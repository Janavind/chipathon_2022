magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< metal1 >>
rect 78 0 114 50560
rect 150 0 186 50560
rect 222 49849 258 50481
rect 222 49059 258 49691
rect 222 48269 258 48901
rect 222 47479 258 48111
rect 222 46689 258 47321
rect 222 45899 258 46531
rect 222 45109 258 45741
rect 222 44319 258 44951
rect 222 43529 258 44161
rect 222 42739 258 43371
rect 222 41949 258 42581
rect 222 41159 258 41791
rect 222 40369 258 41001
rect 222 39579 258 40211
rect 222 38789 258 39421
rect 222 37999 258 38631
rect 222 37209 258 37841
rect 222 36419 258 37051
rect 222 35629 258 36261
rect 222 34839 258 35471
rect 222 34049 258 34681
rect 222 33259 258 33891
rect 222 32469 258 33101
rect 222 31679 258 32311
rect 222 30889 258 31521
rect 222 30099 258 30731
rect 222 29309 258 29941
rect 222 28519 258 29151
rect 222 27729 258 28361
rect 222 26939 258 27571
rect 222 26149 258 26781
rect 222 25359 258 25991
rect 222 24569 258 25201
rect 222 23779 258 24411
rect 222 22989 258 23621
rect 222 22199 258 22831
rect 222 21409 258 22041
rect 222 20619 258 21251
rect 222 19829 258 20461
rect 222 19039 258 19671
rect 222 18249 258 18881
rect 222 17459 258 18091
rect 222 16669 258 17301
rect 222 15879 258 16511
rect 222 15089 258 15721
rect 222 14299 258 14931
rect 222 13509 258 14141
rect 222 12719 258 13351
rect 222 11929 258 12561
rect 222 11139 258 11771
rect 222 10349 258 10981
rect 222 9559 258 10191
rect 222 8769 258 9401
rect 222 7979 258 8611
rect 222 7189 258 7821
rect 222 6399 258 7031
rect 222 5609 258 6241
rect 222 4819 258 5451
rect 222 4029 258 4661
rect 222 3239 258 3871
rect 222 2449 258 3081
rect 222 1659 258 2291
rect 222 869 258 1501
rect 222 79 258 711
rect 294 0 330 50560
rect 366 0 402 50560
rect 846 0 882 50560
rect 918 0 954 50560
rect 990 49849 1026 50481
rect 990 49059 1026 49691
rect 990 48269 1026 48901
rect 990 47479 1026 48111
rect 990 46689 1026 47321
rect 990 45899 1026 46531
rect 990 45109 1026 45741
rect 990 44319 1026 44951
rect 990 43529 1026 44161
rect 990 42739 1026 43371
rect 990 41949 1026 42581
rect 990 41159 1026 41791
rect 990 40369 1026 41001
rect 990 39579 1026 40211
rect 990 38789 1026 39421
rect 990 37999 1026 38631
rect 990 37209 1026 37841
rect 990 36419 1026 37051
rect 990 35629 1026 36261
rect 990 34839 1026 35471
rect 990 34049 1026 34681
rect 990 33259 1026 33891
rect 990 32469 1026 33101
rect 990 31679 1026 32311
rect 990 30889 1026 31521
rect 990 30099 1026 30731
rect 990 29309 1026 29941
rect 990 28519 1026 29151
rect 990 27729 1026 28361
rect 990 26939 1026 27571
rect 990 26149 1026 26781
rect 990 25359 1026 25991
rect 990 24569 1026 25201
rect 990 23779 1026 24411
rect 990 22989 1026 23621
rect 990 22199 1026 22831
rect 990 21409 1026 22041
rect 990 20619 1026 21251
rect 990 19829 1026 20461
rect 990 19039 1026 19671
rect 990 18249 1026 18881
rect 990 17459 1026 18091
rect 990 16669 1026 17301
rect 990 15879 1026 16511
rect 990 15089 1026 15721
rect 990 14299 1026 14931
rect 990 13509 1026 14141
rect 990 12719 1026 13351
rect 990 11929 1026 12561
rect 990 11139 1026 11771
rect 990 10349 1026 10981
rect 990 9559 1026 10191
rect 990 8769 1026 9401
rect 990 7979 1026 8611
rect 990 7189 1026 7821
rect 990 6399 1026 7031
rect 990 5609 1026 6241
rect 990 4819 1026 5451
rect 990 4029 1026 4661
rect 990 3239 1026 3871
rect 990 2449 1026 3081
rect 990 1659 1026 2291
rect 990 869 1026 1501
rect 990 79 1026 711
rect 1062 0 1098 50560
rect 1134 0 1170 50560
rect 1326 0 1362 50560
rect 1398 0 1434 50560
rect 1470 49849 1506 50481
rect 1470 49059 1506 49691
rect 1470 48269 1506 48901
rect 1470 47479 1506 48111
rect 1470 46689 1506 47321
rect 1470 45899 1506 46531
rect 1470 45109 1506 45741
rect 1470 44319 1506 44951
rect 1470 43529 1506 44161
rect 1470 42739 1506 43371
rect 1470 41949 1506 42581
rect 1470 41159 1506 41791
rect 1470 40369 1506 41001
rect 1470 39579 1506 40211
rect 1470 38789 1506 39421
rect 1470 37999 1506 38631
rect 1470 37209 1506 37841
rect 1470 36419 1506 37051
rect 1470 35629 1506 36261
rect 1470 34839 1506 35471
rect 1470 34049 1506 34681
rect 1470 33259 1506 33891
rect 1470 32469 1506 33101
rect 1470 31679 1506 32311
rect 1470 30889 1506 31521
rect 1470 30099 1506 30731
rect 1470 29309 1506 29941
rect 1470 28519 1506 29151
rect 1470 27729 1506 28361
rect 1470 26939 1506 27571
rect 1470 26149 1506 26781
rect 1470 25359 1506 25991
rect 1470 24569 1506 25201
rect 1470 23779 1506 24411
rect 1470 22989 1506 23621
rect 1470 22199 1506 22831
rect 1470 21409 1506 22041
rect 1470 20619 1506 21251
rect 1470 19829 1506 20461
rect 1470 19039 1506 19671
rect 1470 18249 1506 18881
rect 1470 17459 1506 18091
rect 1470 16669 1506 17301
rect 1470 15879 1506 16511
rect 1470 15089 1506 15721
rect 1470 14299 1506 14931
rect 1470 13509 1506 14141
rect 1470 12719 1506 13351
rect 1470 11929 1506 12561
rect 1470 11139 1506 11771
rect 1470 10349 1506 10981
rect 1470 9559 1506 10191
rect 1470 8769 1506 9401
rect 1470 7979 1506 8611
rect 1470 7189 1506 7821
rect 1470 6399 1506 7031
rect 1470 5609 1506 6241
rect 1470 4819 1506 5451
rect 1470 4029 1506 4661
rect 1470 3239 1506 3871
rect 1470 2449 1506 3081
rect 1470 1659 1506 2291
rect 1470 869 1506 1501
rect 1470 79 1506 711
rect 1542 0 1578 50560
rect 1614 0 1650 50560
rect 2094 0 2130 50560
rect 2166 0 2202 50560
rect 2238 49849 2274 50481
rect 2238 49059 2274 49691
rect 2238 48269 2274 48901
rect 2238 47479 2274 48111
rect 2238 46689 2274 47321
rect 2238 45899 2274 46531
rect 2238 45109 2274 45741
rect 2238 44319 2274 44951
rect 2238 43529 2274 44161
rect 2238 42739 2274 43371
rect 2238 41949 2274 42581
rect 2238 41159 2274 41791
rect 2238 40369 2274 41001
rect 2238 39579 2274 40211
rect 2238 38789 2274 39421
rect 2238 37999 2274 38631
rect 2238 37209 2274 37841
rect 2238 36419 2274 37051
rect 2238 35629 2274 36261
rect 2238 34839 2274 35471
rect 2238 34049 2274 34681
rect 2238 33259 2274 33891
rect 2238 32469 2274 33101
rect 2238 31679 2274 32311
rect 2238 30889 2274 31521
rect 2238 30099 2274 30731
rect 2238 29309 2274 29941
rect 2238 28519 2274 29151
rect 2238 27729 2274 28361
rect 2238 26939 2274 27571
rect 2238 26149 2274 26781
rect 2238 25359 2274 25991
rect 2238 24569 2274 25201
rect 2238 23779 2274 24411
rect 2238 22989 2274 23621
rect 2238 22199 2274 22831
rect 2238 21409 2274 22041
rect 2238 20619 2274 21251
rect 2238 19829 2274 20461
rect 2238 19039 2274 19671
rect 2238 18249 2274 18881
rect 2238 17459 2274 18091
rect 2238 16669 2274 17301
rect 2238 15879 2274 16511
rect 2238 15089 2274 15721
rect 2238 14299 2274 14931
rect 2238 13509 2274 14141
rect 2238 12719 2274 13351
rect 2238 11929 2274 12561
rect 2238 11139 2274 11771
rect 2238 10349 2274 10981
rect 2238 9559 2274 10191
rect 2238 8769 2274 9401
rect 2238 7979 2274 8611
rect 2238 7189 2274 7821
rect 2238 6399 2274 7031
rect 2238 5609 2274 6241
rect 2238 4819 2274 5451
rect 2238 4029 2274 4661
rect 2238 3239 2274 3871
rect 2238 2449 2274 3081
rect 2238 1659 2274 2291
rect 2238 869 2274 1501
rect 2238 79 2274 711
rect 2310 0 2346 50560
rect 2382 0 2418 50560
rect 2574 0 2610 50560
rect 2646 0 2682 50560
rect 2718 49849 2754 50481
rect 2718 49059 2754 49691
rect 2718 48269 2754 48901
rect 2718 47479 2754 48111
rect 2718 46689 2754 47321
rect 2718 45899 2754 46531
rect 2718 45109 2754 45741
rect 2718 44319 2754 44951
rect 2718 43529 2754 44161
rect 2718 42739 2754 43371
rect 2718 41949 2754 42581
rect 2718 41159 2754 41791
rect 2718 40369 2754 41001
rect 2718 39579 2754 40211
rect 2718 38789 2754 39421
rect 2718 37999 2754 38631
rect 2718 37209 2754 37841
rect 2718 36419 2754 37051
rect 2718 35629 2754 36261
rect 2718 34839 2754 35471
rect 2718 34049 2754 34681
rect 2718 33259 2754 33891
rect 2718 32469 2754 33101
rect 2718 31679 2754 32311
rect 2718 30889 2754 31521
rect 2718 30099 2754 30731
rect 2718 29309 2754 29941
rect 2718 28519 2754 29151
rect 2718 27729 2754 28361
rect 2718 26939 2754 27571
rect 2718 26149 2754 26781
rect 2718 25359 2754 25991
rect 2718 24569 2754 25201
rect 2718 23779 2754 24411
rect 2718 22989 2754 23621
rect 2718 22199 2754 22831
rect 2718 21409 2754 22041
rect 2718 20619 2754 21251
rect 2718 19829 2754 20461
rect 2718 19039 2754 19671
rect 2718 18249 2754 18881
rect 2718 17459 2754 18091
rect 2718 16669 2754 17301
rect 2718 15879 2754 16511
rect 2718 15089 2754 15721
rect 2718 14299 2754 14931
rect 2718 13509 2754 14141
rect 2718 12719 2754 13351
rect 2718 11929 2754 12561
rect 2718 11139 2754 11771
rect 2718 10349 2754 10981
rect 2718 9559 2754 10191
rect 2718 8769 2754 9401
rect 2718 7979 2754 8611
rect 2718 7189 2754 7821
rect 2718 6399 2754 7031
rect 2718 5609 2754 6241
rect 2718 4819 2754 5451
rect 2718 4029 2754 4661
rect 2718 3239 2754 3871
rect 2718 2449 2754 3081
rect 2718 1659 2754 2291
rect 2718 869 2754 1501
rect 2718 79 2754 711
rect 2790 0 2826 50560
rect 2862 0 2898 50560
rect 3342 0 3378 50560
rect 3414 0 3450 50560
rect 3486 49849 3522 50481
rect 3486 49059 3522 49691
rect 3486 48269 3522 48901
rect 3486 47479 3522 48111
rect 3486 46689 3522 47321
rect 3486 45899 3522 46531
rect 3486 45109 3522 45741
rect 3486 44319 3522 44951
rect 3486 43529 3522 44161
rect 3486 42739 3522 43371
rect 3486 41949 3522 42581
rect 3486 41159 3522 41791
rect 3486 40369 3522 41001
rect 3486 39579 3522 40211
rect 3486 38789 3522 39421
rect 3486 37999 3522 38631
rect 3486 37209 3522 37841
rect 3486 36419 3522 37051
rect 3486 35629 3522 36261
rect 3486 34839 3522 35471
rect 3486 34049 3522 34681
rect 3486 33259 3522 33891
rect 3486 32469 3522 33101
rect 3486 31679 3522 32311
rect 3486 30889 3522 31521
rect 3486 30099 3522 30731
rect 3486 29309 3522 29941
rect 3486 28519 3522 29151
rect 3486 27729 3522 28361
rect 3486 26939 3522 27571
rect 3486 26149 3522 26781
rect 3486 25359 3522 25991
rect 3486 24569 3522 25201
rect 3486 23779 3522 24411
rect 3486 22989 3522 23621
rect 3486 22199 3522 22831
rect 3486 21409 3522 22041
rect 3486 20619 3522 21251
rect 3486 19829 3522 20461
rect 3486 19039 3522 19671
rect 3486 18249 3522 18881
rect 3486 17459 3522 18091
rect 3486 16669 3522 17301
rect 3486 15879 3522 16511
rect 3486 15089 3522 15721
rect 3486 14299 3522 14931
rect 3486 13509 3522 14141
rect 3486 12719 3522 13351
rect 3486 11929 3522 12561
rect 3486 11139 3522 11771
rect 3486 10349 3522 10981
rect 3486 9559 3522 10191
rect 3486 8769 3522 9401
rect 3486 7979 3522 8611
rect 3486 7189 3522 7821
rect 3486 6399 3522 7031
rect 3486 5609 3522 6241
rect 3486 4819 3522 5451
rect 3486 4029 3522 4661
rect 3486 3239 3522 3871
rect 3486 2449 3522 3081
rect 3486 1659 3522 2291
rect 3486 869 3522 1501
rect 3486 79 3522 711
rect 3558 0 3594 50560
rect 3630 0 3666 50560
rect 3822 0 3858 50560
rect 3894 0 3930 50560
rect 3966 49849 4002 50481
rect 3966 49059 4002 49691
rect 3966 48269 4002 48901
rect 3966 47479 4002 48111
rect 3966 46689 4002 47321
rect 3966 45899 4002 46531
rect 3966 45109 4002 45741
rect 3966 44319 4002 44951
rect 3966 43529 4002 44161
rect 3966 42739 4002 43371
rect 3966 41949 4002 42581
rect 3966 41159 4002 41791
rect 3966 40369 4002 41001
rect 3966 39579 4002 40211
rect 3966 38789 4002 39421
rect 3966 37999 4002 38631
rect 3966 37209 4002 37841
rect 3966 36419 4002 37051
rect 3966 35629 4002 36261
rect 3966 34839 4002 35471
rect 3966 34049 4002 34681
rect 3966 33259 4002 33891
rect 3966 32469 4002 33101
rect 3966 31679 4002 32311
rect 3966 30889 4002 31521
rect 3966 30099 4002 30731
rect 3966 29309 4002 29941
rect 3966 28519 4002 29151
rect 3966 27729 4002 28361
rect 3966 26939 4002 27571
rect 3966 26149 4002 26781
rect 3966 25359 4002 25991
rect 3966 24569 4002 25201
rect 3966 23779 4002 24411
rect 3966 22989 4002 23621
rect 3966 22199 4002 22831
rect 3966 21409 4002 22041
rect 3966 20619 4002 21251
rect 3966 19829 4002 20461
rect 3966 19039 4002 19671
rect 3966 18249 4002 18881
rect 3966 17459 4002 18091
rect 3966 16669 4002 17301
rect 3966 15879 4002 16511
rect 3966 15089 4002 15721
rect 3966 14299 4002 14931
rect 3966 13509 4002 14141
rect 3966 12719 4002 13351
rect 3966 11929 4002 12561
rect 3966 11139 4002 11771
rect 3966 10349 4002 10981
rect 3966 9559 4002 10191
rect 3966 8769 4002 9401
rect 3966 7979 4002 8611
rect 3966 7189 4002 7821
rect 3966 6399 4002 7031
rect 3966 5609 4002 6241
rect 3966 4819 4002 5451
rect 3966 4029 4002 4661
rect 3966 3239 4002 3871
rect 3966 2449 4002 3081
rect 3966 1659 4002 2291
rect 3966 869 4002 1501
rect 3966 79 4002 711
rect 4038 0 4074 50560
rect 4110 0 4146 50560
rect 4590 0 4626 50560
rect 4662 0 4698 50560
rect 4734 49849 4770 50481
rect 4734 49059 4770 49691
rect 4734 48269 4770 48901
rect 4734 47479 4770 48111
rect 4734 46689 4770 47321
rect 4734 45899 4770 46531
rect 4734 45109 4770 45741
rect 4734 44319 4770 44951
rect 4734 43529 4770 44161
rect 4734 42739 4770 43371
rect 4734 41949 4770 42581
rect 4734 41159 4770 41791
rect 4734 40369 4770 41001
rect 4734 39579 4770 40211
rect 4734 38789 4770 39421
rect 4734 37999 4770 38631
rect 4734 37209 4770 37841
rect 4734 36419 4770 37051
rect 4734 35629 4770 36261
rect 4734 34839 4770 35471
rect 4734 34049 4770 34681
rect 4734 33259 4770 33891
rect 4734 32469 4770 33101
rect 4734 31679 4770 32311
rect 4734 30889 4770 31521
rect 4734 30099 4770 30731
rect 4734 29309 4770 29941
rect 4734 28519 4770 29151
rect 4734 27729 4770 28361
rect 4734 26939 4770 27571
rect 4734 26149 4770 26781
rect 4734 25359 4770 25991
rect 4734 24569 4770 25201
rect 4734 23779 4770 24411
rect 4734 22989 4770 23621
rect 4734 22199 4770 22831
rect 4734 21409 4770 22041
rect 4734 20619 4770 21251
rect 4734 19829 4770 20461
rect 4734 19039 4770 19671
rect 4734 18249 4770 18881
rect 4734 17459 4770 18091
rect 4734 16669 4770 17301
rect 4734 15879 4770 16511
rect 4734 15089 4770 15721
rect 4734 14299 4770 14931
rect 4734 13509 4770 14141
rect 4734 12719 4770 13351
rect 4734 11929 4770 12561
rect 4734 11139 4770 11771
rect 4734 10349 4770 10981
rect 4734 9559 4770 10191
rect 4734 8769 4770 9401
rect 4734 7979 4770 8611
rect 4734 7189 4770 7821
rect 4734 6399 4770 7031
rect 4734 5609 4770 6241
rect 4734 4819 4770 5451
rect 4734 4029 4770 4661
rect 4734 3239 4770 3871
rect 4734 2449 4770 3081
rect 4734 1659 4770 2291
rect 4734 869 4770 1501
rect 4734 79 4770 711
rect 4806 0 4842 50560
rect 4878 0 4914 50560
rect 5070 0 5106 50560
rect 5142 0 5178 50560
rect 5214 49849 5250 50481
rect 5214 49059 5250 49691
rect 5214 48269 5250 48901
rect 5214 47479 5250 48111
rect 5214 46689 5250 47321
rect 5214 45899 5250 46531
rect 5214 45109 5250 45741
rect 5214 44319 5250 44951
rect 5214 43529 5250 44161
rect 5214 42739 5250 43371
rect 5214 41949 5250 42581
rect 5214 41159 5250 41791
rect 5214 40369 5250 41001
rect 5214 39579 5250 40211
rect 5214 38789 5250 39421
rect 5214 37999 5250 38631
rect 5214 37209 5250 37841
rect 5214 36419 5250 37051
rect 5214 35629 5250 36261
rect 5214 34839 5250 35471
rect 5214 34049 5250 34681
rect 5214 33259 5250 33891
rect 5214 32469 5250 33101
rect 5214 31679 5250 32311
rect 5214 30889 5250 31521
rect 5214 30099 5250 30731
rect 5214 29309 5250 29941
rect 5214 28519 5250 29151
rect 5214 27729 5250 28361
rect 5214 26939 5250 27571
rect 5214 26149 5250 26781
rect 5214 25359 5250 25991
rect 5214 24569 5250 25201
rect 5214 23779 5250 24411
rect 5214 22989 5250 23621
rect 5214 22199 5250 22831
rect 5214 21409 5250 22041
rect 5214 20619 5250 21251
rect 5214 19829 5250 20461
rect 5214 19039 5250 19671
rect 5214 18249 5250 18881
rect 5214 17459 5250 18091
rect 5214 16669 5250 17301
rect 5214 15879 5250 16511
rect 5214 15089 5250 15721
rect 5214 14299 5250 14931
rect 5214 13509 5250 14141
rect 5214 12719 5250 13351
rect 5214 11929 5250 12561
rect 5214 11139 5250 11771
rect 5214 10349 5250 10981
rect 5214 9559 5250 10191
rect 5214 8769 5250 9401
rect 5214 7979 5250 8611
rect 5214 7189 5250 7821
rect 5214 6399 5250 7031
rect 5214 5609 5250 6241
rect 5214 4819 5250 5451
rect 5214 4029 5250 4661
rect 5214 3239 5250 3871
rect 5214 2449 5250 3081
rect 5214 1659 5250 2291
rect 5214 869 5250 1501
rect 5214 79 5250 711
rect 5286 0 5322 50560
rect 5358 0 5394 50560
rect 5838 0 5874 50560
rect 5910 0 5946 50560
rect 5982 49849 6018 50481
rect 5982 49059 6018 49691
rect 5982 48269 6018 48901
rect 5982 47479 6018 48111
rect 5982 46689 6018 47321
rect 5982 45899 6018 46531
rect 5982 45109 6018 45741
rect 5982 44319 6018 44951
rect 5982 43529 6018 44161
rect 5982 42739 6018 43371
rect 5982 41949 6018 42581
rect 5982 41159 6018 41791
rect 5982 40369 6018 41001
rect 5982 39579 6018 40211
rect 5982 38789 6018 39421
rect 5982 37999 6018 38631
rect 5982 37209 6018 37841
rect 5982 36419 6018 37051
rect 5982 35629 6018 36261
rect 5982 34839 6018 35471
rect 5982 34049 6018 34681
rect 5982 33259 6018 33891
rect 5982 32469 6018 33101
rect 5982 31679 6018 32311
rect 5982 30889 6018 31521
rect 5982 30099 6018 30731
rect 5982 29309 6018 29941
rect 5982 28519 6018 29151
rect 5982 27729 6018 28361
rect 5982 26939 6018 27571
rect 5982 26149 6018 26781
rect 5982 25359 6018 25991
rect 5982 24569 6018 25201
rect 5982 23779 6018 24411
rect 5982 22989 6018 23621
rect 5982 22199 6018 22831
rect 5982 21409 6018 22041
rect 5982 20619 6018 21251
rect 5982 19829 6018 20461
rect 5982 19039 6018 19671
rect 5982 18249 6018 18881
rect 5982 17459 6018 18091
rect 5982 16669 6018 17301
rect 5982 15879 6018 16511
rect 5982 15089 6018 15721
rect 5982 14299 6018 14931
rect 5982 13509 6018 14141
rect 5982 12719 6018 13351
rect 5982 11929 6018 12561
rect 5982 11139 6018 11771
rect 5982 10349 6018 10981
rect 5982 9559 6018 10191
rect 5982 8769 6018 9401
rect 5982 7979 6018 8611
rect 5982 7189 6018 7821
rect 5982 6399 6018 7031
rect 5982 5609 6018 6241
rect 5982 4819 6018 5451
rect 5982 4029 6018 4661
rect 5982 3239 6018 3871
rect 5982 2449 6018 3081
rect 5982 1659 6018 2291
rect 5982 869 6018 1501
rect 5982 79 6018 711
rect 6054 0 6090 50560
rect 6126 0 6162 50560
rect 6318 0 6354 50560
rect 6390 0 6426 50560
rect 6462 49849 6498 50481
rect 6462 49059 6498 49691
rect 6462 48269 6498 48901
rect 6462 47479 6498 48111
rect 6462 46689 6498 47321
rect 6462 45899 6498 46531
rect 6462 45109 6498 45741
rect 6462 44319 6498 44951
rect 6462 43529 6498 44161
rect 6462 42739 6498 43371
rect 6462 41949 6498 42581
rect 6462 41159 6498 41791
rect 6462 40369 6498 41001
rect 6462 39579 6498 40211
rect 6462 38789 6498 39421
rect 6462 37999 6498 38631
rect 6462 37209 6498 37841
rect 6462 36419 6498 37051
rect 6462 35629 6498 36261
rect 6462 34839 6498 35471
rect 6462 34049 6498 34681
rect 6462 33259 6498 33891
rect 6462 32469 6498 33101
rect 6462 31679 6498 32311
rect 6462 30889 6498 31521
rect 6462 30099 6498 30731
rect 6462 29309 6498 29941
rect 6462 28519 6498 29151
rect 6462 27729 6498 28361
rect 6462 26939 6498 27571
rect 6462 26149 6498 26781
rect 6462 25359 6498 25991
rect 6462 24569 6498 25201
rect 6462 23779 6498 24411
rect 6462 22989 6498 23621
rect 6462 22199 6498 22831
rect 6462 21409 6498 22041
rect 6462 20619 6498 21251
rect 6462 19829 6498 20461
rect 6462 19039 6498 19671
rect 6462 18249 6498 18881
rect 6462 17459 6498 18091
rect 6462 16669 6498 17301
rect 6462 15879 6498 16511
rect 6462 15089 6498 15721
rect 6462 14299 6498 14931
rect 6462 13509 6498 14141
rect 6462 12719 6498 13351
rect 6462 11929 6498 12561
rect 6462 11139 6498 11771
rect 6462 10349 6498 10981
rect 6462 9559 6498 10191
rect 6462 8769 6498 9401
rect 6462 7979 6498 8611
rect 6462 7189 6498 7821
rect 6462 6399 6498 7031
rect 6462 5609 6498 6241
rect 6462 4819 6498 5451
rect 6462 4029 6498 4661
rect 6462 3239 6498 3871
rect 6462 2449 6498 3081
rect 6462 1659 6498 2291
rect 6462 869 6498 1501
rect 6462 79 6498 711
rect 6534 0 6570 50560
rect 6606 0 6642 50560
rect 7086 0 7122 50560
rect 7158 0 7194 50560
rect 7230 49849 7266 50481
rect 7230 49059 7266 49691
rect 7230 48269 7266 48901
rect 7230 47479 7266 48111
rect 7230 46689 7266 47321
rect 7230 45899 7266 46531
rect 7230 45109 7266 45741
rect 7230 44319 7266 44951
rect 7230 43529 7266 44161
rect 7230 42739 7266 43371
rect 7230 41949 7266 42581
rect 7230 41159 7266 41791
rect 7230 40369 7266 41001
rect 7230 39579 7266 40211
rect 7230 38789 7266 39421
rect 7230 37999 7266 38631
rect 7230 37209 7266 37841
rect 7230 36419 7266 37051
rect 7230 35629 7266 36261
rect 7230 34839 7266 35471
rect 7230 34049 7266 34681
rect 7230 33259 7266 33891
rect 7230 32469 7266 33101
rect 7230 31679 7266 32311
rect 7230 30889 7266 31521
rect 7230 30099 7266 30731
rect 7230 29309 7266 29941
rect 7230 28519 7266 29151
rect 7230 27729 7266 28361
rect 7230 26939 7266 27571
rect 7230 26149 7266 26781
rect 7230 25359 7266 25991
rect 7230 24569 7266 25201
rect 7230 23779 7266 24411
rect 7230 22989 7266 23621
rect 7230 22199 7266 22831
rect 7230 21409 7266 22041
rect 7230 20619 7266 21251
rect 7230 19829 7266 20461
rect 7230 19039 7266 19671
rect 7230 18249 7266 18881
rect 7230 17459 7266 18091
rect 7230 16669 7266 17301
rect 7230 15879 7266 16511
rect 7230 15089 7266 15721
rect 7230 14299 7266 14931
rect 7230 13509 7266 14141
rect 7230 12719 7266 13351
rect 7230 11929 7266 12561
rect 7230 11139 7266 11771
rect 7230 10349 7266 10981
rect 7230 9559 7266 10191
rect 7230 8769 7266 9401
rect 7230 7979 7266 8611
rect 7230 7189 7266 7821
rect 7230 6399 7266 7031
rect 7230 5609 7266 6241
rect 7230 4819 7266 5451
rect 7230 4029 7266 4661
rect 7230 3239 7266 3871
rect 7230 2449 7266 3081
rect 7230 1659 7266 2291
rect 7230 869 7266 1501
rect 7230 79 7266 711
rect 7302 0 7338 50560
rect 7374 0 7410 50560
rect 7566 0 7602 50560
rect 7638 0 7674 50560
rect 7710 49849 7746 50481
rect 7710 49059 7746 49691
rect 7710 48269 7746 48901
rect 7710 47479 7746 48111
rect 7710 46689 7746 47321
rect 7710 45899 7746 46531
rect 7710 45109 7746 45741
rect 7710 44319 7746 44951
rect 7710 43529 7746 44161
rect 7710 42739 7746 43371
rect 7710 41949 7746 42581
rect 7710 41159 7746 41791
rect 7710 40369 7746 41001
rect 7710 39579 7746 40211
rect 7710 38789 7746 39421
rect 7710 37999 7746 38631
rect 7710 37209 7746 37841
rect 7710 36419 7746 37051
rect 7710 35629 7746 36261
rect 7710 34839 7746 35471
rect 7710 34049 7746 34681
rect 7710 33259 7746 33891
rect 7710 32469 7746 33101
rect 7710 31679 7746 32311
rect 7710 30889 7746 31521
rect 7710 30099 7746 30731
rect 7710 29309 7746 29941
rect 7710 28519 7746 29151
rect 7710 27729 7746 28361
rect 7710 26939 7746 27571
rect 7710 26149 7746 26781
rect 7710 25359 7746 25991
rect 7710 24569 7746 25201
rect 7710 23779 7746 24411
rect 7710 22989 7746 23621
rect 7710 22199 7746 22831
rect 7710 21409 7746 22041
rect 7710 20619 7746 21251
rect 7710 19829 7746 20461
rect 7710 19039 7746 19671
rect 7710 18249 7746 18881
rect 7710 17459 7746 18091
rect 7710 16669 7746 17301
rect 7710 15879 7746 16511
rect 7710 15089 7746 15721
rect 7710 14299 7746 14931
rect 7710 13509 7746 14141
rect 7710 12719 7746 13351
rect 7710 11929 7746 12561
rect 7710 11139 7746 11771
rect 7710 10349 7746 10981
rect 7710 9559 7746 10191
rect 7710 8769 7746 9401
rect 7710 7979 7746 8611
rect 7710 7189 7746 7821
rect 7710 6399 7746 7031
rect 7710 5609 7746 6241
rect 7710 4819 7746 5451
rect 7710 4029 7746 4661
rect 7710 3239 7746 3871
rect 7710 2449 7746 3081
rect 7710 1659 7746 2291
rect 7710 869 7746 1501
rect 7710 79 7746 711
rect 7782 0 7818 50560
rect 7854 0 7890 50560
rect 8334 0 8370 50560
rect 8406 0 8442 50560
rect 8478 49849 8514 50481
rect 8478 49059 8514 49691
rect 8478 48269 8514 48901
rect 8478 47479 8514 48111
rect 8478 46689 8514 47321
rect 8478 45899 8514 46531
rect 8478 45109 8514 45741
rect 8478 44319 8514 44951
rect 8478 43529 8514 44161
rect 8478 42739 8514 43371
rect 8478 41949 8514 42581
rect 8478 41159 8514 41791
rect 8478 40369 8514 41001
rect 8478 39579 8514 40211
rect 8478 38789 8514 39421
rect 8478 37999 8514 38631
rect 8478 37209 8514 37841
rect 8478 36419 8514 37051
rect 8478 35629 8514 36261
rect 8478 34839 8514 35471
rect 8478 34049 8514 34681
rect 8478 33259 8514 33891
rect 8478 32469 8514 33101
rect 8478 31679 8514 32311
rect 8478 30889 8514 31521
rect 8478 30099 8514 30731
rect 8478 29309 8514 29941
rect 8478 28519 8514 29151
rect 8478 27729 8514 28361
rect 8478 26939 8514 27571
rect 8478 26149 8514 26781
rect 8478 25359 8514 25991
rect 8478 24569 8514 25201
rect 8478 23779 8514 24411
rect 8478 22989 8514 23621
rect 8478 22199 8514 22831
rect 8478 21409 8514 22041
rect 8478 20619 8514 21251
rect 8478 19829 8514 20461
rect 8478 19039 8514 19671
rect 8478 18249 8514 18881
rect 8478 17459 8514 18091
rect 8478 16669 8514 17301
rect 8478 15879 8514 16511
rect 8478 15089 8514 15721
rect 8478 14299 8514 14931
rect 8478 13509 8514 14141
rect 8478 12719 8514 13351
rect 8478 11929 8514 12561
rect 8478 11139 8514 11771
rect 8478 10349 8514 10981
rect 8478 9559 8514 10191
rect 8478 8769 8514 9401
rect 8478 7979 8514 8611
rect 8478 7189 8514 7821
rect 8478 6399 8514 7031
rect 8478 5609 8514 6241
rect 8478 4819 8514 5451
rect 8478 4029 8514 4661
rect 8478 3239 8514 3871
rect 8478 2449 8514 3081
rect 8478 1659 8514 2291
rect 8478 869 8514 1501
rect 8478 79 8514 711
rect 8550 0 8586 50560
rect 8622 0 8658 50560
rect 8814 0 8850 50560
rect 8886 0 8922 50560
rect 8958 49849 8994 50481
rect 8958 49059 8994 49691
rect 8958 48269 8994 48901
rect 8958 47479 8994 48111
rect 8958 46689 8994 47321
rect 8958 45899 8994 46531
rect 8958 45109 8994 45741
rect 8958 44319 8994 44951
rect 8958 43529 8994 44161
rect 8958 42739 8994 43371
rect 8958 41949 8994 42581
rect 8958 41159 8994 41791
rect 8958 40369 8994 41001
rect 8958 39579 8994 40211
rect 8958 38789 8994 39421
rect 8958 37999 8994 38631
rect 8958 37209 8994 37841
rect 8958 36419 8994 37051
rect 8958 35629 8994 36261
rect 8958 34839 8994 35471
rect 8958 34049 8994 34681
rect 8958 33259 8994 33891
rect 8958 32469 8994 33101
rect 8958 31679 8994 32311
rect 8958 30889 8994 31521
rect 8958 30099 8994 30731
rect 8958 29309 8994 29941
rect 8958 28519 8994 29151
rect 8958 27729 8994 28361
rect 8958 26939 8994 27571
rect 8958 26149 8994 26781
rect 8958 25359 8994 25991
rect 8958 24569 8994 25201
rect 8958 23779 8994 24411
rect 8958 22989 8994 23621
rect 8958 22199 8994 22831
rect 8958 21409 8994 22041
rect 8958 20619 8994 21251
rect 8958 19829 8994 20461
rect 8958 19039 8994 19671
rect 8958 18249 8994 18881
rect 8958 17459 8994 18091
rect 8958 16669 8994 17301
rect 8958 15879 8994 16511
rect 8958 15089 8994 15721
rect 8958 14299 8994 14931
rect 8958 13509 8994 14141
rect 8958 12719 8994 13351
rect 8958 11929 8994 12561
rect 8958 11139 8994 11771
rect 8958 10349 8994 10981
rect 8958 9559 8994 10191
rect 8958 8769 8994 9401
rect 8958 7979 8994 8611
rect 8958 7189 8994 7821
rect 8958 6399 8994 7031
rect 8958 5609 8994 6241
rect 8958 4819 8994 5451
rect 8958 4029 8994 4661
rect 8958 3239 8994 3871
rect 8958 2449 8994 3081
rect 8958 1659 8994 2291
rect 8958 869 8994 1501
rect 8958 79 8994 711
rect 9030 0 9066 50560
rect 9102 0 9138 50560
rect 9582 0 9618 50560
rect 9654 0 9690 50560
rect 9726 49849 9762 50481
rect 9726 49059 9762 49691
rect 9726 48269 9762 48901
rect 9726 47479 9762 48111
rect 9726 46689 9762 47321
rect 9726 45899 9762 46531
rect 9726 45109 9762 45741
rect 9726 44319 9762 44951
rect 9726 43529 9762 44161
rect 9726 42739 9762 43371
rect 9726 41949 9762 42581
rect 9726 41159 9762 41791
rect 9726 40369 9762 41001
rect 9726 39579 9762 40211
rect 9726 38789 9762 39421
rect 9726 37999 9762 38631
rect 9726 37209 9762 37841
rect 9726 36419 9762 37051
rect 9726 35629 9762 36261
rect 9726 34839 9762 35471
rect 9726 34049 9762 34681
rect 9726 33259 9762 33891
rect 9726 32469 9762 33101
rect 9726 31679 9762 32311
rect 9726 30889 9762 31521
rect 9726 30099 9762 30731
rect 9726 29309 9762 29941
rect 9726 28519 9762 29151
rect 9726 27729 9762 28361
rect 9726 26939 9762 27571
rect 9726 26149 9762 26781
rect 9726 25359 9762 25991
rect 9726 24569 9762 25201
rect 9726 23779 9762 24411
rect 9726 22989 9762 23621
rect 9726 22199 9762 22831
rect 9726 21409 9762 22041
rect 9726 20619 9762 21251
rect 9726 19829 9762 20461
rect 9726 19039 9762 19671
rect 9726 18249 9762 18881
rect 9726 17459 9762 18091
rect 9726 16669 9762 17301
rect 9726 15879 9762 16511
rect 9726 15089 9762 15721
rect 9726 14299 9762 14931
rect 9726 13509 9762 14141
rect 9726 12719 9762 13351
rect 9726 11929 9762 12561
rect 9726 11139 9762 11771
rect 9726 10349 9762 10981
rect 9726 9559 9762 10191
rect 9726 8769 9762 9401
rect 9726 7979 9762 8611
rect 9726 7189 9762 7821
rect 9726 6399 9762 7031
rect 9726 5609 9762 6241
rect 9726 4819 9762 5451
rect 9726 4029 9762 4661
rect 9726 3239 9762 3871
rect 9726 2449 9762 3081
rect 9726 1659 9762 2291
rect 9726 869 9762 1501
rect 9726 79 9762 711
rect 9798 0 9834 50560
rect 9870 0 9906 50560
rect 10062 0 10098 50560
rect 10134 0 10170 50560
rect 10206 49849 10242 50481
rect 10206 49059 10242 49691
rect 10206 48269 10242 48901
rect 10206 47479 10242 48111
rect 10206 46689 10242 47321
rect 10206 45899 10242 46531
rect 10206 45109 10242 45741
rect 10206 44319 10242 44951
rect 10206 43529 10242 44161
rect 10206 42739 10242 43371
rect 10206 41949 10242 42581
rect 10206 41159 10242 41791
rect 10206 40369 10242 41001
rect 10206 39579 10242 40211
rect 10206 38789 10242 39421
rect 10206 37999 10242 38631
rect 10206 37209 10242 37841
rect 10206 36419 10242 37051
rect 10206 35629 10242 36261
rect 10206 34839 10242 35471
rect 10206 34049 10242 34681
rect 10206 33259 10242 33891
rect 10206 32469 10242 33101
rect 10206 31679 10242 32311
rect 10206 30889 10242 31521
rect 10206 30099 10242 30731
rect 10206 29309 10242 29941
rect 10206 28519 10242 29151
rect 10206 27729 10242 28361
rect 10206 26939 10242 27571
rect 10206 26149 10242 26781
rect 10206 25359 10242 25991
rect 10206 24569 10242 25201
rect 10206 23779 10242 24411
rect 10206 22989 10242 23621
rect 10206 22199 10242 22831
rect 10206 21409 10242 22041
rect 10206 20619 10242 21251
rect 10206 19829 10242 20461
rect 10206 19039 10242 19671
rect 10206 18249 10242 18881
rect 10206 17459 10242 18091
rect 10206 16669 10242 17301
rect 10206 15879 10242 16511
rect 10206 15089 10242 15721
rect 10206 14299 10242 14931
rect 10206 13509 10242 14141
rect 10206 12719 10242 13351
rect 10206 11929 10242 12561
rect 10206 11139 10242 11771
rect 10206 10349 10242 10981
rect 10206 9559 10242 10191
rect 10206 8769 10242 9401
rect 10206 7979 10242 8611
rect 10206 7189 10242 7821
rect 10206 6399 10242 7031
rect 10206 5609 10242 6241
rect 10206 4819 10242 5451
rect 10206 4029 10242 4661
rect 10206 3239 10242 3871
rect 10206 2449 10242 3081
rect 10206 1659 10242 2291
rect 10206 869 10242 1501
rect 10206 79 10242 711
rect 10278 0 10314 50560
rect 10350 0 10386 50560
rect 10830 0 10866 50560
rect 10902 0 10938 50560
rect 10974 49849 11010 50481
rect 10974 49059 11010 49691
rect 10974 48269 11010 48901
rect 10974 47479 11010 48111
rect 10974 46689 11010 47321
rect 10974 45899 11010 46531
rect 10974 45109 11010 45741
rect 10974 44319 11010 44951
rect 10974 43529 11010 44161
rect 10974 42739 11010 43371
rect 10974 41949 11010 42581
rect 10974 41159 11010 41791
rect 10974 40369 11010 41001
rect 10974 39579 11010 40211
rect 10974 38789 11010 39421
rect 10974 37999 11010 38631
rect 10974 37209 11010 37841
rect 10974 36419 11010 37051
rect 10974 35629 11010 36261
rect 10974 34839 11010 35471
rect 10974 34049 11010 34681
rect 10974 33259 11010 33891
rect 10974 32469 11010 33101
rect 10974 31679 11010 32311
rect 10974 30889 11010 31521
rect 10974 30099 11010 30731
rect 10974 29309 11010 29941
rect 10974 28519 11010 29151
rect 10974 27729 11010 28361
rect 10974 26939 11010 27571
rect 10974 26149 11010 26781
rect 10974 25359 11010 25991
rect 10974 24569 11010 25201
rect 10974 23779 11010 24411
rect 10974 22989 11010 23621
rect 10974 22199 11010 22831
rect 10974 21409 11010 22041
rect 10974 20619 11010 21251
rect 10974 19829 11010 20461
rect 10974 19039 11010 19671
rect 10974 18249 11010 18881
rect 10974 17459 11010 18091
rect 10974 16669 11010 17301
rect 10974 15879 11010 16511
rect 10974 15089 11010 15721
rect 10974 14299 11010 14931
rect 10974 13509 11010 14141
rect 10974 12719 11010 13351
rect 10974 11929 11010 12561
rect 10974 11139 11010 11771
rect 10974 10349 11010 10981
rect 10974 9559 11010 10191
rect 10974 8769 11010 9401
rect 10974 7979 11010 8611
rect 10974 7189 11010 7821
rect 10974 6399 11010 7031
rect 10974 5609 11010 6241
rect 10974 4819 11010 5451
rect 10974 4029 11010 4661
rect 10974 3239 11010 3871
rect 10974 2449 11010 3081
rect 10974 1659 11010 2291
rect 10974 869 11010 1501
rect 10974 79 11010 711
rect 11046 0 11082 50560
rect 11118 0 11154 50560
rect 11310 0 11346 50560
rect 11382 0 11418 50560
rect 11454 49849 11490 50481
rect 11454 49059 11490 49691
rect 11454 48269 11490 48901
rect 11454 47479 11490 48111
rect 11454 46689 11490 47321
rect 11454 45899 11490 46531
rect 11454 45109 11490 45741
rect 11454 44319 11490 44951
rect 11454 43529 11490 44161
rect 11454 42739 11490 43371
rect 11454 41949 11490 42581
rect 11454 41159 11490 41791
rect 11454 40369 11490 41001
rect 11454 39579 11490 40211
rect 11454 38789 11490 39421
rect 11454 37999 11490 38631
rect 11454 37209 11490 37841
rect 11454 36419 11490 37051
rect 11454 35629 11490 36261
rect 11454 34839 11490 35471
rect 11454 34049 11490 34681
rect 11454 33259 11490 33891
rect 11454 32469 11490 33101
rect 11454 31679 11490 32311
rect 11454 30889 11490 31521
rect 11454 30099 11490 30731
rect 11454 29309 11490 29941
rect 11454 28519 11490 29151
rect 11454 27729 11490 28361
rect 11454 26939 11490 27571
rect 11454 26149 11490 26781
rect 11454 25359 11490 25991
rect 11454 24569 11490 25201
rect 11454 23779 11490 24411
rect 11454 22989 11490 23621
rect 11454 22199 11490 22831
rect 11454 21409 11490 22041
rect 11454 20619 11490 21251
rect 11454 19829 11490 20461
rect 11454 19039 11490 19671
rect 11454 18249 11490 18881
rect 11454 17459 11490 18091
rect 11454 16669 11490 17301
rect 11454 15879 11490 16511
rect 11454 15089 11490 15721
rect 11454 14299 11490 14931
rect 11454 13509 11490 14141
rect 11454 12719 11490 13351
rect 11454 11929 11490 12561
rect 11454 11139 11490 11771
rect 11454 10349 11490 10981
rect 11454 9559 11490 10191
rect 11454 8769 11490 9401
rect 11454 7979 11490 8611
rect 11454 7189 11490 7821
rect 11454 6399 11490 7031
rect 11454 5609 11490 6241
rect 11454 4819 11490 5451
rect 11454 4029 11490 4661
rect 11454 3239 11490 3871
rect 11454 2449 11490 3081
rect 11454 1659 11490 2291
rect 11454 869 11490 1501
rect 11454 79 11490 711
rect 11526 0 11562 50560
rect 11598 0 11634 50560
rect 12078 0 12114 50560
rect 12150 0 12186 50560
rect 12222 49849 12258 50481
rect 12222 49059 12258 49691
rect 12222 48269 12258 48901
rect 12222 47479 12258 48111
rect 12222 46689 12258 47321
rect 12222 45899 12258 46531
rect 12222 45109 12258 45741
rect 12222 44319 12258 44951
rect 12222 43529 12258 44161
rect 12222 42739 12258 43371
rect 12222 41949 12258 42581
rect 12222 41159 12258 41791
rect 12222 40369 12258 41001
rect 12222 39579 12258 40211
rect 12222 38789 12258 39421
rect 12222 37999 12258 38631
rect 12222 37209 12258 37841
rect 12222 36419 12258 37051
rect 12222 35629 12258 36261
rect 12222 34839 12258 35471
rect 12222 34049 12258 34681
rect 12222 33259 12258 33891
rect 12222 32469 12258 33101
rect 12222 31679 12258 32311
rect 12222 30889 12258 31521
rect 12222 30099 12258 30731
rect 12222 29309 12258 29941
rect 12222 28519 12258 29151
rect 12222 27729 12258 28361
rect 12222 26939 12258 27571
rect 12222 26149 12258 26781
rect 12222 25359 12258 25991
rect 12222 24569 12258 25201
rect 12222 23779 12258 24411
rect 12222 22989 12258 23621
rect 12222 22199 12258 22831
rect 12222 21409 12258 22041
rect 12222 20619 12258 21251
rect 12222 19829 12258 20461
rect 12222 19039 12258 19671
rect 12222 18249 12258 18881
rect 12222 17459 12258 18091
rect 12222 16669 12258 17301
rect 12222 15879 12258 16511
rect 12222 15089 12258 15721
rect 12222 14299 12258 14931
rect 12222 13509 12258 14141
rect 12222 12719 12258 13351
rect 12222 11929 12258 12561
rect 12222 11139 12258 11771
rect 12222 10349 12258 10981
rect 12222 9559 12258 10191
rect 12222 8769 12258 9401
rect 12222 7979 12258 8611
rect 12222 7189 12258 7821
rect 12222 6399 12258 7031
rect 12222 5609 12258 6241
rect 12222 4819 12258 5451
rect 12222 4029 12258 4661
rect 12222 3239 12258 3871
rect 12222 2449 12258 3081
rect 12222 1659 12258 2291
rect 12222 869 12258 1501
rect 12222 79 12258 711
rect 12294 0 12330 50560
rect 12366 0 12402 50560
rect 12558 0 12594 50560
rect 12630 0 12666 50560
rect 12702 49849 12738 50481
rect 12702 49059 12738 49691
rect 12702 48269 12738 48901
rect 12702 47479 12738 48111
rect 12702 46689 12738 47321
rect 12702 45899 12738 46531
rect 12702 45109 12738 45741
rect 12702 44319 12738 44951
rect 12702 43529 12738 44161
rect 12702 42739 12738 43371
rect 12702 41949 12738 42581
rect 12702 41159 12738 41791
rect 12702 40369 12738 41001
rect 12702 39579 12738 40211
rect 12702 38789 12738 39421
rect 12702 37999 12738 38631
rect 12702 37209 12738 37841
rect 12702 36419 12738 37051
rect 12702 35629 12738 36261
rect 12702 34839 12738 35471
rect 12702 34049 12738 34681
rect 12702 33259 12738 33891
rect 12702 32469 12738 33101
rect 12702 31679 12738 32311
rect 12702 30889 12738 31521
rect 12702 30099 12738 30731
rect 12702 29309 12738 29941
rect 12702 28519 12738 29151
rect 12702 27729 12738 28361
rect 12702 26939 12738 27571
rect 12702 26149 12738 26781
rect 12702 25359 12738 25991
rect 12702 24569 12738 25201
rect 12702 23779 12738 24411
rect 12702 22989 12738 23621
rect 12702 22199 12738 22831
rect 12702 21409 12738 22041
rect 12702 20619 12738 21251
rect 12702 19829 12738 20461
rect 12702 19039 12738 19671
rect 12702 18249 12738 18881
rect 12702 17459 12738 18091
rect 12702 16669 12738 17301
rect 12702 15879 12738 16511
rect 12702 15089 12738 15721
rect 12702 14299 12738 14931
rect 12702 13509 12738 14141
rect 12702 12719 12738 13351
rect 12702 11929 12738 12561
rect 12702 11139 12738 11771
rect 12702 10349 12738 10981
rect 12702 9559 12738 10191
rect 12702 8769 12738 9401
rect 12702 7979 12738 8611
rect 12702 7189 12738 7821
rect 12702 6399 12738 7031
rect 12702 5609 12738 6241
rect 12702 4819 12738 5451
rect 12702 4029 12738 4661
rect 12702 3239 12738 3871
rect 12702 2449 12738 3081
rect 12702 1659 12738 2291
rect 12702 869 12738 1501
rect 12702 79 12738 711
rect 12774 0 12810 50560
rect 12846 0 12882 50560
rect 13326 0 13362 50560
rect 13398 0 13434 50560
rect 13470 49849 13506 50481
rect 13470 49059 13506 49691
rect 13470 48269 13506 48901
rect 13470 47479 13506 48111
rect 13470 46689 13506 47321
rect 13470 45899 13506 46531
rect 13470 45109 13506 45741
rect 13470 44319 13506 44951
rect 13470 43529 13506 44161
rect 13470 42739 13506 43371
rect 13470 41949 13506 42581
rect 13470 41159 13506 41791
rect 13470 40369 13506 41001
rect 13470 39579 13506 40211
rect 13470 38789 13506 39421
rect 13470 37999 13506 38631
rect 13470 37209 13506 37841
rect 13470 36419 13506 37051
rect 13470 35629 13506 36261
rect 13470 34839 13506 35471
rect 13470 34049 13506 34681
rect 13470 33259 13506 33891
rect 13470 32469 13506 33101
rect 13470 31679 13506 32311
rect 13470 30889 13506 31521
rect 13470 30099 13506 30731
rect 13470 29309 13506 29941
rect 13470 28519 13506 29151
rect 13470 27729 13506 28361
rect 13470 26939 13506 27571
rect 13470 26149 13506 26781
rect 13470 25359 13506 25991
rect 13470 24569 13506 25201
rect 13470 23779 13506 24411
rect 13470 22989 13506 23621
rect 13470 22199 13506 22831
rect 13470 21409 13506 22041
rect 13470 20619 13506 21251
rect 13470 19829 13506 20461
rect 13470 19039 13506 19671
rect 13470 18249 13506 18881
rect 13470 17459 13506 18091
rect 13470 16669 13506 17301
rect 13470 15879 13506 16511
rect 13470 15089 13506 15721
rect 13470 14299 13506 14931
rect 13470 13509 13506 14141
rect 13470 12719 13506 13351
rect 13470 11929 13506 12561
rect 13470 11139 13506 11771
rect 13470 10349 13506 10981
rect 13470 9559 13506 10191
rect 13470 8769 13506 9401
rect 13470 7979 13506 8611
rect 13470 7189 13506 7821
rect 13470 6399 13506 7031
rect 13470 5609 13506 6241
rect 13470 4819 13506 5451
rect 13470 4029 13506 4661
rect 13470 3239 13506 3871
rect 13470 2449 13506 3081
rect 13470 1659 13506 2291
rect 13470 869 13506 1501
rect 13470 79 13506 711
rect 13542 0 13578 50560
rect 13614 0 13650 50560
rect 13806 0 13842 50560
rect 13878 0 13914 50560
rect 13950 49849 13986 50481
rect 13950 49059 13986 49691
rect 13950 48269 13986 48901
rect 13950 47479 13986 48111
rect 13950 46689 13986 47321
rect 13950 45899 13986 46531
rect 13950 45109 13986 45741
rect 13950 44319 13986 44951
rect 13950 43529 13986 44161
rect 13950 42739 13986 43371
rect 13950 41949 13986 42581
rect 13950 41159 13986 41791
rect 13950 40369 13986 41001
rect 13950 39579 13986 40211
rect 13950 38789 13986 39421
rect 13950 37999 13986 38631
rect 13950 37209 13986 37841
rect 13950 36419 13986 37051
rect 13950 35629 13986 36261
rect 13950 34839 13986 35471
rect 13950 34049 13986 34681
rect 13950 33259 13986 33891
rect 13950 32469 13986 33101
rect 13950 31679 13986 32311
rect 13950 30889 13986 31521
rect 13950 30099 13986 30731
rect 13950 29309 13986 29941
rect 13950 28519 13986 29151
rect 13950 27729 13986 28361
rect 13950 26939 13986 27571
rect 13950 26149 13986 26781
rect 13950 25359 13986 25991
rect 13950 24569 13986 25201
rect 13950 23779 13986 24411
rect 13950 22989 13986 23621
rect 13950 22199 13986 22831
rect 13950 21409 13986 22041
rect 13950 20619 13986 21251
rect 13950 19829 13986 20461
rect 13950 19039 13986 19671
rect 13950 18249 13986 18881
rect 13950 17459 13986 18091
rect 13950 16669 13986 17301
rect 13950 15879 13986 16511
rect 13950 15089 13986 15721
rect 13950 14299 13986 14931
rect 13950 13509 13986 14141
rect 13950 12719 13986 13351
rect 13950 11929 13986 12561
rect 13950 11139 13986 11771
rect 13950 10349 13986 10981
rect 13950 9559 13986 10191
rect 13950 8769 13986 9401
rect 13950 7979 13986 8611
rect 13950 7189 13986 7821
rect 13950 6399 13986 7031
rect 13950 5609 13986 6241
rect 13950 4819 13986 5451
rect 13950 4029 13986 4661
rect 13950 3239 13986 3871
rect 13950 2449 13986 3081
rect 13950 1659 13986 2291
rect 13950 869 13986 1501
rect 13950 79 13986 711
rect 14022 0 14058 50560
rect 14094 0 14130 50560
rect 14574 0 14610 50560
rect 14646 0 14682 50560
rect 14718 49849 14754 50481
rect 14718 49059 14754 49691
rect 14718 48269 14754 48901
rect 14718 47479 14754 48111
rect 14718 46689 14754 47321
rect 14718 45899 14754 46531
rect 14718 45109 14754 45741
rect 14718 44319 14754 44951
rect 14718 43529 14754 44161
rect 14718 42739 14754 43371
rect 14718 41949 14754 42581
rect 14718 41159 14754 41791
rect 14718 40369 14754 41001
rect 14718 39579 14754 40211
rect 14718 38789 14754 39421
rect 14718 37999 14754 38631
rect 14718 37209 14754 37841
rect 14718 36419 14754 37051
rect 14718 35629 14754 36261
rect 14718 34839 14754 35471
rect 14718 34049 14754 34681
rect 14718 33259 14754 33891
rect 14718 32469 14754 33101
rect 14718 31679 14754 32311
rect 14718 30889 14754 31521
rect 14718 30099 14754 30731
rect 14718 29309 14754 29941
rect 14718 28519 14754 29151
rect 14718 27729 14754 28361
rect 14718 26939 14754 27571
rect 14718 26149 14754 26781
rect 14718 25359 14754 25991
rect 14718 24569 14754 25201
rect 14718 23779 14754 24411
rect 14718 22989 14754 23621
rect 14718 22199 14754 22831
rect 14718 21409 14754 22041
rect 14718 20619 14754 21251
rect 14718 19829 14754 20461
rect 14718 19039 14754 19671
rect 14718 18249 14754 18881
rect 14718 17459 14754 18091
rect 14718 16669 14754 17301
rect 14718 15879 14754 16511
rect 14718 15089 14754 15721
rect 14718 14299 14754 14931
rect 14718 13509 14754 14141
rect 14718 12719 14754 13351
rect 14718 11929 14754 12561
rect 14718 11139 14754 11771
rect 14718 10349 14754 10981
rect 14718 9559 14754 10191
rect 14718 8769 14754 9401
rect 14718 7979 14754 8611
rect 14718 7189 14754 7821
rect 14718 6399 14754 7031
rect 14718 5609 14754 6241
rect 14718 4819 14754 5451
rect 14718 4029 14754 4661
rect 14718 3239 14754 3871
rect 14718 2449 14754 3081
rect 14718 1659 14754 2291
rect 14718 869 14754 1501
rect 14718 79 14754 711
rect 14790 0 14826 50560
rect 14862 0 14898 50560
rect 15054 0 15090 50560
rect 15126 0 15162 50560
rect 15198 49849 15234 50481
rect 15198 49059 15234 49691
rect 15198 48269 15234 48901
rect 15198 47479 15234 48111
rect 15198 46689 15234 47321
rect 15198 45899 15234 46531
rect 15198 45109 15234 45741
rect 15198 44319 15234 44951
rect 15198 43529 15234 44161
rect 15198 42739 15234 43371
rect 15198 41949 15234 42581
rect 15198 41159 15234 41791
rect 15198 40369 15234 41001
rect 15198 39579 15234 40211
rect 15198 38789 15234 39421
rect 15198 37999 15234 38631
rect 15198 37209 15234 37841
rect 15198 36419 15234 37051
rect 15198 35629 15234 36261
rect 15198 34839 15234 35471
rect 15198 34049 15234 34681
rect 15198 33259 15234 33891
rect 15198 32469 15234 33101
rect 15198 31679 15234 32311
rect 15198 30889 15234 31521
rect 15198 30099 15234 30731
rect 15198 29309 15234 29941
rect 15198 28519 15234 29151
rect 15198 27729 15234 28361
rect 15198 26939 15234 27571
rect 15198 26149 15234 26781
rect 15198 25359 15234 25991
rect 15198 24569 15234 25201
rect 15198 23779 15234 24411
rect 15198 22989 15234 23621
rect 15198 22199 15234 22831
rect 15198 21409 15234 22041
rect 15198 20619 15234 21251
rect 15198 19829 15234 20461
rect 15198 19039 15234 19671
rect 15198 18249 15234 18881
rect 15198 17459 15234 18091
rect 15198 16669 15234 17301
rect 15198 15879 15234 16511
rect 15198 15089 15234 15721
rect 15198 14299 15234 14931
rect 15198 13509 15234 14141
rect 15198 12719 15234 13351
rect 15198 11929 15234 12561
rect 15198 11139 15234 11771
rect 15198 10349 15234 10981
rect 15198 9559 15234 10191
rect 15198 8769 15234 9401
rect 15198 7979 15234 8611
rect 15198 7189 15234 7821
rect 15198 6399 15234 7031
rect 15198 5609 15234 6241
rect 15198 4819 15234 5451
rect 15198 4029 15234 4661
rect 15198 3239 15234 3871
rect 15198 2449 15234 3081
rect 15198 1659 15234 2291
rect 15198 869 15234 1501
rect 15198 79 15234 711
rect 15270 0 15306 50560
rect 15342 0 15378 50560
rect 15822 0 15858 50560
rect 15894 0 15930 50560
rect 15966 49849 16002 50481
rect 15966 49059 16002 49691
rect 15966 48269 16002 48901
rect 15966 47479 16002 48111
rect 15966 46689 16002 47321
rect 15966 45899 16002 46531
rect 15966 45109 16002 45741
rect 15966 44319 16002 44951
rect 15966 43529 16002 44161
rect 15966 42739 16002 43371
rect 15966 41949 16002 42581
rect 15966 41159 16002 41791
rect 15966 40369 16002 41001
rect 15966 39579 16002 40211
rect 15966 38789 16002 39421
rect 15966 37999 16002 38631
rect 15966 37209 16002 37841
rect 15966 36419 16002 37051
rect 15966 35629 16002 36261
rect 15966 34839 16002 35471
rect 15966 34049 16002 34681
rect 15966 33259 16002 33891
rect 15966 32469 16002 33101
rect 15966 31679 16002 32311
rect 15966 30889 16002 31521
rect 15966 30099 16002 30731
rect 15966 29309 16002 29941
rect 15966 28519 16002 29151
rect 15966 27729 16002 28361
rect 15966 26939 16002 27571
rect 15966 26149 16002 26781
rect 15966 25359 16002 25991
rect 15966 24569 16002 25201
rect 15966 23779 16002 24411
rect 15966 22989 16002 23621
rect 15966 22199 16002 22831
rect 15966 21409 16002 22041
rect 15966 20619 16002 21251
rect 15966 19829 16002 20461
rect 15966 19039 16002 19671
rect 15966 18249 16002 18881
rect 15966 17459 16002 18091
rect 15966 16669 16002 17301
rect 15966 15879 16002 16511
rect 15966 15089 16002 15721
rect 15966 14299 16002 14931
rect 15966 13509 16002 14141
rect 15966 12719 16002 13351
rect 15966 11929 16002 12561
rect 15966 11139 16002 11771
rect 15966 10349 16002 10981
rect 15966 9559 16002 10191
rect 15966 8769 16002 9401
rect 15966 7979 16002 8611
rect 15966 7189 16002 7821
rect 15966 6399 16002 7031
rect 15966 5609 16002 6241
rect 15966 4819 16002 5451
rect 15966 4029 16002 4661
rect 15966 3239 16002 3871
rect 15966 2449 16002 3081
rect 15966 1659 16002 2291
rect 15966 869 16002 1501
rect 15966 79 16002 711
rect 16038 0 16074 50560
rect 16110 0 16146 50560
rect 16302 0 16338 50560
rect 16374 0 16410 50560
rect 16446 49849 16482 50481
rect 16446 49059 16482 49691
rect 16446 48269 16482 48901
rect 16446 47479 16482 48111
rect 16446 46689 16482 47321
rect 16446 45899 16482 46531
rect 16446 45109 16482 45741
rect 16446 44319 16482 44951
rect 16446 43529 16482 44161
rect 16446 42739 16482 43371
rect 16446 41949 16482 42581
rect 16446 41159 16482 41791
rect 16446 40369 16482 41001
rect 16446 39579 16482 40211
rect 16446 38789 16482 39421
rect 16446 37999 16482 38631
rect 16446 37209 16482 37841
rect 16446 36419 16482 37051
rect 16446 35629 16482 36261
rect 16446 34839 16482 35471
rect 16446 34049 16482 34681
rect 16446 33259 16482 33891
rect 16446 32469 16482 33101
rect 16446 31679 16482 32311
rect 16446 30889 16482 31521
rect 16446 30099 16482 30731
rect 16446 29309 16482 29941
rect 16446 28519 16482 29151
rect 16446 27729 16482 28361
rect 16446 26939 16482 27571
rect 16446 26149 16482 26781
rect 16446 25359 16482 25991
rect 16446 24569 16482 25201
rect 16446 23779 16482 24411
rect 16446 22989 16482 23621
rect 16446 22199 16482 22831
rect 16446 21409 16482 22041
rect 16446 20619 16482 21251
rect 16446 19829 16482 20461
rect 16446 19039 16482 19671
rect 16446 18249 16482 18881
rect 16446 17459 16482 18091
rect 16446 16669 16482 17301
rect 16446 15879 16482 16511
rect 16446 15089 16482 15721
rect 16446 14299 16482 14931
rect 16446 13509 16482 14141
rect 16446 12719 16482 13351
rect 16446 11929 16482 12561
rect 16446 11139 16482 11771
rect 16446 10349 16482 10981
rect 16446 9559 16482 10191
rect 16446 8769 16482 9401
rect 16446 7979 16482 8611
rect 16446 7189 16482 7821
rect 16446 6399 16482 7031
rect 16446 5609 16482 6241
rect 16446 4819 16482 5451
rect 16446 4029 16482 4661
rect 16446 3239 16482 3871
rect 16446 2449 16482 3081
rect 16446 1659 16482 2291
rect 16446 869 16482 1501
rect 16446 79 16482 711
rect 16518 0 16554 50560
rect 16590 0 16626 50560
rect 17070 0 17106 50560
rect 17142 0 17178 50560
rect 17214 49849 17250 50481
rect 17214 49059 17250 49691
rect 17214 48269 17250 48901
rect 17214 47479 17250 48111
rect 17214 46689 17250 47321
rect 17214 45899 17250 46531
rect 17214 45109 17250 45741
rect 17214 44319 17250 44951
rect 17214 43529 17250 44161
rect 17214 42739 17250 43371
rect 17214 41949 17250 42581
rect 17214 41159 17250 41791
rect 17214 40369 17250 41001
rect 17214 39579 17250 40211
rect 17214 38789 17250 39421
rect 17214 37999 17250 38631
rect 17214 37209 17250 37841
rect 17214 36419 17250 37051
rect 17214 35629 17250 36261
rect 17214 34839 17250 35471
rect 17214 34049 17250 34681
rect 17214 33259 17250 33891
rect 17214 32469 17250 33101
rect 17214 31679 17250 32311
rect 17214 30889 17250 31521
rect 17214 30099 17250 30731
rect 17214 29309 17250 29941
rect 17214 28519 17250 29151
rect 17214 27729 17250 28361
rect 17214 26939 17250 27571
rect 17214 26149 17250 26781
rect 17214 25359 17250 25991
rect 17214 24569 17250 25201
rect 17214 23779 17250 24411
rect 17214 22989 17250 23621
rect 17214 22199 17250 22831
rect 17214 21409 17250 22041
rect 17214 20619 17250 21251
rect 17214 19829 17250 20461
rect 17214 19039 17250 19671
rect 17214 18249 17250 18881
rect 17214 17459 17250 18091
rect 17214 16669 17250 17301
rect 17214 15879 17250 16511
rect 17214 15089 17250 15721
rect 17214 14299 17250 14931
rect 17214 13509 17250 14141
rect 17214 12719 17250 13351
rect 17214 11929 17250 12561
rect 17214 11139 17250 11771
rect 17214 10349 17250 10981
rect 17214 9559 17250 10191
rect 17214 8769 17250 9401
rect 17214 7979 17250 8611
rect 17214 7189 17250 7821
rect 17214 6399 17250 7031
rect 17214 5609 17250 6241
rect 17214 4819 17250 5451
rect 17214 4029 17250 4661
rect 17214 3239 17250 3871
rect 17214 2449 17250 3081
rect 17214 1659 17250 2291
rect 17214 869 17250 1501
rect 17214 79 17250 711
rect 17286 0 17322 50560
rect 17358 0 17394 50560
rect 17550 0 17586 50560
rect 17622 0 17658 50560
rect 17694 49849 17730 50481
rect 17694 49059 17730 49691
rect 17694 48269 17730 48901
rect 17694 47479 17730 48111
rect 17694 46689 17730 47321
rect 17694 45899 17730 46531
rect 17694 45109 17730 45741
rect 17694 44319 17730 44951
rect 17694 43529 17730 44161
rect 17694 42739 17730 43371
rect 17694 41949 17730 42581
rect 17694 41159 17730 41791
rect 17694 40369 17730 41001
rect 17694 39579 17730 40211
rect 17694 38789 17730 39421
rect 17694 37999 17730 38631
rect 17694 37209 17730 37841
rect 17694 36419 17730 37051
rect 17694 35629 17730 36261
rect 17694 34839 17730 35471
rect 17694 34049 17730 34681
rect 17694 33259 17730 33891
rect 17694 32469 17730 33101
rect 17694 31679 17730 32311
rect 17694 30889 17730 31521
rect 17694 30099 17730 30731
rect 17694 29309 17730 29941
rect 17694 28519 17730 29151
rect 17694 27729 17730 28361
rect 17694 26939 17730 27571
rect 17694 26149 17730 26781
rect 17694 25359 17730 25991
rect 17694 24569 17730 25201
rect 17694 23779 17730 24411
rect 17694 22989 17730 23621
rect 17694 22199 17730 22831
rect 17694 21409 17730 22041
rect 17694 20619 17730 21251
rect 17694 19829 17730 20461
rect 17694 19039 17730 19671
rect 17694 18249 17730 18881
rect 17694 17459 17730 18091
rect 17694 16669 17730 17301
rect 17694 15879 17730 16511
rect 17694 15089 17730 15721
rect 17694 14299 17730 14931
rect 17694 13509 17730 14141
rect 17694 12719 17730 13351
rect 17694 11929 17730 12561
rect 17694 11139 17730 11771
rect 17694 10349 17730 10981
rect 17694 9559 17730 10191
rect 17694 8769 17730 9401
rect 17694 7979 17730 8611
rect 17694 7189 17730 7821
rect 17694 6399 17730 7031
rect 17694 5609 17730 6241
rect 17694 4819 17730 5451
rect 17694 4029 17730 4661
rect 17694 3239 17730 3871
rect 17694 2449 17730 3081
rect 17694 1659 17730 2291
rect 17694 869 17730 1501
rect 17694 79 17730 711
rect 17766 0 17802 50560
rect 17838 0 17874 50560
rect 18318 0 18354 50560
rect 18390 0 18426 50560
rect 18462 49849 18498 50481
rect 18462 49059 18498 49691
rect 18462 48269 18498 48901
rect 18462 47479 18498 48111
rect 18462 46689 18498 47321
rect 18462 45899 18498 46531
rect 18462 45109 18498 45741
rect 18462 44319 18498 44951
rect 18462 43529 18498 44161
rect 18462 42739 18498 43371
rect 18462 41949 18498 42581
rect 18462 41159 18498 41791
rect 18462 40369 18498 41001
rect 18462 39579 18498 40211
rect 18462 38789 18498 39421
rect 18462 37999 18498 38631
rect 18462 37209 18498 37841
rect 18462 36419 18498 37051
rect 18462 35629 18498 36261
rect 18462 34839 18498 35471
rect 18462 34049 18498 34681
rect 18462 33259 18498 33891
rect 18462 32469 18498 33101
rect 18462 31679 18498 32311
rect 18462 30889 18498 31521
rect 18462 30099 18498 30731
rect 18462 29309 18498 29941
rect 18462 28519 18498 29151
rect 18462 27729 18498 28361
rect 18462 26939 18498 27571
rect 18462 26149 18498 26781
rect 18462 25359 18498 25991
rect 18462 24569 18498 25201
rect 18462 23779 18498 24411
rect 18462 22989 18498 23621
rect 18462 22199 18498 22831
rect 18462 21409 18498 22041
rect 18462 20619 18498 21251
rect 18462 19829 18498 20461
rect 18462 19039 18498 19671
rect 18462 18249 18498 18881
rect 18462 17459 18498 18091
rect 18462 16669 18498 17301
rect 18462 15879 18498 16511
rect 18462 15089 18498 15721
rect 18462 14299 18498 14931
rect 18462 13509 18498 14141
rect 18462 12719 18498 13351
rect 18462 11929 18498 12561
rect 18462 11139 18498 11771
rect 18462 10349 18498 10981
rect 18462 9559 18498 10191
rect 18462 8769 18498 9401
rect 18462 7979 18498 8611
rect 18462 7189 18498 7821
rect 18462 6399 18498 7031
rect 18462 5609 18498 6241
rect 18462 4819 18498 5451
rect 18462 4029 18498 4661
rect 18462 3239 18498 3871
rect 18462 2449 18498 3081
rect 18462 1659 18498 2291
rect 18462 869 18498 1501
rect 18462 79 18498 711
rect 18534 0 18570 50560
rect 18606 0 18642 50560
rect 18798 0 18834 50560
rect 18870 0 18906 50560
rect 18942 49849 18978 50481
rect 18942 49059 18978 49691
rect 18942 48269 18978 48901
rect 18942 47479 18978 48111
rect 18942 46689 18978 47321
rect 18942 45899 18978 46531
rect 18942 45109 18978 45741
rect 18942 44319 18978 44951
rect 18942 43529 18978 44161
rect 18942 42739 18978 43371
rect 18942 41949 18978 42581
rect 18942 41159 18978 41791
rect 18942 40369 18978 41001
rect 18942 39579 18978 40211
rect 18942 38789 18978 39421
rect 18942 37999 18978 38631
rect 18942 37209 18978 37841
rect 18942 36419 18978 37051
rect 18942 35629 18978 36261
rect 18942 34839 18978 35471
rect 18942 34049 18978 34681
rect 18942 33259 18978 33891
rect 18942 32469 18978 33101
rect 18942 31679 18978 32311
rect 18942 30889 18978 31521
rect 18942 30099 18978 30731
rect 18942 29309 18978 29941
rect 18942 28519 18978 29151
rect 18942 27729 18978 28361
rect 18942 26939 18978 27571
rect 18942 26149 18978 26781
rect 18942 25359 18978 25991
rect 18942 24569 18978 25201
rect 18942 23779 18978 24411
rect 18942 22989 18978 23621
rect 18942 22199 18978 22831
rect 18942 21409 18978 22041
rect 18942 20619 18978 21251
rect 18942 19829 18978 20461
rect 18942 19039 18978 19671
rect 18942 18249 18978 18881
rect 18942 17459 18978 18091
rect 18942 16669 18978 17301
rect 18942 15879 18978 16511
rect 18942 15089 18978 15721
rect 18942 14299 18978 14931
rect 18942 13509 18978 14141
rect 18942 12719 18978 13351
rect 18942 11929 18978 12561
rect 18942 11139 18978 11771
rect 18942 10349 18978 10981
rect 18942 9559 18978 10191
rect 18942 8769 18978 9401
rect 18942 7979 18978 8611
rect 18942 7189 18978 7821
rect 18942 6399 18978 7031
rect 18942 5609 18978 6241
rect 18942 4819 18978 5451
rect 18942 4029 18978 4661
rect 18942 3239 18978 3871
rect 18942 2449 18978 3081
rect 18942 1659 18978 2291
rect 18942 869 18978 1501
rect 18942 79 18978 711
rect 19014 0 19050 50560
rect 19086 0 19122 50560
rect 19566 0 19602 50560
rect 19638 0 19674 50560
rect 19710 49849 19746 50481
rect 19710 49059 19746 49691
rect 19710 48269 19746 48901
rect 19710 47479 19746 48111
rect 19710 46689 19746 47321
rect 19710 45899 19746 46531
rect 19710 45109 19746 45741
rect 19710 44319 19746 44951
rect 19710 43529 19746 44161
rect 19710 42739 19746 43371
rect 19710 41949 19746 42581
rect 19710 41159 19746 41791
rect 19710 40369 19746 41001
rect 19710 39579 19746 40211
rect 19710 38789 19746 39421
rect 19710 37999 19746 38631
rect 19710 37209 19746 37841
rect 19710 36419 19746 37051
rect 19710 35629 19746 36261
rect 19710 34839 19746 35471
rect 19710 34049 19746 34681
rect 19710 33259 19746 33891
rect 19710 32469 19746 33101
rect 19710 31679 19746 32311
rect 19710 30889 19746 31521
rect 19710 30099 19746 30731
rect 19710 29309 19746 29941
rect 19710 28519 19746 29151
rect 19710 27729 19746 28361
rect 19710 26939 19746 27571
rect 19710 26149 19746 26781
rect 19710 25359 19746 25991
rect 19710 24569 19746 25201
rect 19710 23779 19746 24411
rect 19710 22989 19746 23621
rect 19710 22199 19746 22831
rect 19710 21409 19746 22041
rect 19710 20619 19746 21251
rect 19710 19829 19746 20461
rect 19710 19039 19746 19671
rect 19710 18249 19746 18881
rect 19710 17459 19746 18091
rect 19710 16669 19746 17301
rect 19710 15879 19746 16511
rect 19710 15089 19746 15721
rect 19710 14299 19746 14931
rect 19710 13509 19746 14141
rect 19710 12719 19746 13351
rect 19710 11929 19746 12561
rect 19710 11139 19746 11771
rect 19710 10349 19746 10981
rect 19710 9559 19746 10191
rect 19710 8769 19746 9401
rect 19710 7979 19746 8611
rect 19710 7189 19746 7821
rect 19710 6399 19746 7031
rect 19710 5609 19746 6241
rect 19710 4819 19746 5451
rect 19710 4029 19746 4661
rect 19710 3239 19746 3871
rect 19710 2449 19746 3081
rect 19710 1659 19746 2291
rect 19710 869 19746 1501
rect 19710 79 19746 711
rect 19782 0 19818 50560
rect 19854 0 19890 50560
rect 20046 0 20082 50560
rect 20118 0 20154 50560
rect 20190 49849 20226 50481
rect 20190 49059 20226 49691
rect 20190 48269 20226 48901
rect 20190 47479 20226 48111
rect 20190 46689 20226 47321
rect 20190 45899 20226 46531
rect 20190 45109 20226 45741
rect 20190 44319 20226 44951
rect 20190 43529 20226 44161
rect 20190 42739 20226 43371
rect 20190 41949 20226 42581
rect 20190 41159 20226 41791
rect 20190 40369 20226 41001
rect 20190 39579 20226 40211
rect 20190 38789 20226 39421
rect 20190 37999 20226 38631
rect 20190 37209 20226 37841
rect 20190 36419 20226 37051
rect 20190 35629 20226 36261
rect 20190 34839 20226 35471
rect 20190 34049 20226 34681
rect 20190 33259 20226 33891
rect 20190 32469 20226 33101
rect 20190 31679 20226 32311
rect 20190 30889 20226 31521
rect 20190 30099 20226 30731
rect 20190 29309 20226 29941
rect 20190 28519 20226 29151
rect 20190 27729 20226 28361
rect 20190 26939 20226 27571
rect 20190 26149 20226 26781
rect 20190 25359 20226 25991
rect 20190 24569 20226 25201
rect 20190 23779 20226 24411
rect 20190 22989 20226 23621
rect 20190 22199 20226 22831
rect 20190 21409 20226 22041
rect 20190 20619 20226 21251
rect 20190 19829 20226 20461
rect 20190 19039 20226 19671
rect 20190 18249 20226 18881
rect 20190 17459 20226 18091
rect 20190 16669 20226 17301
rect 20190 15879 20226 16511
rect 20190 15089 20226 15721
rect 20190 14299 20226 14931
rect 20190 13509 20226 14141
rect 20190 12719 20226 13351
rect 20190 11929 20226 12561
rect 20190 11139 20226 11771
rect 20190 10349 20226 10981
rect 20190 9559 20226 10191
rect 20190 8769 20226 9401
rect 20190 7979 20226 8611
rect 20190 7189 20226 7821
rect 20190 6399 20226 7031
rect 20190 5609 20226 6241
rect 20190 4819 20226 5451
rect 20190 4029 20226 4661
rect 20190 3239 20226 3871
rect 20190 2449 20226 3081
rect 20190 1659 20226 2291
rect 20190 869 20226 1501
rect 20190 79 20226 711
rect 20262 0 20298 50560
rect 20334 0 20370 50560
rect 20814 0 20850 50560
rect 20886 0 20922 50560
rect 20958 49849 20994 50481
rect 20958 49059 20994 49691
rect 20958 48269 20994 48901
rect 20958 47479 20994 48111
rect 20958 46689 20994 47321
rect 20958 45899 20994 46531
rect 20958 45109 20994 45741
rect 20958 44319 20994 44951
rect 20958 43529 20994 44161
rect 20958 42739 20994 43371
rect 20958 41949 20994 42581
rect 20958 41159 20994 41791
rect 20958 40369 20994 41001
rect 20958 39579 20994 40211
rect 20958 38789 20994 39421
rect 20958 37999 20994 38631
rect 20958 37209 20994 37841
rect 20958 36419 20994 37051
rect 20958 35629 20994 36261
rect 20958 34839 20994 35471
rect 20958 34049 20994 34681
rect 20958 33259 20994 33891
rect 20958 32469 20994 33101
rect 20958 31679 20994 32311
rect 20958 30889 20994 31521
rect 20958 30099 20994 30731
rect 20958 29309 20994 29941
rect 20958 28519 20994 29151
rect 20958 27729 20994 28361
rect 20958 26939 20994 27571
rect 20958 26149 20994 26781
rect 20958 25359 20994 25991
rect 20958 24569 20994 25201
rect 20958 23779 20994 24411
rect 20958 22989 20994 23621
rect 20958 22199 20994 22831
rect 20958 21409 20994 22041
rect 20958 20619 20994 21251
rect 20958 19829 20994 20461
rect 20958 19039 20994 19671
rect 20958 18249 20994 18881
rect 20958 17459 20994 18091
rect 20958 16669 20994 17301
rect 20958 15879 20994 16511
rect 20958 15089 20994 15721
rect 20958 14299 20994 14931
rect 20958 13509 20994 14141
rect 20958 12719 20994 13351
rect 20958 11929 20994 12561
rect 20958 11139 20994 11771
rect 20958 10349 20994 10981
rect 20958 9559 20994 10191
rect 20958 8769 20994 9401
rect 20958 7979 20994 8611
rect 20958 7189 20994 7821
rect 20958 6399 20994 7031
rect 20958 5609 20994 6241
rect 20958 4819 20994 5451
rect 20958 4029 20994 4661
rect 20958 3239 20994 3871
rect 20958 2449 20994 3081
rect 20958 1659 20994 2291
rect 20958 869 20994 1501
rect 20958 79 20994 711
rect 21030 0 21066 50560
rect 21102 0 21138 50560
rect 21294 0 21330 50560
rect 21366 0 21402 50560
rect 21438 49849 21474 50481
rect 21438 49059 21474 49691
rect 21438 48269 21474 48901
rect 21438 47479 21474 48111
rect 21438 46689 21474 47321
rect 21438 45899 21474 46531
rect 21438 45109 21474 45741
rect 21438 44319 21474 44951
rect 21438 43529 21474 44161
rect 21438 42739 21474 43371
rect 21438 41949 21474 42581
rect 21438 41159 21474 41791
rect 21438 40369 21474 41001
rect 21438 39579 21474 40211
rect 21438 38789 21474 39421
rect 21438 37999 21474 38631
rect 21438 37209 21474 37841
rect 21438 36419 21474 37051
rect 21438 35629 21474 36261
rect 21438 34839 21474 35471
rect 21438 34049 21474 34681
rect 21438 33259 21474 33891
rect 21438 32469 21474 33101
rect 21438 31679 21474 32311
rect 21438 30889 21474 31521
rect 21438 30099 21474 30731
rect 21438 29309 21474 29941
rect 21438 28519 21474 29151
rect 21438 27729 21474 28361
rect 21438 26939 21474 27571
rect 21438 26149 21474 26781
rect 21438 25359 21474 25991
rect 21438 24569 21474 25201
rect 21438 23779 21474 24411
rect 21438 22989 21474 23621
rect 21438 22199 21474 22831
rect 21438 21409 21474 22041
rect 21438 20619 21474 21251
rect 21438 19829 21474 20461
rect 21438 19039 21474 19671
rect 21438 18249 21474 18881
rect 21438 17459 21474 18091
rect 21438 16669 21474 17301
rect 21438 15879 21474 16511
rect 21438 15089 21474 15721
rect 21438 14299 21474 14931
rect 21438 13509 21474 14141
rect 21438 12719 21474 13351
rect 21438 11929 21474 12561
rect 21438 11139 21474 11771
rect 21438 10349 21474 10981
rect 21438 9559 21474 10191
rect 21438 8769 21474 9401
rect 21438 7979 21474 8611
rect 21438 7189 21474 7821
rect 21438 6399 21474 7031
rect 21438 5609 21474 6241
rect 21438 4819 21474 5451
rect 21438 4029 21474 4661
rect 21438 3239 21474 3871
rect 21438 2449 21474 3081
rect 21438 1659 21474 2291
rect 21438 869 21474 1501
rect 21438 79 21474 711
rect 21510 0 21546 50560
rect 21582 0 21618 50560
rect 22062 0 22098 50560
rect 22134 0 22170 50560
rect 22206 49849 22242 50481
rect 22206 49059 22242 49691
rect 22206 48269 22242 48901
rect 22206 47479 22242 48111
rect 22206 46689 22242 47321
rect 22206 45899 22242 46531
rect 22206 45109 22242 45741
rect 22206 44319 22242 44951
rect 22206 43529 22242 44161
rect 22206 42739 22242 43371
rect 22206 41949 22242 42581
rect 22206 41159 22242 41791
rect 22206 40369 22242 41001
rect 22206 39579 22242 40211
rect 22206 38789 22242 39421
rect 22206 37999 22242 38631
rect 22206 37209 22242 37841
rect 22206 36419 22242 37051
rect 22206 35629 22242 36261
rect 22206 34839 22242 35471
rect 22206 34049 22242 34681
rect 22206 33259 22242 33891
rect 22206 32469 22242 33101
rect 22206 31679 22242 32311
rect 22206 30889 22242 31521
rect 22206 30099 22242 30731
rect 22206 29309 22242 29941
rect 22206 28519 22242 29151
rect 22206 27729 22242 28361
rect 22206 26939 22242 27571
rect 22206 26149 22242 26781
rect 22206 25359 22242 25991
rect 22206 24569 22242 25201
rect 22206 23779 22242 24411
rect 22206 22989 22242 23621
rect 22206 22199 22242 22831
rect 22206 21409 22242 22041
rect 22206 20619 22242 21251
rect 22206 19829 22242 20461
rect 22206 19039 22242 19671
rect 22206 18249 22242 18881
rect 22206 17459 22242 18091
rect 22206 16669 22242 17301
rect 22206 15879 22242 16511
rect 22206 15089 22242 15721
rect 22206 14299 22242 14931
rect 22206 13509 22242 14141
rect 22206 12719 22242 13351
rect 22206 11929 22242 12561
rect 22206 11139 22242 11771
rect 22206 10349 22242 10981
rect 22206 9559 22242 10191
rect 22206 8769 22242 9401
rect 22206 7979 22242 8611
rect 22206 7189 22242 7821
rect 22206 6399 22242 7031
rect 22206 5609 22242 6241
rect 22206 4819 22242 5451
rect 22206 4029 22242 4661
rect 22206 3239 22242 3871
rect 22206 2449 22242 3081
rect 22206 1659 22242 2291
rect 22206 869 22242 1501
rect 22206 79 22242 711
rect 22278 0 22314 50560
rect 22350 0 22386 50560
rect 22542 0 22578 50560
rect 22614 0 22650 50560
rect 22686 49849 22722 50481
rect 22686 49059 22722 49691
rect 22686 48269 22722 48901
rect 22686 47479 22722 48111
rect 22686 46689 22722 47321
rect 22686 45899 22722 46531
rect 22686 45109 22722 45741
rect 22686 44319 22722 44951
rect 22686 43529 22722 44161
rect 22686 42739 22722 43371
rect 22686 41949 22722 42581
rect 22686 41159 22722 41791
rect 22686 40369 22722 41001
rect 22686 39579 22722 40211
rect 22686 38789 22722 39421
rect 22686 37999 22722 38631
rect 22686 37209 22722 37841
rect 22686 36419 22722 37051
rect 22686 35629 22722 36261
rect 22686 34839 22722 35471
rect 22686 34049 22722 34681
rect 22686 33259 22722 33891
rect 22686 32469 22722 33101
rect 22686 31679 22722 32311
rect 22686 30889 22722 31521
rect 22686 30099 22722 30731
rect 22686 29309 22722 29941
rect 22686 28519 22722 29151
rect 22686 27729 22722 28361
rect 22686 26939 22722 27571
rect 22686 26149 22722 26781
rect 22686 25359 22722 25991
rect 22686 24569 22722 25201
rect 22686 23779 22722 24411
rect 22686 22989 22722 23621
rect 22686 22199 22722 22831
rect 22686 21409 22722 22041
rect 22686 20619 22722 21251
rect 22686 19829 22722 20461
rect 22686 19039 22722 19671
rect 22686 18249 22722 18881
rect 22686 17459 22722 18091
rect 22686 16669 22722 17301
rect 22686 15879 22722 16511
rect 22686 15089 22722 15721
rect 22686 14299 22722 14931
rect 22686 13509 22722 14141
rect 22686 12719 22722 13351
rect 22686 11929 22722 12561
rect 22686 11139 22722 11771
rect 22686 10349 22722 10981
rect 22686 9559 22722 10191
rect 22686 8769 22722 9401
rect 22686 7979 22722 8611
rect 22686 7189 22722 7821
rect 22686 6399 22722 7031
rect 22686 5609 22722 6241
rect 22686 4819 22722 5451
rect 22686 4029 22722 4661
rect 22686 3239 22722 3871
rect 22686 2449 22722 3081
rect 22686 1659 22722 2291
rect 22686 869 22722 1501
rect 22686 79 22722 711
rect 22758 0 22794 50560
rect 22830 0 22866 50560
rect 23310 0 23346 50560
rect 23382 0 23418 50560
rect 23454 49849 23490 50481
rect 23454 49059 23490 49691
rect 23454 48269 23490 48901
rect 23454 47479 23490 48111
rect 23454 46689 23490 47321
rect 23454 45899 23490 46531
rect 23454 45109 23490 45741
rect 23454 44319 23490 44951
rect 23454 43529 23490 44161
rect 23454 42739 23490 43371
rect 23454 41949 23490 42581
rect 23454 41159 23490 41791
rect 23454 40369 23490 41001
rect 23454 39579 23490 40211
rect 23454 38789 23490 39421
rect 23454 37999 23490 38631
rect 23454 37209 23490 37841
rect 23454 36419 23490 37051
rect 23454 35629 23490 36261
rect 23454 34839 23490 35471
rect 23454 34049 23490 34681
rect 23454 33259 23490 33891
rect 23454 32469 23490 33101
rect 23454 31679 23490 32311
rect 23454 30889 23490 31521
rect 23454 30099 23490 30731
rect 23454 29309 23490 29941
rect 23454 28519 23490 29151
rect 23454 27729 23490 28361
rect 23454 26939 23490 27571
rect 23454 26149 23490 26781
rect 23454 25359 23490 25991
rect 23454 24569 23490 25201
rect 23454 23779 23490 24411
rect 23454 22989 23490 23621
rect 23454 22199 23490 22831
rect 23454 21409 23490 22041
rect 23454 20619 23490 21251
rect 23454 19829 23490 20461
rect 23454 19039 23490 19671
rect 23454 18249 23490 18881
rect 23454 17459 23490 18091
rect 23454 16669 23490 17301
rect 23454 15879 23490 16511
rect 23454 15089 23490 15721
rect 23454 14299 23490 14931
rect 23454 13509 23490 14141
rect 23454 12719 23490 13351
rect 23454 11929 23490 12561
rect 23454 11139 23490 11771
rect 23454 10349 23490 10981
rect 23454 9559 23490 10191
rect 23454 8769 23490 9401
rect 23454 7979 23490 8611
rect 23454 7189 23490 7821
rect 23454 6399 23490 7031
rect 23454 5609 23490 6241
rect 23454 4819 23490 5451
rect 23454 4029 23490 4661
rect 23454 3239 23490 3871
rect 23454 2449 23490 3081
rect 23454 1659 23490 2291
rect 23454 869 23490 1501
rect 23454 79 23490 711
rect 23526 0 23562 50560
rect 23598 0 23634 50560
rect 23790 0 23826 50560
rect 23862 0 23898 50560
rect 23934 49849 23970 50481
rect 23934 49059 23970 49691
rect 23934 48269 23970 48901
rect 23934 47479 23970 48111
rect 23934 46689 23970 47321
rect 23934 45899 23970 46531
rect 23934 45109 23970 45741
rect 23934 44319 23970 44951
rect 23934 43529 23970 44161
rect 23934 42739 23970 43371
rect 23934 41949 23970 42581
rect 23934 41159 23970 41791
rect 23934 40369 23970 41001
rect 23934 39579 23970 40211
rect 23934 38789 23970 39421
rect 23934 37999 23970 38631
rect 23934 37209 23970 37841
rect 23934 36419 23970 37051
rect 23934 35629 23970 36261
rect 23934 34839 23970 35471
rect 23934 34049 23970 34681
rect 23934 33259 23970 33891
rect 23934 32469 23970 33101
rect 23934 31679 23970 32311
rect 23934 30889 23970 31521
rect 23934 30099 23970 30731
rect 23934 29309 23970 29941
rect 23934 28519 23970 29151
rect 23934 27729 23970 28361
rect 23934 26939 23970 27571
rect 23934 26149 23970 26781
rect 23934 25359 23970 25991
rect 23934 24569 23970 25201
rect 23934 23779 23970 24411
rect 23934 22989 23970 23621
rect 23934 22199 23970 22831
rect 23934 21409 23970 22041
rect 23934 20619 23970 21251
rect 23934 19829 23970 20461
rect 23934 19039 23970 19671
rect 23934 18249 23970 18881
rect 23934 17459 23970 18091
rect 23934 16669 23970 17301
rect 23934 15879 23970 16511
rect 23934 15089 23970 15721
rect 23934 14299 23970 14931
rect 23934 13509 23970 14141
rect 23934 12719 23970 13351
rect 23934 11929 23970 12561
rect 23934 11139 23970 11771
rect 23934 10349 23970 10981
rect 23934 9559 23970 10191
rect 23934 8769 23970 9401
rect 23934 7979 23970 8611
rect 23934 7189 23970 7821
rect 23934 6399 23970 7031
rect 23934 5609 23970 6241
rect 23934 4819 23970 5451
rect 23934 4029 23970 4661
rect 23934 3239 23970 3871
rect 23934 2449 23970 3081
rect 23934 1659 23970 2291
rect 23934 869 23970 1501
rect 23934 79 23970 711
rect 24006 0 24042 50560
rect 24078 0 24114 50560
rect 24558 0 24594 50560
rect 24630 0 24666 50560
rect 24702 49849 24738 50481
rect 24702 49059 24738 49691
rect 24702 48269 24738 48901
rect 24702 47479 24738 48111
rect 24702 46689 24738 47321
rect 24702 45899 24738 46531
rect 24702 45109 24738 45741
rect 24702 44319 24738 44951
rect 24702 43529 24738 44161
rect 24702 42739 24738 43371
rect 24702 41949 24738 42581
rect 24702 41159 24738 41791
rect 24702 40369 24738 41001
rect 24702 39579 24738 40211
rect 24702 38789 24738 39421
rect 24702 37999 24738 38631
rect 24702 37209 24738 37841
rect 24702 36419 24738 37051
rect 24702 35629 24738 36261
rect 24702 34839 24738 35471
rect 24702 34049 24738 34681
rect 24702 33259 24738 33891
rect 24702 32469 24738 33101
rect 24702 31679 24738 32311
rect 24702 30889 24738 31521
rect 24702 30099 24738 30731
rect 24702 29309 24738 29941
rect 24702 28519 24738 29151
rect 24702 27729 24738 28361
rect 24702 26939 24738 27571
rect 24702 26149 24738 26781
rect 24702 25359 24738 25991
rect 24702 24569 24738 25201
rect 24702 23779 24738 24411
rect 24702 22989 24738 23621
rect 24702 22199 24738 22831
rect 24702 21409 24738 22041
rect 24702 20619 24738 21251
rect 24702 19829 24738 20461
rect 24702 19039 24738 19671
rect 24702 18249 24738 18881
rect 24702 17459 24738 18091
rect 24702 16669 24738 17301
rect 24702 15879 24738 16511
rect 24702 15089 24738 15721
rect 24702 14299 24738 14931
rect 24702 13509 24738 14141
rect 24702 12719 24738 13351
rect 24702 11929 24738 12561
rect 24702 11139 24738 11771
rect 24702 10349 24738 10981
rect 24702 9559 24738 10191
rect 24702 8769 24738 9401
rect 24702 7979 24738 8611
rect 24702 7189 24738 7821
rect 24702 6399 24738 7031
rect 24702 5609 24738 6241
rect 24702 4819 24738 5451
rect 24702 4029 24738 4661
rect 24702 3239 24738 3871
rect 24702 2449 24738 3081
rect 24702 1659 24738 2291
rect 24702 869 24738 1501
rect 24702 79 24738 711
rect 24774 0 24810 50560
rect 24846 0 24882 50560
rect 25038 0 25074 50560
rect 25110 0 25146 50560
rect 25182 49849 25218 50481
rect 25182 49059 25218 49691
rect 25182 48269 25218 48901
rect 25182 47479 25218 48111
rect 25182 46689 25218 47321
rect 25182 45899 25218 46531
rect 25182 45109 25218 45741
rect 25182 44319 25218 44951
rect 25182 43529 25218 44161
rect 25182 42739 25218 43371
rect 25182 41949 25218 42581
rect 25182 41159 25218 41791
rect 25182 40369 25218 41001
rect 25182 39579 25218 40211
rect 25182 38789 25218 39421
rect 25182 37999 25218 38631
rect 25182 37209 25218 37841
rect 25182 36419 25218 37051
rect 25182 35629 25218 36261
rect 25182 34839 25218 35471
rect 25182 34049 25218 34681
rect 25182 33259 25218 33891
rect 25182 32469 25218 33101
rect 25182 31679 25218 32311
rect 25182 30889 25218 31521
rect 25182 30099 25218 30731
rect 25182 29309 25218 29941
rect 25182 28519 25218 29151
rect 25182 27729 25218 28361
rect 25182 26939 25218 27571
rect 25182 26149 25218 26781
rect 25182 25359 25218 25991
rect 25182 24569 25218 25201
rect 25182 23779 25218 24411
rect 25182 22989 25218 23621
rect 25182 22199 25218 22831
rect 25182 21409 25218 22041
rect 25182 20619 25218 21251
rect 25182 19829 25218 20461
rect 25182 19039 25218 19671
rect 25182 18249 25218 18881
rect 25182 17459 25218 18091
rect 25182 16669 25218 17301
rect 25182 15879 25218 16511
rect 25182 15089 25218 15721
rect 25182 14299 25218 14931
rect 25182 13509 25218 14141
rect 25182 12719 25218 13351
rect 25182 11929 25218 12561
rect 25182 11139 25218 11771
rect 25182 10349 25218 10981
rect 25182 9559 25218 10191
rect 25182 8769 25218 9401
rect 25182 7979 25218 8611
rect 25182 7189 25218 7821
rect 25182 6399 25218 7031
rect 25182 5609 25218 6241
rect 25182 4819 25218 5451
rect 25182 4029 25218 4661
rect 25182 3239 25218 3871
rect 25182 2449 25218 3081
rect 25182 1659 25218 2291
rect 25182 869 25218 1501
rect 25182 79 25218 711
rect 25254 0 25290 50560
rect 25326 0 25362 50560
rect 25806 0 25842 50560
rect 25878 0 25914 50560
rect 25950 49849 25986 50481
rect 25950 49059 25986 49691
rect 25950 48269 25986 48901
rect 25950 47479 25986 48111
rect 25950 46689 25986 47321
rect 25950 45899 25986 46531
rect 25950 45109 25986 45741
rect 25950 44319 25986 44951
rect 25950 43529 25986 44161
rect 25950 42739 25986 43371
rect 25950 41949 25986 42581
rect 25950 41159 25986 41791
rect 25950 40369 25986 41001
rect 25950 39579 25986 40211
rect 25950 38789 25986 39421
rect 25950 37999 25986 38631
rect 25950 37209 25986 37841
rect 25950 36419 25986 37051
rect 25950 35629 25986 36261
rect 25950 34839 25986 35471
rect 25950 34049 25986 34681
rect 25950 33259 25986 33891
rect 25950 32469 25986 33101
rect 25950 31679 25986 32311
rect 25950 30889 25986 31521
rect 25950 30099 25986 30731
rect 25950 29309 25986 29941
rect 25950 28519 25986 29151
rect 25950 27729 25986 28361
rect 25950 26939 25986 27571
rect 25950 26149 25986 26781
rect 25950 25359 25986 25991
rect 25950 24569 25986 25201
rect 25950 23779 25986 24411
rect 25950 22989 25986 23621
rect 25950 22199 25986 22831
rect 25950 21409 25986 22041
rect 25950 20619 25986 21251
rect 25950 19829 25986 20461
rect 25950 19039 25986 19671
rect 25950 18249 25986 18881
rect 25950 17459 25986 18091
rect 25950 16669 25986 17301
rect 25950 15879 25986 16511
rect 25950 15089 25986 15721
rect 25950 14299 25986 14931
rect 25950 13509 25986 14141
rect 25950 12719 25986 13351
rect 25950 11929 25986 12561
rect 25950 11139 25986 11771
rect 25950 10349 25986 10981
rect 25950 9559 25986 10191
rect 25950 8769 25986 9401
rect 25950 7979 25986 8611
rect 25950 7189 25986 7821
rect 25950 6399 25986 7031
rect 25950 5609 25986 6241
rect 25950 4819 25986 5451
rect 25950 4029 25986 4661
rect 25950 3239 25986 3871
rect 25950 2449 25986 3081
rect 25950 1659 25986 2291
rect 25950 869 25986 1501
rect 25950 79 25986 711
rect 26022 0 26058 50560
rect 26094 0 26130 50560
rect 26286 0 26322 50560
rect 26358 0 26394 50560
rect 26430 49849 26466 50481
rect 26430 49059 26466 49691
rect 26430 48269 26466 48901
rect 26430 47479 26466 48111
rect 26430 46689 26466 47321
rect 26430 45899 26466 46531
rect 26430 45109 26466 45741
rect 26430 44319 26466 44951
rect 26430 43529 26466 44161
rect 26430 42739 26466 43371
rect 26430 41949 26466 42581
rect 26430 41159 26466 41791
rect 26430 40369 26466 41001
rect 26430 39579 26466 40211
rect 26430 38789 26466 39421
rect 26430 37999 26466 38631
rect 26430 37209 26466 37841
rect 26430 36419 26466 37051
rect 26430 35629 26466 36261
rect 26430 34839 26466 35471
rect 26430 34049 26466 34681
rect 26430 33259 26466 33891
rect 26430 32469 26466 33101
rect 26430 31679 26466 32311
rect 26430 30889 26466 31521
rect 26430 30099 26466 30731
rect 26430 29309 26466 29941
rect 26430 28519 26466 29151
rect 26430 27729 26466 28361
rect 26430 26939 26466 27571
rect 26430 26149 26466 26781
rect 26430 25359 26466 25991
rect 26430 24569 26466 25201
rect 26430 23779 26466 24411
rect 26430 22989 26466 23621
rect 26430 22199 26466 22831
rect 26430 21409 26466 22041
rect 26430 20619 26466 21251
rect 26430 19829 26466 20461
rect 26430 19039 26466 19671
rect 26430 18249 26466 18881
rect 26430 17459 26466 18091
rect 26430 16669 26466 17301
rect 26430 15879 26466 16511
rect 26430 15089 26466 15721
rect 26430 14299 26466 14931
rect 26430 13509 26466 14141
rect 26430 12719 26466 13351
rect 26430 11929 26466 12561
rect 26430 11139 26466 11771
rect 26430 10349 26466 10981
rect 26430 9559 26466 10191
rect 26430 8769 26466 9401
rect 26430 7979 26466 8611
rect 26430 7189 26466 7821
rect 26430 6399 26466 7031
rect 26430 5609 26466 6241
rect 26430 4819 26466 5451
rect 26430 4029 26466 4661
rect 26430 3239 26466 3871
rect 26430 2449 26466 3081
rect 26430 1659 26466 2291
rect 26430 869 26466 1501
rect 26430 79 26466 711
rect 26502 0 26538 50560
rect 26574 0 26610 50560
rect 27054 0 27090 50560
rect 27126 0 27162 50560
rect 27198 49849 27234 50481
rect 27198 49059 27234 49691
rect 27198 48269 27234 48901
rect 27198 47479 27234 48111
rect 27198 46689 27234 47321
rect 27198 45899 27234 46531
rect 27198 45109 27234 45741
rect 27198 44319 27234 44951
rect 27198 43529 27234 44161
rect 27198 42739 27234 43371
rect 27198 41949 27234 42581
rect 27198 41159 27234 41791
rect 27198 40369 27234 41001
rect 27198 39579 27234 40211
rect 27198 38789 27234 39421
rect 27198 37999 27234 38631
rect 27198 37209 27234 37841
rect 27198 36419 27234 37051
rect 27198 35629 27234 36261
rect 27198 34839 27234 35471
rect 27198 34049 27234 34681
rect 27198 33259 27234 33891
rect 27198 32469 27234 33101
rect 27198 31679 27234 32311
rect 27198 30889 27234 31521
rect 27198 30099 27234 30731
rect 27198 29309 27234 29941
rect 27198 28519 27234 29151
rect 27198 27729 27234 28361
rect 27198 26939 27234 27571
rect 27198 26149 27234 26781
rect 27198 25359 27234 25991
rect 27198 24569 27234 25201
rect 27198 23779 27234 24411
rect 27198 22989 27234 23621
rect 27198 22199 27234 22831
rect 27198 21409 27234 22041
rect 27198 20619 27234 21251
rect 27198 19829 27234 20461
rect 27198 19039 27234 19671
rect 27198 18249 27234 18881
rect 27198 17459 27234 18091
rect 27198 16669 27234 17301
rect 27198 15879 27234 16511
rect 27198 15089 27234 15721
rect 27198 14299 27234 14931
rect 27198 13509 27234 14141
rect 27198 12719 27234 13351
rect 27198 11929 27234 12561
rect 27198 11139 27234 11771
rect 27198 10349 27234 10981
rect 27198 9559 27234 10191
rect 27198 8769 27234 9401
rect 27198 7979 27234 8611
rect 27198 7189 27234 7821
rect 27198 6399 27234 7031
rect 27198 5609 27234 6241
rect 27198 4819 27234 5451
rect 27198 4029 27234 4661
rect 27198 3239 27234 3871
rect 27198 2449 27234 3081
rect 27198 1659 27234 2291
rect 27198 869 27234 1501
rect 27198 79 27234 711
rect 27270 0 27306 50560
rect 27342 0 27378 50560
rect 27534 0 27570 50560
rect 27606 0 27642 50560
rect 27678 49849 27714 50481
rect 27678 49059 27714 49691
rect 27678 48269 27714 48901
rect 27678 47479 27714 48111
rect 27678 46689 27714 47321
rect 27678 45899 27714 46531
rect 27678 45109 27714 45741
rect 27678 44319 27714 44951
rect 27678 43529 27714 44161
rect 27678 42739 27714 43371
rect 27678 41949 27714 42581
rect 27678 41159 27714 41791
rect 27678 40369 27714 41001
rect 27678 39579 27714 40211
rect 27678 38789 27714 39421
rect 27678 37999 27714 38631
rect 27678 37209 27714 37841
rect 27678 36419 27714 37051
rect 27678 35629 27714 36261
rect 27678 34839 27714 35471
rect 27678 34049 27714 34681
rect 27678 33259 27714 33891
rect 27678 32469 27714 33101
rect 27678 31679 27714 32311
rect 27678 30889 27714 31521
rect 27678 30099 27714 30731
rect 27678 29309 27714 29941
rect 27678 28519 27714 29151
rect 27678 27729 27714 28361
rect 27678 26939 27714 27571
rect 27678 26149 27714 26781
rect 27678 25359 27714 25991
rect 27678 24569 27714 25201
rect 27678 23779 27714 24411
rect 27678 22989 27714 23621
rect 27678 22199 27714 22831
rect 27678 21409 27714 22041
rect 27678 20619 27714 21251
rect 27678 19829 27714 20461
rect 27678 19039 27714 19671
rect 27678 18249 27714 18881
rect 27678 17459 27714 18091
rect 27678 16669 27714 17301
rect 27678 15879 27714 16511
rect 27678 15089 27714 15721
rect 27678 14299 27714 14931
rect 27678 13509 27714 14141
rect 27678 12719 27714 13351
rect 27678 11929 27714 12561
rect 27678 11139 27714 11771
rect 27678 10349 27714 10981
rect 27678 9559 27714 10191
rect 27678 8769 27714 9401
rect 27678 7979 27714 8611
rect 27678 7189 27714 7821
rect 27678 6399 27714 7031
rect 27678 5609 27714 6241
rect 27678 4819 27714 5451
rect 27678 4029 27714 4661
rect 27678 3239 27714 3871
rect 27678 2449 27714 3081
rect 27678 1659 27714 2291
rect 27678 869 27714 1501
rect 27678 79 27714 711
rect 27750 0 27786 50560
rect 27822 0 27858 50560
rect 28302 0 28338 50560
rect 28374 0 28410 50560
rect 28446 49849 28482 50481
rect 28446 49059 28482 49691
rect 28446 48269 28482 48901
rect 28446 47479 28482 48111
rect 28446 46689 28482 47321
rect 28446 45899 28482 46531
rect 28446 45109 28482 45741
rect 28446 44319 28482 44951
rect 28446 43529 28482 44161
rect 28446 42739 28482 43371
rect 28446 41949 28482 42581
rect 28446 41159 28482 41791
rect 28446 40369 28482 41001
rect 28446 39579 28482 40211
rect 28446 38789 28482 39421
rect 28446 37999 28482 38631
rect 28446 37209 28482 37841
rect 28446 36419 28482 37051
rect 28446 35629 28482 36261
rect 28446 34839 28482 35471
rect 28446 34049 28482 34681
rect 28446 33259 28482 33891
rect 28446 32469 28482 33101
rect 28446 31679 28482 32311
rect 28446 30889 28482 31521
rect 28446 30099 28482 30731
rect 28446 29309 28482 29941
rect 28446 28519 28482 29151
rect 28446 27729 28482 28361
rect 28446 26939 28482 27571
rect 28446 26149 28482 26781
rect 28446 25359 28482 25991
rect 28446 24569 28482 25201
rect 28446 23779 28482 24411
rect 28446 22989 28482 23621
rect 28446 22199 28482 22831
rect 28446 21409 28482 22041
rect 28446 20619 28482 21251
rect 28446 19829 28482 20461
rect 28446 19039 28482 19671
rect 28446 18249 28482 18881
rect 28446 17459 28482 18091
rect 28446 16669 28482 17301
rect 28446 15879 28482 16511
rect 28446 15089 28482 15721
rect 28446 14299 28482 14931
rect 28446 13509 28482 14141
rect 28446 12719 28482 13351
rect 28446 11929 28482 12561
rect 28446 11139 28482 11771
rect 28446 10349 28482 10981
rect 28446 9559 28482 10191
rect 28446 8769 28482 9401
rect 28446 7979 28482 8611
rect 28446 7189 28482 7821
rect 28446 6399 28482 7031
rect 28446 5609 28482 6241
rect 28446 4819 28482 5451
rect 28446 4029 28482 4661
rect 28446 3239 28482 3871
rect 28446 2449 28482 3081
rect 28446 1659 28482 2291
rect 28446 869 28482 1501
rect 28446 79 28482 711
rect 28518 0 28554 50560
rect 28590 0 28626 50560
rect 28782 0 28818 50560
rect 28854 0 28890 50560
rect 28926 49849 28962 50481
rect 28926 49059 28962 49691
rect 28926 48269 28962 48901
rect 28926 47479 28962 48111
rect 28926 46689 28962 47321
rect 28926 45899 28962 46531
rect 28926 45109 28962 45741
rect 28926 44319 28962 44951
rect 28926 43529 28962 44161
rect 28926 42739 28962 43371
rect 28926 41949 28962 42581
rect 28926 41159 28962 41791
rect 28926 40369 28962 41001
rect 28926 39579 28962 40211
rect 28926 38789 28962 39421
rect 28926 37999 28962 38631
rect 28926 37209 28962 37841
rect 28926 36419 28962 37051
rect 28926 35629 28962 36261
rect 28926 34839 28962 35471
rect 28926 34049 28962 34681
rect 28926 33259 28962 33891
rect 28926 32469 28962 33101
rect 28926 31679 28962 32311
rect 28926 30889 28962 31521
rect 28926 30099 28962 30731
rect 28926 29309 28962 29941
rect 28926 28519 28962 29151
rect 28926 27729 28962 28361
rect 28926 26939 28962 27571
rect 28926 26149 28962 26781
rect 28926 25359 28962 25991
rect 28926 24569 28962 25201
rect 28926 23779 28962 24411
rect 28926 22989 28962 23621
rect 28926 22199 28962 22831
rect 28926 21409 28962 22041
rect 28926 20619 28962 21251
rect 28926 19829 28962 20461
rect 28926 19039 28962 19671
rect 28926 18249 28962 18881
rect 28926 17459 28962 18091
rect 28926 16669 28962 17301
rect 28926 15879 28962 16511
rect 28926 15089 28962 15721
rect 28926 14299 28962 14931
rect 28926 13509 28962 14141
rect 28926 12719 28962 13351
rect 28926 11929 28962 12561
rect 28926 11139 28962 11771
rect 28926 10349 28962 10981
rect 28926 9559 28962 10191
rect 28926 8769 28962 9401
rect 28926 7979 28962 8611
rect 28926 7189 28962 7821
rect 28926 6399 28962 7031
rect 28926 5609 28962 6241
rect 28926 4819 28962 5451
rect 28926 4029 28962 4661
rect 28926 3239 28962 3871
rect 28926 2449 28962 3081
rect 28926 1659 28962 2291
rect 28926 869 28962 1501
rect 28926 79 28962 711
rect 28998 0 29034 50560
rect 29070 0 29106 50560
rect 29550 0 29586 50560
rect 29622 0 29658 50560
rect 29694 49849 29730 50481
rect 29694 49059 29730 49691
rect 29694 48269 29730 48901
rect 29694 47479 29730 48111
rect 29694 46689 29730 47321
rect 29694 45899 29730 46531
rect 29694 45109 29730 45741
rect 29694 44319 29730 44951
rect 29694 43529 29730 44161
rect 29694 42739 29730 43371
rect 29694 41949 29730 42581
rect 29694 41159 29730 41791
rect 29694 40369 29730 41001
rect 29694 39579 29730 40211
rect 29694 38789 29730 39421
rect 29694 37999 29730 38631
rect 29694 37209 29730 37841
rect 29694 36419 29730 37051
rect 29694 35629 29730 36261
rect 29694 34839 29730 35471
rect 29694 34049 29730 34681
rect 29694 33259 29730 33891
rect 29694 32469 29730 33101
rect 29694 31679 29730 32311
rect 29694 30889 29730 31521
rect 29694 30099 29730 30731
rect 29694 29309 29730 29941
rect 29694 28519 29730 29151
rect 29694 27729 29730 28361
rect 29694 26939 29730 27571
rect 29694 26149 29730 26781
rect 29694 25359 29730 25991
rect 29694 24569 29730 25201
rect 29694 23779 29730 24411
rect 29694 22989 29730 23621
rect 29694 22199 29730 22831
rect 29694 21409 29730 22041
rect 29694 20619 29730 21251
rect 29694 19829 29730 20461
rect 29694 19039 29730 19671
rect 29694 18249 29730 18881
rect 29694 17459 29730 18091
rect 29694 16669 29730 17301
rect 29694 15879 29730 16511
rect 29694 15089 29730 15721
rect 29694 14299 29730 14931
rect 29694 13509 29730 14141
rect 29694 12719 29730 13351
rect 29694 11929 29730 12561
rect 29694 11139 29730 11771
rect 29694 10349 29730 10981
rect 29694 9559 29730 10191
rect 29694 8769 29730 9401
rect 29694 7979 29730 8611
rect 29694 7189 29730 7821
rect 29694 6399 29730 7031
rect 29694 5609 29730 6241
rect 29694 4819 29730 5451
rect 29694 4029 29730 4661
rect 29694 3239 29730 3871
rect 29694 2449 29730 3081
rect 29694 1659 29730 2291
rect 29694 869 29730 1501
rect 29694 79 29730 711
rect 29766 0 29802 50560
rect 29838 0 29874 50560
rect 30030 0 30066 50560
rect 30102 0 30138 50560
rect 30174 49849 30210 50481
rect 30174 49059 30210 49691
rect 30174 48269 30210 48901
rect 30174 47479 30210 48111
rect 30174 46689 30210 47321
rect 30174 45899 30210 46531
rect 30174 45109 30210 45741
rect 30174 44319 30210 44951
rect 30174 43529 30210 44161
rect 30174 42739 30210 43371
rect 30174 41949 30210 42581
rect 30174 41159 30210 41791
rect 30174 40369 30210 41001
rect 30174 39579 30210 40211
rect 30174 38789 30210 39421
rect 30174 37999 30210 38631
rect 30174 37209 30210 37841
rect 30174 36419 30210 37051
rect 30174 35629 30210 36261
rect 30174 34839 30210 35471
rect 30174 34049 30210 34681
rect 30174 33259 30210 33891
rect 30174 32469 30210 33101
rect 30174 31679 30210 32311
rect 30174 30889 30210 31521
rect 30174 30099 30210 30731
rect 30174 29309 30210 29941
rect 30174 28519 30210 29151
rect 30174 27729 30210 28361
rect 30174 26939 30210 27571
rect 30174 26149 30210 26781
rect 30174 25359 30210 25991
rect 30174 24569 30210 25201
rect 30174 23779 30210 24411
rect 30174 22989 30210 23621
rect 30174 22199 30210 22831
rect 30174 21409 30210 22041
rect 30174 20619 30210 21251
rect 30174 19829 30210 20461
rect 30174 19039 30210 19671
rect 30174 18249 30210 18881
rect 30174 17459 30210 18091
rect 30174 16669 30210 17301
rect 30174 15879 30210 16511
rect 30174 15089 30210 15721
rect 30174 14299 30210 14931
rect 30174 13509 30210 14141
rect 30174 12719 30210 13351
rect 30174 11929 30210 12561
rect 30174 11139 30210 11771
rect 30174 10349 30210 10981
rect 30174 9559 30210 10191
rect 30174 8769 30210 9401
rect 30174 7979 30210 8611
rect 30174 7189 30210 7821
rect 30174 6399 30210 7031
rect 30174 5609 30210 6241
rect 30174 4819 30210 5451
rect 30174 4029 30210 4661
rect 30174 3239 30210 3871
rect 30174 2449 30210 3081
rect 30174 1659 30210 2291
rect 30174 869 30210 1501
rect 30174 79 30210 711
rect 30246 0 30282 50560
rect 30318 0 30354 50560
rect 30798 0 30834 50560
rect 30870 0 30906 50560
rect 30942 49849 30978 50481
rect 30942 49059 30978 49691
rect 30942 48269 30978 48901
rect 30942 47479 30978 48111
rect 30942 46689 30978 47321
rect 30942 45899 30978 46531
rect 30942 45109 30978 45741
rect 30942 44319 30978 44951
rect 30942 43529 30978 44161
rect 30942 42739 30978 43371
rect 30942 41949 30978 42581
rect 30942 41159 30978 41791
rect 30942 40369 30978 41001
rect 30942 39579 30978 40211
rect 30942 38789 30978 39421
rect 30942 37999 30978 38631
rect 30942 37209 30978 37841
rect 30942 36419 30978 37051
rect 30942 35629 30978 36261
rect 30942 34839 30978 35471
rect 30942 34049 30978 34681
rect 30942 33259 30978 33891
rect 30942 32469 30978 33101
rect 30942 31679 30978 32311
rect 30942 30889 30978 31521
rect 30942 30099 30978 30731
rect 30942 29309 30978 29941
rect 30942 28519 30978 29151
rect 30942 27729 30978 28361
rect 30942 26939 30978 27571
rect 30942 26149 30978 26781
rect 30942 25359 30978 25991
rect 30942 24569 30978 25201
rect 30942 23779 30978 24411
rect 30942 22989 30978 23621
rect 30942 22199 30978 22831
rect 30942 21409 30978 22041
rect 30942 20619 30978 21251
rect 30942 19829 30978 20461
rect 30942 19039 30978 19671
rect 30942 18249 30978 18881
rect 30942 17459 30978 18091
rect 30942 16669 30978 17301
rect 30942 15879 30978 16511
rect 30942 15089 30978 15721
rect 30942 14299 30978 14931
rect 30942 13509 30978 14141
rect 30942 12719 30978 13351
rect 30942 11929 30978 12561
rect 30942 11139 30978 11771
rect 30942 10349 30978 10981
rect 30942 9559 30978 10191
rect 30942 8769 30978 9401
rect 30942 7979 30978 8611
rect 30942 7189 30978 7821
rect 30942 6399 30978 7031
rect 30942 5609 30978 6241
rect 30942 4819 30978 5451
rect 30942 4029 30978 4661
rect 30942 3239 30978 3871
rect 30942 2449 30978 3081
rect 30942 1659 30978 2291
rect 30942 869 30978 1501
rect 30942 79 30978 711
rect 31014 0 31050 50560
rect 31086 0 31122 50560
rect 31278 0 31314 50560
rect 31350 0 31386 50560
rect 31422 49849 31458 50481
rect 31422 49059 31458 49691
rect 31422 48269 31458 48901
rect 31422 47479 31458 48111
rect 31422 46689 31458 47321
rect 31422 45899 31458 46531
rect 31422 45109 31458 45741
rect 31422 44319 31458 44951
rect 31422 43529 31458 44161
rect 31422 42739 31458 43371
rect 31422 41949 31458 42581
rect 31422 41159 31458 41791
rect 31422 40369 31458 41001
rect 31422 39579 31458 40211
rect 31422 38789 31458 39421
rect 31422 37999 31458 38631
rect 31422 37209 31458 37841
rect 31422 36419 31458 37051
rect 31422 35629 31458 36261
rect 31422 34839 31458 35471
rect 31422 34049 31458 34681
rect 31422 33259 31458 33891
rect 31422 32469 31458 33101
rect 31422 31679 31458 32311
rect 31422 30889 31458 31521
rect 31422 30099 31458 30731
rect 31422 29309 31458 29941
rect 31422 28519 31458 29151
rect 31422 27729 31458 28361
rect 31422 26939 31458 27571
rect 31422 26149 31458 26781
rect 31422 25359 31458 25991
rect 31422 24569 31458 25201
rect 31422 23779 31458 24411
rect 31422 22989 31458 23621
rect 31422 22199 31458 22831
rect 31422 21409 31458 22041
rect 31422 20619 31458 21251
rect 31422 19829 31458 20461
rect 31422 19039 31458 19671
rect 31422 18249 31458 18881
rect 31422 17459 31458 18091
rect 31422 16669 31458 17301
rect 31422 15879 31458 16511
rect 31422 15089 31458 15721
rect 31422 14299 31458 14931
rect 31422 13509 31458 14141
rect 31422 12719 31458 13351
rect 31422 11929 31458 12561
rect 31422 11139 31458 11771
rect 31422 10349 31458 10981
rect 31422 9559 31458 10191
rect 31422 8769 31458 9401
rect 31422 7979 31458 8611
rect 31422 7189 31458 7821
rect 31422 6399 31458 7031
rect 31422 5609 31458 6241
rect 31422 4819 31458 5451
rect 31422 4029 31458 4661
rect 31422 3239 31458 3871
rect 31422 2449 31458 3081
rect 31422 1659 31458 2291
rect 31422 869 31458 1501
rect 31422 79 31458 711
rect 31494 0 31530 50560
rect 31566 0 31602 50560
rect 32046 0 32082 50560
rect 32118 0 32154 50560
rect 32190 49849 32226 50481
rect 32190 49059 32226 49691
rect 32190 48269 32226 48901
rect 32190 47479 32226 48111
rect 32190 46689 32226 47321
rect 32190 45899 32226 46531
rect 32190 45109 32226 45741
rect 32190 44319 32226 44951
rect 32190 43529 32226 44161
rect 32190 42739 32226 43371
rect 32190 41949 32226 42581
rect 32190 41159 32226 41791
rect 32190 40369 32226 41001
rect 32190 39579 32226 40211
rect 32190 38789 32226 39421
rect 32190 37999 32226 38631
rect 32190 37209 32226 37841
rect 32190 36419 32226 37051
rect 32190 35629 32226 36261
rect 32190 34839 32226 35471
rect 32190 34049 32226 34681
rect 32190 33259 32226 33891
rect 32190 32469 32226 33101
rect 32190 31679 32226 32311
rect 32190 30889 32226 31521
rect 32190 30099 32226 30731
rect 32190 29309 32226 29941
rect 32190 28519 32226 29151
rect 32190 27729 32226 28361
rect 32190 26939 32226 27571
rect 32190 26149 32226 26781
rect 32190 25359 32226 25991
rect 32190 24569 32226 25201
rect 32190 23779 32226 24411
rect 32190 22989 32226 23621
rect 32190 22199 32226 22831
rect 32190 21409 32226 22041
rect 32190 20619 32226 21251
rect 32190 19829 32226 20461
rect 32190 19039 32226 19671
rect 32190 18249 32226 18881
rect 32190 17459 32226 18091
rect 32190 16669 32226 17301
rect 32190 15879 32226 16511
rect 32190 15089 32226 15721
rect 32190 14299 32226 14931
rect 32190 13509 32226 14141
rect 32190 12719 32226 13351
rect 32190 11929 32226 12561
rect 32190 11139 32226 11771
rect 32190 10349 32226 10981
rect 32190 9559 32226 10191
rect 32190 8769 32226 9401
rect 32190 7979 32226 8611
rect 32190 7189 32226 7821
rect 32190 6399 32226 7031
rect 32190 5609 32226 6241
rect 32190 4819 32226 5451
rect 32190 4029 32226 4661
rect 32190 3239 32226 3871
rect 32190 2449 32226 3081
rect 32190 1659 32226 2291
rect 32190 869 32226 1501
rect 32190 79 32226 711
rect 32262 0 32298 50560
rect 32334 0 32370 50560
rect 32526 0 32562 50560
rect 32598 0 32634 50560
rect 32670 49849 32706 50481
rect 32670 49059 32706 49691
rect 32670 48269 32706 48901
rect 32670 47479 32706 48111
rect 32670 46689 32706 47321
rect 32670 45899 32706 46531
rect 32670 45109 32706 45741
rect 32670 44319 32706 44951
rect 32670 43529 32706 44161
rect 32670 42739 32706 43371
rect 32670 41949 32706 42581
rect 32670 41159 32706 41791
rect 32670 40369 32706 41001
rect 32670 39579 32706 40211
rect 32670 38789 32706 39421
rect 32670 37999 32706 38631
rect 32670 37209 32706 37841
rect 32670 36419 32706 37051
rect 32670 35629 32706 36261
rect 32670 34839 32706 35471
rect 32670 34049 32706 34681
rect 32670 33259 32706 33891
rect 32670 32469 32706 33101
rect 32670 31679 32706 32311
rect 32670 30889 32706 31521
rect 32670 30099 32706 30731
rect 32670 29309 32706 29941
rect 32670 28519 32706 29151
rect 32670 27729 32706 28361
rect 32670 26939 32706 27571
rect 32670 26149 32706 26781
rect 32670 25359 32706 25991
rect 32670 24569 32706 25201
rect 32670 23779 32706 24411
rect 32670 22989 32706 23621
rect 32670 22199 32706 22831
rect 32670 21409 32706 22041
rect 32670 20619 32706 21251
rect 32670 19829 32706 20461
rect 32670 19039 32706 19671
rect 32670 18249 32706 18881
rect 32670 17459 32706 18091
rect 32670 16669 32706 17301
rect 32670 15879 32706 16511
rect 32670 15089 32706 15721
rect 32670 14299 32706 14931
rect 32670 13509 32706 14141
rect 32670 12719 32706 13351
rect 32670 11929 32706 12561
rect 32670 11139 32706 11771
rect 32670 10349 32706 10981
rect 32670 9559 32706 10191
rect 32670 8769 32706 9401
rect 32670 7979 32706 8611
rect 32670 7189 32706 7821
rect 32670 6399 32706 7031
rect 32670 5609 32706 6241
rect 32670 4819 32706 5451
rect 32670 4029 32706 4661
rect 32670 3239 32706 3871
rect 32670 2449 32706 3081
rect 32670 1659 32706 2291
rect 32670 869 32706 1501
rect 32670 79 32706 711
rect 32742 0 32778 50560
rect 32814 0 32850 50560
rect 33294 0 33330 50560
rect 33366 0 33402 50560
rect 33438 49849 33474 50481
rect 33438 49059 33474 49691
rect 33438 48269 33474 48901
rect 33438 47479 33474 48111
rect 33438 46689 33474 47321
rect 33438 45899 33474 46531
rect 33438 45109 33474 45741
rect 33438 44319 33474 44951
rect 33438 43529 33474 44161
rect 33438 42739 33474 43371
rect 33438 41949 33474 42581
rect 33438 41159 33474 41791
rect 33438 40369 33474 41001
rect 33438 39579 33474 40211
rect 33438 38789 33474 39421
rect 33438 37999 33474 38631
rect 33438 37209 33474 37841
rect 33438 36419 33474 37051
rect 33438 35629 33474 36261
rect 33438 34839 33474 35471
rect 33438 34049 33474 34681
rect 33438 33259 33474 33891
rect 33438 32469 33474 33101
rect 33438 31679 33474 32311
rect 33438 30889 33474 31521
rect 33438 30099 33474 30731
rect 33438 29309 33474 29941
rect 33438 28519 33474 29151
rect 33438 27729 33474 28361
rect 33438 26939 33474 27571
rect 33438 26149 33474 26781
rect 33438 25359 33474 25991
rect 33438 24569 33474 25201
rect 33438 23779 33474 24411
rect 33438 22989 33474 23621
rect 33438 22199 33474 22831
rect 33438 21409 33474 22041
rect 33438 20619 33474 21251
rect 33438 19829 33474 20461
rect 33438 19039 33474 19671
rect 33438 18249 33474 18881
rect 33438 17459 33474 18091
rect 33438 16669 33474 17301
rect 33438 15879 33474 16511
rect 33438 15089 33474 15721
rect 33438 14299 33474 14931
rect 33438 13509 33474 14141
rect 33438 12719 33474 13351
rect 33438 11929 33474 12561
rect 33438 11139 33474 11771
rect 33438 10349 33474 10981
rect 33438 9559 33474 10191
rect 33438 8769 33474 9401
rect 33438 7979 33474 8611
rect 33438 7189 33474 7821
rect 33438 6399 33474 7031
rect 33438 5609 33474 6241
rect 33438 4819 33474 5451
rect 33438 4029 33474 4661
rect 33438 3239 33474 3871
rect 33438 2449 33474 3081
rect 33438 1659 33474 2291
rect 33438 869 33474 1501
rect 33438 79 33474 711
rect 33510 0 33546 50560
rect 33582 0 33618 50560
rect 33774 0 33810 50560
rect 33846 0 33882 50560
rect 33918 49849 33954 50481
rect 33918 49059 33954 49691
rect 33918 48269 33954 48901
rect 33918 47479 33954 48111
rect 33918 46689 33954 47321
rect 33918 45899 33954 46531
rect 33918 45109 33954 45741
rect 33918 44319 33954 44951
rect 33918 43529 33954 44161
rect 33918 42739 33954 43371
rect 33918 41949 33954 42581
rect 33918 41159 33954 41791
rect 33918 40369 33954 41001
rect 33918 39579 33954 40211
rect 33918 38789 33954 39421
rect 33918 37999 33954 38631
rect 33918 37209 33954 37841
rect 33918 36419 33954 37051
rect 33918 35629 33954 36261
rect 33918 34839 33954 35471
rect 33918 34049 33954 34681
rect 33918 33259 33954 33891
rect 33918 32469 33954 33101
rect 33918 31679 33954 32311
rect 33918 30889 33954 31521
rect 33918 30099 33954 30731
rect 33918 29309 33954 29941
rect 33918 28519 33954 29151
rect 33918 27729 33954 28361
rect 33918 26939 33954 27571
rect 33918 26149 33954 26781
rect 33918 25359 33954 25991
rect 33918 24569 33954 25201
rect 33918 23779 33954 24411
rect 33918 22989 33954 23621
rect 33918 22199 33954 22831
rect 33918 21409 33954 22041
rect 33918 20619 33954 21251
rect 33918 19829 33954 20461
rect 33918 19039 33954 19671
rect 33918 18249 33954 18881
rect 33918 17459 33954 18091
rect 33918 16669 33954 17301
rect 33918 15879 33954 16511
rect 33918 15089 33954 15721
rect 33918 14299 33954 14931
rect 33918 13509 33954 14141
rect 33918 12719 33954 13351
rect 33918 11929 33954 12561
rect 33918 11139 33954 11771
rect 33918 10349 33954 10981
rect 33918 9559 33954 10191
rect 33918 8769 33954 9401
rect 33918 7979 33954 8611
rect 33918 7189 33954 7821
rect 33918 6399 33954 7031
rect 33918 5609 33954 6241
rect 33918 4819 33954 5451
rect 33918 4029 33954 4661
rect 33918 3239 33954 3871
rect 33918 2449 33954 3081
rect 33918 1659 33954 2291
rect 33918 869 33954 1501
rect 33918 79 33954 711
rect 33990 0 34026 50560
rect 34062 0 34098 50560
rect 34542 0 34578 50560
rect 34614 0 34650 50560
rect 34686 49849 34722 50481
rect 34686 49059 34722 49691
rect 34686 48269 34722 48901
rect 34686 47479 34722 48111
rect 34686 46689 34722 47321
rect 34686 45899 34722 46531
rect 34686 45109 34722 45741
rect 34686 44319 34722 44951
rect 34686 43529 34722 44161
rect 34686 42739 34722 43371
rect 34686 41949 34722 42581
rect 34686 41159 34722 41791
rect 34686 40369 34722 41001
rect 34686 39579 34722 40211
rect 34686 38789 34722 39421
rect 34686 37999 34722 38631
rect 34686 37209 34722 37841
rect 34686 36419 34722 37051
rect 34686 35629 34722 36261
rect 34686 34839 34722 35471
rect 34686 34049 34722 34681
rect 34686 33259 34722 33891
rect 34686 32469 34722 33101
rect 34686 31679 34722 32311
rect 34686 30889 34722 31521
rect 34686 30099 34722 30731
rect 34686 29309 34722 29941
rect 34686 28519 34722 29151
rect 34686 27729 34722 28361
rect 34686 26939 34722 27571
rect 34686 26149 34722 26781
rect 34686 25359 34722 25991
rect 34686 24569 34722 25201
rect 34686 23779 34722 24411
rect 34686 22989 34722 23621
rect 34686 22199 34722 22831
rect 34686 21409 34722 22041
rect 34686 20619 34722 21251
rect 34686 19829 34722 20461
rect 34686 19039 34722 19671
rect 34686 18249 34722 18881
rect 34686 17459 34722 18091
rect 34686 16669 34722 17301
rect 34686 15879 34722 16511
rect 34686 15089 34722 15721
rect 34686 14299 34722 14931
rect 34686 13509 34722 14141
rect 34686 12719 34722 13351
rect 34686 11929 34722 12561
rect 34686 11139 34722 11771
rect 34686 10349 34722 10981
rect 34686 9559 34722 10191
rect 34686 8769 34722 9401
rect 34686 7979 34722 8611
rect 34686 7189 34722 7821
rect 34686 6399 34722 7031
rect 34686 5609 34722 6241
rect 34686 4819 34722 5451
rect 34686 4029 34722 4661
rect 34686 3239 34722 3871
rect 34686 2449 34722 3081
rect 34686 1659 34722 2291
rect 34686 869 34722 1501
rect 34686 79 34722 711
rect 34758 0 34794 50560
rect 34830 0 34866 50560
rect 35022 0 35058 50560
rect 35094 0 35130 50560
rect 35166 49849 35202 50481
rect 35166 49059 35202 49691
rect 35166 48269 35202 48901
rect 35166 47479 35202 48111
rect 35166 46689 35202 47321
rect 35166 45899 35202 46531
rect 35166 45109 35202 45741
rect 35166 44319 35202 44951
rect 35166 43529 35202 44161
rect 35166 42739 35202 43371
rect 35166 41949 35202 42581
rect 35166 41159 35202 41791
rect 35166 40369 35202 41001
rect 35166 39579 35202 40211
rect 35166 38789 35202 39421
rect 35166 37999 35202 38631
rect 35166 37209 35202 37841
rect 35166 36419 35202 37051
rect 35166 35629 35202 36261
rect 35166 34839 35202 35471
rect 35166 34049 35202 34681
rect 35166 33259 35202 33891
rect 35166 32469 35202 33101
rect 35166 31679 35202 32311
rect 35166 30889 35202 31521
rect 35166 30099 35202 30731
rect 35166 29309 35202 29941
rect 35166 28519 35202 29151
rect 35166 27729 35202 28361
rect 35166 26939 35202 27571
rect 35166 26149 35202 26781
rect 35166 25359 35202 25991
rect 35166 24569 35202 25201
rect 35166 23779 35202 24411
rect 35166 22989 35202 23621
rect 35166 22199 35202 22831
rect 35166 21409 35202 22041
rect 35166 20619 35202 21251
rect 35166 19829 35202 20461
rect 35166 19039 35202 19671
rect 35166 18249 35202 18881
rect 35166 17459 35202 18091
rect 35166 16669 35202 17301
rect 35166 15879 35202 16511
rect 35166 15089 35202 15721
rect 35166 14299 35202 14931
rect 35166 13509 35202 14141
rect 35166 12719 35202 13351
rect 35166 11929 35202 12561
rect 35166 11139 35202 11771
rect 35166 10349 35202 10981
rect 35166 9559 35202 10191
rect 35166 8769 35202 9401
rect 35166 7979 35202 8611
rect 35166 7189 35202 7821
rect 35166 6399 35202 7031
rect 35166 5609 35202 6241
rect 35166 4819 35202 5451
rect 35166 4029 35202 4661
rect 35166 3239 35202 3871
rect 35166 2449 35202 3081
rect 35166 1659 35202 2291
rect 35166 869 35202 1501
rect 35166 79 35202 711
rect 35238 0 35274 50560
rect 35310 0 35346 50560
rect 35790 0 35826 50560
rect 35862 0 35898 50560
rect 35934 49849 35970 50481
rect 35934 49059 35970 49691
rect 35934 48269 35970 48901
rect 35934 47479 35970 48111
rect 35934 46689 35970 47321
rect 35934 45899 35970 46531
rect 35934 45109 35970 45741
rect 35934 44319 35970 44951
rect 35934 43529 35970 44161
rect 35934 42739 35970 43371
rect 35934 41949 35970 42581
rect 35934 41159 35970 41791
rect 35934 40369 35970 41001
rect 35934 39579 35970 40211
rect 35934 38789 35970 39421
rect 35934 37999 35970 38631
rect 35934 37209 35970 37841
rect 35934 36419 35970 37051
rect 35934 35629 35970 36261
rect 35934 34839 35970 35471
rect 35934 34049 35970 34681
rect 35934 33259 35970 33891
rect 35934 32469 35970 33101
rect 35934 31679 35970 32311
rect 35934 30889 35970 31521
rect 35934 30099 35970 30731
rect 35934 29309 35970 29941
rect 35934 28519 35970 29151
rect 35934 27729 35970 28361
rect 35934 26939 35970 27571
rect 35934 26149 35970 26781
rect 35934 25359 35970 25991
rect 35934 24569 35970 25201
rect 35934 23779 35970 24411
rect 35934 22989 35970 23621
rect 35934 22199 35970 22831
rect 35934 21409 35970 22041
rect 35934 20619 35970 21251
rect 35934 19829 35970 20461
rect 35934 19039 35970 19671
rect 35934 18249 35970 18881
rect 35934 17459 35970 18091
rect 35934 16669 35970 17301
rect 35934 15879 35970 16511
rect 35934 15089 35970 15721
rect 35934 14299 35970 14931
rect 35934 13509 35970 14141
rect 35934 12719 35970 13351
rect 35934 11929 35970 12561
rect 35934 11139 35970 11771
rect 35934 10349 35970 10981
rect 35934 9559 35970 10191
rect 35934 8769 35970 9401
rect 35934 7979 35970 8611
rect 35934 7189 35970 7821
rect 35934 6399 35970 7031
rect 35934 5609 35970 6241
rect 35934 4819 35970 5451
rect 35934 4029 35970 4661
rect 35934 3239 35970 3871
rect 35934 2449 35970 3081
rect 35934 1659 35970 2291
rect 35934 869 35970 1501
rect 35934 79 35970 711
rect 36006 0 36042 50560
rect 36078 0 36114 50560
rect 36270 0 36306 50560
rect 36342 0 36378 50560
rect 36414 49849 36450 50481
rect 36414 49059 36450 49691
rect 36414 48269 36450 48901
rect 36414 47479 36450 48111
rect 36414 46689 36450 47321
rect 36414 45899 36450 46531
rect 36414 45109 36450 45741
rect 36414 44319 36450 44951
rect 36414 43529 36450 44161
rect 36414 42739 36450 43371
rect 36414 41949 36450 42581
rect 36414 41159 36450 41791
rect 36414 40369 36450 41001
rect 36414 39579 36450 40211
rect 36414 38789 36450 39421
rect 36414 37999 36450 38631
rect 36414 37209 36450 37841
rect 36414 36419 36450 37051
rect 36414 35629 36450 36261
rect 36414 34839 36450 35471
rect 36414 34049 36450 34681
rect 36414 33259 36450 33891
rect 36414 32469 36450 33101
rect 36414 31679 36450 32311
rect 36414 30889 36450 31521
rect 36414 30099 36450 30731
rect 36414 29309 36450 29941
rect 36414 28519 36450 29151
rect 36414 27729 36450 28361
rect 36414 26939 36450 27571
rect 36414 26149 36450 26781
rect 36414 25359 36450 25991
rect 36414 24569 36450 25201
rect 36414 23779 36450 24411
rect 36414 22989 36450 23621
rect 36414 22199 36450 22831
rect 36414 21409 36450 22041
rect 36414 20619 36450 21251
rect 36414 19829 36450 20461
rect 36414 19039 36450 19671
rect 36414 18249 36450 18881
rect 36414 17459 36450 18091
rect 36414 16669 36450 17301
rect 36414 15879 36450 16511
rect 36414 15089 36450 15721
rect 36414 14299 36450 14931
rect 36414 13509 36450 14141
rect 36414 12719 36450 13351
rect 36414 11929 36450 12561
rect 36414 11139 36450 11771
rect 36414 10349 36450 10981
rect 36414 9559 36450 10191
rect 36414 8769 36450 9401
rect 36414 7979 36450 8611
rect 36414 7189 36450 7821
rect 36414 6399 36450 7031
rect 36414 5609 36450 6241
rect 36414 4819 36450 5451
rect 36414 4029 36450 4661
rect 36414 3239 36450 3871
rect 36414 2449 36450 3081
rect 36414 1659 36450 2291
rect 36414 869 36450 1501
rect 36414 79 36450 711
rect 36486 0 36522 50560
rect 36558 0 36594 50560
rect 37038 0 37074 50560
rect 37110 0 37146 50560
rect 37182 49849 37218 50481
rect 37182 49059 37218 49691
rect 37182 48269 37218 48901
rect 37182 47479 37218 48111
rect 37182 46689 37218 47321
rect 37182 45899 37218 46531
rect 37182 45109 37218 45741
rect 37182 44319 37218 44951
rect 37182 43529 37218 44161
rect 37182 42739 37218 43371
rect 37182 41949 37218 42581
rect 37182 41159 37218 41791
rect 37182 40369 37218 41001
rect 37182 39579 37218 40211
rect 37182 38789 37218 39421
rect 37182 37999 37218 38631
rect 37182 37209 37218 37841
rect 37182 36419 37218 37051
rect 37182 35629 37218 36261
rect 37182 34839 37218 35471
rect 37182 34049 37218 34681
rect 37182 33259 37218 33891
rect 37182 32469 37218 33101
rect 37182 31679 37218 32311
rect 37182 30889 37218 31521
rect 37182 30099 37218 30731
rect 37182 29309 37218 29941
rect 37182 28519 37218 29151
rect 37182 27729 37218 28361
rect 37182 26939 37218 27571
rect 37182 26149 37218 26781
rect 37182 25359 37218 25991
rect 37182 24569 37218 25201
rect 37182 23779 37218 24411
rect 37182 22989 37218 23621
rect 37182 22199 37218 22831
rect 37182 21409 37218 22041
rect 37182 20619 37218 21251
rect 37182 19829 37218 20461
rect 37182 19039 37218 19671
rect 37182 18249 37218 18881
rect 37182 17459 37218 18091
rect 37182 16669 37218 17301
rect 37182 15879 37218 16511
rect 37182 15089 37218 15721
rect 37182 14299 37218 14931
rect 37182 13509 37218 14141
rect 37182 12719 37218 13351
rect 37182 11929 37218 12561
rect 37182 11139 37218 11771
rect 37182 10349 37218 10981
rect 37182 9559 37218 10191
rect 37182 8769 37218 9401
rect 37182 7979 37218 8611
rect 37182 7189 37218 7821
rect 37182 6399 37218 7031
rect 37182 5609 37218 6241
rect 37182 4819 37218 5451
rect 37182 4029 37218 4661
rect 37182 3239 37218 3871
rect 37182 2449 37218 3081
rect 37182 1659 37218 2291
rect 37182 869 37218 1501
rect 37182 79 37218 711
rect 37254 0 37290 50560
rect 37326 0 37362 50560
rect 37518 0 37554 50560
rect 37590 0 37626 50560
rect 37662 49849 37698 50481
rect 37662 49059 37698 49691
rect 37662 48269 37698 48901
rect 37662 47479 37698 48111
rect 37662 46689 37698 47321
rect 37662 45899 37698 46531
rect 37662 45109 37698 45741
rect 37662 44319 37698 44951
rect 37662 43529 37698 44161
rect 37662 42739 37698 43371
rect 37662 41949 37698 42581
rect 37662 41159 37698 41791
rect 37662 40369 37698 41001
rect 37662 39579 37698 40211
rect 37662 38789 37698 39421
rect 37662 37999 37698 38631
rect 37662 37209 37698 37841
rect 37662 36419 37698 37051
rect 37662 35629 37698 36261
rect 37662 34839 37698 35471
rect 37662 34049 37698 34681
rect 37662 33259 37698 33891
rect 37662 32469 37698 33101
rect 37662 31679 37698 32311
rect 37662 30889 37698 31521
rect 37662 30099 37698 30731
rect 37662 29309 37698 29941
rect 37662 28519 37698 29151
rect 37662 27729 37698 28361
rect 37662 26939 37698 27571
rect 37662 26149 37698 26781
rect 37662 25359 37698 25991
rect 37662 24569 37698 25201
rect 37662 23779 37698 24411
rect 37662 22989 37698 23621
rect 37662 22199 37698 22831
rect 37662 21409 37698 22041
rect 37662 20619 37698 21251
rect 37662 19829 37698 20461
rect 37662 19039 37698 19671
rect 37662 18249 37698 18881
rect 37662 17459 37698 18091
rect 37662 16669 37698 17301
rect 37662 15879 37698 16511
rect 37662 15089 37698 15721
rect 37662 14299 37698 14931
rect 37662 13509 37698 14141
rect 37662 12719 37698 13351
rect 37662 11929 37698 12561
rect 37662 11139 37698 11771
rect 37662 10349 37698 10981
rect 37662 9559 37698 10191
rect 37662 8769 37698 9401
rect 37662 7979 37698 8611
rect 37662 7189 37698 7821
rect 37662 6399 37698 7031
rect 37662 5609 37698 6241
rect 37662 4819 37698 5451
rect 37662 4029 37698 4661
rect 37662 3239 37698 3871
rect 37662 2449 37698 3081
rect 37662 1659 37698 2291
rect 37662 869 37698 1501
rect 37662 79 37698 711
rect 37734 0 37770 50560
rect 37806 0 37842 50560
rect 38286 0 38322 50560
rect 38358 0 38394 50560
rect 38430 49849 38466 50481
rect 38430 49059 38466 49691
rect 38430 48269 38466 48901
rect 38430 47479 38466 48111
rect 38430 46689 38466 47321
rect 38430 45899 38466 46531
rect 38430 45109 38466 45741
rect 38430 44319 38466 44951
rect 38430 43529 38466 44161
rect 38430 42739 38466 43371
rect 38430 41949 38466 42581
rect 38430 41159 38466 41791
rect 38430 40369 38466 41001
rect 38430 39579 38466 40211
rect 38430 38789 38466 39421
rect 38430 37999 38466 38631
rect 38430 37209 38466 37841
rect 38430 36419 38466 37051
rect 38430 35629 38466 36261
rect 38430 34839 38466 35471
rect 38430 34049 38466 34681
rect 38430 33259 38466 33891
rect 38430 32469 38466 33101
rect 38430 31679 38466 32311
rect 38430 30889 38466 31521
rect 38430 30099 38466 30731
rect 38430 29309 38466 29941
rect 38430 28519 38466 29151
rect 38430 27729 38466 28361
rect 38430 26939 38466 27571
rect 38430 26149 38466 26781
rect 38430 25359 38466 25991
rect 38430 24569 38466 25201
rect 38430 23779 38466 24411
rect 38430 22989 38466 23621
rect 38430 22199 38466 22831
rect 38430 21409 38466 22041
rect 38430 20619 38466 21251
rect 38430 19829 38466 20461
rect 38430 19039 38466 19671
rect 38430 18249 38466 18881
rect 38430 17459 38466 18091
rect 38430 16669 38466 17301
rect 38430 15879 38466 16511
rect 38430 15089 38466 15721
rect 38430 14299 38466 14931
rect 38430 13509 38466 14141
rect 38430 12719 38466 13351
rect 38430 11929 38466 12561
rect 38430 11139 38466 11771
rect 38430 10349 38466 10981
rect 38430 9559 38466 10191
rect 38430 8769 38466 9401
rect 38430 7979 38466 8611
rect 38430 7189 38466 7821
rect 38430 6399 38466 7031
rect 38430 5609 38466 6241
rect 38430 4819 38466 5451
rect 38430 4029 38466 4661
rect 38430 3239 38466 3871
rect 38430 2449 38466 3081
rect 38430 1659 38466 2291
rect 38430 869 38466 1501
rect 38430 79 38466 711
rect 38502 0 38538 50560
rect 38574 0 38610 50560
rect 38766 0 38802 50560
rect 38838 0 38874 50560
rect 38910 49849 38946 50481
rect 38910 49059 38946 49691
rect 38910 48269 38946 48901
rect 38910 47479 38946 48111
rect 38910 46689 38946 47321
rect 38910 45899 38946 46531
rect 38910 45109 38946 45741
rect 38910 44319 38946 44951
rect 38910 43529 38946 44161
rect 38910 42739 38946 43371
rect 38910 41949 38946 42581
rect 38910 41159 38946 41791
rect 38910 40369 38946 41001
rect 38910 39579 38946 40211
rect 38910 38789 38946 39421
rect 38910 37999 38946 38631
rect 38910 37209 38946 37841
rect 38910 36419 38946 37051
rect 38910 35629 38946 36261
rect 38910 34839 38946 35471
rect 38910 34049 38946 34681
rect 38910 33259 38946 33891
rect 38910 32469 38946 33101
rect 38910 31679 38946 32311
rect 38910 30889 38946 31521
rect 38910 30099 38946 30731
rect 38910 29309 38946 29941
rect 38910 28519 38946 29151
rect 38910 27729 38946 28361
rect 38910 26939 38946 27571
rect 38910 26149 38946 26781
rect 38910 25359 38946 25991
rect 38910 24569 38946 25201
rect 38910 23779 38946 24411
rect 38910 22989 38946 23621
rect 38910 22199 38946 22831
rect 38910 21409 38946 22041
rect 38910 20619 38946 21251
rect 38910 19829 38946 20461
rect 38910 19039 38946 19671
rect 38910 18249 38946 18881
rect 38910 17459 38946 18091
rect 38910 16669 38946 17301
rect 38910 15879 38946 16511
rect 38910 15089 38946 15721
rect 38910 14299 38946 14931
rect 38910 13509 38946 14141
rect 38910 12719 38946 13351
rect 38910 11929 38946 12561
rect 38910 11139 38946 11771
rect 38910 10349 38946 10981
rect 38910 9559 38946 10191
rect 38910 8769 38946 9401
rect 38910 7979 38946 8611
rect 38910 7189 38946 7821
rect 38910 6399 38946 7031
rect 38910 5609 38946 6241
rect 38910 4819 38946 5451
rect 38910 4029 38946 4661
rect 38910 3239 38946 3871
rect 38910 2449 38946 3081
rect 38910 1659 38946 2291
rect 38910 869 38946 1501
rect 38910 79 38946 711
rect 38982 0 39018 50560
rect 39054 0 39090 50560
rect 39534 0 39570 50560
rect 39606 0 39642 50560
rect 39678 49849 39714 50481
rect 39678 49059 39714 49691
rect 39678 48269 39714 48901
rect 39678 47479 39714 48111
rect 39678 46689 39714 47321
rect 39678 45899 39714 46531
rect 39678 45109 39714 45741
rect 39678 44319 39714 44951
rect 39678 43529 39714 44161
rect 39678 42739 39714 43371
rect 39678 41949 39714 42581
rect 39678 41159 39714 41791
rect 39678 40369 39714 41001
rect 39678 39579 39714 40211
rect 39678 38789 39714 39421
rect 39678 37999 39714 38631
rect 39678 37209 39714 37841
rect 39678 36419 39714 37051
rect 39678 35629 39714 36261
rect 39678 34839 39714 35471
rect 39678 34049 39714 34681
rect 39678 33259 39714 33891
rect 39678 32469 39714 33101
rect 39678 31679 39714 32311
rect 39678 30889 39714 31521
rect 39678 30099 39714 30731
rect 39678 29309 39714 29941
rect 39678 28519 39714 29151
rect 39678 27729 39714 28361
rect 39678 26939 39714 27571
rect 39678 26149 39714 26781
rect 39678 25359 39714 25991
rect 39678 24569 39714 25201
rect 39678 23779 39714 24411
rect 39678 22989 39714 23621
rect 39678 22199 39714 22831
rect 39678 21409 39714 22041
rect 39678 20619 39714 21251
rect 39678 19829 39714 20461
rect 39678 19039 39714 19671
rect 39678 18249 39714 18881
rect 39678 17459 39714 18091
rect 39678 16669 39714 17301
rect 39678 15879 39714 16511
rect 39678 15089 39714 15721
rect 39678 14299 39714 14931
rect 39678 13509 39714 14141
rect 39678 12719 39714 13351
rect 39678 11929 39714 12561
rect 39678 11139 39714 11771
rect 39678 10349 39714 10981
rect 39678 9559 39714 10191
rect 39678 8769 39714 9401
rect 39678 7979 39714 8611
rect 39678 7189 39714 7821
rect 39678 6399 39714 7031
rect 39678 5609 39714 6241
rect 39678 4819 39714 5451
rect 39678 4029 39714 4661
rect 39678 3239 39714 3871
rect 39678 2449 39714 3081
rect 39678 1659 39714 2291
rect 39678 869 39714 1501
rect 39678 79 39714 711
rect 39750 0 39786 50560
rect 39822 0 39858 50560
<< metal2 >>
rect 186 50505 294 50615
rect 954 50505 1062 50615
rect 1434 50505 1542 50615
rect 2202 50505 2310 50615
rect 2682 50505 2790 50615
rect 3450 50505 3558 50615
rect 3930 50505 4038 50615
rect 4698 50505 4806 50615
rect 5178 50505 5286 50615
rect 5946 50505 6054 50615
rect 6426 50505 6534 50615
rect 7194 50505 7302 50615
rect 7674 50505 7782 50615
rect 8442 50505 8550 50615
rect 8922 50505 9030 50615
rect 9690 50505 9798 50615
rect 10170 50505 10278 50615
rect 10938 50505 11046 50615
rect 11418 50505 11526 50615
rect 12186 50505 12294 50615
rect 12666 50505 12774 50615
rect 13434 50505 13542 50615
rect 13914 50505 14022 50615
rect 14682 50505 14790 50615
rect 15162 50505 15270 50615
rect 15930 50505 16038 50615
rect 16410 50505 16518 50615
rect 17178 50505 17286 50615
rect 17658 50505 17766 50615
rect 18426 50505 18534 50615
rect 18906 50505 19014 50615
rect 19674 50505 19782 50615
rect 20154 50505 20262 50615
rect 20922 50505 21030 50615
rect 21402 50505 21510 50615
rect 22170 50505 22278 50615
rect 22650 50505 22758 50615
rect 23418 50505 23526 50615
rect 23898 50505 24006 50615
rect 24666 50505 24774 50615
rect 25146 50505 25254 50615
rect 25914 50505 26022 50615
rect 26394 50505 26502 50615
rect 27162 50505 27270 50615
rect 27642 50505 27750 50615
rect 28410 50505 28518 50615
rect 28890 50505 28998 50615
rect 29658 50505 29766 50615
rect 30138 50505 30246 50615
rect 30906 50505 31014 50615
rect 31386 50505 31494 50615
rect 32154 50505 32262 50615
rect 32634 50505 32742 50615
rect 33402 50505 33510 50615
rect 33882 50505 33990 50615
rect 34650 50505 34758 50615
rect 35130 50505 35238 50615
rect 35898 50505 36006 50615
rect 36378 50505 36486 50615
rect 37146 50505 37254 50615
rect 37626 50505 37734 50615
rect 38394 50505 38502 50615
rect 38874 50505 38982 50615
rect 39642 50505 39750 50615
rect 0 50409 39936 50457
rect 186 50285 294 50361
rect 954 50285 1062 50361
rect 1434 50285 1542 50361
rect 2202 50285 2310 50361
rect 2682 50285 2790 50361
rect 3450 50285 3558 50361
rect 3930 50285 4038 50361
rect 4698 50285 4806 50361
rect 5178 50285 5286 50361
rect 5946 50285 6054 50361
rect 6426 50285 6534 50361
rect 7194 50285 7302 50361
rect 7674 50285 7782 50361
rect 8442 50285 8550 50361
rect 8922 50285 9030 50361
rect 9690 50285 9798 50361
rect 10170 50285 10278 50361
rect 10938 50285 11046 50361
rect 11418 50285 11526 50361
rect 12186 50285 12294 50361
rect 12666 50285 12774 50361
rect 13434 50285 13542 50361
rect 13914 50285 14022 50361
rect 14682 50285 14790 50361
rect 15162 50285 15270 50361
rect 15930 50285 16038 50361
rect 16410 50285 16518 50361
rect 17178 50285 17286 50361
rect 17658 50285 17766 50361
rect 18426 50285 18534 50361
rect 18906 50285 19014 50361
rect 19674 50285 19782 50361
rect 20154 50285 20262 50361
rect 20922 50285 21030 50361
rect 21402 50285 21510 50361
rect 22170 50285 22278 50361
rect 22650 50285 22758 50361
rect 23418 50285 23526 50361
rect 23898 50285 24006 50361
rect 24666 50285 24774 50361
rect 25146 50285 25254 50361
rect 25914 50285 26022 50361
rect 26394 50285 26502 50361
rect 27162 50285 27270 50361
rect 27642 50285 27750 50361
rect 28410 50285 28518 50361
rect 28890 50285 28998 50361
rect 29658 50285 29766 50361
rect 30138 50285 30246 50361
rect 30906 50285 31014 50361
rect 31386 50285 31494 50361
rect 32154 50285 32262 50361
rect 32634 50285 32742 50361
rect 33402 50285 33510 50361
rect 33882 50285 33990 50361
rect 34650 50285 34758 50361
rect 35130 50285 35238 50361
rect 35898 50285 36006 50361
rect 36378 50285 36486 50361
rect 37146 50285 37254 50361
rect 37626 50285 37734 50361
rect 38394 50285 38502 50361
rect 38874 50285 38982 50361
rect 39642 50285 39750 50361
rect 0 50189 39936 50237
rect 0 50093 39936 50141
rect 186 49969 294 50045
rect 954 49969 1062 50045
rect 1434 49969 1542 50045
rect 2202 49969 2310 50045
rect 2682 49969 2790 50045
rect 3450 49969 3558 50045
rect 3930 49969 4038 50045
rect 4698 49969 4806 50045
rect 5178 49969 5286 50045
rect 5946 49969 6054 50045
rect 6426 49969 6534 50045
rect 7194 49969 7302 50045
rect 7674 49969 7782 50045
rect 8442 49969 8550 50045
rect 8922 49969 9030 50045
rect 9690 49969 9798 50045
rect 10170 49969 10278 50045
rect 10938 49969 11046 50045
rect 11418 49969 11526 50045
rect 12186 49969 12294 50045
rect 12666 49969 12774 50045
rect 13434 49969 13542 50045
rect 13914 49969 14022 50045
rect 14682 49969 14790 50045
rect 15162 49969 15270 50045
rect 15930 49969 16038 50045
rect 16410 49969 16518 50045
rect 17178 49969 17286 50045
rect 17658 49969 17766 50045
rect 18426 49969 18534 50045
rect 18906 49969 19014 50045
rect 19674 49969 19782 50045
rect 20154 49969 20262 50045
rect 20922 49969 21030 50045
rect 21402 49969 21510 50045
rect 22170 49969 22278 50045
rect 22650 49969 22758 50045
rect 23418 49969 23526 50045
rect 23898 49969 24006 50045
rect 24666 49969 24774 50045
rect 25146 49969 25254 50045
rect 25914 49969 26022 50045
rect 26394 49969 26502 50045
rect 27162 49969 27270 50045
rect 27642 49969 27750 50045
rect 28410 49969 28518 50045
rect 28890 49969 28998 50045
rect 29658 49969 29766 50045
rect 30138 49969 30246 50045
rect 30906 49969 31014 50045
rect 31386 49969 31494 50045
rect 32154 49969 32262 50045
rect 32634 49969 32742 50045
rect 33402 49969 33510 50045
rect 33882 49969 33990 50045
rect 34650 49969 34758 50045
rect 35130 49969 35238 50045
rect 35898 49969 36006 50045
rect 36378 49969 36486 50045
rect 37146 49969 37254 50045
rect 37626 49969 37734 50045
rect 38394 49969 38502 50045
rect 38874 49969 38982 50045
rect 39642 49969 39750 50045
rect 0 49873 39936 49921
rect 186 49715 294 49825
rect 954 49715 1062 49825
rect 1434 49715 1542 49825
rect 2202 49715 2310 49825
rect 2682 49715 2790 49825
rect 3450 49715 3558 49825
rect 3930 49715 4038 49825
rect 4698 49715 4806 49825
rect 5178 49715 5286 49825
rect 5946 49715 6054 49825
rect 6426 49715 6534 49825
rect 7194 49715 7302 49825
rect 7674 49715 7782 49825
rect 8442 49715 8550 49825
rect 8922 49715 9030 49825
rect 9690 49715 9798 49825
rect 10170 49715 10278 49825
rect 10938 49715 11046 49825
rect 11418 49715 11526 49825
rect 12186 49715 12294 49825
rect 12666 49715 12774 49825
rect 13434 49715 13542 49825
rect 13914 49715 14022 49825
rect 14682 49715 14790 49825
rect 15162 49715 15270 49825
rect 15930 49715 16038 49825
rect 16410 49715 16518 49825
rect 17178 49715 17286 49825
rect 17658 49715 17766 49825
rect 18426 49715 18534 49825
rect 18906 49715 19014 49825
rect 19674 49715 19782 49825
rect 20154 49715 20262 49825
rect 20922 49715 21030 49825
rect 21402 49715 21510 49825
rect 22170 49715 22278 49825
rect 22650 49715 22758 49825
rect 23418 49715 23526 49825
rect 23898 49715 24006 49825
rect 24666 49715 24774 49825
rect 25146 49715 25254 49825
rect 25914 49715 26022 49825
rect 26394 49715 26502 49825
rect 27162 49715 27270 49825
rect 27642 49715 27750 49825
rect 28410 49715 28518 49825
rect 28890 49715 28998 49825
rect 29658 49715 29766 49825
rect 30138 49715 30246 49825
rect 30906 49715 31014 49825
rect 31386 49715 31494 49825
rect 32154 49715 32262 49825
rect 32634 49715 32742 49825
rect 33402 49715 33510 49825
rect 33882 49715 33990 49825
rect 34650 49715 34758 49825
rect 35130 49715 35238 49825
rect 35898 49715 36006 49825
rect 36378 49715 36486 49825
rect 37146 49715 37254 49825
rect 37626 49715 37734 49825
rect 38394 49715 38502 49825
rect 38874 49715 38982 49825
rect 39642 49715 39750 49825
rect 0 49619 39936 49667
rect 186 49495 294 49571
rect 954 49495 1062 49571
rect 1434 49495 1542 49571
rect 2202 49495 2310 49571
rect 2682 49495 2790 49571
rect 3450 49495 3558 49571
rect 3930 49495 4038 49571
rect 4698 49495 4806 49571
rect 5178 49495 5286 49571
rect 5946 49495 6054 49571
rect 6426 49495 6534 49571
rect 7194 49495 7302 49571
rect 7674 49495 7782 49571
rect 8442 49495 8550 49571
rect 8922 49495 9030 49571
rect 9690 49495 9798 49571
rect 10170 49495 10278 49571
rect 10938 49495 11046 49571
rect 11418 49495 11526 49571
rect 12186 49495 12294 49571
rect 12666 49495 12774 49571
rect 13434 49495 13542 49571
rect 13914 49495 14022 49571
rect 14682 49495 14790 49571
rect 15162 49495 15270 49571
rect 15930 49495 16038 49571
rect 16410 49495 16518 49571
rect 17178 49495 17286 49571
rect 17658 49495 17766 49571
rect 18426 49495 18534 49571
rect 18906 49495 19014 49571
rect 19674 49495 19782 49571
rect 20154 49495 20262 49571
rect 20922 49495 21030 49571
rect 21402 49495 21510 49571
rect 22170 49495 22278 49571
rect 22650 49495 22758 49571
rect 23418 49495 23526 49571
rect 23898 49495 24006 49571
rect 24666 49495 24774 49571
rect 25146 49495 25254 49571
rect 25914 49495 26022 49571
rect 26394 49495 26502 49571
rect 27162 49495 27270 49571
rect 27642 49495 27750 49571
rect 28410 49495 28518 49571
rect 28890 49495 28998 49571
rect 29658 49495 29766 49571
rect 30138 49495 30246 49571
rect 30906 49495 31014 49571
rect 31386 49495 31494 49571
rect 32154 49495 32262 49571
rect 32634 49495 32742 49571
rect 33402 49495 33510 49571
rect 33882 49495 33990 49571
rect 34650 49495 34758 49571
rect 35130 49495 35238 49571
rect 35898 49495 36006 49571
rect 36378 49495 36486 49571
rect 37146 49495 37254 49571
rect 37626 49495 37734 49571
rect 38394 49495 38502 49571
rect 38874 49495 38982 49571
rect 39642 49495 39750 49571
rect 0 49399 39936 49447
rect 0 49303 39936 49351
rect 186 49179 294 49255
rect 954 49179 1062 49255
rect 1434 49179 1542 49255
rect 2202 49179 2310 49255
rect 2682 49179 2790 49255
rect 3450 49179 3558 49255
rect 3930 49179 4038 49255
rect 4698 49179 4806 49255
rect 5178 49179 5286 49255
rect 5946 49179 6054 49255
rect 6426 49179 6534 49255
rect 7194 49179 7302 49255
rect 7674 49179 7782 49255
rect 8442 49179 8550 49255
rect 8922 49179 9030 49255
rect 9690 49179 9798 49255
rect 10170 49179 10278 49255
rect 10938 49179 11046 49255
rect 11418 49179 11526 49255
rect 12186 49179 12294 49255
rect 12666 49179 12774 49255
rect 13434 49179 13542 49255
rect 13914 49179 14022 49255
rect 14682 49179 14790 49255
rect 15162 49179 15270 49255
rect 15930 49179 16038 49255
rect 16410 49179 16518 49255
rect 17178 49179 17286 49255
rect 17658 49179 17766 49255
rect 18426 49179 18534 49255
rect 18906 49179 19014 49255
rect 19674 49179 19782 49255
rect 20154 49179 20262 49255
rect 20922 49179 21030 49255
rect 21402 49179 21510 49255
rect 22170 49179 22278 49255
rect 22650 49179 22758 49255
rect 23418 49179 23526 49255
rect 23898 49179 24006 49255
rect 24666 49179 24774 49255
rect 25146 49179 25254 49255
rect 25914 49179 26022 49255
rect 26394 49179 26502 49255
rect 27162 49179 27270 49255
rect 27642 49179 27750 49255
rect 28410 49179 28518 49255
rect 28890 49179 28998 49255
rect 29658 49179 29766 49255
rect 30138 49179 30246 49255
rect 30906 49179 31014 49255
rect 31386 49179 31494 49255
rect 32154 49179 32262 49255
rect 32634 49179 32742 49255
rect 33402 49179 33510 49255
rect 33882 49179 33990 49255
rect 34650 49179 34758 49255
rect 35130 49179 35238 49255
rect 35898 49179 36006 49255
rect 36378 49179 36486 49255
rect 37146 49179 37254 49255
rect 37626 49179 37734 49255
rect 38394 49179 38502 49255
rect 38874 49179 38982 49255
rect 39642 49179 39750 49255
rect 0 49083 39936 49131
rect 186 48925 294 49035
rect 954 48925 1062 49035
rect 1434 48925 1542 49035
rect 2202 48925 2310 49035
rect 2682 48925 2790 49035
rect 3450 48925 3558 49035
rect 3930 48925 4038 49035
rect 4698 48925 4806 49035
rect 5178 48925 5286 49035
rect 5946 48925 6054 49035
rect 6426 48925 6534 49035
rect 7194 48925 7302 49035
rect 7674 48925 7782 49035
rect 8442 48925 8550 49035
rect 8922 48925 9030 49035
rect 9690 48925 9798 49035
rect 10170 48925 10278 49035
rect 10938 48925 11046 49035
rect 11418 48925 11526 49035
rect 12186 48925 12294 49035
rect 12666 48925 12774 49035
rect 13434 48925 13542 49035
rect 13914 48925 14022 49035
rect 14682 48925 14790 49035
rect 15162 48925 15270 49035
rect 15930 48925 16038 49035
rect 16410 48925 16518 49035
rect 17178 48925 17286 49035
rect 17658 48925 17766 49035
rect 18426 48925 18534 49035
rect 18906 48925 19014 49035
rect 19674 48925 19782 49035
rect 20154 48925 20262 49035
rect 20922 48925 21030 49035
rect 21402 48925 21510 49035
rect 22170 48925 22278 49035
rect 22650 48925 22758 49035
rect 23418 48925 23526 49035
rect 23898 48925 24006 49035
rect 24666 48925 24774 49035
rect 25146 48925 25254 49035
rect 25914 48925 26022 49035
rect 26394 48925 26502 49035
rect 27162 48925 27270 49035
rect 27642 48925 27750 49035
rect 28410 48925 28518 49035
rect 28890 48925 28998 49035
rect 29658 48925 29766 49035
rect 30138 48925 30246 49035
rect 30906 48925 31014 49035
rect 31386 48925 31494 49035
rect 32154 48925 32262 49035
rect 32634 48925 32742 49035
rect 33402 48925 33510 49035
rect 33882 48925 33990 49035
rect 34650 48925 34758 49035
rect 35130 48925 35238 49035
rect 35898 48925 36006 49035
rect 36378 48925 36486 49035
rect 37146 48925 37254 49035
rect 37626 48925 37734 49035
rect 38394 48925 38502 49035
rect 38874 48925 38982 49035
rect 39642 48925 39750 49035
rect 0 48829 39936 48877
rect 186 48705 294 48781
rect 954 48705 1062 48781
rect 1434 48705 1542 48781
rect 2202 48705 2310 48781
rect 2682 48705 2790 48781
rect 3450 48705 3558 48781
rect 3930 48705 4038 48781
rect 4698 48705 4806 48781
rect 5178 48705 5286 48781
rect 5946 48705 6054 48781
rect 6426 48705 6534 48781
rect 7194 48705 7302 48781
rect 7674 48705 7782 48781
rect 8442 48705 8550 48781
rect 8922 48705 9030 48781
rect 9690 48705 9798 48781
rect 10170 48705 10278 48781
rect 10938 48705 11046 48781
rect 11418 48705 11526 48781
rect 12186 48705 12294 48781
rect 12666 48705 12774 48781
rect 13434 48705 13542 48781
rect 13914 48705 14022 48781
rect 14682 48705 14790 48781
rect 15162 48705 15270 48781
rect 15930 48705 16038 48781
rect 16410 48705 16518 48781
rect 17178 48705 17286 48781
rect 17658 48705 17766 48781
rect 18426 48705 18534 48781
rect 18906 48705 19014 48781
rect 19674 48705 19782 48781
rect 20154 48705 20262 48781
rect 20922 48705 21030 48781
rect 21402 48705 21510 48781
rect 22170 48705 22278 48781
rect 22650 48705 22758 48781
rect 23418 48705 23526 48781
rect 23898 48705 24006 48781
rect 24666 48705 24774 48781
rect 25146 48705 25254 48781
rect 25914 48705 26022 48781
rect 26394 48705 26502 48781
rect 27162 48705 27270 48781
rect 27642 48705 27750 48781
rect 28410 48705 28518 48781
rect 28890 48705 28998 48781
rect 29658 48705 29766 48781
rect 30138 48705 30246 48781
rect 30906 48705 31014 48781
rect 31386 48705 31494 48781
rect 32154 48705 32262 48781
rect 32634 48705 32742 48781
rect 33402 48705 33510 48781
rect 33882 48705 33990 48781
rect 34650 48705 34758 48781
rect 35130 48705 35238 48781
rect 35898 48705 36006 48781
rect 36378 48705 36486 48781
rect 37146 48705 37254 48781
rect 37626 48705 37734 48781
rect 38394 48705 38502 48781
rect 38874 48705 38982 48781
rect 39642 48705 39750 48781
rect 0 48609 39936 48657
rect 0 48513 39936 48561
rect 186 48389 294 48465
rect 954 48389 1062 48465
rect 1434 48389 1542 48465
rect 2202 48389 2310 48465
rect 2682 48389 2790 48465
rect 3450 48389 3558 48465
rect 3930 48389 4038 48465
rect 4698 48389 4806 48465
rect 5178 48389 5286 48465
rect 5946 48389 6054 48465
rect 6426 48389 6534 48465
rect 7194 48389 7302 48465
rect 7674 48389 7782 48465
rect 8442 48389 8550 48465
rect 8922 48389 9030 48465
rect 9690 48389 9798 48465
rect 10170 48389 10278 48465
rect 10938 48389 11046 48465
rect 11418 48389 11526 48465
rect 12186 48389 12294 48465
rect 12666 48389 12774 48465
rect 13434 48389 13542 48465
rect 13914 48389 14022 48465
rect 14682 48389 14790 48465
rect 15162 48389 15270 48465
rect 15930 48389 16038 48465
rect 16410 48389 16518 48465
rect 17178 48389 17286 48465
rect 17658 48389 17766 48465
rect 18426 48389 18534 48465
rect 18906 48389 19014 48465
rect 19674 48389 19782 48465
rect 20154 48389 20262 48465
rect 20922 48389 21030 48465
rect 21402 48389 21510 48465
rect 22170 48389 22278 48465
rect 22650 48389 22758 48465
rect 23418 48389 23526 48465
rect 23898 48389 24006 48465
rect 24666 48389 24774 48465
rect 25146 48389 25254 48465
rect 25914 48389 26022 48465
rect 26394 48389 26502 48465
rect 27162 48389 27270 48465
rect 27642 48389 27750 48465
rect 28410 48389 28518 48465
rect 28890 48389 28998 48465
rect 29658 48389 29766 48465
rect 30138 48389 30246 48465
rect 30906 48389 31014 48465
rect 31386 48389 31494 48465
rect 32154 48389 32262 48465
rect 32634 48389 32742 48465
rect 33402 48389 33510 48465
rect 33882 48389 33990 48465
rect 34650 48389 34758 48465
rect 35130 48389 35238 48465
rect 35898 48389 36006 48465
rect 36378 48389 36486 48465
rect 37146 48389 37254 48465
rect 37626 48389 37734 48465
rect 38394 48389 38502 48465
rect 38874 48389 38982 48465
rect 39642 48389 39750 48465
rect 0 48293 39936 48341
rect 186 48135 294 48245
rect 954 48135 1062 48245
rect 1434 48135 1542 48245
rect 2202 48135 2310 48245
rect 2682 48135 2790 48245
rect 3450 48135 3558 48245
rect 3930 48135 4038 48245
rect 4698 48135 4806 48245
rect 5178 48135 5286 48245
rect 5946 48135 6054 48245
rect 6426 48135 6534 48245
rect 7194 48135 7302 48245
rect 7674 48135 7782 48245
rect 8442 48135 8550 48245
rect 8922 48135 9030 48245
rect 9690 48135 9798 48245
rect 10170 48135 10278 48245
rect 10938 48135 11046 48245
rect 11418 48135 11526 48245
rect 12186 48135 12294 48245
rect 12666 48135 12774 48245
rect 13434 48135 13542 48245
rect 13914 48135 14022 48245
rect 14682 48135 14790 48245
rect 15162 48135 15270 48245
rect 15930 48135 16038 48245
rect 16410 48135 16518 48245
rect 17178 48135 17286 48245
rect 17658 48135 17766 48245
rect 18426 48135 18534 48245
rect 18906 48135 19014 48245
rect 19674 48135 19782 48245
rect 20154 48135 20262 48245
rect 20922 48135 21030 48245
rect 21402 48135 21510 48245
rect 22170 48135 22278 48245
rect 22650 48135 22758 48245
rect 23418 48135 23526 48245
rect 23898 48135 24006 48245
rect 24666 48135 24774 48245
rect 25146 48135 25254 48245
rect 25914 48135 26022 48245
rect 26394 48135 26502 48245
rect 27162 48135 27270 48245
rect 27642 48135 27750 48245
rect 28410 48135 28518 48245
rect 28890 48135 28998 48245
rect 29658 48135 29766 48245
rect 30138 48135 30246 48245
rect 30906 48135 31014 48245
rect 31386 48135 31494 48245
rect 32154 48135 32262 48245
rect 32634 48135 32742 48245
rect 33402 48135 33510 48245
rect 33882 48135 33990 48245
rect 34650 48135 34758 48245
rect 35130 48135 35238 48245
rect 35898 48135 36006 48245
rect 36378 48135 36486 48245
rect 37146 48135 37254 48245
rect 37626 48135 37734 48245
rect 38394 48135 38502 48245
rect 38874 48135 38982 48245
rect 39642 48135 39750 48245
rect 0 48039 39936 48087
rect 186 47915 294 47991
rect 954 47915 1062 47991
rect 1434 47915 1542 47991
rect 2202 47915 2310 47991
rect 2682 47915 2790 47991
rect 3450 47915 3558 47991
rect 3930 47915 4038 47991
rect 4698 47915 4806 47991
rect 5178 47915 5286 47991
rect 5946 47915 6054 47991
rect 6426 47915 6534 47991
rect 7194 47915 7302 47991
rect 7674 47915 7782 47991
rect 8442 47915 8550 47991
rect 8922 47915 9030 47991
rect 9690 47915 9798 47991
rect 10170 47915 10278 47991
rect 10938 47915 11046 47991
rect 11418 47915 11526 47991
rect 12186 47915 12294 47991
rect 12666 47915 12774 47991
rect 13434 47915 13542 47991
rect 13914 47915 14022 47991
rect 14682 47915 14790 47991
rect 15162 47915 15270 47991
rect 15930 47915 16038 47991
rect 16410 47915 16518 47991
rect 17178 47915 17286 47991
rect 17658 47915 17766 47991
rect 18426 47915 18534 47991
rect 18906 47915 19014 47991
rect 19674 47915 19782 47991
rect 20154 47915 20262 47991
rect 20922 47915 21030 47991
rect 21402 47915 21510 47991
rect 22170 47915 22278 47991
rect 22650 47915 22758 47991
rect 23418 47915 23526 47991
rect 23898 47915 24006 47991
rect 24666 47915 24774 47991
rect 25146 47915 25254 47991
rect 25914 47915 26022 47991
rect 26394 47915 26502 47991
rect 27162 47915 27270 47991
rect 27642 47915 27750 47991
rect 28410 47915 28518 47991
rect 28890 47915 28998 47991
rect 29658 47915 29766 47991
rect 30138 47915 30246 47991
rect 30906 47915 31014 47991
rect 31386 47915 31494 47991
rect 32154 47915 32262 47991
rect 32634 47915 32742 47991
rect 33402 47915 33510 47991
rect 33882 47915 33990 47991
rect 34650 47915 34758 47991
rect 35130 47915 35238 47991
rect 35898 47915 36006 47991
rect 36378 47915 36486 47991
rect 37146 47915 37254 47991
rect 37626 47915 37734 47991
rect 38394 47915 38502 47991
rect 38874 47915 38982 47991
rect 39642 47915 39750 47991
rect 0 47819 39936 47867
rect 0 47723 39936 47771
rect 186 47599 294 47675
rect 954 47599 1062 47675
rect 1434 47599 1542 47675
rect 2202 47599 2310 47675
rect 2682 47599 2790 47675
rect 3450 47599 3558 47675
rect 3930 47599 4038 47675
rect 4698 47599 4806 47675
rect 5178 47599 5286 47675
rect 5946 47599 6054 47675
rect 6426 47599 6534 47675
rect 7194 47599 7302 47675
rect 7674 47599 7782 47675
rect 8442 47599 8550 47675
rect 8922 47599 9030 47675
rect 9690 47599 9798 47675
rect 10170 47599 10278 47675
rect 10938 47599 11046 47675
rect 11418 47599 11526 47675
rect 12186 47599 12294 47675
rect 12666 47599 12774 47675
rect 13434 47599 13542 47675
rect 13914 47599 14022 47675
rect 14682 47599 14790 47675
rect 15162 47599 15270 47675
rect 15930 47599 16038 47675
rect 16410 47599 16518 47675
rect 17178 47599 17286 47675
rect 17658 47599 17766 47675
rect 18426 47599 18534 47675
rect 18906 47599 19014 47675
rect 19674 47599 19782 47675
rect 20154 47599 20262 47675
rect 20922 47599 21030 47675
rect 21402 47599 21510 47675
rect 22170 47599 22278 47675
rect 22650 47599 22758 47675
rect 23418 47599 23526 47675
rect 23898 47599 24006 47675
rect 24666 47599 24774 47675
rect 25146 47599 25254 47675
rect 25914 47599 26022 47675
rect 26394 47599 26502 47675
rect 27162 47599 27270 47675
rect 27642 47599 27750 47675
rect 28410 47599 28518 47675
rect 28890 47599 28998 47675
rect 29658 47599 29766 47675
rect 30138 47599 30246 47675
rect 30906 47599 31014 47675
rect 31386 47599 31494 47675
rect 32154 47599 32262 47675
rect 32634 47599 32742 47675
rect 33402 47599 33510 47675
rect 33882 47599 33990 47675
rect 34650 47599 34758 47675
rect 35130 47599 35238 47675
rect 35898 47599 36006 47675
rect 36378 47599 36486 47675
rect 37146 47599 37254 47675
rect 37626 47599 37734 47675
rect 38394 47599 38502 47675
rect 38874 47599 38982 47675
rect 39642 47599 39750 47675
rect 0 47503 39936 47551
rect 186 47345 294 47455
rect 954 47345 1062 47455
rect 1434 47345 1542 47455
rect 2202 47345 2310 47455
rect 2682 47345 2790 47455
rect 3450 47345 3558 47455
rect 3930 47345 4038 47455
rect 4698 47345 4806 47455
rect 5178 47345 5286 47455
rect 5946 47345 6054 47455
rect 6426 47345 6534 47455
rect 7194 47345 7302 47455
rect 7674 47345 7782 47455
rect 8442 47345 8550 47455
rect 8922 47345 9030 47455
rect 9690 47345 9798 47455
rect 10170 47345 10278 47455
rect 10938 47345 11046 47455
rect 11418 47345 11526 47455
rect 12186 47345 12294 47455
rect 12666 47345 12774 47455
rect 13434 47345 13542 47455
rect 13914 47345 14022 47455
rect 14682 47345 14790 47455
rect 15162 47345 15270 47455
rect 15930 47345 16038 47455
rect 16410 47345 16518 47455
rect 17178 47345 17286 47455
rect 17658 47345 17766 47455
rect 18426 47345 18534 47455
rect 18906 47345 19014 47455
rect 19674 47345 19782 47455
rect 20154 47345 20262 47455
rect 20922 47345 21030 47455
rect 21402 47345 21510 47455
rect 22170 47345 22278 47455
rect 22650 47345 22758 47455
rect 23418 47345 23526 47455
rect 23898 47345 24006 47455
rect 24666 47345 24774 47455
rect 25146 47345 25254 47455
rect 25914 47345 26022 47455
rect 26394 47345 26502 47455
rect 27162 47345 27270 47455
rect 27642 47345 27750 47455
rect 28410 47345 28518 47455
rect 28890 47345 28998 47455
rect 29658 47345 29766 47455
rect 30138 47345 30246 47455
rect 30906 47345 31014 47455
rect 31386 47345 31494 47455
rect 32154 47345 32262 47455
rect 32634 47345 32742 47455
rect 33402 47345 33510 47455
rect 33882 47345 33990 47455
rect 34650 47345 34758 47455
rect 35130 47345 35238 47455
rect 35898 47345 36006 47455
rect 36378 47345 36486 47455
rect 37146 47345 37254 47455
rect 37626 47345 37734 47455
rect 38394 47345 38502 47455
rect 38874 47345 38982 47455
rect 39642 47345 39750 47455
rect 0 47249 39936 47297
rect 186 47125 294 47201
rect 954 47125 1062 47201
rect 1434 47125 1542 47201
rect 2202 47125 2310 47201
rect 2682 47125 2790 47201
rect 3450 47125 3558 47201
rect 3930 47125 4038 47201
rect 4698 47125 4806 47201
rect 5178 47125 5286 47201
rect 5946 47125 6054 47201
rect 6426 47125 6534 47201
rect 7194 47125 7302 47201
rect 7674 47125 7782 47201
rect 8442 47125 8550 47201
rect 8922 47125 9030 47201
rect 9690 47125 9798 47201
rect 10170 47125 10278 47201
rect 10938 47125 11046 47201
rect 11418 47125 11526 47201
rect 12186 47125 12294 47201
rect 12666 47125 12774 47201
rect 13434 47125 13542 47201
rect 13914 47125 14022 47201
rect 14682 47125 14790 47201
rect 15162 47125 15270 47201
rect 15930 47125 16038 47201
rect 16410 47125 16518 47201
rect 17178 47125 17286 47201
rect 17658 47125 17766 47201
rect 18426 47125 18534 47201
rect 18906 47125 19014 47201
rect 19674 47125 19782 47201
rect 20154 47125 20262 47201
rect 20922 47125 21030 47201
rect 21402 47125 21510 47201
rect 22170 47125 22278 47201
rect 22650 47125 22758 47201
rect 23418 47125 23526 47201
rect 23898 47125 24006 47201
rect 24666 47125 24774 47201
rect 25146 47125 25254 47201
rect 25914 47125 26022 47201
rect 26394 47125 26502 47201
rect 27162 47125 27270 47201
rect 27642 47125 27750 47201
rect 28410 47125 28518 47201
rect 28890 47125 28998 47201
rect 29658 47125 29766 47201
rect 30138 47125 30246 47201
rect 30906 47125 31014 47201
rect 31386 47125 31494 47201
rect 32154 47125 32262 47201
rect 32634 47125 32742 47201
rect 33402 47125 33510 47201
rect 33882 47125 33990 47201
rect 34650 47125 34758 47201
rect 35130 47125 35238 47201
rect 35898 47125 36006 47201
rect 36378 47125 36486 47201
rect 37146 47125 37254 47201
rect 37626 47125 37734 47201
rect 38394 47125 38502 47201
rect 38874 47125 38982 47201
rect 39642 47125 39750 47201
rect 0 47029 39936 47077
rect 0 46933 39936 46981
rect 186 46809 294 46885
rect 954 46809 1062 46885
rect 1434 46809 1542 46885
rect 2202 46809 2310 46885
rect 2682 46809 2790 46885
rect 3450 46809 3558 46885
rect 3930 46809 4038 46885
rect 4698 46809 4806 46885
rect 5178 46809 5286 46885
rect 5946 46809 6054 46885
rect 6426 46809 6534 46885
rect 7194 46809 7302 46885
rect 7674 46809 7782 46885
rect 8442 46809 8550 46885
rect 8922 46809 9030 46885
rect 9690 46809 9798 46885
rect 10170 46809 10278 46885
rect 10938 46809 11046 46885
rect 11418 46809 11526 46885
rect 12186 46809 12294 46885
rect 12666 46809 12774 46885
rect 13434 46809 13542 46885
rect 13914 46809 14022 46885
rect 14682 46809 14790 46885
rect 15162 46809 15270 46885
rect 15930 46809 16038 46885
rect 16410 46809 16518 46885
rect 17178 46809 17286 46885
rect 17658 46809 17766 46885
rect 18426 46809 18534 46885
rect 18906 46809 19014 46885
rect 19674 46809 19782 46885
rect 20154 46809 20262 46885
rect 20922 46809 21030 46885
rect 21402 46809 21510 46885
rect 22170 46809 22278 46885
rect 22650 46809 22758 46885
rect 23418 46809 23526 46885
rect 23898 46809 24006 46885
rect 24666 46809 24774 46885
rect 25146 46809 25254 46885
rect 25914 46809 26022 46885
rect 26394 46809 26502 46885
rect 27162 46809 27270 46885
rect 27642 46809 27750 46885
rect 28410 46809 28518 46885
rect 28890 46809 28998 46885
rect 29658 46809 29766 46885
rect 30138 46809 30246 46885
rect 30906 46809 31014 46885
rect 31386 46809 31494 46885
rect 32154 46809 32262 46885
rect 32634 46809 32742 46885
rect 33402 46809 33510 46885
rect 33882 46809 33990 46885
rect 34650 46809 34758 46885
rect 35130 46809 35238 46885
rect 35898 46809 36006 46885
rect 36378 46809 36486 46885
rect 37146 46809 37254 46885
rect 37626 46809 37734 46885
rect 38394 46809 38502 46885
rect 38874 46809 38982 46885
rect 39642 46809 39750 46885
rect 0 46713 39936 46761
rect 186 46555 294 46665
rect 954 46555 1062 46665
rect 1434 46555 1542 46665
rect 2202 46555 2310 46665
rect 2682 46555 2790 46665
rect 3450 46555 3558 46665
rect 3930 46555 4038 46665
rect 4698 46555 4806 46665
rect 5178 46555 5286 46665
rect 5946 46555 6054 46665
rect 6426 46555 6534 46665
rect 7194 46555 7302 46665
rect 7674 46555 7782 46665
rect 8442 46555 8550 46665
rect 8922 46555 9030 46665
rect 9690 46555 9798 46665
rect 10170 46555 10278 46665
rect 10938 46555 11046 46665
rect 11418 46555 11526 46665
rect 12186 46555 12294 46665
rect 12666 46555 12774 46665
rect 13434 46555 13542 46665
rect 13914 46555 14022 46665
rect 14682 46555 14790 46665
rect 15162 46555 15270 46665
rect 15930 46555 16038 46665
rect 16410 46555 16518 46665
rect 17178 46555 17286 46665
rect 17658 46555 17766 46665
rect 18426 46555 18534 46665
rect 18906 46555 19014 46665
rect 19674 46555 19782 46665
rect 20154 46555 20262 46665
rect 20922 46555 21030 46665
rect 21402 46555 21510 46665
rect 22170 46555 22278 46665
rect 22650 46555 22758 46665
rect 23418 46555 23526 46665
rect 23898 46555 24006 46665
rect 24666 46555 24774 46665
rect 25146 46555 25254 46665
rect 25914 46555 26022 46665
rect 26394 46555 26502 46665
rect 27162 46555 27270 46665
rect 27642 46555 27750 46665
rect 28410 46555 28518 46665
rect 28890 46555 28998 46665
rect 29658 46555 29766 46665
rect 30138 46555 30246 46665
rect 30906 46555 31014 46665
rect 31386 46555 31494 46665
rect 32154 46555 32262 46665
rect 32634 46555 32742 46665
rect 33402 46555 33510 46665
rect 33882 46555 33990 46665
rect 34650 46555 34758 46665
rect 35130 46555 35238 46665
rect 35898 46555 36006 46665
rect 36378 46555 36486 46665
rect 37146 46555 37254 46665
rect 37626 46555 37734 46665
rect 38394 46555 38502 46665
rect 38874 46555 38982 46665
rect 39642 46555 39750 46665
rect 0 46459 39936 46507
rect 186 46335 294 46411
rect 954 46335 1062 46411
rect 1434 46335 1542 46411
rect 2202 46335 2310 46411
rect 2682 46335 2790 46411
rect 3450 46335 3558 46411
rect 3930 46335 4038 46411
rect 4698 46335 4806 46411
rect 5178 46335 5286 46411
rect 5946 46335 6054 46411
rect 6426 46335 6534 46411
rect 7194 46335 7302 46411
rect 7674 46335 7782 46411
rect 8442 46335 8550 46411
rect 8922 46335 9030 46411
rect 9690 46335 9798 46411
rect 10170 46335 10278 46411
rect 10938 46335 11046 46411
rect 11418 46335 11526 46411
rect 12186 46335 12294 46411
rect 12666 46335 12774 46411
rect 13434 46335 13542 46411
rect 13914 46335 14022 46411
rect 14682 46335 14790 46411
rect 15162 46335 15270 46411
rect 15930 46335 16038 46411
rect 16410 46335 16518 46411
rect 17178 46335 17286 46411
rect 17658 46335 17766 46411
rect 18426 46335 18534 46411
rect 18906 46335 19014 46411
rect 19674 46335 19782 46411
rect 20154 46335 20262 46411
rect 20922 46335 21030 46411
rect 21402 46335 21510 46411
rect 22170 46335 22278 46411
rect 22650 46335 22758 46411
rect 23418 46335 23526 46411
rect 23898 46335 24006 46411
rect 24666 46335 24774 46411
rect 25146 46335 25254 46411
rect 25914 46335 26022 46411
rect 26394 46335 26502 46411
rect 27162 46335 27270 46411
rect 27642 46335 27750 46411
rect 28410 46335 28518 46411
rect 28890 46335 28998 46411
rect 29658 46335 29766 46411
rect 30138 46335 30246 46411
rect 30906 46335 31014 46411
rect 31386 46335 31494 46411
rect 32154 46335 32262 46411
rect 32634 46335 32742 46411
rect 33402 46335 33510 46411
rect 33882 46335 33990 46411
rect 34650 46335 34758 46411
rect 35130 46335 35238 46411
rect 35898 46335 36006 46411
rect 36378 46335 36486 46411
rect 37146 46335 37254 46411
rect 37626 46335 37734 46411
rect 38394 46335 38502 46411
rect 38874 46335 38982 46411
rect 39642 46335 39750 46411
rect 0 46239 39936 46287
rect 0 46143 39936 46191
rect 186 46019 294 46095
rect 954 46019 1062 46095
rect 1434 46019 1542 46095
rect 2202 46019 2310 46095
rect 2682 46019 2790 46095
rect 3450 46019 3558 46095
rect 3930 46019 4038 46095
rect 4698 46019 4806 46095
rect 5178 46019 5286 46095
rect 5946 46019 6054 46095
rect 6426 46019 6534 46095
rect 7194 46019 7302 46095
rect 7674 46019 7782 46095
rect 8442 46019 8550 46095
rect 8922 46019 9030 46095
rect 9690 46019 9798 46095
rect 10170 46019 10278 46095
rect 10938 46019 11046 46095
rect 11418 46019 11526 46095
rect 12186 46019 12294 46095
rect 12666 46019 12774 46095
rect 13434 46019 13542 46095
rect 13914 46019 14022 46095
rect 14682 46019 14790 46095
rect 15162 46019 15270 46095
rect 15930 46019 16038 46095
rect 16410 46019 16518 46095
rect 17178 46019 17286 46095
rect 17658 46019 17766 46095
rect 18426 46019 18534 46095
rect 18906 46019 19014 46095
rect 19674 46019 19782 46095
rect 20154 46019 20262 46095
rect 20922 46019 21030 46095
rect 21402 46019 21510 46095
rect 22170 46019 22278 46095
rect 22650 46019 22758 46095
rect 23418 46019 23526 46095
rect 23898 46019 24006 46095
rect 24666 46019 24774 46095
rect 25146 46019 25254 46095
rect 25914 46019 26022 46095
rect 26394 46019 26502 46095
rect 27162 46019 27270 46095
rect 27642 46019 27750 46095
rect 28410 46019 28518 46095
rect 28890 46019 28998 46095
rect 29658 46019 29766 46095
rect 30138 46019 30246 46095
rect 30906 46019 31014 46095
rect 31386 46019 31494 46095
rect 32154 46019 32262 46095
rect 32634 46019 32742 46095
rect 33402 46019 33510 46095
rect 33882 46019 33990 46095
rect 34650 46019 34758 46095
rect 35130 46019 35238 46095
rect 35898 46019 36006 46095
rect 36378 46019 36486 46095
rect 37146 46019 37254 46095
rect 37626 46019 37734 46095
rect 38394 46019 38502 46095
rect 38874 46019 38982 46095
rect 39642 46019 39750 46095
rect 0 45923 39936 45971
rect 186 45765 294 45875
rect 954 45765 1062 45875
rect 1434 45765 1542 45875
rect 2202 45765 2310 45875
rect 2682 45765 2790 45875
rect 3450 45765 3558 45875
rect 3930 45765 4038 45875
rect 4698 45765 4806 45875
rect 5178 45765 5286 45875
rect 5946 45765 6054 45875
rect 6426 45765 6534 45875
rect 7194 45765 7302 45875
rect 7674 45765 7782 45875
rect 8442 45765 8550 45875
rect 8922 45765 9030 45875
rect 9690 45765 9798 45875
rect 10170 45765 10278 45875
rect 10938 45765 11046 45875
rect 11418 45765 11526 45875
rect 12186 45765 12294 45875
rect 12666 45765 12774 45875
rect 13434 45765 13542 45875
rect 13914 45765 14022 45875
rect 14682 45765 14790 45875
rect 15162 45765 15270 45875
rect 15930 45765 16038 45875
rect 16410 45765 16518 45875
rect 17178 45765 17286 45875
rect 17658 45765 17766 45875
rect 18426 45765 18534 45875
rect 18906 45765 19014 45875
rect 19674 45765 19782 45875
rect 20154 45765 20262 45875
rect 20922 45765 21030 45875
rect 21402 45765 21510 45875
rect 22170 45765 22278 45875
rect 22650 45765 22758 45875
rect 23418 45765 23526 45875
rect 23898 45765 24006 45875
rect 24666 45765 24774 45875
rect 25146 45765 25254 45875
rect 25914 45765 26022 45875
rect 26394 45765 26502 45875
rect 27162 45765 27270 45875
rect 27642 45765 27750 45875
rect 28410 45765 28518 45875
rect 28890 45765 28998 45875
rect 29658 45765 29766 45875
rect 30138 45765 30246 45875
rect 30906 45765 31014 45875
rect 31386 45765 31494 45875
rect 32154 45765 32262 45875
rect 32634 45765 32742 45875
rect 33402 45765 33510 45875
rect 33882 45765 33990 45875
rect 34650 45765 34758 45875
rect 35130 45765 35238 45875
rect 35898 45765 36006 45875
rect 36378 45765 36486 45875
rect 37146 45765 37254 45875
rect 37626 45765 37734 45875
rect 38394 45765 38502 45875
rect 38874 45765 38982 45875
rect 39642 45765 39750 45875
rect 0 45669 39936 45717
rect 186 45545 294 45621
rect 954 45545 1062 45621
rect 1434 45545 1542 45621
rect 2202 45545 2310 45621
rect 2682 45545 2790 45621
rect 3450 45545 3558 45621
rect 3930 45545 4038 45621
rect 4698 45545 4806 45621
rect 5178 45545 5286 45621
rect 5946 45545 6054 45621
rect 6426 45545 6534 45621
rect 7194 45545 7302 45621
rect 7674 45545 7782 45621
rect 8442 45545 8550 45621
rect 8922 45545 9030 45621
rect 9690 45545 9798 45621
rect 10170 45545 10278 45621
rect 10938 45545 11046 45621
rect 11418 45545 11526 45621
rect 12186 45545 12294 45621
rect 12666 45545 12774 45621
rect 13434 45545 13542 45621
rect 13914 45545 14022 45621
rect 14682 45545 14790 45621
rect 15162 45545 15270 45621
rect 15930 45545 16038 45621
rect 16410 45545 16518 45621
rect 17178 45545 17286 45621
rect 17658 45545 17766 45621
rect 18426 45545 18534 45621
rect 18906 45545 19014 45621
rect 19674 45545 19782 45621
rect 20154 45545 20262 45621
rect 20922 45545 21030 45621
rect 21402 45545 21510 45621
rect 22170 45545 22278 45621
rect 22650 45545 22758 45621
rect 23418 45545 23526 45621
rect 23898 45545 24006 45621
rect 24666 45545 24774 45621
rect 25146 45545 25254 45621
rect 25914 45545 26022 45621
rect 26394 45545 26502 45621
rect 27162 45545 27270 45621
rect 27642 45545 27750 45621
rect 28410 45545 28518 45621
rect 28890 45545 28998 45621
rect 29658 45545 29766 45621
rect 30138 45545 30246 45621
rect 30906 45545 31014 45621
rect 31386 45545 31494 45621
rect 32154 45545 32262 45621
rect 32634 45545 32742 45621
rect 33402 45545 33510 45621
rect 33882 45545 33990 45621
rect 34650 45545 34758 45621
rect 35130 45545 35238 45621
rect 35898 45545 36006 45621
rect 36378 45545 36486 45621
rect 37146 45545 37254 45621
rect 37626 45545 37734 45621
rect 38394 45545 38502 45621
rect 38874 45545 38982 45621
rect 39642 45545 39750 45621
rect 0 45449 39936 45497
rect 0 45353 39936 45401
rect 186 45229 294 45305
rect 954 45229 1062 45305
rect 1434 45229 1542 45305
rect 2202 45229 2310 45305
rect 2682 45229 2790 45305
rect 3450 45229 3558 45305
rect 3930 45229 4038 45305
rect 4698 45229 4806 45305
rect 5178 45229 5286 45305
rect 5946 45229 6054 45305
rect 6426 45229 6534 45305
rect 7194 45229 7302 45305
rect 7674 45229 7782 45305
rect 8442 45229 8550 45305
rect 8922 45229 9030 45305
rect 9690 45229 9798 45305
rect 10170 45229 10278 45305
rect 10938 45229 11046 45305
rect 11418 45229 11526 45305
rect 12186 45229 12294 45305
rect 12666 45229 12774 45305
rect 13434 45229 13542 45305
rect 13914 45229 14022 45305
rect 14682 45229 14790 45305
rect 15162 45229 15270 45305
rect 15930 45229 16038 45305
rect 16410 45229 16518 45305
rect 17178 45229 17286 45305
rect 17658 45229 17766 45305
rect 18426 45229 18534 45305
rect 18906 45229 19014 45305
rect 19674 45229 19782 45305
rect 20154 45229 20262 45305
rect 20922 45229 21030 45305
rect 21402 45229 21510 45305
rect 22170 45229 22278 45305
rect 22650 45229 22758 45305
rect 23418 45229 23526 45305
rect 23898 45229 24006 45305
rect 24666 45229 24774 45305
rect 25146 45229 25254 45305
rect 25914 45229 26022 45305
rect 26394 45229 26502 45305
rect 27162 45229 27270 45305
rect 27642 45229 27750 45305
rect 28410 45229 28518 45305
rect 28890 45229 28998 45305
rect 29658 45229 29766 45305
rect 30138 45229 30246 45305
rect 30906 45229 31014 45305
rect 31386 45229 31494 45305
rect 32154 45229 32262 45305
rect 32634 45229 32742 45305
rect 33402 45229 33510 45305
rect 33882 45229 33990 45305
rect 34650 45229 34758 45305
rect 35130 45229 35238 45305
rect 35898 45229 36006 45305
rect 36378 45229 36486 45305
rect 37146 45229 37254 45305
rect 37626 45229 37734 45305
rect 38394 45229 38502 45305
rect 38874 45229 38982 45305
rect 39642 45229 39750 45305
rect 0 45133 39936 45181
rect 186 44975 294 45085
rect 954 44975 1062 45085
rect 1434 44975 1542 45085
rect 2202 44975 2310 45085
rect 2682 44975 2790 45085
rect 3450 44975 3558 45085
rect 3930 44975 4038 45085
rect 4698 44975 4806 45085
rect 5178 44975 5286 45085
rect 5946 44975 6054 45085
rect 6426 44975 6534 45085
rect 7194 44975 7302 45085
rect 7674 44975 7782 45085
rect 8442 44975 8550 45085
rect 8922 44975 9030 45085
rect 9690 44975 9798 45085
rect 10170 44975 10278 45085
rect 10938 44975 11046 45085
rect 11418 44975 11526 45085
rect 12186 44975 12294 45085
rect 12666 44975 12774 45085
rect 13434 44975 13542 45085
rect 13914 44975 14022 45085
rect 14682 44975 14790 45085
rect 15162 44975 15270 45085
rect 15930 44975 16038 45085
rect 16410 44975 16518 45085
rect 17178 44975 17286 45085
rect 17658 44975 17766 45085
rect 18426 44975 18534 45085
rect 18906 44975 19014 45085
rect 19674 44975 19782 45085
rect 20154 44975 20262 45085
rect 20922 44975 21030 45085
rect 21402 44975 21510 45085
rect 22170 44975 22278 45085
rect 22650 44975 22758 45085
rect 23418 44975 23526 45085
rect 23898 44975 24006 45085
rect 24666 44975 24774 45085
rect 25146 44975 25254 45085
rect 25914 44975 26022 45085
rect 26394 44975 26502 45085
rect 27162 44975 27270 45085
rect 27642 44975 27750 45085
rect 28410 44975 28518 45085
rect 28890 44975 28998 45085
rect 29658 44975 29766 45085
rect 30138 44975 30246 45085
rect 30906 44975 31014 45085
rect 31386 44975 31494 45085
rect 32154 44975 32262 45085
rect 32634 44975 32742 45085
rect 33402 44975 33510 45085
rect 33882 44975 33990 45085
rect 34650 44975 34758 45085
rect 35130 44975 35238 45085
rect 35898 44975 36006 45085
rect 36378 44975 36486 45085
rect 37146 44975 37254 45085
rect 37626 44975 37734 45085
rect 38394 44975 38502 45085
rect 38874 44975 38982 45085
rect 39642 44975 39750 45085
rect 0 44879 39936 44927
rect 186 44755 294 44831
rect 954 44755 1062 44831
rect 1434 44755 1542 44831
rect 2202 44755 2310 44831
rect 2682 44755 2790 44831
rect 3450 44755 3558 44831
rect 3930 44755 4038 44831
rect 4698 44755 4806 44831
rect 5178 44755 5286 44831
rect 5946 44755 6054 44831
rect 6426 44755 6534 44831
rect 7194 44755 7302 44831
rect 7674 44755 7782 44831
rect 8442 44755 8550 44831
rect 8922 44755 9030 44831
rect 9690 44755 9798 44831
rect 10170 44755 10278 44831
rect 10938 44755 11046 44831
rect 11418 44755 11526 44831
rect 12186 44755 12294 44831
rect 12666 44755 12774 44831
rect 13434 44755 13542 44831
rect 13914 44755 14022 44831
rect 14682 44755 14790 44831
rect 15162 44755 15270 44831
rect 15930 44755 16038 44831
rect 16410 44755 16518 44831
rect 17178 44755 17286 44831
rect 17658 44755 17766 44831
rect 18426 44755 18534 44831
rect 18906 44755 19014 44831
rect 19674 44755 19782 44831
rect 20154 44755 20262 44831
rect 20922 44755 21030 44831
rect 21402 44755 21510 44831
rect 22170 44755 22278 44831
rect 22650 44755 22758 44831
rect 23418 44755 23526 44831
rect 23898 44755 24006 44831
rect 24666 44755 24774 44831
rect 25146 44755 25254 44831
rect 25914 44755 26022 44831
rect 26394 44755 26502 44831
rect 27162 44755 27270 44831
rect 27642 44755 27750 44831
rect 28410 44755 28518 44831
rect 28890 44755 28998 44831
rect 29658 44755 29766 44831
rect 30138 44755 30246 44831
rect 30906 44755 31014 44831
rect 31386 44755 31494 44831
rect 32154 44755 32262 44831
rect 32634 44755 32742 44831
rect 33402 44755 33510 44831
rect 33882 44755 33990 44831
rect 34650 44755 34758 44831
rect 35130 44755 35238 44831
rect 35898 44755 36006 44831
rect 36378 44755 36486 44831
rect 37146 44755 37254 44831
rect 37626 44755 37734 44831
rect 38394 44755 38502 44831
rect 38874 44755 38982 44831
rect 39642 44755 39750 44831
rect 0 44659 39936 44707
rect 0 44563 39936 44611
rect 186 44439 294 44515
rect 954 44439 1062 44515
rect 1434 44439 1542 44515
rect 2202 44439 2310 44515
rect 2682 44439 2790 44515
rect 3450 44439 3558 44515
rect 3930 44439 4038 44515
rect 4698 44439 4806 44515
rect 5178 44439 5286 44515
rect 5946 44439 6054 44515
rect 6426 44439 6534 44515
rect 7194 44439 7302 44515
rect 7674 44439 7782 44515
rect 8442 44439 8550 44515
rect 8922 44439 9030 44515
rect 9690 44439 9798 44515
rect 10170 44439 10278 44515
rect 10938 44439 11046 44515
rect 11418 44439 11526 44515
rect 12186 44439 12294 44515
rect 12666 44439 12774 44515
rect 13434 44439 13542 44515
rect 13914 44439 14022 44515
rect 14682 44439 14790 44515
rect 15162 44439 15270 44515
rect 15930 44439 16038 44515
rect 16410 44439 16518 44515
rect 17178 44439 17286 44515
rect 17658 44439 17766 44515
rect 18426 44439 18534 44515
rect 18906 44439 19014 44515
rect 19674 44439 19782 44515
rect 20154 44439 20262 44515
rect 20922 44439 21030 44515
rect 21402 44439 21510 44515
rect 22170 44439 22278 44515
rect 22650 44439 22758 44515
rect 23418 44439 23526 44515
rect 23898 44439 24006 44515
rect 24666 44439 24774 44515
rect 25146 44439 25254 44515
rect 25914 44439 26022 44515
rect 26394 44439 26502 44515
rect 27162 44439 27270 44515
rect 27642 44439 27750 44515
rect 28410 44439 28518 44515
rect 28890 44439 28998 44515
rect 29658 44439 29766 44515
rect 30138 44439 30246 44515
rect 30906 44439 31014 44515
rect 31386 44439 31494 44515
rect 32154 44439 32262 44515
rect 32634 44439 32742 44515
rect 33402 44439 33510 44515
rect 33882 44439 33990 44515
rect 34650 44439 34758 44515
rect 35130 44439 35238 44515
rect 35898 44439 36006 44515
rect 36378 44439 36486 44515
rect 37146 44439 37254 44515
rect 37626 44439 37734 44515
rect 38394 44439 38502 44515
rect 38874 44439 38982 44515
rect 39642 44439 39750 44515
rect 0 44343 39936 44391
rect 186 44185 294 44295
rect 954 44185 1062 44295
rect 1434 44185 1542 44295
rect 2202 44185 2310 44295
rect 2682 44185 2790 44295
rect 3450 44185 3558 44295
rect 3930 44185 4038 44295
rect 4698 44185 4806 44295
rect 5178 44185 5286 44295
rect 5946 44185 6054 44295
rect 6426 44185 6534 44295
rect 7194 44185 7302 44295
rect 7674 44185 7782 44295
rect 8442 44185 8550 44295
rect 8922 44185 9030 44295
rect 9690 44185 9798 44295
rect 10170 44185 10278 44295
rect 10938 44185 11046 44295
rect 11418 44185 11526 44295
rect 12186 44185 12294 44295
rect 12666 44185 12774 44295
rect 13434 44185 13542 44295
rect 13914 44185 14022 44295
rect 14682 44185 14790 44295
rect 15162 44185 15270 44295
rect 15930 44185 16038 44295
rect 16410 44185 16518 44295
rect 17178 44185 17286 44295
rect 17658 44185 17766 44295
rect 18426 44185 18534 44295
rect 18906 44185 19014 44295
rect 19674 44185 19782 44295
rect 20154 44185 20262 44295
rect 20922 44185 21030 44295
rect 21402 44185 21510 44295
rect 22170 44185 22278 44295
rect 22650 44185 22758 44295
rect 23418 44185 23526 44295
rect 23898 44185 24006 44295
rect 24666 44185 24774 44295
rect 25146 44185 25254 44295
rect 25914 44185 26022 44295
rect 26394 44185 26502 44295
rect 27162 44185 27270 44295
rect 27642 44185 27750 44295
rect 28410 44185 28518 44295
rect 28890 44185 28998 44295
rect 29658 44185 29766 44295
rect 30138 44185 30246 44295
rect 30906 44185 31014 44295
rect 31386 44185 31494 44295
rect 32154 44185 32262 44295
rect 32634 44185 32742 44295
rect 33402 44185 33510 44295
rect 33882 44185 33990 44295
rect 34650 44185 34758 44295
rect 35130 44185 35238 44295
rect 35898 44185 36006 44295
rect 36378 44185 36486 44295
rect 37146 44185 37254 44295
rect 37626 44185 37734 44295
rect 38394 44185 38502 44295
rect 38874 44185 38982 44295
rect 39642 44185 39750 44295
rect 0 44089 39936 44137
rect 186 43965 294 44041
rect 954 43965 1062 44041
rect 1434 43965 1542 44041
rect 2202 43965 2310 44041
rect 2682 43965 2790 44041
rect 3450 43965 3558 44041
rect 3930 43965 4038 44041
rect 4698 43965 4806 44041
rect 5178 43965 5286 44041
rect 5946 43965 6054 44041
rect 6426 43965 6534 44041
rect 7194 43965 7302 44041
rect 7674 43965 7782 44041
rect 8442 43965 8550 44041
rect 8922 43965 9030 44041
rect 9690 43965 9798 44041
rect 10170 43965 10278 44041
rect 10938 43965 11046 44041
rect 11418 43965 11526 44041
rect 12186 43965 12294 44041
rect 12666 43965 12774 44041
rect 13434 43965 13542 44041
rect 13914 43965 14022 44041
rect 14682 43965 14790 44041
rect 15162 43965 15270 44041
rect 15930 43965 16038 44041
rect 16410 43965 16518 44041
rect 17178 43965 17286 44041
rect 17658 43965 17766 44041
rect 18426 43965 18534 44041
rect 18906 43965 19014 44041
rect 19674 43965 19782 44041
rect 20154 43965 20262 44041
rect 20922 43965 21030 44041
rect 21402 43965 21510 44041
rect 22170 43965 22278 44041
rect 22650 43965 22758 44041
rect 23418 43965 23526 44041
rect 23898 43965 24006 44041
rect 24666 43965 24774 44041
rect 25146 43965 25254 44041
rect 25914 43965 26022 44041
rect 26394 43965 26502 44041
rect 27162 43965 27270 44041
rect 27642 43965 27750 44041
rect 28410 43965 28518 44041
rect 28890 43965 28998 44041
rect 29658 43965 29766 44041
rect 30138 43965 30246 44041
rect 30906 43965 31014 44041
rect 31386 43965 31494 44041
rect 32154 43965 32262 44041
rect 32634 43965 32742 44041
rect 33402 43965 33510 44041
rect 33882 43965 33990 44041
rect 34650 43965 34758 44041
rect 35130 43965 35238 44041
rect 35898 43965 36006 44041
rect 36378 43965 36486 44041
rect 37146 43965 37254 44041
rect 37626 43965 37734 44041
rect 38394 43965 38502 44041
rect 38874 43965 38982 44041
rect 39642 43965 39750 44041
rect 0 43869 39936 43917
rect 0 43773 39936 43821
rect 186 43649 294 43725
rect 954 43649 1062 43725
rect 1434 43649 1542 43725
rect 2202 43649 2310 43725
rect 2682 43649 2790 43725
rect 3450 43649 3558 43725
rect 3930 43649 4038 43725
rect 4698 43649 4806 43725
rect 5178 43649 5286 43725
rect 5946 43649 6054 43725
rect 6426 43649 6534 43725
rect 7194 43649 7302 43725
rect 7674 43649 7782 43725
rect 8442 43649 8550 43725
rect 8922 43649 9030 43725
rect 9690 43649 9798 43725
rect 10170 43649 10278 43725
rect 10938 43649 11046 43725
rect 11418 43649 11526 43725
rect 12186 43649 12294 43725
rect 12666 43649 12774 43725
rect 13434 43649 13542 43725
rect 13914 43649 14022 43725
rect 14682 43649 14790 43725
rect 15162 43649 15270 43725
rect 15930 43649 16038 43725
rect 16410 43649 16518 43725
rect 17178 43649 17286 43725
rect 17658 43649 17766 43725
rect 18426 43649 18534 43725
rect 18906 43649 19014 43725
rect 19674 43649 19782 43725
rect 20154 43649 20262 43725
rect 20922 43649 21030 43725
rect 21402 43649 21510 43725
rect 22170 43649 22278 43725
rect 22650 43649 22758 43725
rect 23418 43649 23526 43725
rect 23898 43649 24006 43725
rect 24666 43649 24774 43725
rect 25146 43649 25254 43725
rect 25914 43649 26022 43725
rect 26394 43649 26502 43725
rect 27162 43649 27270 43725
rect 27642 43649 27750 43725
rect 28410 43649 28518 43725
rect 28890 43649 28998 43725
rect 29658 43649 29766 43725
rect 30138 43649 30246 43725
rect 30906 43649 31014 43725
rect 31386 43649 31494 43725
rect 32154 43649 32262 43725
rect 32634 43649 32742 43725
rect 33402 43649 33510 43725
rect 33882 43649 33990 43725
rect 34650 43649 34758 43725
rect 35130 43649 35238 43725
rect 35898 43649 36006 43725
rect 36378 43649 36486 43725
rect 37146 43649 37254 43725
rect 37626 43649 37734 43725
rect 38394 43649 38502 43725
rect 38874 43649 38982 43725
rect 39642 43649 39750 43725
rect 0 43553 39936 43601
rect 186 43395 294 43505
rect 954 43395 1062 43505
rect 1434 43395 1542 43505
rect 2202 43395 2310 43505
rect 2682 43395 2790 43505
rect 3450 43395 3558 43505
rect 3930 43395 4038 43505
rect 4698 43395 4806 43505
rect 5178 43395 5286 43505
rect 5946 43395 6054 43505
rect 6426 43395 6534 43505
rect 7194 43395 7302 43505
rect 7674 43395 7782 43505
rect 8442 43395 8550 43505
rect 8922 43395 9030 43505
rect 9690 43395 9798 43505
rect 10170 43395 10278 43505
rect 10938 43395 11046 43505
rect 11418 43395 11526 43505
rect 12186 43395 12294 43505
rect 12666 43395 12774 43505
rect 13434 43395 13542 43505
rect 13914 43395 14022 43505
rect 14682 43395 14790 43505
rect 15162 43395 15270 43505
rect 15930 43395 16038 43505
rect 16410 43395 16518 43505
rect 17178 43395 17286 43505
rect 17658 43395 17766 43505
rect 18426 43395 18534 43505
rect 18906 43395 19014 43505
rect 19674 43395 19782 43505
rect 20154 43395 20262 43505
rect 20922 43395 21030 43505
rect 21402 43395 21510 43505
rect 22170 43395 22278 43505
rect 22650 43395 22758 43505
rect 23418 43395 23526 43505
rect 23898 43395 24006 43505
rect 24666 43395 24774 43505
rect 25146 43395 25254 43505
rect 25914 43395 26022 43505
rect 26394 43395 26502 43505
rect 27162 43395 27270 43505
rect 27642 43395 27750 43505
rect 28410 43395 28518 43505
rect 28890 43395 28998 43505
rect 29658 43395 29766 43505
rect 30138 43395 30246 43505
rect 30906 43395 31014 43505
rect 31386 43395 31494 43505
rect 32154 43395 32262 43505
rect 32634 43395 32742 43505
rect 33402 43395 33510 43505
rect 33882 43395 33990 43505
rect 34650 43395 34758 43505
rect 35130 43395 35238 43505
rect 35898 43395 36006 43505
rect 36378 43395 36486 43505
rect 37146 43395 37254 43505
rect 37626 43395 37734 43505
rect 38394 43395 38502 43505
rect 38874 43395 38982 43505
rect 39642 43395 39750 43505
rect 0 43299 39936 43347
rect 186 43175 294 43251
rect 954 43175 1062 43251
rect 1434 43175 1542 43251
rect 2202 43175 2310 43251
rect 2682 43175 2790 43251
rect 3450 43175 3558 43251
rect 3930 43175 4038 43251
rect 4698 43175 4806 43251
rect 5178 43175 5286 43251
rect 5946 43175 6054 43251
rect 6426 43175 6534 43251
rect 7194 43175 7302 43251
rect 7674 43175 7782 43251
rect 8442 43175 8550 43251
rect 8922 43175 9030 43251
rect 9690 43175 9798 43251
rect 10170 43175 10278 43251
rect 10938 43175 11046 43251
rect 11418 43175 11526 43251
rect 12186 43175 12294 43251
rect 12666 43175 12774 43251
rect 13434 43175 13542 43251
rect 13914 43175 14022 43251
rect 14682 43175 14790 43251
rect 15162 43175 15270 43251
rect 15930 43175 16038 43251
rect 16410 43175 16518 43251
rect 17178 43175 17286 43251
rect 17658 43175 17766 43251
rect 18426 43175 18534 43251
rect 18906 43175 19014 43251
rect 19674 43175 19782 43251
rect 20154 43175 20262 43251
rect 20922 43175 21030 43251
rect 21402 43175 21510 43251
rect 22170 43175 22278 43251
rect 22650 43175 22758 43251
rect 23418 43175 23526 43251
rect 23898 43175 24006 43251
rect 24666 43175 24774 43251
rect 25146 43175 25254 43251
rect 25914 43175 26022 43251
rect 26394 43175 26502 43251
rect 27162 43175 27270 43251
rect 27642 43175 27750 43251
rect 28410 43175 28518 43251
rect 28890 43175 28998 43251
rect 29658 43175 29766 43251
rect 30138 43175 30246 43251
rect 30906 43175 31014 43251
rect 31386 43175 31494 43251
rect 32154 43175 32262 43251
rect 32634 43175 32742 43251
rect 33402 43175 33510 43251
rect 33882 43175 33990 43251
rect 34650 43175 34758 43251
rect 35130 43175 35238 43251
rect 35898 43175 36006 43251
rect 36378 43175 36486 43251
rect 37146 43175 37254 43251
rect 37626 43175 37734 43251
rect 38394 43175 38502 43251
rect 38874 43175 38982 43251
rect 39642 43175 39750 43251
rect 0 43079 39936 43127
rect 0 42983 39936 43031
rect 186 42859 294 42935
rect 954 42859 1062 42935
rect 1434 42859 1542 42935
rect 2202 42859 2310 42935
rect 2682 42859 2790 42935
rect 3450 42859 3558 42935
rect 3930 42859 4038 42935
rect 4698 42859 4806 42935
rect 5178 42859 5286 42935
rect 5946 42859 6054 42935
rect 6426 42859 6534 42935
rect 7194 42859 7302 42935
rect 7674 42859 7782 42935
rect 8442 42859 8550 42935
rect 8922 42859 9030 42935
rect 9690 42859 9798 42935
rect 10170 42859 10278 42935
rect 10938 42859 11046 42935
rect 11418 42859 11526 42935
rect 12186 42859 12294 42935
rect 12666 42859 12774 42935
rect 13434 42859 13542 42935
rect 13914 42859 14022 42935
rect 14682 42859 14790 42935
rect 15162 42859 15270 42935
rect 15930 42859 16038 42935
rect 16410 42859 16518 42935
rect 17178 42859 17286 42935
rect 17658 42859 17766 42935
rect 18426 42859 18534 42935
rect 18906 42859 19014 42935
rect 19674 42859 19782 42935
rect 20154 42859 20262 42935
rect 20922 42859 21030 42935
rect 21402 42859 21510 42935
rect 22170 42859 22278 42935
rect 22650 42859 22758 42935
rect 23418 42859 23526 42935
rect 23898 42859 24006 42935
rect 24666 42859 24774 42935
rect 25146 42859 25254 42935
rect 25914 42859 26022 42935
rect 26394 42859 26502 42935
rect 27162 42859 27270 42935
rect 27642 42859 27750 42935
rect 28410 42859 28518 42935
rect 28890 42859 28998 42935
rect 29658 42859 29766 42935
rect 30138 42859 30246 42935
rect 30906 42859 31014 42935
rect 31386 42859 31494 42935
rect 32154 42859 32262 42935
rect 32634 42859 32742 42935
rect 33402 42859 33510 42935
rect 33882 42859 33990 42935
rect 34650 42859 34758 42935
rect 35130 42859 35238 42935
rect 35898 42859 36006 42935
rect 36378 42859 36486 42935
rect 37146 42859 37254 42935
rect 37626 42859 37734 42935
rect 38394 42859 38502 42935
rect 38874 42859 38982 42935
rect 39642 42859 39750 42935
rect 0 42763 39936 42811
rect 186 42605 294 42715
rect 954 42605 1062 42715
rect 1434 42605 1542 42715
rect 2202 42605 2310 42715
rect 2682 42605 2790 42715
rect 3450 42605 3558 42715
rect 3930 42605 4038 42715
rect 4698 42605 4806 42715
rect 5178 42605 5286 42715
rect 5946 42605 6054 42715
rect 6426 42605 6534 42715
rect 7194 42605 7302 42715
rect 7674 42605 7782 42715
rect 8442 42605 8550 42715
rect 8922 42605 9030 42715
rect 9690 42605 9798 42715
rect 10170 42605 10278 42715
rect 10938 42605 11046 42715
rect 11418 42605 11526 42715
rect 12186 42605 12294 42715
rect 12666 42605 12774 42715
rect 13434 42605 13542 42715
rect 13914 42605 14022 42715
rect 14682 42605 14790 42715
rect 15162 42605 15270 42715
rect 15930 42605 16038 42715
rect 16410 42605 16518 42715
rect 17178 42605 17286 42715
rect 17658 42605 17766 42715
rect 18426 42605 18534 42715
rect 18906 42605 19014 42715
rect 19674 42605 19782 42715
rect 20154 42605 20262 42715
rect 20922 42605 21030 42715
rect 21402 42605 21510 42715
rect 22170 42605 22278 42715
rect 22650 42605 22758 42715
rect 23418 42605 23526 42715
rect 23898 42605 24006 42715
rect 24666 42605 24774 42715
rect 25146 42605 25254 42715
rect 25914 42605 26022 42715
rect 26394 42605 26502 42715
rect 27162 42605 27270 42715
rect 27642 42605 27750 42715
rect 28410 42605 28518 42715
rect 28890 42605 28998 42715
rect 29658 42605 29766 42715
rect 30138 42605 30246 42715
rect 30906 42605 31014 42715
rect 31386 42605 31494 42715
rect 32154 42605 32262 42715
rect 32634 42605 32742 42715
rect 33402 42605 33510 42715
rect 33882 42605 33990 42715
rect 34650 42605 34758 42715
rect 35130 42605 35238 42715
rect 35898 42605 36006 42715
rect 36378 42605 36486 42715
rect 37146 42605 37254 42715
rect 37626 42605 37734 42715
rect 38394 42605 38502 42715
rect 38874 42605 38982 42715
rect 39642 42605 39750 42715
rect 0 42509 39936 42557
rect 186 42385 294 42461
rect 954 42385 1062 42461
rect 1434 42385 1542 42461
rect 2202 42385 2310 42461
rect 2682 42385 2790 42461
rect 3450 42385 3558 42461
rect 3930 42385 4038 42461
rect 4698 42385 4806 42461
rect 5178 42385 5286 42461
rect 5946 42385 6054 42461
rect 6426 42385 6534 42461
rect 7194 42385 7302 42461
rect 7674 42385 7782 42461
rect 8442 42385 8550 42461
rect 8922 42385 9030 42461
rect 9690 42385 9798 42461
rect 10170 42385 10278 42461
rect 10938 42385 11046 42461
rect 11418 42385 11526 42461
rect 12186 42385 12294 42461
rect 12666 42385 12774 42461
rect 13434 42385 13542 42461
rect 13914 42385 14022 42461
rect 14682 42385 14790 42461
rect 15162 42385 15270 42461
rect 15930 42385 16038 42461
rect 16410 42385 16518 42461
rect 17178 42385 17286 42461
rect 17658 42385 17766 42461
rect 18426 42385 18534 42461
rect 18906 42385 19014 42461
rect 19674 42385 19782 42461
rect 20154 42385 20262 42461
rect 20922 42385 21030 42461
rect 21402 42385 21510 42461
rect 22170 42385 22278 42461
rect 22650 42385 22758 42461
rect 23418 42385 23526 42461
rect 23898 42385 24006 42461
rect 24666 42385 24774 42461
rect 25146 42385 25254 42461
rect 25914 42385 26022 42461
rect 26394 42385 26502 42461
rect 27162 42385 27270 42461
rect 27642 42385 27750 42461
rect 28410 42385 28518 42461
rect 28890 42385 28998 42461
rect 29658 42385 29766 42461
rect 30138 42385 30246 42461
rect 30906 42385 31014 42461
rect 31386 42385 31494 42461
rect 32154 42385 32262 42461
rect 32634 42385 32742 42461
rect 33402 42385 33510 42461
rect 33882 42385 33990 42461
rect 34650 42385 34758 42461
rect 35130 42385 35238 42461
rect 35898 42385 36006 42461
rect 36378 42385 36486 42461
rect 37146 42385 37254 42461
rect 37626 42385 37734 42461
rect 38394 42385 38502 42461
rect 38874 42385 38982 42461
rect 39642 42385 39750 42461
rect 0 42289 39936 42337
rect 0 42193 39936 42241
rect 186 42069 294 42145
rect 954 42069 1062 42145
rect 1434 42069 1542 42145
rect 2202 42069 2310 42145
rect 2682 42069 2790 42145
rect 3450 42069 3558 42145
rect 3930 42069 4038 42145
rect 4698 42069 4806 42145
rect 5178 42069 5286 42145
rect 5946 42069 6054 42145
rect 6426 42069 6534 42145
rect 7194 42069 7302 42145
rect 7674 42069 7782 42145
rect 8442 42069 8550 42145
rect 8922 42069 9030 42145
rect 9690 42069 9798 42145
rect 10170 42069 10278 42145
rect 10938 42069 11046 42145
rect 11418 42069 11526 42145
rect 12186 42069 12294 42145
rect 12666 42069 12774 42145
rect 13434 42069 13542 42145
rect 13914 42069 14022 42145
rect 14682 42069 14790 42145
rect 15162 42069 15270 42145
rect 15930 42069 16038 42145
rect 16410 42069 16518 42145
rect 17178 42069 17286 42145
rect 17658 42069 17766 42145
rect 18426 42069 18534 42145
rect 18906 42069 19014 42145
rect 19674 42069 19782 42145
rect 20154 42069 20262 42145
rect 20922 42069 21030 42145
rect 21402 42069 21510 42145
rect 22170 42069 22278 42145
rect 22650 42069 22758 42145
rect 23418 42069 23526 42145
rect 23898 42069 24006 42145
rect 24666 42069 24774 42145
rect 25146 42069 25254 42145
rect 25914 42069 26022 42145
rect 26394 42069 26502 42145
rect 27162 42069 27270 42145
rect 27642 42069 27750 42145
rect 28410 42069 28518 42145
rect 28890 42069 28998 42145
rect 29658 42069 29766 42145
rect 30138 42069 30246 42145
rect 30906 42069 31014 42145
rect 31386 42069 31494 42145
rect 32154 42069 32262 42145
rect 32634 42069 32742 42145
rect 33402 42069 33510 42145
rect 33882 42069 33990 42145
rect 34650 42069 34758 42145
rect 35130 42069 35238 42145
rect 35898 42069 36006 42145
rect 36378 42069 36486 42145
rect 37146 42069 37254 42145
rect 37626 42069 37734 42145
rect 38394 42069 38502 42145
rect 38874 42069 38982 42145
rect 39642 42069 39750 42145
rect 0 41973 39936 42021
rect 186 41815 294 41925
rect 954 41815 1062 41925
rect 1434 41815 1542 41925
rect 2202 41815 2310 41925
rect 2682 41815 2790 41925
rect 3450 41815 3558 41925
rect 3930 41815 4038 41925
rect 4698 41815 4806 41925
rect 5178 41815 5286 41925
rect 5946 41815 6054 41925
rect 6426 41815 6534 41925
rect 7194 41815 7302 41925
rect 7674 41815 7782 41925
rect 8442 41815 8550 41925
rect 8922 41815 9030 41925
rect 9690 41815 9798 41925
rect 10170 41815 10278 41925
rect 10938 41815 11046 41925
rect 11418 41815 11526 41925
rect 12186 41815 12294 41925
rect 12666 41815 12774 41925
rect 13434 41815 13542 41925
rect 13914 41815 14022 41925
rect 14682 41815 14790 41925
rect 15162 41815 15270 41925
rect 15930 41815 16038 41925
rect 16410 41815 16518 41925
rect 17178 41815 17286 41925
rect 17658 41815 17766 41925
rect 18426 41815 18534 41925
rect 18906 41815 19014 41925
rect 19674 41815 19782 41925
rect 20154 41815 20262 41925
rect 20922 41815 21030 41925
rect 21402 41815 21510 41925
rect 22170 41815 22278 41925
rect 22650 41815 22758 41925
rect 23418 41815 23526 41925
rect 23898 41815 24006 41925
rect 24666 41815 24774 41925
rect 25146 41815 25254 41925
rect 25914 41815 26022 41925
rect 26394 41815 26502 41925
rect 27162 41815 27270 41925
rect 27642 41815 27750 41925
rect 28410 41815 28518 41925
rect 28890 41815 28998 41925
rect 29658 41815 29766 41925
rect 30138 41815 30246 41925
rect 30906 41815 31014 41925
rect 31386 41815 31494 41925
rect 32154 41815 32262 41925
rect 32634 41815 32742 41925
rect 33402 41815 33510 41925
rect 33882 41815 33990 41925
rect 34650 41815 34758 41925
rect 35130 41815 35238 41925
rect 35898 41815 36006 41925
rect 36378 41815 36486 41925
rect 37146 41815 37254 41925
rect 37626 41815 37734 41925
rect 38394 41815 38502 41925
rect 38874 41815 38982 41925
rect 39642 41815 39750 41925
rect 0 41719 39936 41767
rect 186 41595 294 41671
rect 954 41595 1062 41671
rect 1434 41595 1542 41671
rect 2202 41595 2310 41671
rect 2682 41595 2790 41671
rect 3450 41595 3558 41671
rect 3930 41595 4038 41671
rect 4698 41595 4806 41671
rect 5178 41595 5286 41671
rect 5946 41595 6054 41671
rect 6426 41595 6534 41671
rect 7194 41595 7302 41671
rect 7674 41595 7782 41671
rect 8442 41595 8550 41671
rect 8922 41595 9030 41671
rect 9690 41595 9798 41671
rect 10170 41595 10278 41671
rect 10938 41595 11046 41671
rect 11418 41595 11526 41671
rect 12186 41595 12294 41671
rect 12666 41595 12774 41671
rect 13434 41595 13542 41671
rect 13914 41595 14022 41671
rect 14682 41595 14790 41671
rect 15162 41595 15270 41671
rect 15930 41595 16038 41671
rect 16410 41595 16518 41671
rect 17178 41595 17286 41671
rect 17658 41595 17766 41671
rect 18426 41595 18534 41671
rect 18906 41595 19014 41671
rect 19674 41595 19782 41671
rect 20154 41595 20262 41671
rect 20922 41595 21030 41671
rect 21402 41595 21510 41671
rect 22170 41595 22278 41671
rect 22650 41595 22758 41671
rect 23418 41595 23526 41671
rect 23898 41595 24006 41671
rect 24666 41595 24774 41671
rect 25146 41595 25254 41671
rect 25914 41595 26022 41671
rect 26394 41595 26502 41671
rect 27162 41595 27270 41671
rect 27642 41595 27750 41671
rect 28410 41595 28518 41671
rect 28890 41595 28998 41671
rect 29658 41595 29766 41671
rect 30138 41595 30246 41671
rect 30906 41595 31014 41671
rect 31386 41595 31494 41671
rect 32154 41595 32262 41671
rect 32634 41595 32742 41671
rect 33402 41595 33510 41671
rect 33882 41595 33990 41671
rect 34650 41595 34758 41671
rect 35130 41595 35238 41671
rect 35898 41595 36006 41671
rect 36378 41595 36486 41671
rect 37146 41595 37254 41671
rect 37626 41595 37734 41671
rect 38394 41595 38502 41671
rect 38874 41595 38982 41671
rect 39642 41595 39750 41671
rect 0 41499 39936 41547
rect 0 41403 39936 41451
rect 186 41279 294 41355
rect 954 41279 1062 41355
rect 1434 41279 1542 41355
rect 2202 41279 2310 41355
rect 2682 41279 2790 41355
rect 3450 41279 3558 41355
rect 3930 41279 4038 41355
rect 4698 41279 4806 41355
rect 5178 41279 5286 41355
rect 5946 41279 6054 41355
rect 6426 41279 6534 41355
rect 7194 41279 7302 41355
rect 7674 41279 7782 41355
rect 8442 41279 8550 41355
rect 8922 41279 9030 41355
rect 9690 41279 9798 41355
rect 10170 41279 10278 41355
rect 10938 41279 11046 41355
rect 11418 41279 11526 41355
rect 12186 41279 12294 41355
rect 12666 41279 12774 41355
rect 13434 41279 13542 41355
rect 13914 41279 14022 41355
rect 14682 41279 14790 41355
rect 15162 41279 15270 41355
rect 15930 41279 16038 41355
rect 16410 41279 16518 41355
rect 17178 41279 17286 41355
rect 17658 41279 17766 41355
rect 18426 41279 18534 41355
rect 18906 41279 19014 41355
rect 19674 41279 19782 41355
rect 20154 41279 20262 41355
rect 20922 41279 21030 41355
rect 21402 41279 21510 41355
rect 22170 41279 22278 41355
rect 22650 41279 22758 41355
rect 23418 41279 23526 41355
rect 23898 41279 24006 41355
rect 24666 41279 24774 41355
rect 25146 41279 25254 41355
rect 25914 41279 26022 41355
rect 26394 41279 26502 41355
rect 27162 41279 27270 41355
rect 27642 41279 27750 41355
rect 28410 41279 28518 41355
rect 28890 41279 28998 41355
rect 29658 41279 29766 41355
rect 30138 41279 30246 41355
rect 30906 41279 31014 41355
rect 31386 41279 31494 41355
rect 32154 41279 32262 41355
rect 32634 41279 32742 41355
rect 33402 41279 33510 41355
rect 33882 41279 33990 41355
rect 34650 41279 34758 41355
rect 35130 41279 35238 41355
rect 35898 41279 36006 41355
rect 36378 41279 36486 41355
rect 37146 41279 37254 41355
rect 37626 41279 37734 41355
rect 38394 41279 38502 41355
rect 38874 41279 38982 41355
rect 39642 41279 39750 41355
rect 0 41183 39936 41231
rect 186 41025 294 41135
rect 954 41025 1062 41135
rect 1434 41025 1542 41135
rect 2202 41025 2310 41135
rect 2682 41025 2790 41135
rect 3450 41025 3558 41135
rect 3930 41025 4038 41135
rect 4698 41025 4806 41135
rect 5178 41025 5286 41135
rect 5946 41025 6054 41135
rect 6426 41025 6534 41135
rect 7194 41025 7302 41135
rect 7674 41025 7782 41135
rect 8442 41025 8550 41135
rect 8922 41025 9030 41135
rect 9690 41025 9798 41135
rect 10170 41025 10278 41135
rect 10938 41025 11046 41135
rect 11418 41025 11526 41135
rect 12186 41025 12294 41135
rect 12666 41025 12774 41135
rect 13434 41025 13542 41135
rect 13914 41025 14022 41135
rect 14682 41025 14790 41135
rect 15162 41025 15270 41135
rect 15930 41025 16038 41135
rect 16410 41025 16518 41135
rect 17178 41025 17286 41135
rect 17658 41025 17766 41135
rect 18426 41025 18534 41135
rect 18906 41025 19014 41135
rect 19674 41025 19782 41135
rect 20154 41025 20262 41135
rect 20922 41025 21030 41135
rect 21402 41025 21510 41135
rect 22170 41025 22278 41135
rect 22650 41025 22758 41135
rect 23418 41025 23526 41135
rect 23898 41025 24006 41135
rect 24666 41025 24774 41135
rect 25146 41025 25254 41135
rect 25914 41025 26022 41135
rect 26394 41025 26502 41135
rect 27162 41025 27270 41135
rect 27642 41025 27750 41135
rect 28410 41025 28518 41135
rect 28890 41025 28998 41135
rect 29658 41025 29766 41135
rect 30138 41025 30246 41135
rect 30906 41025 31014 41135
rect 31386 41025 31494 41135
rect 32154 41025 32262 41135
rect 32634 41025 32742 41135
rect 33402 41025 33510 41135
rect 33882 41025 33990 41135
rect 34650 41025 34758 41135
rect 35130 41025 35238 41135
rect 35898 41025 36006 41135
rect 36378 41025 36486 41135
rect 37146 41025 37254 41135
rect 37626 41025 37734 41135
rect 38394 41025 38502 41135
rect 38874 41025 38982 41135
rect 39642 41025 39750 41135
rect 0 40929 39936 40977
rect 186 40805 294 40881
rect 954 40805 1062 40881
rect 1434 40805 1542 40881
rect 2202 40805 2310 40881
rect 2682 40805 2790 40881
rect 3450 40805 3558 40881
rect 3930 40805 4038 40881
rect 4698 40805 4806 40881
rect 5178 40805 5286 40881
rect 5946 40805 6054 40881
rect 6426 40805 6534 40881
rect 7194 40805 7302 40881
rect 7674 40805 7782 40881
rect 8442 40805 8550 40881
rect 8922 40805 9030 40881
rect 9690 40805 9798 40881
rect 10170 40805 10278 40881
rect 10938 40805 11046 40881
rect 11418 40805 11526 40881
rect 12186 40805 12294 40881
rect 12666 40805 12774 40881
rect 13434 40805 13542 40881
rect 13914 40805 14022 40881
rect 14682 40805 14790 40881
rect 15162 40805 15270 40881
rect 15930 40805 16038 40881
rect 16410 40805 16518 40881
rect 17178 40805 17286 40881
rect 17658 40805 17766 40881
rect 18426 40805 18534 40881
rect 18906 40805 19014 40881
rect 19674 40805 19782 40881
rect 20154 40805 20262 40881
rect 20922 40805 21030 40881
rect 21402 40805 21510 40881
rect 22170 40805 22278 40881
rect 22650 40805 22758 40881
rect 23418 40805 23526 40881
rect 23898 40805 24006 40881
rect 24666 40805 24774 40881
rect 25146 40805 25254 40881
rect 25914 40805 26022 40881
rect 26394 40805 26502 40881
rect 27162 40805 27270 40881
rect 27642 40805 27750 40881
rect 28410 40805 28518 40881
rect 28890 40805 28998 40881
rect 29658 40805 29766 40881
rect 30138 40805 30246 40881
rect 30906 40805 31014 40881
rect 31386 40805 31494 40881
rect 32154 40805 32262 40881
rect 32634 40805 32742 40881
rect 33402 40805 33510 40881
rect 33882 40805 33990 40881
rect 34650 40805 34758 40881
rect 35130 40805 35238 40881
rect 35898 40805 36006 40881
rect 36378 40805 36486 40881
rect 37146 40805 37254 40881
rect 37626 40805 37734 40881
rect 38394 40805 38502 40881
rect 38874 40805 38982 40881
rect 39642 40805 39750 40881
rect 0 40709 39936 40757
rect 0 40613 39936 40661
rect 186 40489 294 40565
rect 954 40489 1062 40565
rect 1434 40489 1542 40565
rect 2202 40489 2310 40565
rect 2682 40489 2790 40565
rect 3450 40489 3558 40565
rect 3930 40489 4038 40565
rect 4698 40489 4806 40565
rect 5178 40489 5286 40565
rect 5946 40489 6054 40565
rect 6426 40489 6534 40565
rect 7194 40489 7302 40565
rect 7674 40489 7782 40565
rect 8442 40489 8550 40565
rect 8922 40489 9030 40565
rect 9690 40489 9798 40565
rect 10170 40489 10278 40565
rect 10938 40489 11046 40565
rect 11418 40489 11526 40565
rect 12186 40489 12294 40565
rect 12666 40489 12774 40565
rect 13434 40489 13542 40565
rect 13914 40489 14022 40565
rect 14682 40489 14790 40565
rect 15162 40489 15270 40565
rect 15930 40489 16038 40565
rect 16410 40489 16518 40565
rect 17178 40489 17286 40565
rect 17658 40489 17766 40565
rect 18426 40489 18534 40565
rect 18906 40489 19014 40565
rect 19674 40489 19782 40565
rect 20154 40489 20262 40565
rect 20922 40489 21030 40565
rect 21402 40489 21510 40565
rect 22170 40489 22278 40565
rect 22650 40489 22758 40565
rect 23418 40489 23526 40565
rect 23898 40489 24006 40565
rect 24666 40489 24774 40565
rect 25146 40489 25254 40565
rect 25914 40489 26022 40565
rect 26394 40489 26502 40565
rect 27162 40489 27270 40565
rect 27642 40489 27750 40565
rect 28410 40489 28518 40565
rect 28890 40489 28998 40565
rect 29658 40489 29766 40565
rect 30138 40489 30246 40565
rect 30906 40489 31014 40565
rect 31386 40489 31494 40565
rect 32154 40489 32262 40565
rect 32634 40489 32742 40565
rect 33402 40489 33510 40565
rect 33882 40489 33990 40565
rect 34650 40489 34758 40565
rect 35130 40489 35238 40565
rect 35898 40489 36006 40565
rect 36378 40489 36486 40565
rect 37146 40489 37254 40565
rect 37626 40489 37734 40565
rect 38394 40489 38502 40565
rect 38874 40489 38982 40565
rect 39642 40489 39750 40565
rect 0 40393 39936 40441
rect 186 40235 294 40345
rect 954 40235 1062 40345
rect 1434 40235 1542 40345
rect 2202 40235 2310 40345
rect 2682 40235 2790 40345
rect 3450 40235 3558 40345
rect 3930 40235 4038 40345
rect 4698 40235 4806 40345
rect 5178 40235 5286 40345
rect 5946 40235 6054 40345
rect 6426 40235 6534 40345
rect 7194 40235 7302 40345
rect 7674 40235 7782 40345
rect 8442 40235 8550 40345
rect 8922 40235 9030 40345
rect 9690 40235 9798 40345
rect 10170 40235 10278 40345
rect 10938 40235 11046 40345
rect 11418 40235 11526 40345
rect 12186 40235 12294 40345
rect 12666 40235 12774 40345
rect 13434 40235 13542 40345
rect 13914 40235 14022 40345
rect 14682 40235 14790 40345
rect 15162 40235 15270 40345
rect 15930 40235 16038 40345
rect 16410 40235 16518 40345
rect 17178 40235 17286 40345
rect 17658 40235 17766 40345
rect 18426 40235 18534 40345
rect 18906 40235 19014 40345
rect 19674 40235 19782 40345
rect 20154 40235 20262 40345
rect 20922 40235 21030 40345
rect 21402 40235 21510 40345
rect 22170 40235 22278 40345
rect 22650 40235 22758 40345
rect 23418 40235 23526 40345
rect 23898 40235 24006 40345
rect 24666 40235 24774 40345
rect 25146 40235 25254 40345
rect 25914 40235 26022 40345
rect 26394 40235 26502 40345
rect 27162 40235 27270 40345
rect 27642 40235 27750 40345
rect 28410 40235 28518 40345
rect 28890 40235 28998 40345
rect 29658 40235 29766 40345
rect 30138 40235 30246 40345
rect 30906 40235 31014 40345
rect 31386 40235 31494 40345
rect 32154 40235 32262 40345
rect 32634 40235 32742 40345
rect 33402 40235 33510 40345
rect 33882 40235 33990 40345
rect 34650 40235 34758 40345
rect 35130 40235 35238 40345
rect 35898 40235 36006 40345
rect 36378 40235 36486 40345
rect 37146 40235 37254 40345
rect 37626 40235 37734 40345
rect 38394 40235 38502 40345
rect 38874 40235 38982 40345
rect 39642 40235 39750 40345
rect 0 40139 39936 40187
rect 186 40015 294 40091
rect 954 40015 1062 40091
rect 1434 40015 1542 40091
rect 2202 40015 2310 40091
rect 2682 40015 2790 40091
rect 3450 40015 3558 40091
rect 3930 40015 4038 40091
rect 4698 40015 4806 40091
rect 5178 40015 5286 40091
rect 5946 40015 6054 40091
rect 6426 40015 6534 40091
rect 7194 40015 7302 40091
rect 7674 40015 7782 40091
rect 8442 40015 8550 40091
rect 8922 40015 9030 40091
rect 9690 40015 9798 40091
rect 10170 40015 10278 40091
rect 10938 40015 11046 40091
rect 11418 40015 11526 40091
rect 12186 40015 12294 40091
rect 12666 40015 12774 40091
rect 13434 40015 13542 40091
rect 13914 40015 14022 40091
rect 14682 40015 14790 40091
rect 15162 40015 15270 40091
rect 15930 40015 16038 40091
rect 16410 40015 16518 40091
rect 17178 40015 17286 40091
rect 17658 40015 17766 40091
rect 18426 40015 18534 40091
rect 18906 40015 19014 40091
rect 19674 40015 19782 40091
rect 20154 40015 20262 40091
rect 20922 40015 21030 40091
rect 21402 40015 21510 40091
rect 22170 40015 22278 40091
rect 22650 40015 22758 40091
rect 23418 40015 23526 40091
rect 23898 40015 24006 40091
rect 24666 40015 24774 40091
rect 25146 40015 25254 40091
rect 25914 40015 26022 40091
rect 26394 40015 26502 40091
rect 27162 40015 27270 40091
rect 27642 40015 27750 40091
rect 28410 40015 28518 40091
rect 28890 40015 28998 40091
rect 29658 40015 29766 40091
rect 30138 40015 30246 40091
rect 30906 40015 31014 40091
rect 31386 40015 31494 40091
rect 32154 40015 32262 40091
rect 32634 40015 32742 40091
rect 33402 40015 33510 40091
rect 33882 40015 33990 40091
rect 34650 40015 34758 40091
rect 35130 40015 35238 40091
rect 35898 40015 36006 40091
rect 36378 40015 36486 40091
rect 37146 40015 37254 40091
rect 37626 40015 37734 40091
rect 38394 40015 38502 40091
rect 38874 40015 38982 40091
rect 39642 40015 39750 40091
rect 0 39919 39936 39967
rect 0 39823 39936 39871
rect 186 39699 294 39775
rect 954 39699 1062 39775
rect 1434 39699 1542 39775
rect 2202 39699 2310 39775
rect 2682 39699 2790 39775
rect 3450 39699 3558 39775
rect 3930 39699 4038 39775
rect 4698 39699 4806 39775
rect 5178 39699 5286 39775
rect 5946 39699 6054 39775
rect 6426 39699 6534 39775
rect 7194 39699 7302 39775
rect 7674 39699 7782 39775
rect 8442 39699 8550 39775
rect 8922 39699 9030 39775
rect 9690 39699 9798 39775
rect 10170 39699 10278 39775
rect 10938 39699 11046 39775
rect 11418 39699 11526 39775
rect 12186 39699 12294 39775
rect 12666 39699 12774 39775
rect 13434 39699 13542 39775
rect 13914 39699 14022 39775
rect 14682 39699 14790 39775
rect 15162 39699 15270 39775
rect 15930 39699 16038 39775
rect 16410 39699 16518 39775
rect 17178 39699 17286 39775
rect 17658 39699 17766 39775
rect 18426 39699 18534 39775
rect 18906 39699 19014 39775
rect 19674 39699 19782 39775
rect 20154 39699 20262 39775
rect 20922 39699 21030 39775
rect 21402 39699 21510 39775
rect 22170 39699 22278 39775
rect 22650 39699 22758 39775
rect 23418 39699 23526 39775
rect 23898 39699 24006 39775
rect 24666 39699 24774 39775
rect 25146 39699 25254 39775
rect 25914 39699 26022 39775
rect 26394 39699 26502 39775
rect 27162 39699 27270 39775
rect 27642 39699 27750 39775
rect 28410 39699 28518 39775
rect 28890 39699 28998 39775
rect 29658 39699 29766 39775
rect 30138 39699 30246 39775
rect 30906 39699 31014 39775
rect 31386 39699 31494 39775
rect 32154 39699 32262 39775
rect 32634 39699 32742 39775
rect 33402 39699 33510 39775
rect 33882 39699 33990 39775
rect 34650 39699 34758 39775
rect 35130 39699 35238 39775
rect 35898 39699 36006 39775
rect 36378 39699 36486 39775
rect 37146 39699 37254 39775
rect 37626 39699 37734 39775
rect 38394 39699 38502 39775
rect 38874 39699 38982 39775
rect 39642 39699 39750 39775
rect 0 39603 39936 39651
rect 186 39445 294 39555
rect 954 39445 1062 39555
rect 1434 39445 1542 39555
rect 2202 39445 2310 39555
rect 2682 39445 2790 39555
rect 3450 39445 3558 39555
rect 3930 39445 4038 39555
rect 4698 39445 4806 39555
rect 5178 39445 5286 39555
rect 5946 39445 6054 39555
rect 6426 39445 6534 39555
rect 7194 39445 7302 39555
rect 7674 39445 7782 39555
rect 8442 39445 8550 39555
rect 8922 39445 9030 39555
rect 9690 39445 9798 39555
rect 10170 39445 10278 39555
rect 10938 39445 11046 39555
rect 11418 39445 11526 39555
rect 12186 39445 12294 39555
rect 12666 39445 12774 39555
rect 13434 39445 13542 39555
rect 13914 39445 14022 39555
rect 14682 39445 14790 39555
rect 15162 39445 15270 39555
rect 15930 39445 16038 39555
rect 16410 39445 16518 39555
rect 17178 39445 17286 39555
rect 17658 39445 17766 39555
rect 18426 39445 18534 39555
rect 18906 39445 19014 39555
rect 19674 39445 19782 39555
rect 20154 39445 20262 39555
rect 20922 39445 21030 39555
rect 21402 39445 21510 39555
rect 22170 39445 22278 39555
rect 22650 39445 22758 39555
rect 23418 39445 23526 39555
rect 23898 39445 24006 39555
rect 24666 39445 24774 39555
rect 25146 39445 25254 39555
rect 25914 39445 26022 39555
rect 26394 39445 26502 39555
rect 27162 39445 27270 39555
rect 27642 39445 27750 39555
rect 28410 39445 28518 39555
rect 28890 39445 28998 39555
rect 29658 39445 29766 39555
rect 30138 39445 30246 39555
rect 30906 39445 31014 39555
rect 31386 39445 31494 39555
rect 32154 39445 32262 39555
rect 32634 39445 32742 39555
rect 33402 39445 33510 39555
rect 33882 39445 33990 39555
rect 34650 39445 34758 39555
rect 35130 39445 35238 39555
rect 35898 39445 36006 39555
rect 36378 39445 36486 39555
rect 37146 39445 37254 39555
rect 37626 39445 37734 39555
rect 38394 39445 38502 39555
rect 38874 39445 38982 39555
rect 39642 39445 39750 39555
rect 0 39349 39936 39397
rect 186 39225 294 39301
rect 954 39225 1062 39301
rect 1434 39225 1542 39301
rect 2202 39225 2310 39301
rect 2682 39225 2790 39301
rect 3450 39225 3558 39301
rect 3930 39225 4038 39301
rect 4698 39225 4806 39301
rect 5178 39225 5286 39301
rect 5946 39225 6054 39301
rect 6426 39225 6534 39301
rect 7194 39225 7302 39301
rect 7674 39225 7782 39301
rect 8442 39225 8550 39301
rect 8922 39225 9030 39301
rect 9690 39225 9798 39301
rect 10170 39225 10278 39301
rect 10938 39225 11046 39301
rect 11418 39225 11526 39301
rect 12186 39225 12294 39301
rect 12666 39225 12774 39301
rect 13434 39225 13542 39301
rect 13914 39225 14022 39301
rect 14682 39225 14790 39301
rect 15162 39225 15270 39301
rect 15930 39225 16038 39301
rect 16410 39225 16518 39301
rect 17178 39225 17286 39301
rect 17658 39225 17766 39301
rect 18426 39225 18534 39301
rect 18906 39225 19014 39301
rect 19674 39225 19782 39301
rect 20154 39225 20262 39301
rect 20922 39225 21030 39301
rect 21402 39225 21510 39301
rect 22170 39225 22278 39301
rect 22650 39225 22758 39301
rect 23418 39225 23526 39301
rect 23898 39225 24006 39301
rect 24666 39225 24774 39301
rect 25146 39225 25254 39301
rect 25914 39225 26022 39301
rect 26394 39225 26502 39301
rect 27162 39225 27270 39301
rect 27642 39225 27750 39301
rect 28410 39225 28518 39301
rect 28890 39225 28998 39301
rect 29658 39225 29766 39301
rect 30138 39225 30246 39301
rect 30906 39225 31014 39301
rect 31386 39225 31494 39301
rect 32154 39225 32262 39301
rect 32634 39225 32742 39301
rect 33402 39225 33510 39301
rect 33882 39225 33990 39301
rect 34650 39225 34758 39301
rect 35130 39225 35238 39301
rect 35898 39225 36006 39301
rect 36378 39225 36486 39301
rect 37146 39225 37254 39301
rect 37626 39225 37734 39301
rect 38394 39225 38502 39301
rect 38874 39225 38982 39301
rect 39642 39225 39750 39301
rect 0 39129 39936 39177
rect 0 39033 39936 39081
rect 186 38909 294 38985
rect 954 38909 1062 38985
rect 1434 38909 1542 38985
rect 2202 38909 2310 38985
rect 2682 38909 2790 38985
rect 3450 38909 3558 38985
rect 3930 38909 4038 38985
rect 4698 38909 4806 38985
rect 5178 38909 5286 38985
rect 5946 38909 6054 38985
rect 6426 38909 6534 38985
rect 7194 38909 7302 38985
rect 7674 38909 7782 38985
rect 8442 38909 8550 38985
rect 8922 38909 9030 38985
rect 9690 38909 9798 38985
rect 10170 38909 10278 38985
rect 10938 38909 11046 38985
rect 11418 38909 11526 38985
rect 12186 38909 12294 38985
rect 12666 38909 12774 38985
rect 13434 38909 13542 38985
rect 13914 38909 14022 38985
rect 14682 38909 14790 38985
rect 15162 38909 15270 38985
rect 15930 38909 16038 38985
rect 16410 38909 16518 38985
rect 17178 38909 17286 38985
rect 17658 38909 17766 38985
rect 18426 38909 18534 38985
rect 18906 38909 19014 38985
rect 19674 38909 19782 38985
rect 20154 38909 20262 38985
rect 20922 38909 21030 38985
rect 21402 38909 21510 38985
rect 22170 38909 22278 38985
rect 22650 38909 22758 38985
rect 23418 38909 23526 38985
rect 23898 38909 24006 38985
rect 24666 38909 24774 38985
rect 25146 38909 25254 38985
rect 25914 38909 26022 38985
rect 26394 38909 26502 38985
rect 27162 38909 27270 38985
rect 27642 38909 27750 38985
rect 28410 38909 28518 38985
rect 28890 38909 28998 38985
rect 29658 38909 29766 38985
rect 30138 38909 30246 38985
rect 30906 38909 31014 38985
rect 31386 38909 31494 38985
rect 32154 38909 32262 38985
rect 32634 38909 32742 38985
rect 33402 38909 33510 38985
rect 33882 38909 33990 38985
rect 34650 38909 34758 38985
rect 35130 38909 35238 38985
rect 35898 38909 36006 38985
rect 36378 38909 36486 38985
rect 37146 38909 37254 38985
rect 37626 38909 37734 38985
rect 38394 38909 38502 38985
rect 38874 38909 38982 38985
rect 39642 38909 39750 38985
rect 0 38813 39936 38861
rect 186 38655 294 38765
rect 954 38655 1062 38765
rect 1434 38655 1542 38765
rect 2202 38655 2310 38765
rect 2682 38655 2790 38765
rect 3450 38655 3558 38765
rect 3930 38655 4038 38765
rect 4698 38655 4806 38765
rect 5178 38655 5286 38765
rect 5946 38655 6054 38765
rect 6426 38655 6534 38765
rect 7194 38655 7302 38765
rect 7674 38655 7782 38765
rect 8442 38655 8550 38765
rect 8922 38655 9030 38765
rect 9690 38655 9798 38765
rect 10170 38655 10278 38765
rect 10938 38655 11046 38765
rect 11418 38655 11526 38765
rect 12186 38655 12294 38765
rect 12666 38655 12774 38765
rect 13434 38655 13542 38765
rect 13914 38655 14022 38765
rect 14682 38655 14790 38765
rect 15162 38655 15270 38765
rect 15930 38655 16038 38765
rect 16410 38655 16518 38765
rect 17178 38655 17286 38765
rect 17658 38655 17766 38765
rect 18426 38655 18534 38765
rect 18906 38655 19014 38765
rect 19674 38655 19782 38765
rect 20154 38655 20262 38765
rect 20922 38655 21030 38765
rect 21402 38655 21510 38765
rect 22170 38655 22278 38765
rect 22650 38655 22758 38765
rect 23418 38655 23526 38765
rect 23898 38655 24006 38765
rect 24666 38655 24774 38765
rect 25146 38655 25254 38765
rect 25914 38655 26022 38765
rect 26394 38655 26502 38765
rect 27162 38655 27270 38765
rect 27642 38655 27750 38765
rect 28410 38655 28518 38765
rect 28890 38655 28998 38765
rect 29658 38655 29766 38765
rect 30138 38655 30246 38765
rect 30906 38655 31014 38765
rect 31386 38655 31494 38765
rect 32154 38655 32262 38765
rect 32634 38655 32742 38765
rect 33402 38655 33510 38765
rect 33882 38655 33990 38765
rect 34650 38655 34758 38765
rect 35130 38655 35238 38765
rect 35898 38655 36006 38765
rect 36378 38655 36486 38765
rect 37146 38655 37254 38765
rect 37626 38655 37734 38765
rect 38394 38655 38502 38765
rect 38874 38655 38982 38765
rect 39642 38655 39750 38765
rect 0 38559 39936 38607
rect 186 38435 294 38511
rect 954 38435 1062 38511
rect 1434 38435 1542 38511
rect 2202 38435 2310 38511
rect 2682 38435 2790 38511
rect 3450 38435 3558 38511
rect 3930 38435 4038 38511
rect 4698 38435 4806 38511
rect 5178 38435 5286 38511
rect 5946 38435 6054 38511
rect 6426 38435 6534 38511
rect 7194 38435 7302 38511
rect 7674 38435 7782 38511
rect 8442 38435 8550 38511
rect 8922 38435 9030 38511
rect 9690 38435 9798 38511
rect 10170 38435 10278 38511
rect 10938 38435 11046 38511
rect 11418 38435 11526 38511
rect 12186 38435 12294 38511
rect 12666 38435 12774 38511
rect 13434 38435 13542 38511
rect 13914 38435 14022 38511
rect 14682 38435 14790 38511
rect 15162 38435 15270 38511
rect 15930 38435 16038 38511
rect 16410 38435 16518 38511
rect 17178 38435 17286 38511
rect 17658 38435 17766 38511
rect 18426 38435 18534 38511
rect 18906 38435 19014 38511
rect 19674 38435 19782 38511
rect 20154 38435 20262 38511
rect 20922 38435 21030 38511
rect 21402 38435 21510 38511
rect 22170 38435 22278 38511
rect 22650 38435 22758 38511
rect 23418 38435 23526 38511
rect 23898 38435 24006 38511
rect 24666 38435 24774 38511
rect 25146 38435 25254 38511
rect 25914 38435 26022 38511
rect 26394 38435 26502 38511
rect 27162 38435 27270 38511
rect 27642 38435 27750 38511
rect 28410 38435 28518 38511
rect 28890 38435 28998 38511
rect 29658 38435 29766 38511
rect 30138 38435 30246 38511
rect 30906 38435 31014 38511
rect 31386 38435 31494 38511
rect 32154 38435 32262 38511
rect 32634 38435 32742 38511
rect 33402 38435 33510 38511
rect 33882 38435 33990 38511
rect 34650 38435 34758 38511
rect 35130 38435 35238 38511
rect 35898 38435 36006 38511
rect 36378 38435 36486 38511
rect 37146 38435 37254 38511
rect 37626 38435 37734 38511
rect 38394 38435 38502 38511
rect 38874 38435 38982 38511
rect 39642 38435 39750 38511
rect 0 38339 39936 38387
rect 0 38243 39936 38291
rect 186 38119 294 38195
rect 954 38119 1062 38195
rect 1434 38119 1542 38195
rect 2202 38119 2310 38195
rect 2682 38119 2790 38195
rect 3450 38119 3558 38195
rect 3930 38119 4038 38195
rect 4698 38119 4806 38195
rect 5178 38119 5286 38195
rect 5946 38119 6054 38195
rect 6426 38119 6534 38195
rect 7194 38119 7302 38195
rect 7674 38119 7782 38195
rect 8442 38119 8550 38195
rect 8922 38119 9030 38195
rect 9690 38119 9798 38195
rect 10170 38119 10278 38195
rect 10938 38119 11046 38195
rect 11418 38119 11526 38195
rect 12186 38119 12294 38195
rect 12666 38119 12774 38195
rect 13434 38119 13542 38195
rect 13914 38119 14022 38195
rect 14682 38119 14790 38195
rect 15162 38119 15270 38195
rect 15930 38119 16038 38195
rect 16410 38119 16518 38195
rect 17178 38119 17286 38195
rect 17658 38119 17766 38195
rect 18426 38119 18534 38195
rect 18906 38119 19014 38195
rect 19674 38119 19782 38195
rect 20154 38119 20262 38195
rect 20922 38119 21030 38195
rect 21402 38119 21510 38195
rect 22170 38119 22278 38195
rect 22650 38119 22758 38195
rect 23418 38119 23526 38195
rect 23898 38119 24006 38195
rect 24666 38119 24774 38195
rect 25146 38119 25254 38195
rect 25914 38119 26022 38195
rect 26394 38119 26502 38195
rect 27162 38119 27270 38195
rect 27642 38119 27750 38195
rect 28410 38119 28518 38195
rect 28890 38119 28998 38195
rect 29658 38119 29766 38195
rect 30138 38119 30246 38195
rect 30906 38119 31014 38195
rect 31386 38119 31494 38195
rect 32154 38119 32262 38195
rect 32634 38119 32742 38195
rect 33402 38119 33510 38195
rect 33882 38119 33990 38195
rect 34650 38119 34758 38195
rect 35130 38119 35238 38195
rect 35898 38119 36006 38195
rect 36378 38119 36486 38195
rect 37146 38119 37254 38195
rect 37626 38119 37734 38195
rect 38394 38119 38502 38195
rect 38874 38119 38982 38195
rect 39642 38119 39750 38195
rect 0 38023 39936 38071
rect 186 37865 294 37975
rect 954 37865 1062 37975
rect 1434 37865 1542 37975
rect 2202 37865 2310 37975
rect 2682 37865 2790 37975
rect 3450 37865 3558 37975
rect 3930 37865 4038 37975
rect 4698 37865 4806 37975
rect 5178 37865 5286 37975
rect 5946 37865 6054 37975
rect 6426 37865 6534 37975
rect 7194 37865 7302 37975
rect 7674 37865 7782 37975
rect 8442 37865 8550 37975
rect 8922 37865 9030 37975
rect 9690 37865 9798 37975
rect 10170 37865 10278 37975
rect 10938 37865 11046 37975
rect 11418 37865 11526 37975
rect 12186 37865 12294 37975
rect 12666 37865 12774 37975
rect 13434 37865 13542 37975
rect 13914 37865 14022 37975
rect 14682 37865 14790 37975
rect 15162 37865 15270 37975
rect 15930 37865 16038 37975
rect 16410 37865 16518 37975
rect 17178 37865 17286 37975
rect 17658 37865 17766 37975
rect 18426 37865 18534 37975
rect 18906 37865 19014 37975
rect 19674 37865 19782 37975
rect 20154 37865 20262 37975
rect 20922 37865 21030 37975
rect 21402 37865 21510 37975
rect 22170 37865 22278 37975
rect 22650 37865 22758 37975
rect 23418 37865 23526 37975
rect 23898 37865 24006 37975
rect 24666 37865 24774 37975
rect 25146 37865 25254 37975
rect 25914 37865 26022 37975
rect 26394 37865 26502 37975
rect 27162 37865 27270 37975
rect 27642 37865 27750 37975
rect 28410 37865 28518 37975
rect 28890 37865 28998 37975
rect 29658 37865 29766 37975
rect 30138 37865 30246 37975
rect 30906 37865 31014 37975
rect 31386 37865 31494 37975
rect 32154 37865 32262 37975
rect 32634 37865 32742 37975
rect 33402 37865 33510 37975
rect 33882 37865 33990 37975
rect 34650 37865 34758 37975
rect 35130 37865 35238 37975
rect 35898 37865 36006 37975
rect 36378 37865 36486 37975
rect 37146 37865 37254 37975
rect 37626 37865 37734 37975
rect 38394 37865 38502 37975
rect 38874 37865 38982 37975
rect 39642 37865 39750 37975
rect 0 37769 39936 37817
rect 186 37645 294 37721
rect 954 37645 1062 37721
rect 1434 37645 1542 37721
rect 2202 37645 2310 37721
rect 2682 37645 2790 37721
rect 3450 37645 3558 37721
rect 3930 37645 4038 37721
rect 4698 37645 4806 37721
rect 5178 37645 5286 37721
rect 5946 37645 6054 37721
rect 6426 37645 6534 37721
rect 7194 37645 7302 37721
rect 7674 37645 7782 37721
rect 8442 37645 8550 37721
rect 8922 37645 9030 37721
rect 9690 37645 9798 37721
rect 10170 37645 10278 37721
rect 10938 37645 11046 37721
rect 11418 37645 11526 37721
rect 12186 37645 12294 37721
rect 12666 37645 12774 37721
rect 13434 37645 13542 37721
rect 13914 37645 14022 37721
rect 14682 37645 14790 37721
rect 15162 37645 15270 37721
rect 15930 37645 16038 37721
rect 16410 37645 16518 37721
rect 17178 37645 17286 37721
rect 17658 37645 17766 37721
rect 18426 37645 18534 37721
rect 18906 37645 19014 37721
rect 19674 37645 19782 37721
rect 20154 37645 20262 37721
rect 20922 37645 21030 37721
rect 21402 37645 21510 37721
rect 22170 37645 22278 37721
rect 22650 37645 22758 37721
rect 23418 37645 23526 37721
rect 23898 37645 24006 37721
rect 24666 37645 24774 37721
rect 25146 37645 25254 37721
rect 25914 37645 26022 37721
rect 26394 37645 26502 37721
rect 27162 37645 27270 37721
rect 27642 37645 27750 37721
rect 28410 37645 28518 37721
rect 28890 37645 28998 37721
rect 29658 37645 29766 37721
rect 30138 37645 30246 37721
rect 30906 37645 31014 37721
rect 31386 37645 31494 37721
rect 32154 37645 32262 37721
rect 32634 37645 32742 37721
rect 33402 37645 33510 37721
rect 33882 37645 33990 37721
rect 34650 37645 34758 37721
rect 35130 37645 35238 37721
rect 35898 37645 36006 37721
rect 36378 37645 36486 37721
rect 37146 37645 37254 37721
rect 37626 37645 37734 37721
rect 38394 37645 38502 37721
rect 38874 37645 38982 37721
rect 39642 37645 39750 37721
rect 0 37549 39936 37597
rect 0 37453 39936 37501
rect 186 37329 294 37405
rect 954 37329 1062 37405
rect 1434 37329 1542 37405
rect 2202 37329 2310 37405
rect 2682 37329 2790 37405
rect 3450 37329 3558 37405
rect 3930 37329 4038 37405
rect 4698 37329 4806 37405
rect 5178 37329 5286 37405
rect 5946 37329 6054 37405
rect 6426 37329 6534 37405
rect 7194 37329 7302 37405
rect 7674 37329 7782 37405
rect 8442 37329 8550 37405
rect 8922 37329 9030 37405
rect 9690 37329 9798 37405
rect 10170 37329 10278 37405
rect 10938 37329 11046 37405
rect 11418 37329 11526 37405
rect 12186 37329 12294 37405
rect 12666 37329 12774 37405
rect 13434 37329 13542 37405
rect 13914 37329 14022 37405
rect 14682 37329 14790 37405
rect 15162 37329 15270 37405
rect 15930 37329 16038 37405
rect 16410 37329 16518 37405
rect 17178 37329 17286 37405
rect 17658 37329 17766 37405
rect 18426 37329 18534 37405
rect 18906 37329 19014 37405
rect 19674 37329 19782 37405
rect 20154 37329 20262 37405
rect 20922 37329 21030 37405
rect 21402 37329 21510 37405
rect 22170 37329 22278 37405
rect 22650 37329 22758 37405
rect 23418 37329 23526 37405
rect 23898 37329 24006 37405
rect 24666 37329 24774 37405
rect 25146 37329 25254 37405
rect 25914 37329 26022 37405
rect 26394 37329 26502 37405
rect 27162 37329 27270 37405
rect 27642 37329 27750 37405
rect 28410 37329 28518 37405
rect 28890 37329 28998 37405
rect 29658 37329 29766 37405
rect 30138 37329 30246 37405
rect 30906 37329 31014 37405
rect 31386 37329 31494 37405
rect 32154 37329 32262 37405
rect 32634 37329 32742 37405
rect 33402 37329 33510 37405
rect 33882 37329 33990 37405
rect 34650 37329 34758 37405
rect 35130 37329 35238 37405
rect 35898 37329 36006 37405
rect 36378 37329 36486 37405
rect 37146 37329 37254 37405
rect 37626 37329 37734 37405
rect 38394 37329 38502 37405
rect 38874 37329 38982 37405
rect 39642 37329 39750 37405
rect 0 37233 39936 37281
rect 186 37075 294 37185
rect 954 37075 1062 37185
rect 1434 37075 1542 37185
rect 2202 37075 2310 37185
rect 2682 37075 2790 37185
rect 3450 37075 3558 37185
rect 3930 37075 4038 37185
rect 4698 37075 4806 37185
rect 5178 37075 5286 37185
rect 5946 37075 6054 37185
rect 6426 37075 6534 37185
rect 7194 37075 7302 37185
rect 7674 37075 7782 37185
rect 8442 37075 8550 37185
rect 8922 37075 9030 37185
rect 9690 37075 9798 37185
rect 10170 37075 10278 37185
rect 10938 37075 11046 37185
rect 11418 37075 11526 37185
rect 12186 37075 12294 37185
rect 12666 37075 12774 37185
rect 13434 37075 13542 37185
rect 13914 37075 14022 37185
rect 14682 37075 14790 37185
rect 15162 37075 15270 37185
rect 15930 37075 16038 37185
rect 16410 37075 16518 37185
rect 17178 37075 17286 37185
rect 17658 37075 17766 37185
rect 18426 37075 18534 37185
rect 18906 37075 19014 37185
rect 19674 37075 19782 37185
rect 20154 37075 20262 37185
rect 20922 37075 21030 37185
rect 21402 37075 21510 37185
rect 22170 37075 22278 37185
rect 22650 37075 22758 37185
rect 23418 37075 23526 37185
rect 23898 37075 24006 37185
rect 24666 37075 24774 37185
rect 25146 37075 25254 37185
rect 25914 37075 26022 37185
rect 26394 37075 26502 37185
rect 27162 37075 27270 37185
rect 27642 37075 27750 37185
rect 28410 37075 28518 37185
rect 28890 37075 28998 37185
rect 29658 37075 29766 37185
rect 30138 37075 30246 37185
rect 30906 37075 31014 37185
rect 31386 37075 31494 37185
rect 32154 37075 32262 37185
rect 32634 37075 32742 37185
rect 33402 37075 33510 37185
rect 33882 37075 33990 37185
rect 34650 37075 34758 37185
rect 35130 37075 35238 37185
rect 35898 37075 36006 37185
rect 36378 37075 36486 37185
rect 37146 37075 37254 37185
rect 37626 37075 37734 37185
rect 38394 37075 38502 37185
rect 38874 37075 38982 37185
rect 39642 37075 39750 37185
rect 0 36979 39936 37027
rect 186 36855 294 36931
rect 954 36855 1062 36931
rect 1434 36855 1542 36931
rect 2202 36855 2310 36931
rect 2682 36855 2790 36931
rect 3450 36855 3558 36931
rect 3930 36855 4038 36931
rect 4698 36855 4806 36931
rect 5178 36855 5286 36931
rect 5946 36855 6054 36931
rect 6426 36855 6534 36931
rect 7194 36855 7302 36931
rect 7674 36855 7782 36931
rect 8442 36855 8550 36931
rect 8922 36855 9030 36931
rect 9690 36855 9798 36931
rect 10170 36855 10278 36931
rect 10938 36855 11046 36931
rect 11418 36855 11526 36931
rect 12186 36855 12294 36931
rect 12666 36855 12774 36931
rect 13434 36855 13542 36931
rect 13914 36855 14022 36931
rect 14682 36855 14790 36931
rect 15162 36855 15270 36931
rect 15930 36855 16038 36931
rect 16410 36855 16518 36931
rect 17178 36855 17286 36931
rect 17658 36855 17766 36931
rect 18426 36855 18534 36931
rect 18906 36855 19014 36931
rect 19674 36855 19782 36931
rect 20154 36855 20262 36931
rect 20922 36855 21030 36931
rect 21402 36855 21510 36931
rect 22170 36855 22278 36931
rect 22650 36855 22758 36931
rect 23418 36855 23526 36931
rect 23898 36855 24006 36931
rect 24666 36855 24774 36931
rect 25146 36855 25254 36931
rect 25914 36855 26022 36931
rect 26394 36855 26502 36931
rect 27162 36855 27270 36931
rect 27642 36855 27750 36931
rect 28410 36855 28518 36931
rect 28890 36855 28998 36931
rect 29658 36855 29766 36931
rect 30138 36855 30246 36931
rect 30906 36855 31014 36931
rect 31386 36855 31494 36931
rect 32154 36855 32262 36931
rect 32634 36855 32742 36931
rect 33402 36855 33510 36931
rect 33882 36855 33990 36931
rect 34650 36855 34758 36931
rect 35130 36855 35238 36931
rect 35898 36855 36006 36931
rect 36378 36855 36486 36931
rect 37146 36855 37254 36931
rect 37626 36855 37734 36931
rect 38394 36855 38502 36931
rect 38874 36855 38982 36931
rect 39642 36855 39750 36931
rect 0 36759 39936 36807
rect 0 36663 39936 36711
rect 186 36539 294 36615
rect 954 36539 1062 36615
rect 1434 36539 1542 36615
rect 2202 36539 2310 36615
rect 2682 36539 2790 36615
rect 3450 36539 3558 36615
rect 3930 36539 4038 36615
rect 4698 36539 4806 36615
rect 5178 36539 5286 36615
rect 5946 36539 6054 36615
rect 6426 36539 6534 36615
rect 7194 36539 7302 36615
rect 7674 36539 7782 36615
rect 8442 36539 8550 36615
rect 8922 36539 9030 36615
rect 9690 36539 9798 36615
rect 10170 36539 10278 36615
rect 10938 36539 11046 36615
rect 11418 36539 11526 36615
rect 12186 36539 12294 36615
rect 12666 36539 12774 36615
rect 13434 36539 13542 36615
rect 13914 36539 14022 36615
rect 14682 36539 14790 36615
rect 15162 36539 15270 36615
rect 15930 36539 16038 36615
rect 16410 36539 16518 36615
rect 17178 36539 17286 36615
rect 17658 36539 17766 36615
rect 18426 36539 18534 36615
rect 18906 36539 19014 36615
rect 19674 36539 19782 36615
rect 20154 36539 20262 36615
rect 20922 36539 21030 36615
rect 21402 36539 21510 36615
rect 22170 36539 22278 36615
rect 22650 36539 22758 36615
rect 23418 36539 23526 36615
rect 23898 36539 24006 36615
rect 24666 36539 24774 36615
rect 25146 36539 25254 36615
rect 25914 36539 26022 36615
rect 26394 36539 26502 36615
rect 27162 36539 27270 36615
rect 27642 36539 27750 36615
rect 28410 36539 28518 36615
rect 28890 36539 28998 36615
rect 29658 36539 29766 36615
rect 30138 36539 30246 36615
rect 30906 36539 31014 36615
rect 31386 36539 31494 36615
rect 32154 36539 32262 36615
rect 32634 36539 32742 36615
rect 33402 36539 33510 36615
rect 33882 36539 33990 36615
rect 34650 36539 34758 36615
rect 35130 36539 35238 36615
rect 35898 36539 36006 36615
rect 36378 36539 36486 36615
rect 37146 36539 37254 36615
rect 37626 36539 37734 36615
rect 38394 36539 38502 36615
rect 38874 36539 38982 36615
rect 39642 36539 39750 36615
rect 0 36443 39936 36491
rect 186 36285 294 36395
rect 954 36285 1062 36395
rect 1434 36285 1542 36395
rect 2202 36285 2310 36395
rect 2682 36285 2790 36395
rect 3450 36285 3558 36395
rect 3930 36285 4038 36395
rect 4698 36285 4806 36395
rect 5178 36285 5286 36395
rect 5946 36285 6054 36395
rect 6426 36285 6534 36395
rect 7194 36285 7302 36395
rect 7674 36285 7782 36395
rect 8442 36285 8550 36395
rect 8922 36285 9030 36395
rect 9690 36285 9798 36395
rect 10170 36285 10278 36395
rect 10938 36285 11046 36395
rect 11418 36285 11526 36395
rect 12186 36285 12294 36395
rect 12666 36285 12774 36395
rect 13434 36285 13542 36395
rect 13914 36285 14022 36395
rect 14682 36285 14790 36395
rect 15162 36285 15270 36395
rect 15930 36285 16038 36395
rect 16410 36285 16518 36395
rect 17178 36285 17286 36395
rect 17658 36285 17766 36395
rect 18426 36285 18534 36395
rect 18906 36285 19014 36395
rect 19674 36285 19782 36395
rect 20154 36285 20262 36395
rect 20922 36285 21030 36395
rect 21402 36285 21510 36395
rect 22170 36285 22278 36395
rect 22650 36285 22758 36395
rect 23418 36285 23526 36395
rect 23898 36285 24006 36395
rect 24666 36285 24774 36395
rect 25146 36285 25254 36395
rect 25914 36285 26022 36395
rect 26394 36285 26502 36395
rect 27162 36285 27270 36395
rect 27642 36285 27750 36395
rect 28410 36285 28518 36395
rect 28890 36285 28998 36395
rect 29658 36285 29766 36395
rect 30138 36285 30246 36395
rect 30906 36285 31014 36395
rect 31386 36285 31494 36395
rect 32154 36285 32262 36395
rect 32634 36285 32742 36395
rect 33402 36285 33510 36395
rect 33882 36285 33990 36395
rect 34650 36285 34758 36395
rect 35130 36285 35238 36395
rect 35898 36285 36006 36395
rect 36378 36285 36486 36395
rect 37146 36285 37254 36395
rect 37626 36285 37734 36395
rect 38394 36285 38502 36395
rect 38874 36285 38982 36395
rect 39642 36285 39750 36395
rect 0 36189 39936 36237
rect 186 36065 294 36141
rect 954 36065 1062 36141
rect 1434 36065 1542 36141
rect 2202 36065 2310 36141
rect 2682 36065 2790 36141
rect 3450 36065 3558 36141
rect 3930 36065 4038 36141
rect 4698 36065 4806 36141
rect 5178 36065 5286 36141
rect 5946 36065 6054 36141
rect 6426 36065 6534 36141
rect 7194 36065 7302 36141
rect 7674 36065 7782 36141
rect 8442 36065 8550 36141
rect 8922 36065 9030 36141
rect 9690 36065 9798 36141
rect 10170 36065 10278 36141
rect 10938 36065 11046 36141
rect 11418 36065 11526 36141
rect 12186 36065 12294 36141
rect 12666 36065 12774 36141
rect 13434 36065 13542 36141
rect 13914 36065 14022 36141
rect 14682 36065 14790 36141
rect 15162 36065 15270 36141
rect 15930 36065 16038 36141
rect 16410 36065 16518 36141
rect 17178 36065 17286 36141
rect 17658 36065 17766 36141
rect 18426 36065 18534 36141
rect 18906 36065 19014 36141
rect 19674 36065 19782 36141
rect 20154 36065 20262 36141
rect 20922 36065 21030 36141
rect 21402 36065 21510 36141
rect 22170 36065 22278 36141
rect 22650 36065 22758 36141
rect 23418 36065 23526 36141
rect 23898 36065 24006 36141
rect 24666 36065 24774 36141
rect 25146 36065 25254 36141
rect 25914 36065 26022 36141
rect 26394 36065 26502 36141
rect 27162 36065 27270 36141
rect 27642 36065 27750 36141
rect 28410 36065 28518 36141
rect 28890 36065 28998 36141
rect 29658 36065 29766 36141
rect 30138 36065 30246 36141
rect 30906 36065 31014 36141
rect 31386 36065 31494 36141
rect 32154 36065 32262 36141
rect 32634 36065 32742 36141
rect 33402 36065 33510 36141
rect 33882 36065 33990 36141
rect 34650 36065 34758 36141
rect 35130 36065 35238 36141
rect 35898 36065 36006 36141
rect 36378 36065 36486 36141
rect 37146 36065 37254 36141
rect 37626 36065 37734 36141
rect 38394 36065 38502 36141
rect 38874 36065 38982 36141
rect 39642 36065 39750 36141
rect 0 35969 39936 36017
rect 0 35873 39936 35921
rect 186 35749 294 35825
rect 954 35749 1062 35825
rect 1434 35749 1542 35825
rect 2202 35749 2310 35825
rect 2682 35749 2790 35825
rect 3450 35749 3558 35825
rect 3930 35749 4038 35825
rect 4698 35749 4806 35825
rect 5178 35749 5286 35825
rect 5946 35749 6054 35825
rect 6426 35749 6534 35825
rect 7194 35749 7302 35825
rect 7674 35749 7782 35825
rect 8442 35749 8550 35825
rect 8922 35749 9030 35825
rect 9690 35749 9798 35825
rect 10170 35749 10278 35825
rect 10938 35749 11046 35825
rect 11418 35749 11526 35825
rect 12186 35749 12294 35825
rect 12666 35749 12774 35825
rect 13434 35749 13542 35825
rect 13914 35749 14022 35825
rect 14682 35749 14790 35825
rect 15162 35749 15270 35825
rect 15930 35749 16038 35825
rect 16410 35749 16518 35825
rect 17178 35749 17286 35825
rect 17658 35749 17766 35825
rect 18426 35749 18534 35825
rect 18906 35749 19014 35825
rect 19674 35749 19782 35825
rect 20154 35749 20262 35825
rect 20922 35749 21030 35825
rect 21402 35749 21510 35825
rect 22170 35749 22278 35825
rect 22650 35749 22758 35825
rect 23418 35749 23526 35825
rect 23898 35749 24006 35825
rect 24666 35749 24774 35825
rect 25146 35749 25254 35825
rect 25914 35749 26022 35825
rect 26394 35749 26502 35825
rect 27162 35749 27270 35825
rect 27642 35749 27750 35825
rect 28410 35749 28518 35825
rect 28890 35749 28998 35825
rect 29658 35749 29766 35825
rect 30138 35749 30246 35825
rect 30906 35749 31014 35825
rect 31386 35749 31494 35825
rect 32154 35749 32262 35825
rect 32634 35749 32742 35825
rect 33402 35749 33510 35825
rect 33882 35749 33990 35825
rect 34650 35749 34758 35825
rect 35130 35749 35238 35825
rect 35898 35749 36006 35825
rect 36378 35749 36486 35825
rect 37146 35749 37254 35825
rect 37626 35749 37734 35825
rect 38394 35749 38502 35825
rect 38874 35749 38982 35825
rect 39642 35749 39750 35825
rect 0 35653 39936 35701
rect 186 35495 294 35605
rect 954 35495 1062 35605
rect 1434 35495 1542 35605
rect 2202 35495 2310 35605
rect 2682 35495 2790 35605
rect 3450 35495 3558 35605
rect 3930 35495 4038 35605
rect 4698 35495 4806 35605
rect 5178 35495 5286 35605
rect 5946 35495 6054 35605
rect 6426 35495 6534 35605
rect 7194 35495 7302 35605
rect 7674 35495 7782 35605
rect 8442 35495 8550 35605
rect 8922 35495 9030 35605
rect 9690 35495 9798 35605
rect 10170 35495 10278 35605
rect 10938 35495 11046 35605
rect 11418 35495 11526 35605
rect 12186 35495 12294 35605
rect 12666 35495 12774 35605
rect 13434 35495 13542 35605
rect 13914 35495 14022 35605
rect 14682 35495 14790 35605
rect 15162 35495 15270 35605
rect 15930 35495 16038 35605
rect 16410 35495 16518 35605
rect 17178 35495 17286 35605
rect 17658 35495 17766 35605
rect 18426 35495 18534 35605
rect 18906 35495 19014 35605
rect 19674 35495 19782 35605
rect 20154 35495 20262 35605
rect 20922 35495 21030 35605
rect 21402 35495 21510 35605
rect 22170 35495 22278 35605
rect 22650 35495 22758 35605
rect 23418 35495 23526 35605
rect 23898 35495 24006 35605
rect 24666 35495 24774 35605
rect 25146 35495 25254 35605
rect 25914 35495 26022 35605
rect 26394 35495 26502 35605
rect 27162 35495 27270 35605
rect 27642 35495 27750 35605
rect 28410 35495 28518 35605
rect 28890 35495 28998 35605
rect 29658 35495 29766 35605
rect 30138 35495 30246 35605
rect 30906 35495 31014 35605
rect 31386 35495 31494 35605
rect 32154 35495 32262 35605
rect 32634 35495 32742 35605
rect 33402 35495 33510 35605
rect 33882 35495 33990 35605
rect 34650 35495 34758 35605
rect 35130 35495 35238 35605
rect 35898 35495 36006 35605
rect 36378 35495 36486 35605
rect 37146 35495 37254 35605
rect 37626 35495 37734 35605
rect 38394 35495 38502 35605
rect 38874 35495 38982 35605
rect 39642 35495 39750 35605
rect 0 35399 39936 35447
rect 186 35275 294 35351
rect 954 35275 1062 35351
rect 1434 35275 1542 35351
rect 2202 35275 2310 35351
rect 2682 35275 2790 35351
rect 3450 35275 3558 35351
rect 3930 35275 4038 35351
rect 4698 35275 4806 35351
rect 5178 35275 5286 35351
rect 5946 35275 6054 35351
rect 6426 35275 6534 35351
rect 7194 35275 7302 35351
rect 7674 35275 7782 35351
rect 8442 35275 8550 35351
rect 8922 35275 9030 35351
rect 9690 35275 9798 35351
rect 10170 35275 10278 35351
rect 10938 35275 11046 35351
rect 11418 35275 11526 35351
rect 12186 35275 12294 35351
rect 12666 35275 12774 35351
rect 13434 35275 13542 35351
rect 13914 35275 14022 35351
rect 14682 35275 14790 35351
rect 15162 35275 15270 35351
rect 15930 35275 16038 35351
rect 16410 35275 16518 35351
rect 17178 35275 17286 35351
rect 17658 35275 17766 35351
rect 18426 35275 18534 35351
rect 18906 35275 19014 35351
rect 19674 35275 19782 35351
rect 20154 35275 20262 35351
rect 20922 35275 21030 35351
rect 21402 35275 21510 35351
rect 22170 35275 22278 35351
rect 22650 35275 22758 35351
rect 23418 35275 23526 35351
rect 23898 35275 24006 35351
rect 24666 35275 24774 35351
rect 25146 35275 25254 35351
rect 25914 35275 26022 35351
rect 26394 35275 26502 35351
rect 27162 35275 27270 35351
rect 27642 35275 27750 35351
rect 28410 35275 28518 35351
rect 28890 35275 28998 35351
rect 29658 35275 29766 35351
rect 30138 35275 30246 35351
rect 30906 35275 31014 35351
rect 31386 35275 31494 35351
rect 32154 35275 32262 35351
rect 32634 35275 32742 35351
rect 33402 35275 33510 35351
rect 33882 35275 33990 35351
rect 34650 35275 34758 35351
rect 35130 35275 35238 35351
rect 35898 35275 36006 35351
rect 36378 35275 36486 35351
rect 37146 35275 37254 35351
rect 37626 35275 37734 35351
rect 38394 35275 38502 35351
rect 38874 35275 38982 35351
rect 39642 35275 39750 35351
rect 0 35179 39936 35227
rect 0 35083 39936 35131
rect 186 34959 294 35035
rect 954 34959 1062 35035
rect 1434 34959 1542 35035
rect 2202 34959 2310 35035
rect 2682 34959 2790 35035
rect 3450 34959 3558 35035
rect 3930 34959 4038 35035
rect 4698 34959 4806 35035
rect 5178 34959 5286 35035
rect 5946 34959 6054 35035
rect 6426 34959 6534 35035
rect 7194 34959 7302 35035
rect 7674 34959 7782 35035
rect 8442 34959 8550 35035
rect 8922 34959 9030 35035
rect 9690 34959 9798 35035
rect 10170 34959 10278 35035
rect 10938 34959 11046 35035
rect 11418 34959 11526 35035
rect 12186 34959 12294 35035
rect 12666 34959 12774 35035
rect 13434 34959 13542 35035
rect 13914 34959 14022 35035
rect 14682 34959 14790 35035
rect 15162 34959 15270 35035
rect 15930 34959 16038 35035
rect 16410 34959 16518 35035
rect 17178 34959 17286 35035
rect 17658 34959 17766 35035
rect 18426 34959 18534 35035
rect 18906 34959 19014 35035
rect 19674 34959 19782 35035
rect 20154 34959 20262 35035
rect 20922 34959 21030 35035
rect 21402 34959 21510 35035
rect 22170 34959 22278 35035
rect 22650 34959 22758 35035
rect 23418 34959 23526 35035
rect 23898 34959 24006 35035
rect 24666 34959 24774 35035
rect 25146 34959 25254 35035
rect 25914 34959 26022 35035
rect 26394 34959 26502 35035
rect 27162 34959 27270 35035
rect 27642 34959 27750 35035
rect 28410 34959 28518 35035
rect 28890 34959 28998 35035
rect 29658 34959 29766 35035
rect 30138 34959 30246 35035
rect 30906 34959 31014 35035
rect 31386 34959 31494 35035
rect 32154 34959 32262 35035
rect 32634 34959 32742 35035
rect 33402 34959 33510 35035
rect 33882 34959 33990 35035
rect 34650 34959 34758 35035
rect 35130 34959 35238 35035
rect 35898 34959 36006 35035
rect 36378 34959 36486 35035
rect 37146 34959 37254 35035
rect 37626 34959 37734 35035
rect 38394 34959 38502 35035
rect 38874 34959 38982 35035
rect 39642 34959 39750 35035
rect 0 34863 39936 34911
rect 186 34705 294 34815
rect 954 34705 1062 34815
rect 1434 34705 1542 34815
rect 2202 34705 2310 34815
rect 2682 34705 2790 34815
rect 3450 34705 3558 34815
rect 3930 34705 4038 34815
rect 4698 34705 4806 34815
rect 5178 34705 5286 34815
rect 5946 34705 6054 34815
rect 6426 34705 6534 34815
rect 7194 34705 7302 34815
rect 7674 34705 7782 34815
rect 8442 34705 8550 34815
rect 8922 34705 9030 34815
rect 9690 34705 9798 34815
rect 10170 34705 10278 34815
rect 10938 34705 11046 34815
rect 11418 34705 11526 34815
rect 12186 34705 12294 34815
rect 12666 34705 12774 34815
rect 13434 34705 13542 34815
rect 13914 34705 14022 34815
rect 14682 34705 14790 34815
rect 15162 34705 15270 34815
rect 15930 34705 16038 34815
rect 16410 34705 16518 34815
rect 17178 34705 17286 34815
rect 17658 34705 17766 34815
rect 18426 34705 18534 34815
rect 18906 34705 19014 34815
rect 19674 34705 19782 34815
rect 20154 34705 20262 34815
rect 20922 34705 21030 34815
rect 21402 34705 21510 34815
rect 22170 34705 22278 34815
rect 22650 34705 22758 34815
rect 23418 34705 23526 34815
rect 23898 34705 24006 34815
rect 24666 34705 24774 34815
rect 25146 34705 25254 34815
rect 25914 34705 26022 34815
rect 26394 34705 26502 34815
rect 27162 34705 27270 34815
rect 27642 34705 27750 34815
rect 28410 34705 28518 34815
rect 28890 34705 28998 34815
rect 29658 34705 29766 34815
rect 30138 34705 30246 34815
rect 30906 34705 31014 34815
rect 31386 34705 31494 34815
rect 32154 34705 32262 34815
rect 32634 34705 32742 34815
rect 33402 34705 33510 34815
rect 33882 34705 33990 34815
rect 34650 34705 34758 34815
rect 35130 34705 35238 34815
rect 35898 34705 36006 34815
rect 36378 34705 36486 34815
rect 37146 34705 37254 34815
rect 37626 34705 37734 34815
rect 38394 34705 38502 34815
rect 38874 34705 38982 34815
rect 39642 34705 39750 34815
rect 0 34609 39936 34657
rect 186 34485 294 34561
rect 954 34485 1062 34561
rect 1434 34485 1542 34561
rect 2202 34485 2310 34561
rect 2682 34485 2790 34561
rect 3450 34485 3558 34561
rect 3930 34485 4038 34561
rect 4698 34485 4806 34561
rect 5178 34485 5286 34561
rect 5946 34485 6054 34561
rect 6426 34485 6534 34561
rect 7194 34485 7302 34561
rect 7674 34485 7782 34561
rect 8442 34485 8550 34561
rect 8922 34485 9030 34561
rect 9690 34485 9798 34561
rect 10170 34485 10278 34561
rect 10938 34485 11046 34561
rect 11418 34485 11526 34561
rect 12186 34485 12294 34561
rect 12666 34485 12774 34561
rect 13434 34485 13542 34561
rect 13914 34485 14022 34561
rect 14682 34485 14790 34561
rect 15162 34485 15270 34561
rect 15930 34485 16038 34561
rect 16410 34485 16518 34561
rect 17178 34485 17286 34561
rect 17658 34485 17766 34561
rect 18426 34485 18534 34561
rect 18906 34485 19014 34561
rect 19674 34485 19782 34561
rect 20154 34485 20262 34561
rect 20922 34485 21030 34561
rect 21402 34485 21510 34561
rect 22170 34485 22278 34561
rect 22650 34485 22758 34561
rect 23418 34485 23526 34561
rect 23898 34485 24006 34561
rect 24666 34485 24774 34561
rect 25146 34485 25254 34561
rect 25914 34485 26022 34561
rect 26394 34485 26502 34561
rect 27162 34485 27270 34561
rect 27642 34485 27750 34561
rect 28410 34485 28518 34561
rect 28890 34485 28998 34561
rect 29658 34485 29766 34561
rect 30138 34485 30246 34561
rect 30906 34485 31014 34561
rect 31386 34485 31494 34561
rect 32154 34485 32262 34561
rect 32634 34485 32742 34561
rect 33402 34485 33510 34561
rect 33882 34485 33990 34561
rect 34650 34485 34758 34561
rect 35130 34485 35238 34561
rect 35898 34485 36006 34561
rect 36378 34485 36486 34561
rect 37146 34485 37254 34561
rect 37626 34485 37734 34561
rect 38394 34485 38502 34561
rect 38874 34485 38982 34561
rect 39642 34485 39750 34561
rect 0 34389 39936 34437
rect 0 34293 39936 34341
rect 186 34169 294 34245
rect 954 34169 1062 34245
rect 1434 34169 1542 34245
rect 2202 34169 2310 34245
rect 2682 34169 2790 34245
rect 3450 34169 3558 34245
rect 3930 34169 4038 34245
rect 4698 34169 4806 34245
rect 5178 34169 5286 34245
rect 5946 34169 6054 34245
rect 6426 34169 6534 34245
rect 7194 34169 7302 34245
rect 7674 34169 7782 34245
rect 8442 34169 8550 34245
rect 8922 34169 9030 34245
rect 9690 34169 9798 34245
rect 10170 34169 10278 34245
rect 10938 34169 11046 34245
rect 11418 34169 11526 34245
rect 12186 34169 12294 34245
rect 12666 34169 12774 34245
rect 13434 34169 13542 34245
rect 13914 34169 14022 34245
rect 14682 34169 14790 34245
rect 15162 34169 15270 34245
rect 15930 34169 16038 34245
rect 16410 34169 16518 34245
rect 17178 34169 17286 34245
rect 17658 34169 17766 34245
rect 18426 34169 18534 34245
rect 18906 34169 19014 34245
rect 19674 34169 19782 34245
rect 20154 34169 20262 34245
rect 20922 34169 21030 34245
rect 21402 34169 21510 34245
rect 22170 34169 22278 34245
rect 22650 34169 22758 34245
rect 23418 34169 23526 34245
rect 23898 34169 24006 34245
rect 24666 34169 24774 34245
rect 25146 34169 25254 34245
rect 25914 34169 26022 34245
rect 26394 34169 26502 34245
rect 27162 34169 27270 34245
rect 27642 34169 27750 34245
rect 28410 34169 28518 34245
rect 28890 34169 28998 34245
rect 29658 34169 29766 34245
rect 30138 34169 30246 34245
rect 30906 34169 31014 34245
rect 31386 34169 31494 34245
rect 32154 34169 32262 34245
rect 32634 34169 32742 34245
rect 33402 34169 33510 34245
rect 33882 34169 33990 34245
rect 34650 34169 34758 34245
rect 35130 34169 35238 34245
rect 35898 34169 36006 34245
rect 36378 34169 36486 34245
rect 37146 34169 37254 34245
rect 37626 34169 37734 34245
rect 38394 34169 38502 34245
rect 38874 34169 38982 34245
rect 39642 34169 39750 34245
rect 0 34073 39936 34121
rect 186 33915 294 34025
rect 954 33915 1062 34025
rect 1434 33915 1542 34025
rect 2202 33915 2310 34025
rect 2682 33915 2790 34025
rect 3450 33915 3558 34025
rect 3930 33915 4038 34025
rect 4698 33915 4806 34025
rect 5178 33915 5286 34025
rect 5946 33915 6054 34025
rect 6426 33915 6534 34025
rect 7194 33915 7302 34025
rect 7674 33915 7782 34025
rect 8442 33915 8550 34025
rect 8922 33915 9030 34025
rect 9690 33915 9798 34025
rect 10170 33915 10278 34025
rect 10938 33915 11046 34025
rect 11418 33915 11526 34025
rect 12186 33915 12294 34025
rect 12666 33915 12774 34025
rect 13434 33915 13542 34025
rect 13914 33915 14022 34025
rect 14682 33915 14790 34025
rect 15162 33915 15270 34025
rect 15930 33915 16038 34025
rect 16410 33915 16518 34025
rect 17178 33915 17286 34025
rect 17658 33915 17766 34025
rect 18426 33915 18534 34025
rect 18906 33915 19014 34025
rect 19674 33915 19782 34025
rect 20154 33915 20262 34025
rect 20922 33915 21030 34025
rect 21402 33915 21510 34025
rect 22170 33915 22278 34025
rect 22650 33915 22758 34025
rect 23418 33915 23526 34025
rect 23898 33915 24006 34025
rect 24666 33915 24774 34025
rect 25146 33915 25254 34025
rect 25914 33915 26022 34025
rect 26394 33915 26502 34025
rect 27162 33915 27270 34025
rect 27642 33915 27750 34025
rect 28410 33915 28518 34025
rect 28890 33915 28998 34025
rect 29658 33915 29766 34025
rect 30138 33915 30246 34025
rect 30906 33915 31014 34025
rect 31386 33915 31494 34025
rect 32154 33915 32262 34025
rect 32634 33915 32742 34025
rect 33402 33915 33510 34025
rect 33882 33915 33990 34025
rect 34650 33915 34758 34025
rect 35130 33915 35238 34025
rect 35898 33915 36006 34025
rect 36378 33915 36486 34025
rect 37146 33915 37254 34025
rect 37626 33915 37734 34025
rect 38394 33915 38502 34025
rect 38874 33915 38982 34025
rect 39642 33915 39750 34025
rect 0 33819 39936 33867
rect 186 33695 294 33771
rect 954 33695 1062 33771
rect 1434 33695 1542 33771
rect 2202 33695 2310 33771
rect 2682 33695 2790 33771
rect 3450 33695 3558 33771
rect 3930 33695 4038 33771
rect 4698 33695 4806 33771
rect 5178 33695 5286 33771
rect 5946 33695 6054 33771
rect 6426 33695 6534 33771
rect 7194 33695 7302 33771
rect 7674 33695 7782 33771
rect 8442 33695 8550 33771
rect 8922 33695 9030 33771
rect 9690 33695 9798 33771
rect 10170 33695 10278 33771
rect 10938 33695 11046 33771
rect 11418 33695 11526 33771
rect 12186 33695 12294 33771
rect 12666 33695 12774 33771
rect 13434 33695 13542 33771
rect 13914 33695 14022 33771
rect 14682 33695 14790 33771
rect 15162 33695 15270 33771
rect 15930 33695 16038 33771
rect 16410 33695 16518 33771
rect 17178 33695 17286 33771
rect 17658 33695 17766 33771
rect 18426 33695 18534 33771
rect 18906 33695 19014 33771
rect 19674 33695 19782 33771
rect 20154 33695 20262 33771
rect 20922 33695 21030 33771
rect 21402 33695 21510 33771
rect 22170 33695 22278 33771
rect 22650 33695 22758 33771
rect 23418 33695 23526 33771
rect 23898 33695 24006 33771
rect 24666 33695 24774 33771
rect 25146 33695 25254 33771
rect 25914 33695 26022 33771
rect 26394 33695 26502 33771
rect 27162 33695 27270 33771
rect 27642 33695 27750 33771
rect 28410 33695 28518 33771
rect 28890 33695 28998 33771
rect 29658 33695 29766 33771
rect 30138 33695 30246 33771
rect 30906 33695 31014 33771
rect 31386 33695 31494 33771
rect 32154 33695 32262 33771
rect 32634 33695 32742 33771
rect 33402 33695 33510 33771
rect 33882 33695 33990 33771
rect 34650 33695 34758 33771
rect 35130 33695 35238 33771
rect 35898 33695 36006 33771
rect 36378 33695 36486 33771
rect 37146 33695 37254 33771
rect 37626 33695 37734 33771
rect 38394 33695 38502 33771
rect 38874 33695 38982 33771
rect 39642 33695 39750 33771
rect 0 33599 39936 33647
rect 0 33503 39936 33551
rect 186 33379 294 33455
rect 954 33379 1062 33455
rect 1434 33379 1542 33455
rect 2202 33379 2310 33455
rect 2682 33379 2790 33455
rect 3450 33379 3558 33455
rect 3930 33379 4038 33455
rect 4698 33379 4806 33455
rect 5178 33379 5286 33455
rect 5946 33379 6054 33455
rect 6426 33379 6534 33455
rect 7194 33379 7302 33455
rect 7674 33379 7782 33455
rect 8442 33379 8550 33455
rect 8922 33379 9030 33455
rect 9690 33379 9798 33455
rect 10170 33379 10278 33455
rect 10938 33379 11046 33455
rect 11418 33379 11526 33455
rect 12186 33379 12294 33455
rect 12666 33379 12774 33455
rect 13434 33379 13542 33455
rect 13914 33379 14022 33455
rect 14682 33379 14790 33455
rect 15162 33379 15270 33455
rect 15930 33379 16038 33455
rect 16410 33379 16518 33455
rect 17178 33379 17286 33455
rect 17658 33379 17766 33455
rect 18426 33379 18534 33455
rect 18906 33379 19014 33455
rect 19674 33379 19782 33455
rect 20154 33379 20262 33455
rect 20922 33379 21030 33455
rect 21402 33379 21510 33455
rect 22170 33379 22278 33455
rect 22650 33379 22758 33455
rect 23418 33379 23526 33455
rect 23898 33379 24006 33455
rect 24666 33379 24774 33455
rect 25146 33379 25254 33455
rect 25914 33379 26022 33455
rect 26394 33379 26502 33455
rect 27162 33379 27270 33455
rect 27642 33379 27750 33455
rect 28410 33379 28518 33455
rect 28890 33379 28998 33455
rect 29658 33379 29766 33455
rect 30138 33379 30246 33455
rect 30906 33379 31014 33455
rect 31386 33379 31494 33455
rect 32154 33379 32262 33455
rect 32634 33379 32742 33455
rect 33402 33379 33510 33455
rect 33882 33379 33990 33455
rect 34650 33379 34758 33455
rect 35130 33379 35238 33455
rect 35898 33379 36006 33455
rect 36378 33379 36486 33455
rect 37146 33379 37254 33455
rect 37626 33379 37734 33455
rect 38394 33379 38502 33455
rect 38874 33379 38982 33455
rect 39642 33379 39750 33455
rect 0 33283 39936 33331
rect 186 33125 294 33235
rect 954 33125 1062 33235
rect 1434 33125 1542 33235
rect 2202 33125 2310 33235
rect 2682 33125 2790 33235
rect 3450 33125 3558 33235
rect 3930 33125 4038 33235
rect 4698 33125 4806 33235
rect 5178 33125 5286 33235
rect 5946 33125 6054 33235
rect 6426 33125 6534 33235
rect 7194 33125 7302 33235
rect 7674 33125 7782 33235
rect 8442 33125 8550 33235
rect 8922 33125 9030 33235
rect 9690 33125 9798 33235
rect 10170 33125 10278 33235
rect 10938 33125 11046 33235
rect 11418 33125 11526 33235
rect 12186 33125 12294 33235
rect 12666 33125 12774 33235
rect 13434 33125 13542 33235
rect 13914 33125 14022 33235
rect 14682 33125 14790 33235
rect 15162 33125 15270 33235
rect 15930 33125 16038 33235
rect 16410 33125 16518 33235
rect 17178 33125 17286 33235
rect 17658 33125 17766 33235
rect 18426 33125 18534 33235
rect 18906 33125 19014 33235
rect 19674 33125 19782 33235
rect 20154 33125 20262 33235
rect 20922 33125 21030 33235
rect 21402 33125 21510 33235
rect 22170 33125 22278 33235
rect 22650 33125 22758 33235
rect 23418 33125 23526 33235
rect 23898 33125 24006 33235
rect 24666 33125 24774 33235
rect 25146 33125 25254 33235
rect 25914 33125 26022 33235
rect 26394 33125 26502 33235
rect 27162 33125 27270 33235
rect 27642 33125 27750 33235
rect 28410 33125 28518 33235
rect 28890 33125 28998 33235
rect 29658 33125 29766 33235
rect 30138 33125 30246 33235
rect 30906 33125 31014 33235
rect 31386 33125 31494 33235
rect 32154 33125 32262 33235
rect 32634 33125 32742 33235
rect 33402 33125 33510 33235
rect 33882 33125 33990 33235
rect 34650 33125 34758 33235
rect 35130 33125 35238 33235
rect 35898 33125 36006 33235
rect 36378 33125 36486 33235
rect 37146 33125 37254 33235
rect 37626 33125 37734 33235
rect 38394 33125 38502 33235
rect 38874 33125 38982 33235
rect 39642 33125 39750 33235
rect 0 33029 39936 33077
rect 186 32905 294 32981
rect 954 32905 1062 32981
rect 1434 32905 1542 32981
rect 2202 32905 2310 32981
rect 2682 32905 2790 32981
rect 3450 32905 3558 32981
rect 3930 32905 4038 32981
rect 4698 32905 4806 32981
rect 5178 32905 5286 32981
rect 5946 32905 6054 32981
rect 6426 32905 6534 32981
rect 7194 32905 7302 32981
rect 7674 32905 7782 32981
rect 8442 32905 8550 32981
rect 8922 32905 9030 32981
rect 9690 32905 9798 32981
rect 10170 32905 10278 32981
rect 10938 32905 11046 32981
rect 11418 32905 11526 32981
rect 12186 32905 12294 32981
rect 12666 32905 12774 32981
rect 13434 32905 13542 32981
rect 13914 32905 14022 32981
rect 14682 32905 14790 32981
rect 15162 32905 15270 32981
rect 15930 32905 16038 32981
rect 16410 32905 16518 32981
rect 17178 32905 17286 32981
rect 17658 32905 17766 32981
rect 18426 32905 18534 32981
rect 18906 32905 19014 32981
rect 19674 32905 19782 32981
rect 20154 32905 20262 32981
rect 20922 32905 21030 32981
rect 21402 32905 21510 32981
rect 22170 32905 22278 32981
rect 22650 32905 22758 32981
rect 23418 32905 23526 32981
rect 23898 32905 24006 32981
rect 24666 32905 24774 32981
rect 25146 32905 25254 32981
rect 25914 32905 26022 32981
rect 26394 32905 26502 32981
rect 27162 32905 27270 32981
rect 27642 32905 27750 32981
rect 28410 32905 28518 32981
rect 28890 32905 28998 32981
rect 29658 32905 29766 32981
rect 30138 32905 30246 32981
rect 30906 32905 31014 32981
rect 31386 32905 31494 32981
rect 32154 32905 32262 32981
rect 32634 32905 32742 32981
rect 33402 32905 33510 32981
rect 33882 32905 33990 32981
rect 34650 32905 34758 32981
rect 35130 32905 35238 32981
rect 35898 32905 36006 32981
rect 36378 32905 36486 32981
rect 37146 32905 37254 32981
rect 37626 32905 37734 32981
rect 38394 32905 38502 32981
rect 38874 32905 38982 32981
rect 39642 32905 39750 32981
rect 0 32809 39936 32857
rect 0 32713 39936 32761
rect 186 32589 294 32665
rect 954 32589 1062 32665
rect 1434 32589 1542 32665
rect 2202 32589 2310 32665
rect 2682 32589 2790 32665
rect 3450 32589 3558 32665
rect 3930 32589 4038 32665
rect 4698 32589 4806 32665
rect 5178 32589 5286 32665
rect 5946 32589 6054 32665
rect 6426 32589 6534 32665
rect 7194 32589 7302 32665
rect 7674 32589 7782 32665
rect 8442 32589 8550 32665
rect 8922 32589 9030 32665
rect 9690 32589 9798 32665
rect 10170 32589 10278 32665
rect 10938 32589 11046 32665
rect 11418 32589 11526 32665
rect 12186 32589 12294 32665
rect 12666 32589 12774 32665
rect 13434 32589 13542 32665
rect 13914 32589 14022 32665
rect 14682 32589 14790 32665
rect 15162 32589 15270 32665
rect 15930 32589 16038 32665
rect 16410 32589 16518 32665
rect 17178 32589 17286 32665
rect 17658 32589 17766 32665
rect 18426 32589 18534 32665
rect 18906 32589 19014 32665
rect 19674 32589 19782 32665
rect 20154 32589 20262 32665
rect 20922 32589 21030 32665
rect 21402 32589 21510 32665
rect 22170 32589 22278 32665
rect 22650 32589 22758 32665
rect 23418 32589 23526 32665
rect 23898 32589 24006 32665
rect 24666 32589 24774 32665
rect 25146 32589 25254 32665
rect 25914 32589 26022 32665
rect 26394 32589 26502 32665
rect 27162 32589 27270 32665
rect 27642 32589 27750 32665
rect 28410 32589 28518 32665
rect 28890 32589 28998 32665
rect 29658 32589 29766 32665
rect 30138 32589 30246 32665
rect 30906 32589 31014 32665
rect 31386 32589 31494 32665
rect 32154 32589 32262 32665
rect 32634 32589 32742 32665
rect 33402 32589 33510 32665
rect 33882 32589 33990 32665
rect 34650 32589 34758 32665
rect 35130 32589 35238 32665
rect 35898 32589 36006 32665
rect 36378 32589 36486 32665
rect 37146 32589 37254 32665
rect 37626 32589 37734 32665
rect 38394 32589 38502 32665
rect 38874 32589 38982 32665
rect 39642 32589 39750 32665
rect 0 32493 39936 32541
rect 186 32335 294 32445
rect 954 32335 1062 32445
rect 1434 32335 1542 32445
rect 2202 32335 2310 32445
rect 2682 32335 2790 32445
rect 3450 32335 3558 32445
rect 3930 32335 4038 32445
rect 4698 32335 4806 32445
rect 5178 32335 5286 32445
rect 5946 32335 6054 32445
rect 6426 32335 6534 32445
rect 7194 32335 7302 32445
rect 7674 32335 7782 32445
rect 8442 32335 8550 32445
rect 8922 32335 9030 32445
rect 9690 32335 9798 32445
rect 10170 32335 10278 32445
rect 10938 32335 11046 32445
rect 11418 32335 11526 32445
rect 12186 32335 12294 32445
rect 12666 32335 12774 32445
rect 13434 32335 13542 32445
rect 13914 32335 14022 32445
rect 14682 32335 14790 32445
rect 15162 32335 15270 32445
rect 15930 32335 16038 32445
rect 16410 32335 16518 32445
rect 17178 32335 17286 32445
rect 17658 32335 17766 32445
rect 18426 32335 18534 32445
rect 18906 32335 19014 32445
rect 19674 32335 19782 32445
rect 20154 32335 20262 32445
rect 20922 32335 21030 32445
rect 21402 32335 21510 32445
rect 22170 32335 22278 32445
rect 22650 32335 22758 32445
rect 23418 32335 23526 32445
rect 23898 32335 24006 32445
rect 24666 32335 24774 32445
rect 25146 32335 25254 32445
rect 25914 32335 26022 32445
rect 26394 32335 26502 32445
rect 27162 32335 27270 32445
rect 27642 32335 27750 32445
rect 28410 32335 28518 32445
rect 28890 32335 28998 32445
rect 29658 32335 29766 32445
rect 30138 32335 30246 32445
rect 30906 32335 31014 32445
rect 31386 32335 31494 32445
rect 32154 32335 32262 32445
rect 32634 32335 32742 32445
rect 33402 32335 33510 32445
rect 33882 32335 33990 32445
rect 34650 32335 34758 32445
rect 35130 32335 35238 32445
rect 35898 32335 36006 32445
rect 36378 32335 36486 32445
rect 37146 32335 37254 32445
rect 37626 32335 37734 32445
rect 38394 32335 38502 32445
rect 38874 32335 38982 32445
rect 39642 32335 39750 32445
rect 0 32239 39936 32287
rect 186 32115 294 32191
rect 954 32115 1062 32191
rect 1434 32115 1542 32191
rect 2202 32115 2310 32191
rect 2682 32115 2790 32191
rect 3450 32115 3558 32191
rect 3930 32115 4038 32191
rect 4698 32115 4806 32191
rect 5178 32115 5286 32191
rect 5946 32115 6054 32191
rect 6426 32115 6534 32191
rect 7194 32115 7302 32191
rect 7674 32115 7782 32191
rect 8442 32115 8550 32191
rect 8922 32115 9030 32191
rect 9690 32115 9798 32191
rect 10170 32115 10278 32191
rect 10938 32115 11046 32191
rect 11418 32115 11526 32191
rect 12186 32115 12294 32191
rect 12666 32115 12774 32191
rect 13434 32115 13542 32191
rect 13914 32115 14022 32191
rect 14682 32115 14790 32191
rect 15162 32115 15270 32191
rect 15930 32115 16038 32191
rect 16410 32115 16518 32191
rect 17178 32115 17286 32191
rect 17658 32115 17766 32191
rect 18426 32115 18534 32191
rect 18906 32115 19014 32191
rect 19674 32115 19782 32191
rect 20154 32115 20262 32191
rect 20922 32115 21030 32191
rect 21402 32115 21510 32191
rect 22170 32115 22278 32191
rect 22650 32115 22758 32191
rect 23418 32115 23526 32191
rect 23898 32115 24006 32191
rect 24666 32115 24774 32191
rect 25146 32115 25254 32191
rect 25914 32115 26022 32191
rect 26394 32115 26502 32191
rect 27162 32115 27270 32191
rect 27642 32115 27750 32191
rect 28410 32115 28518 32191
rect 28890 32115 28998 32191
rect 29658 32115 29766 32191
rect 30138 32115 30246 32191
rect 30906 32115 31014 32191
rect 31386 32115 31494 32191
rect 32154 32115 32262 32191
rect 32634 32115 32742 32191
rect 33402 32115 33510 32191
rect 33882 32115 33990 32191
rect 34650 32115 34758 32191
rect 35130 32115 35238 32191
rect 35898 32115 36006 32191
rect 36378 32115 36486 32191
rect 37146 32115 37254 32191
rect 37626 32115 37734 32191
rect 38394 32115 38502 32191
rect 38874 32115 38982 32191
rect 39642 32115 39750 32191
rect 0 32019 39936 32067
rect 0 31923 39936 31971
rect 186 31799 294 31875
rect 954 31799 1062 31875
rect 1434 31799 1542 31875
rect 2202 31799 2310 31875
rect 2682 31799 2790 31875
rect 3450 31799 3558 31875
rect 3930 31799 4038 31875
rect 4698 31799 4806 31875
rect 5178 31799 5286 31875
rect 5946 31799 6054 31875
rect 6426 31799 6534 31875
rect 7194 31799 7302 31875
rect 7674 31799 7782 31875
rect 8442 31799 8550 31875
rect 8922 31799 9030 31875
rect 9690 31799 9798 31875
rect 10170 31799 10278 31875
rect 10938 31799 11046 31875
rect 11418 31799 11526 31875
rect 12186 31799 12294 31875
rect 12666 31799 12774 31875
rect 13434 31799 13542 31875
rect 13914 31799 14022 31875
rect 14682 31799 14790 31875
rect 15162 31799 15270 31875
rect 15930 31799 16038 31875
rect 16410 31799 16518 31875
rect 17178 31799 17286 31875
rect 17658 31799 17766 31875
rect 18426 31799 18534 31875
rect 18906 31799 19014 31875
rect 19674 31799 19782 31875
rect 20154 31799 20262 31875
rect 20922 31799 21030 31875
rect 21402 31799 21510 31875
rect 22170 31799 22278 31875
rect 22650 31799 22758 31875
rect 23418 31799 23526 31875
rect 23898 31799 24006 31875
rect 24666 31799 24774 31875
rect 25146 31799 25254 31875
rect 25914 31799 26022 31875
rect 26394 31799 26502 31875
rect 27162 31799 27270 31875
rect 27642 31799 27750 31875
rect 28410 31799 28518 31875
rect 28890 31799 28998 31875
rect 29658 31799 29766 31875
rect 30138 31799 30246 31875
rect 30906 31799 31014 31875
rect 31386 31799 31494 31875
rect 32154 31799 32262 31875
rect 32634 31799 32742 31875
rect 33402 31799 33510 31875
rect 33882 31799 33990 31875
rect 34650 31799 34758 31875
rect 35130 31799 35238 31875
rect 35898 31799 36006 31875
rect 36378 31799 36486 31875
rect 37146 31799 37254 31875
rect 37626 31799 37734 31875
rect 38394 31799 38502 31875
rect 38874 31799 38982 31875
rect 39642 31799 39750 31875
rect 0 31703 39936 31751
rect 186 31545 294 31655
rect 954 31545 1062 31655
rect 1434 31545 1542 31655
rect 2202 31545 2310 31655
rect 2682 31545 2790 31655
rect 3450 31545 3558 31655
rect 3930 31545 4038 31655
rect 4698 31545 4806 31655
rect 5178 31545 5286 31655
rect 5946 31545 6054 31655
rect 6426 31545 6534 31655
rect 7194 31545 7302 31655
rect 7674 31545 7782 31655
rect 8442 31545 8550 31655
rect 8922 31545 9030 31655
rect 9690 31545 9798 31655
rect 10170 31545 10278 31655
rect 10938 31545 11046 31655
rect 11418 31545 11526 31655
rect 12186 31545 12294 31655
rect 12666 31545 12774 31655
rect 13434 31545 13542 31655
rect 13914 31545 14022 31655
rect 14682 31545 14790 31655
rect 15162 31545 15270 31655
rect 15930 31545 16038 31655
rect 16410 31545 16518 31655
rect 17178 31545 17286 31655
rect 17658 31545 17766 31655
rect 18426 31545 18534 31655
rect 18906 31545 19014 31655
rect 19674 31545 19782 31655
rect 20154 31545 20262 31655
rect 20922 31545 21030 31655
rect 21402 31545 21510 31655
rect 22170 31545 22278 31655
rect 22650 31545 22758 31655
rect 23418 31545 23526 31655
rect 23898 31545 24006 31655
rect 24666 31545 24774 31655
rect 25146 31545 25254 31655
rect 25914 31545 26022 31655
rect 26394 31545 26502 31655
rect 27162 31545 27270 31655
rect 27642 31545 27750 31655
rect 28410 31545 28518 31655
rect 28890 31545 28998 31655
rect 29658 31545 29766 31655
rect 30138 31545 30246 31655
rect 30906 31545 31014 31655
rect 31386 31545 31494 31655
rect 32154 31545 32262 31655
rect 32634 31545 32742 31655
rect 33402 31545 33510 31655
rect 33882 31545 33990 31655
rect 34650 31545 34758 31655
rect 35130 31545 35238 31655
rect 35898 31545 36006 31655
rect 36378 31545 36486 31655
rect 37146 31545 37254 31655
rect 37626 31545 37734 31655
rect 38394 31545 38502 31655
rect 38874 31545 38982 31655
rect 39642 31545 39750 31655
rect 0 31449 39936 31497
rect 186 31325 294 31401
rect 954 31325 1062 31401
rect 1434 31325 1542 31401
rect 2202 31325 2310 31401
rect 2682 31325 2790 31401
rect 3450 31325 3558 31401
rect 3930 31325 4038 31401
rect 4698 31325 4806 31401
rect 5178 31325 5286 31401
rect 5946 31325 6054 31401
rect 6426 31325 6534 31401
rect 7194 31325 7302 31401
rect 7674 31325 7782 31401
rect 8442 31325 8550 31401
rect 8922 31325 9030 31401
rect 9690 31325 9798 31401
rect 10170 31325 10278 31401
rect 10938 31325 11046 31401
rect 11418 31325 11526 31401
rect 12186 31325 12294 31401
rect 12666 31325 12774 31401
rect 13434 31325 13542 31401
rect 13914 31325 14022 31401
rect 14682 31325 14790 31401
rect 15162 31325 15270 31401
rect 15930 31325 16038 31401
rect 16410 31325 16518 31401
rect 17178 31325 17286 31401
rect 17658 31325 17766 31401
rect 18426 31325 18534 31401
rect 18906 31325 19014 31401
rect 19674 31325 19782 31401
rect 20154 31325 20262 31401
rect 20922 31325 21030 31401
rect 21402 31325 21510 31401
rect 22170 31325 22278 31401
rect 22650 31325 22758 31401
rect 23418 31325 23526 31401
rect 23898 31325 24006 31401
rect 24666 31325 24774 31401
rect 25146 31325 25254 31401
rect 25914 31325 26022 31401
rect 26394 31325 26502 31401
rect 27162 31325 27270 31401
rect 27642 31325 27750 31401
rect 28410 31325 28518 31401
rect 28890 31325 28998 31401
rect 29658 31325 29766 31401
rect 30138 31325 30246 31401
rect 30906 31325 31014 31401
rect 31386 31325 31494 31401
rect 32154 31325 32262 31401
rect 32634 31325 32742 31401
rect 33402 31325 33510 31401
rect 33882 31325 33990 31401
rect 34650 31325 34758 31401
rect 35130 31325 35238 31401
rect 35898 31325 36006 31401
rect 36378 31325 36486 31401
rect 37146 31325 37254 31401
rect 37626 31325 37734 31401
rect 38394 31325 38502 31401
rect 38874 31325 38982 31401
rect 39642 31325 39750 31401
rect 0 31229 39936 31277
rect 0 31133 39936 31181
rect 186 31009 294 31085
rect 954 31009 1062 31085
rect 1434 31009 1542 31085
rect 2202 31009 2310 31085
rect 2682 31009 2790 31085
rect 3450 31009 3558 31085
rect 3930 31009 4038 31085
rect 4698 31009 4806 31085
rect 5178 31009 5286 31085
rect 5946 31009 6054 31085
rect 6426 31009 6534 31085
rect 7194 31009 7302 31085
rect 7674 31009 7782 31085
rect 8442 31009 8550 31085
rect 8922 31009 9030 31085
rect 9690 31009 9798 31085
rect 10170 31009 10278 31085
rect 10938 31009 11046 31085
rect 11418 31009 11526 31085
rect 12186 31009 12294 31085
rect 12666 31009 12774 31085
rect 13434 31009 13542 31085
rect 13914 31009 14022 31085
rect 14682 31009 14790 31085
rect 15162 31009 15270 31085
rect 15930 31009 16038 31085
rect 16410 31009 16518 31085
rect 17178 31009 17286 31085
rect 17658 31009 17766 31085
rect 18426 31009 18534 31085
rect 18906 31009 19014 31085
rect 19674 31009 19782 31085
rect 20154 31009 20262 31085
rect 20922 31009 21030 31085
rect 21402 31009 21510 31085
rect 22170 31009 22278 31085
rect 22650 31009 22758 31085
rect 23418 31009 23526 31085
rect 23898 31009 24006 31085
rect 24666 31009 24774 31085
rect 25146 31009 25254 31085
rect 25914 31009 26022 31085
rect 26394 31009 26502 31085
rect 27162 31009 27270 31085
rect 27642 31009 27750 31085
rect 28410 31009 28518 31085
rect 28890 31009 28998 31085
rect 29658 31009 29766 31085
rect 30138 31009 30246 31085
rect 30906 31009 31014 31085
rect 31386 31009 31494 31085
rect 32154 31009 32262 31085
rect 32634 31009 32742 31085
rect 33402 31009 33510 31085
rect 33882 31009 33990 31085
rect 34650 31009 34758 31085
rect 35130 31009 35238 31085
rect 35898 31009 36006 31085
rect 36378 31009 36486 31085
rect 37146 31009 37254 31085
rect 37626 31009 37734 31085
rect 38394 31009 38502 31085
rect 38874 31009 38982 31085
rect 39642 31009 39750 31085
rect 0 30913 39936 30961
rect 186 30755 294 30865
rect 954 30755 1062 30865
rect 1434 30755 1542 30865
rect 2202 30755 2310 30865
rect 2682 30755 2790 30865
rect 3450 30755 3558 30865
rect 3930 30755 4038 30865
rect 4698 30755 4806 30865
rect 5178 30755 5286 30865
rect 5946 30755 6054 30865
rect 6426 30755 6534 30865
rect 7194 30755 7302 30865
rect 7674 30755 7782 30865
rect 8442 30755 8550 30865
rect 8922 30755 9030 30865
rect 9690 30755 9798 30865
rect 10170 30755 10278 30865
rect 10938 30755 11046 30865
rect 11418 30755 11526 30865
rect 12186 30755 12294 30865
rect 12666 30755 12774 30865
rect 13434 30755 13542 30865
rect 13914 30755 14022 30865
rect 14682 30755 14790 30865
rect 15162 30755 15270 30865
rect 15930 30755 16038 30865
rect 16410 30755 16518 30865
rect 17178 30755 17286 30865
rect 17658 30755 17766 30865
rect 18426 30755 18534 30865
rect 18906 30755 19014 30865
rect 19674 30755 19782 30865
rect 20154 30755 20262 30865
rect 20922 30755 21030 30865
rect 21402 30755 21510 30865
rect 22170 30755 22278 30865
rect 22650 30755 22758 30865
rect 23418 30755 23526 30865
rect 23898 30755 24006 30865
rect 24666 30755 24774 30865
rect 25146 30755 25254 30865
rect 25914 30755 26022 30865
rect 26394 30755 26502 30865
rect 27162 30755 27270 30865
rect 27642 30755 27750 30865
rect 28410 30755 28518 30865
rect 28890 30755 28998 30865
rect 29658 30755 29766 30865
rect 30138 30755 30246 30865
rect 30906 30755 31014 30865
rect 31386 30755 31494 30865
rect 32154 30755 32262 30865
rect 32634 30755 32742 30865
rect 33402 30755 33510 30865
rect 33882 30755 33990 30865
rect 34650 30755 34758 30865
rect 35130 30755 35238 30865
rect 35898 30755 36006 30865
rect 36378 30755 36486 30865
rect 37146 30755 37254 30865
rect 37626 30755 37734 30865
rect 38394 30755 38502 30865
rect 38874 30755 38982 30865
rect 39642 30755 39750 30865
rect 0 30659 39936 30707
rect 186 30535 294 30611
rect 954 30535 1062 30611
rect 1434 30535 1542 30611
rect 2202 30535 2310 30611
rect 2682 30535 2790 30611
rect 3450 30535 3558 30611
rect 3930 30535 4038 30611
rect 4698 30535 4806 30611
rect 5178 30535 5286 30611
rect 5946 30535 6054 30611
rect 6426 30535 6534 30611
rect 7194 30535 7302 30611
rect 7674 30535 7782 30611
rect 8442 30535 8550 30611
rect 8922 30535 9030 30611
rect 9690 30535 9798 30611
rect 10170 30535 10278 30611
rect 10938 30535 11046 30611
rect 11418 30535 11526 30611
rect 12186 30535 12294 30611
rect 12666 30535 12774 30611
rect 13434 30535 13542 30611
rect 13914 30535 14022 30611
rect 14682 30535 14790 30611
rect 15162 30535 15270 30611
rect 15930 30535 16038 30611
rect 16410 30535 16518 30611
rect 17178 30535 17286 30611
rect 17658 30535 17766 30611
rect 18426 30535 18534 30611
rect 18906 30535 19014 30611
rect 19674 30535 19782 30611
rect 20154 30535 20262 30611
rect 20922 30535 21030 30611
rect 21402 30535 21510 30611
rect 22170 30535 22278 30611
rect 22650 30535 22758 30611
rect 23418 30535 23526 30611
rect 23898 30535 24006 30611
rect 24666 30535 24774 30611
rect 25146 30535 25254 30611
rect 25914 30535 26022 30611
rect 26394 30535 26502 30611
rect 27162 30535 27270 30611
rect 27642 30535 27750 30611
rect 28410 30535 28518 30611
rect 28890 30535 28998 30611
rect 29658 30535 29766 30611
rect 30138 30535 30246 30611
rect 30906 30535 31014 30611
rect 31386 30535 31494 30611
rect 32154 30535 32262 30611
rect 32634 30535 32742 30611
rect 33402 30535 33510 30611
rect 33882 30535 33990 30611
rect 34650 30535 34758 30611
rect 35130 30535 35238 30611
rect 35898 30535 36006 30611
rect 36378 30535 36486 30611
rect 37146 30535 37254 30611
rect 37626 30535 37734 30611
rect 38394 30535 38502 30611
rect 38874 30535 38982 30611
rect 39642 30535 39750 30611
rect 0 30439 39936 30487
rect 0 30343 39936 30391
rect 186 30219 294 30295
rect 954 30219 1062 30295
rect 1434 30219 1542 30295
rect 2202 30219 2310 30295
rect 2682 30219 2790 30295
rect 3450 30219 3558 30295
rect 3930 30219 4038 30295
rect 4698 30219 4806 30295
rect 5178 30219 5286 30295
rect 5946 30219 6054 30295
rect 6426 30219 6534 30295
rect 7194 30219 7302 30295
rect 7674 30219 7782 30295
rect 8442 30219 8550 30295
rect 8922 30219 9030 30295
rect 9690 30219 9798 30295
rect 10170 30219 10278 30295
rect 10938 30219 11046 30295
rect 11418 30219 11526 30295
rect 12186 30219 12294 30295
rect 12666 30219 12774 30295
rect 13434 30219 13542 30295
rect 13914 30219 14022 30295
rect 14682 30219 14790 30295
rect 15162 30219 15270 30295
rect 15930 30219 16038 30295
rect 16410 30219 16518 30295
rect 17178 30219 17286 30295
rect 17658 30219 17766 30295
rect 18426 30219 18534 30295
rect 18906 30219 19014 30295
rect 19674 30219 19782 30295
rect 20154 30219 20262 30295
rect 20922 30219 21030 30295
rect 21402 30219 21510 30295
rect 22170 30219 22278 30295
rect 22650 30219 22758 30295
rect 23418 30219 23526 30295
rect 23898 30219 24006 30295
rect 24666 30219 24774 30295
rect 25146 30219 25254 30295
rect 25914 30219 26022 30295
rect 26394 30219 26502 30295
rect 27162 30219 27270 30295
rect 27642 30219 27750 30295
rect 28410 30219 28518 30295
rect 28890 30219 28998 30295
rect 29658 30219 29766 30295
rect 30138 30219 30246 30295
rect 30906 30219 31014 30295
rect 31386 30219 31494 30295
rect 32154 30219 32262 30295
rect 32634 30219 32742 30295
rect 33402 30219 33510 30295
rect 33882 30219 33990 30295
rect 34650 30219 34758 30295
rect 35130 30219 35238 30295
rect 35898 30219 36006 30295
rect 36378 30219 36486 30295
rect 37146 30219 37254 30295
rect 37626 30219 37734 30295
rect 38394 30219 38502 30295
rect 38874 30219 38982 30295
rect 39642 30219 39750 30295
rect 0 30123 39936 30171
rect 186 29965 294 30075
rect 954 29965 1062 30075
rect 1434 29965 1542 30075
rect 2202 29965 2310 30075
rect 2682 29965 2790 30075
rect 3450 29965 3558 30075
rect 3930 29965 4038 30075
rect 4698 29965 4806 30075
rect 5178 29965 5286 30075
rect 5946 29965 6054 30075
rect 6426 29965 6534 30075
rect 7194 29965 7302 30075
rect 7674 29965 7782 30075
rect 8442 29965 8550 30075
rect 8922 29965 9030 30075
rect 9690 29965 9798 30075
rect 10170 29965 10278 30075
rect 10938 29965 11046 30075
rect 11418 29965 11526 30075
rect 12186 29965 12294 30075
rect 12666 29965 12774 30075
rect 13434 29965 13542 30075
rect 13914 29965 14022 30075
rect 14682 29965 14790 30075
rect 15162 29965 15270 30075
rect 15930 29965 16038 30075
rect 16410 29965 16518 30075
rect 17178 29965 17286 30075
rect 17658 29965 17766 30075
rect 18426 29965 18534 30075
rect 18906 29965 19014 30075
rect 19674 29965 19782 30075
rect 20154 29965 20262 30075
rect 20922 29965 21030 30075
rect 21402 29965 21510 30075
rect 22170 29965 22278 30075
rect 22650 29965 22758 30075
rect 23418 29965 23526 30075
rect 23898 29965 24006 30075
rect 24666 29965 24774 30075
rect 25146 29965 25254 30075
rect 25914 29965 26022 30075
rect 26394 29965 26502 30075
rect 27162 29965 27270 30075
rect 27642 29965 27750 30075
rect 28410 29965 28518 30075
rect 28890 29965 28998 30075
rect 29658 29965 29766 30075
rect 30138 29965 30246 30075
rect 30906 29965 31014 30075
rect 31386 29965 31494 30075
rect 32154 29965 32262 30075
rect 32634 29965 32742 30075
rect 33402 29965 33510 30075
rect 33882 29965 33990 30075
rect 34650 29965 34758 30075
rect 35130 29965 35238 30075
rect 35898 29965 36006 30075
rect 36378 29965 36486 30075
rect 37146 29965 37254 30075
rect 37626 29965 37734 30075
rect 38394 29965 38502 30075
rect 38874 29965 38982 30075
rect 39642 29965 39750 30075
rect 0 29869 39936 29917
rect 186 29745 294 29821
rect 954 29745 1062 29821
rect 1434 29745 1542 29821
rect 2202 29745 2310 29821
rect 2682 29745 2790 29821
rect 3450 29745 3558 29821
rect 3930 29745 4038 29821
rect 4698 29745 4806 29821
rect 5178 29745 5286 29821
rect 5946 29745 6054 29821
rect 6426 29745 6534 29821
rect 7194 29745 7302 29821
rect 7674 29745 7782 29821
rect 8442 29745 8550 29821
rect 8922 29745 9030 29821
rect 9690 29745 9798 29821
rect 10170 29745 10278 29821
rect 10938 29745 11046 29821
rect 11418 29745 11526 29821
rect 12186 29745 12294 29821
rect 12666 29745 12774 29821
rect 13434 29745 13542 29821
rect 13914 29745 14022 29821
rect 14682 29745 14790 29821
rect 15162 29745 15270 29821
rect 15930 29745 16038 29821
rect 16410 29745 16518 29821
rect 17178 29745 17286 29821
rect 17658 29745 17766 29821
rect 18426 29745 18534 29821
rect 18906 29745 19014 29821
rect 19674 29745 19782 29821
rect 20154 29745 20262 29821
rect 20922 29745 21030 29821
rect 21402 29745 21510 29821
rect 22170 29745 22278 29821
rect 22650 29745 22758 29821
rect 23418 29745 23526 29821
rect 23898 29745 24006 29821
rect 24666 29745 24774 29821
rect 25146 29745 25254 29821
rect 25914 29745 26022 29821
rect 26394 29745 26502 29821
rect 27162 29745 27270 29821
rect 27642 29745 27750 29821
rect 28410 29745 28518 29821
rect 28890 29745 28998 29821
rect 29658 29745 29766 29821
rect 30138 29745 30246 29821
rect 30906 29745 31014 29821
rect 31386 29745 31494 29821
rect 32154 29745 32262 29821
rect 32634 29745 32742 29821
rect 33402 29745 33510 29821
rect 33882 29745 33990 29821
rect 34650 29745 34758 29821
rect 35130 29745 35238 29821
rect 35898 29745 36006 29821
rect 36378 29745 36486 29821
rect 37146 29745 37254 29821
rect 37626 29745 37734 29821
rect 38394 29745 38502 29821
rect 38874 29745 38982 29821
rect 39642 29745 39750 29821
rect 0 29649 39936 29697
rect 0 29553 39936 29601
rect 186 29429 294 29505
rect 954 29429 1062 29505
rect 1434 29429 1542 29505
rect 2202 29429 2310 29505
rect 2682 29429 2790 29505
rect 3450 29429 3558 29505
rect 3930 29429 4038 29505
rect 4698 29429 4806 29505
rect 5178 29429 5286 29505
rect 5946 29429 6054 29505
rect 6426 29429 6534 29505
rect 7194 29429 7302 29505
rect 7674 29429 7782 29505
rect 8442 29429 8550 29505
rect 8922 29429 9030 29505
rect 9690 29429 9798 29505
rect 10170 29429 10278 29505
rect 10938 29429 11046 29505
rect 11418 29429 11526 29505
rect 12186 29429 12294 29505
rect 12666 29429 12774 29505
rect 13434 29429 13542 29505
rect 13914 29429 14022 29505
rect 14682 29429 14790 29505
rect 15162 29429 15270 29505
rect 15930 29429 16038 29505
rect 16410 29429 16518 29505
rect 17178 29429 17286 29505
rect 17658 29429 17766 29505
rect 18426 29429 18534 29505
rect 18906 29429 19014 29505
rect 19674 29429 19782 29505
rect 20154 29429 20262 29505
rect 20922 29429 21030 29505
rect 21402 29429 21510 29505
rect 22170 29429 22278 29505
rect 22650 29429 22758 29505
rect 23418 29429 23526 29505
rect 23898 29429 24006 29505
rect 24666 29429 24774 29505
rect 25146 29429 25254 29505
rect 25914 29429 26022 29505
rect 26394 29429 26502 29505
rect 27162 29429 27270 29505
rect 27642 29429 27750 29505
rect 28410 29429 28518 29505
rect 28890 29429 28998 29505
rect 29658 29429 29766 29505
rect 30138 29429 30246 29505
rect 30906 29429 31014 29505
rect 31386 29429 31494 29505
rect 32154 29429 32262 29505
rect 32634 29429 32742 29505
rect 33402 29429 33510 29505
rect 33882 29429 33990 29505
rect 34650 29429 34758 29505
rect 35130 29429 35238 29505
rect 35898 29429 36006 29505
rect 36378 29429 36486 29505
rect 37146 29429 37254 29505
rect 37626 29429 37734 29505
rect 38394 29429 38502 29505
rect 38874 29429 38982 29505
rect 39642 29429 39750 29505
rect 0 29333 39936 29381
rect 186 29175 294 29285
rect 954 29175 1062 29285
rect 1434 29175 1542 29285
rect 2202 29175 2310 29285
rect 2682 29175 2790 29285
rect 3450 29175 3558 29285
rect 3930 29175 4038 29285
rect 4698 29175 4806 29285
rect 5178 29175 5286 29285
rect 5946 29175 6054 29285
rect 6426 29175 6534 29285
rect 7194 29175 7302 29285
rect 7674 29175 7782 29285
rect 8442 29175 8550 29285
rect 8922 29175 9030 29285
rect 9690 29175 9798 29285
rect 10170 29175 10278 29285
rect 10938 29175 11046 29285
rect 11418 29175 11526 29285
rect 12186 29175 12294 29285
rect 12666 29175 12774 29285
rect 13434 29175 13542 29285
rect 13914 29175 14022 29285
rect 14682 29175 14790 29285
rect 15162 29175 15270 29285
rect 15930 29175 16038 29285
rect 16410 29175 16518 29285
rect 17178 29175 17286 29285
rect 17658 29175 17766 29285
rect 18426 29175 18534 29285
rect 18906 29175 19014 29285
rect 19674 29175 19782 29285
rect 20154 29175 20262 29285
rect 20922 29175 21030 29285
rect 21402 29175 21510 29285
rect 22170 29175 22278 29285
rect 22650 29175 22758 29285
rect 23418 29175 23526 29285
rect 23898 29175 24006 29285
rect 24666 29175 24774 29285
rect 25146 29175 25254 29285
rect 25914 29175 26022 29285
rect 26394 29175 26502 29285
rect 27162 29175 27270 29285
rect 27642 29175 27750 29285
rect 28410 29175 28518 29285
rect 28890 29175 28998 29285
rect 29658 29175 29766 29285
rect 30138 29175 30246 29285
rect 30906 29175 31014 29285
rect 31386 29175 31494 29285
rect 32154 29175 32262 29285
rect 32634 29175 32742 29285
rect 33402 29175 33510 29285
rect 33882 29175 33990 29285
rect 34650 29175 34758 29285
rect 35130 29175 35238 29285
rect 35898 29175 36006 29285
rect 36378 29175 36486 29285
rect 37146 29175 37254 29285
rect 37626 29175 37734 29285
rect 38394 29175 38502 29285
rect 38874 29175 38982 29285
rect 39642 29175 39750 29285
rect 0 29079 39936 29127
rect 186 28955 294 29031
rect 954 28955 1062 29031
rect 1434 28955 1542 29031
rect 2202 28955 2310 29031
rect 2682 28955 2790 29031
rect 3450 28955 3558 29031
rect 3930 28955 4038 29031
rect 4698 28955 4806 29031
rect 5178 28955 5286 29031
rect 5946 28955 6054 29031
rect 6426 28955 6534 29031
rect 7194 28955 7302 29031
rect 7674 28955 7782 29031
rect 8442 28955 8550 29031
rect 8922 28955 9030 29031
rect 9690 28955 9798 29031
rect 10170 28955 10278 29031
rect 10938 28955 11046 29031
rect 11418 28955 11526 29031
rect 12186 28955 12294 29031
rect 12666 28955 12774 29031
rect 13434 28955 13542 29031
rect 13914 28955 14022 29031
rect 14682 28955 14790 29031
rect 15162 28955 15270 29031
rect 15930 28955 16038 29031
rect 16410 28955 16518 29031
rect 17178 28955 17286 29031
rect 17658 28955 17766 29031
rect 18426 28955 18534 29031
rect 18906 28955 19014 29031
rect 19674 28955 19782 29031
rect 20154 28955 20262 29031
rect 20922 28955 21030 29031
rect 21402 28955 21510 29031
rect 22170 28955 22278 29031
rect 22650 28955 22758 29031
rect 23418 28955 23526 29031
rect 23898 28955 24006 29031
rect 24666 28955 24774 29031
rect 25146 28955 25254 29031
rect 25914 28955 26022 29031
rect 26394 28955 26502 29031
rect 27162 28955 27270 29031
rect 27642 28955 27750 29031
rect 28410 28955 28518 29031
rect 28890 28955 28998 29031
rect 29658 28955 29766 29031
rect 30138 28955 30246 29031
rect 30906 28955 31014 29031
rect 31386 28955 31494 29031
rect 32154 28955 32262 29031
rect 32634 28955 32742 29031
rect 33402 28955 33510 29031
rect 33882 28955 33990 29031
rect 34650 28955 34758 29031
rect 35130 28955 35238 29031
rect 35898 28955 36006 29031
rect 36378 28955 36486 29031
rect 37146 28955 37254 29031
rect 37626 28955 37734 29031
rect 38394 28955 38502 29031
rect 38874 28955 38982 29031
rect 39642 28955 39750 29031
rect 0 28859 39936 28907
rect 0 28763 39936 28811
rect 186 28639 294 28715
rect 954 28639 1062 28715
rect 1434 28639 1542 28715
rect 2202 28639 2310 28715
rect 2682 28639 2790 28715
rect 3450 28639 3558 28715
rect 3930 28639 4038 28715
rect 4698 28639 4806 28715
rect 5178 28639 5286 28715
rect 5946 28639 6054 28715
rect 6426 28639 6534 28715
rect 7194 28639 7302 28715
rect 7674 28639 7782 28715
rect 8442 28639 8550 28715
rect 8922 28639 9030 28715
rect 9690 28639 9798 28715
rect 10170 28639 10278 28715
rect 10938 28639 11046 28715
rect 11418 28639 11526 28715
rect 12186 28639 12294 28715
rect 12666 28639 12774 28715
rect 13434 28639 13542 28715
rect 13914 28639 14022 28715
rect 14682 28639 14790 28715
rect 15162 28639 15270 28715
rect 15930 28639 16038 28715
rect 16410 28639 16518 28715
rect 17178 28639 17286 28715
rect 17658 28639 17766 28715
rect 18426 28639 18534 28715
rect 18906 28639 19014 28715
rect 19674 28639 19782 28715
rect 20154 28639 20262 28715
rect 20922 28639 21030 28715
rect 21402 28639 21510 28715
rect 22170 28639 22278 28715
rect 22650 28639 22758 28715
rect 23418 28639 23526 28715
rect 23898 28639 24006 28715
rect 24666 28639 24774 28715
rect 25146 28639 25254 28715
rect 25914 28639 26022 28715
rect 26394 28639 26502 28715
rect 27162 28639 27270 28715
rect 27642 28639 27750 28715
rect 28410 28639 28518 28715
rect 28890 28639 28998 28715
rect 29658 28639 29766 28715
rect 30138 28639 30246 28715
rect 30906 28639 31014 28715
rect 31386 28639 31494 28715
rect 32154 28639 32262 28715
rect 32634 28639 32742 28715
rect 33402 28639 33510 28715
rect 33882 28639 33990 28715
rect 34650 28639 34758 28715
rect 35130 28639 35238 28715
rect 35898 28639 36006 28715
rect 36378 28639 36486 28715
rect 37146 28639 37254 28715
rect 37626 28639 37734 28715
rect 38394 28639 38502 28715
rect 38874 28639 38982 28715
rect 39642 28639 39750 28715
rect 0 28543 39936 28591
rect 186 28385 294 28495
rect 954 28385 1062 28495
rect 1434 28385 1542 28495
rect 2202 28385 2310 28495
rect 2682 28385 2790 28495
rect 3450 28385 3558 28495
rect 3930 28385 4038 28495
rect 4698 28385 4806 28495
rect 5178 28385 5286 28495
rect 5946 28385 6054 28495
rect 6426 28385 6534 28495
rect 7194 28385 7302 28495
rect 7674 28385 7782 28495
rect 8442 28385 8550 28495
rect 8922 28385 9030 28495
rect 9690 28385 9798 28495
rect 10170 28385 10278 28495
rect 10938 28385 11046 28495
rect 11418 28385 11526 28495
rect 12186 28385 12294 28495
rect 12666 28385 12774 28495
rect 13434 28385 13542 28495
rect 13914 28385 14022 28495
rect 14682 28385 14790 28495
rect 15162 28385 15270 28495
rect 15930 28385 16038 28495
rect 16410 28385 16518 28495
rect 17178 28385 17286 28495
rect 17658 28385 17766 28495
rect 18426 28385 18534 28495
rect 18906 28385 19014 28495
rect 19674 28385 19782 28495
rect 20154 28385 20262 28495
rect 20922 28385 21030 28495
rect 21402 28385 21510 28495
rect 22170 28385 22278 28495
rect 22650 28385 22758 28495
rect 23418 28385 23526 28495
rect 23898 28385 24006 28495
rect 24666 28385 24774 28495
rect 25146 28385 25254 28495
rect 25914 28385 26022 28495
rect 26394 28385 26502 28495
rect 27162 28385 27270 28495
rect 27642 28385 27750 28495
rect 28410 28385 28518 28495
rect 28890 28385 28998 28495
rect 29658 28385 29766 28495
rect 30138 28385 30246 28495
rect 30906 28385 31014 28495
rect 31386 28385 31494 28495
rect 32154 28385 32262 28495
rect 32634 28385 32742 28495
rect 33402 28385 33510 28495
rect 33882 28385 33990 28495
rect 34650 28385 34758 28495
rect 35130 28385 35238 28495
rect 35898 28385 36006 28495
rect 36378 28385 36486 28495
rect 37146 28385 37254 28495
rect 37626 28385 37734 28495
rect 38394 28385 38502 28495
rect 38874 28385 38982 28495
rect 39642 28385 39750 28495
rect 0 28289 39936 28337
rect 186 28165 294 28241
rect 954 28165 1062 28241
rect 1434 28165 1542 28241
rect 2202 28165 2310 28241
rect 2682 28165 2790 28241
rect 3450 28165 3558 28241
rect 3930 28165 4038 28241
rect 4698 28165 4806 28241
rect 5178 28165 5286 28241
rect 5946 28165 6054 28241
rect 6426 28165 6534 28241
rect 7194 28165 7302 28241
rect 7674 28165 7782 28241
rect 8442 28165 8550 28241
rect 8922 28165 9030 28241
rect 9690 28165 9798 28241
rect 10170 28165 10278 28241
rect 10938 28165 11046 28241
rect 11418 28165 11526 28241
rect 12186 28165 12294 28241
rect 12666 28165 12774 28241
rect 13434 28165 13542 28241
rect 13914 28165 14022 28241
rect 14682 28165 14790 28241
rect 15162 28165 15270 28241
rect 15930 28165 16038 28241
rect 16410 28165 16518 28241
rect 17178 28165 17286 28241
rect 17658 28165 17766 28241
rect 18426 28165 18534 28241
rect 18906 28165 19014 28241
rect 19674 28165 19782 28241
rect 20154 28165 20262 28241
rect 20922 28165 21030 28241
rect 21402 28165 21510 28241
rect 22170 28165 22278 28241
rect 22650 28165 22758 28241
rect 23418 28165 23526 28241
rect 23898 28165 24006 28241
rect 24666 28165 24774 28241
rect 25146 28165 25254 28241
rect 25914 28165 26022 28241
rect 26394 28165 26502 28241
rect 27162 28165 27270 28241
rect 27642 28165 27750 28241
rect 28410 28165 28518 28241
rect 28890 28165 28998 28241
rect 29658 28165 29766 28241
rect 30138 28165 30246 28241
rect 30906 28165 31014 28241
rect 31386 28165 31494 28241
rect 32154 28165 32262 28241
rect 32634 28165 32742 28241
rect 33402 28165 33510 28241
rect 33882 28165 33990 28241
rect 34650 28165 34758 28241
rect 35130 28165 35238 28241
rect 35898 28165 36006 28241
rect 36378 28165 36486 28241
rect 37146 28165 37254 28241
rect 37626 28165 37734 28241
rect 38394 28165 38502 28241
rect 38874 28165 38982 28241
rect 39642 28165 39750 28241
rect 0 28069 39936 28117
rect 0 27973 39936 28021
rect 186 27849 294 27925
rect 954 27849 1062 27925
rect 1434 27849 1542 27925
rect 2202 27849 2310 27925
rect 2682 27849 2790 27925
rect 3450 27849 3558 27925
rect 3930 27849 4038 27925
rect 4698 27849 4806 27925
rect 5178 27849 5286 27925
rect 5946 27849 6054 27925
rect 6426 27849 6534 27925
rect 7194 27849 7302 27925
rect 7674 27849 7782 27925
rect 8442 27849 8550 27925
rect 8922 27849 9030 27925
rect 9690 27849 9798 27925
rect 10170 27849 10278 27925
rect 10938 27849 11046 27925
rect 11418 27849 11526 27925
rect 12186 27849 12294 27925
rect 12666 27849 12774 27925
rect 13434 27849 13542 27925
rect 13914 27849 14022 27925
rect 14682 27849 14790 27925
rect 15162 27849 15270 27925
rect 15930 27849 16038 27925
rect 16410 27849 16518 27925
rect 17178 27849 17286 27925
rect 17658 27849 17766 27925
rect 18426 27849 18534 27925
rect 18906 27849 19014 27925
rect 19674 27849 19782 27925
rect 20154 27849 20262 27925
rect 20922 27849 21030 27925
rect 21402 27849 21510 27925
rect 22170 27849 22278 27925
rect 22650 27849 22758 27925
rect 23418 27849 23526 27925
rect 23898 27849 24006 27925
rect 24666 27849 24774 27925
rect 25146 27849 25254 27925
rect 25914 27849 26022 27925
rect 26394 27849 26502 27925
rect 27162 27849 27270 27925
rect 27642 27849 27750 27925
rect 28410 27849 28518 27925
rect 28890 27849 28998 27925
rect 29658 27849 29766 27925
rect 30138 27849 30246 27925
rect 30906 27849 31014 27925
rect 31386 27849 31494 27925
rect 32154 27849 32262 27925
rect 32634 27849 32742 27925
rect 33402 27849 33510 27925
rect 33882 27849 33990 27925
rect 34650 27849 34758 27925
rect 35130 27849 35238 27925
rect 35898 27849 36006 27925
rect 36378 27849 36486 27925
rect 37146 27849 37254 27925
rect 37626 27849 37734 27925
rect 38394 27849 38502 27925
rect 38874 27849 38982 27925
rect 39642 27849 39750 27925
rect 0 27753 39936 27801
rect 186 27595 294 27705
rect 954 27595 1062 27705
rect 1434 27595 1542 27705
rect 2202 27595 2310 27705
rect 2682 27595 2790 27705
rect 3450 27595 3558 27705
rect 3930 27595 4038 27705
rect 4698 27595 4806 27705
rect 5178 27595 5286 27705
rect 5946 27595 6054 27705
rect 6426 27595 6534 27705
rect 7194 27595 7302 27705
rect 7674 27595 7782 27705
rect 8442 27595 8550 27705
rect 8922 27595 9030 27705
rect 9690 27595 9798 27705
rect 10170 27595 10278 27705
rect 10938 27595 11046 27705
rect 11418 27595 11526 27705
rect 12186 27595 12294 27705
rect 12666 27595 12774 27705
rect 13434 27595 13542 27705
rect 13914 27595 14022 27705
rect 14682 27595 14790 27705
rect 15162 27595 15270 27705
rect 15930 27595 16038 27705
rect 16410 27595 16518 27705
rect 17178 27595 17286 27705
rect 17658 27595 17766 27705
rect 18426 27595 18534 27705
rect 18906 27595 19014 27705
rect 19674 27595 19782 27705
rect 20154 27595 20262 27705
rect 20922 27595 21030 27705
rect 21402 27595 21510 27705
rect 22170 27595 22278 27705
rect 22650 27595 22758 27705
rect 23418 27595 23526 27705
rect 23898 27595 24006 27705
rect 24666 27595 24774 27705
rect 25146 27595 25254 27705
rect 25914 27595 26022 27705
rect 26394 27595 26502 27705
rect 27162 27595 27270 27705
rect 27642 27595 27750 27705
rect 28410 27595 28518 27705
rect 28890 27595 28998 27705
rect 29658 27595 29766 27705
rect 30138 27595 30246 27705
rect 30906 27595 31014 27705
rect 31386 27595 31494 27705
rect 32154 27595 32262 27705
rect 32634 27595 32742 27705
rect 33402 27595 33510 27705
rect 33882 27595 33990 27705
rect 34650 27595 34758 27705
rect 35130 27595 35238 27705
rect 35898 27595 36006 27705
rect 36378 27595 36486 27705
rect 37146 27595 37254 27705
rect 37626 27595 37734 27705
rect 38394 27595 38502 27705
rect 38874 27595 38982 27705
rect 39642 27595 39750 27705
rect 0 27499 39936 27547
rect 186 27375 294 27451
rect 954 27375 1062 27451
rect 1434 27375 1542 27451
rect 2202 27375 2310 27451
rect 2682 27375 2790 27451
rect 3450 27375 3558 27451
rect 3930 27375 4038 27451
rect 4698 27375 4806 27451
rect 5178 27375 5286 27451
rect 5946 27375 6054 27451
rect 6426 27375 6534 27451
rect 7194 27375 7302 27451
rect 7674 27375 7782 27451
rect 8442 27375 8550 27451
rect 8922 27375 9030 27451
rect 9690 27375 9798 27451
rect 10170 27375 10278 27451
rect 10938 27375 11046 27451
rect 11418 27375 11526 27451
rect 12186 27375 12294 27451
rect 12666 27375 12774 27451
rect 13434 27375 13542 27451
rect 13914 27375 14022 27451
rect 14682 27375 14790 27451
rect 15162 27375 15270 27451
rect 15930 27375 16038 27451
rect 16410 27375 16518 27451
rect 17178 27375 17286 27451
rect 17658 27375 17766 27451
rect 18426 27375 18534 27451
rect 18906 27375 19014 27451
rect 19674 27375 19782 27451
rect 20154 27375 20262 27451
rect 20922 27375 21030 27451
rect 21402 27375 21510 27451
rect 22170 27375 22278 27451
rect 22650 27375 22758 27451
rect 23418 27375 23526 27451
rect 23898 27375 24006 27451
rect 24666 27375 24774 27451
rect 25146 27375 25254 27451
rect 25914 27375 26022 27451
rect 26394 27375 26502 27451
rect 27162 27375 27270 27451
rect 27642 27375 27750 27451
rect 28410 27375 28518 27451
rect 28890 27375 28998 27451
rect 29658 27375 29766 27451
rect 30138 27375 30246 27451
rect 30906 27375 31014 27451
rect 31386 27375 31494 27451
rect 32154 27375 32262 27451
rect 32634 27375 32742 27451
rect 33402 27375 33510 27451
rect 33882 27375 33990 27451
rect 34650 27375 34758 27451
rect 35130 27375 35238 27451
rect 35898 27375 36006 27451
rect 36378 27375 36486 27451
rect 37146 27375 37254 27451
rect 37626 27375 37734 27451
rect 38394 27375 38502 27451
rect 38874 27375 38982 27451
rect 39642 27375 39750 27451
rect 0 27279 39936 27327
rect 0 27183 39936 27231
rect 186 27059 294 27135
rect 954 27059 1062 27135
rect 1434 27059 1542 27135
rect 2202 27059 2310 27135
rect 2682 27059 2790 27135
rect 3450 27059 3558 27135
rect 3930 27059 4038 27135
rect 4698 27059 4806 27135
rect 5178 27059 5286 27135
rect 5946 27059 6054 27135
rect 6426 27059 6534 27135
rect 7194 27059 7302 27135
rect 7674 27059 7782 27135
rect 8442 27059 8550 27135
rect 8922 27059 9030 27135
rect 9690 27059 9798 27135
rect 10170 27059 10278 27135
rect 10938 27059 11046 27135
rect 11418 27059 11526 27135
rect 12186 27059 12294 27135
rect 12666 27059 12774 27135
rect 13434 27059 13542 27135
rect 13914 27059 14022 27135
rect 14682 27059 14790 27135
rect 15162 27059 15270 27135
rect 15930 27059 16038 27135
rect 16410 27059 16518 27135
rect 17178 27059 17286 27135
rect 17658 27059 17766 27135
rect 18426 27059 18534 27135
rect 18906 27059 19014 27135
rect 19674 27059 19782 27135
rect 20154 27059 20262 27135
rect 20922 27059 21030 27135
rect 21402 27059 21510 27135
rect 22170 27059 22278 27135
rect 22650 27059 22758 27135
rect 23418 27059 23526 27135
rect 23898 27059 24006 27135
rect 24666 27059 24774 27135
rect 25146 27059 25254 27135
rect 25914 27059 26022 27135
rect 26394 27059 26502 27135
rect 27162 27059 27270 27135
rect 27642 27059 27750 27135
rect 28410 27059 28518 27135
rect 28890 27059 28998 27135
rect 29658 27059 29766 27135
rect 30138 27059 30246 27135
rect 30906 27059 31014 27135
rect 31386 27059 31494 27135
rect 32154 27059 32262 27135
rect 32634 27059 32742 27135
rect 33402 27059 33510 27135
rect 33882 27059 33990 27135
rect 34650 27059 34758 27135
rect 35130 27059 35238 27135
rect 35898 27059 36006 27135
rect 36378 27059 36486 27135
rect 37146 27059 37254 27135
rect 37626 27059 37734 27135
rect 38394 27059 38502 27135
rect 38874 27059 38982 27135
rect 39642 27059 39750 27135
rect 0 26963 39936 27011
rect 186 26805 294 26915
rect 954 26805 1062 26915
rect 1434 26805 1542 26915
rect 2202 26805 2310 26915
rect 2682 26805 2790 26915
rect 3450 26805 3558 26915
rect 3930 26805 4038 26915
rect 4698 26805 4806 26915
rect 5178 26805 5286 26915
rect 5946 26805 6054 26915
rect 6426 26805 6534 26915
rect 7194 26805 7302 26915
rect 7674 26805 7782 26915
rect 8442 26805 8550 26915
rect 8922 26805 9030 26915
rect 9690 26805 9798 26915
rect 10170 26805 10278 26915
rect 10938 26805 11046 26915
rect 11418 26805 11526 26915
rect 12186 26805 12294 26915
rect 12666 26805 12774 26915
rect 13434 26805 13542 26915
rect 13914 26805 14022 26915
rect 14682 26805 14790 26915
rect 15162 26805 15270 26915
rect 15930 26805 16038 26915
rect 16410 26805 16518 26915
rect 17178 26805 17286 26915
rect 17658 26805 17766 26915
rect 18426 26805 18534 26915
rect 18906 26805 19014 26915
rect 19674 26805 19782 26915
rect 20154 26805 20262 26915
rect 20922 26805 21030 26915
rect 21402 26805 21510 26915
rect 22170 26805 22278 26915
rect 22650 26805 22758 26915
rect 23418 26805 23526 26915
rect 23898 26805 24006 26915
rect 24666 26805 24774 26915
rect 25146 26805 25254 26915
rect 25914 26805 26022 26915
rect 26394 26805 26502 26915
rect 27162 26805 27270 26915
rect 27642 26805 27750 26915
rect 28410 26805 28518 26915
rect 28890 26805 28998 26915
rect 29658 26805 29766 26915
rect 30138 26805 30246 26915
rect 30906 26805 31014 26915
rect 31386 26805 31494 26915
rect 32154 26805 32262 26915
rect 32634 26805 32742 26915
rect 33402 26805 33510 26915
rect 33882 26805 33990 26915
rect 34650 26805 34758 26915
rect 35130 26805 35238 26915
rect 35898 26805 36006 26915
rect 36378 26805 36486 26915
rect 37146 26805 37254 26915
rect 37626 26805 37734 26915
rect 38394 26805 38502 26915
rect 38874 26805 38982 26915
rect 39642 26805 39750 26915
rect 0 26709 39936 26757
rect 186 26585 294 26661
rect 954 26585 1062 26661
rect 1434 26585 1542 26661
rect 2202 26585 2310 26661
rect 2682 26585 2790 26661
rect 3450 26585 3558 26661
rect 3930 26585 4038 26661
rect 4698 26585 4806 26661
rect 5178 26585 5286 26661
rect 5946 26585 6054 26661
rect 6426 26585 6534 26661
rect 7194 26585 7302 26661
rect 7674 26585 7782 26661
rect 8442 26585 8550 26661
rect 8922 26585 9030 26661
rect 9690 26585 9798 26661
rect 10170 26585 10278 26661
rect 10938 26585 11046 26661
rect 11418 26585 11526 26661
rect 12186 26585 12294 26661
rect 12666 26585 12774 26661
rect 13434 26585 13542 26661
rect 13914 26585 14022 26661
rect 14682 26585 14790 26661
rect 15162 26585 15270 26661
rect 15930 26585 16038 26661
rect 16410 26585 16518 26661
rect 17178 26585 17286 26661
rect 17658 26585 17766 26661
rect 18426 26585 18534 26661
rect 18906 26585 19014 26661
rect 19674 26585 19782 26661
rect 20154 26585 20262 26661
rect 20922 26585 21030 26661
rect 21402 26585 21510 26661
rect 22170 26585 22278 26661
rect 22650 26585 22758 26661
rect 23418 26585 23526 26661
rect 23898 26585 24006 26661
rect 24666 26585 24774 26661
rect 25146 26585 25254 26661
rect 25914 26585 26022 26661
rect 26394 26585 26502 26661
rect 27162 26585 27270 26661
rect 27642 26585 27750 26661
rect 28410 26585 28518 26661
rect 28890 26585 28998 26661
rect 29658 26585 29766 26661
rect 30138 26585 30246 26661
rect 30906 26585 31014 26661
rect 31386 26585 31494 26661
rect 32154 26585 32262 26661
rect 32634 26585 32742 26661
rect 33402 26585 33510 26661
rect 33882 26585 33990 26661
rect 34650 26585 34758 26661
rect 35130 26585 35238 26661
rect 35898 26585 36006 26661
rect 36378 26585 36486 26661
rect 37146 26585 37254 26661
rect 37626 26585 37734 26661
rect 38394 26585 38502 26661
rect 38874 26585 38982 26661
rect 39642 26585 39750 26661
rect 0 26489 39936 26537
rect 0 26393 39936 26441
rect 186 26269 294 26345
rect 954 26269 1062 26345
rect 1434 26269 1542 26345
rect 2202 26269 2310 26345
rect 2682 26269 2790 26345
rect 3450 26269 3558 26345
rect 3930 26269 4038 26345
rect 4698 26269 4806 26345
rect 5178 26269 5286 26345
rect 5946 26269 6054 26345
rect 6426 26269 6534 26345
rect 7194 26269 7302 26345
rect 7674 26269 7782 26345
rect 8442 26269 8550 26345
rect 8922 26269 9030 26345
rect 9690 26269 9798 26345
rect 10170 26269 10278 26345
rect 10938 26269 11046 26345
rect 11418 26269 11526 26345
rect 12186 26269 12294 26345
rect 12666 26269 12774 26345
rect 13434 26269 13542 26345
rect 13914 26269 14022 26345
rect 14682 26269 14790 26345
rect 15162 26269 15270 26345
rect 15930 26269 16038 26345
rect 16410 26269 16518 26345
rect 17178 26269 17286 26345
rect 17658 26269 17766 26345
rect 18426 26269 18534 26345
rect 18906 26269 19014 26345
rect 19674 26269 19782 26345
rect 20154 26269 20262 26345
rect 20922 26269 21030 26345
rect 21402 26269 21510 26345
rect 22170 26269 22278 26345
rect 22650 26269 22758 26345
rect 23418 26269 23526 26345
rect 23898 26269 24006 26345
rect 24666 26269 24774 26345
rect 25146 26269 25254 26345
rect 25914 26269 26022 26345
rect 26394 26269 26502 26345
rect 27162 26269 27270 26345
rect 27642 26269 27750 26345
rect 28410 26269 28518 26345
rect 28890 26269 28998 26345
rect 29658 26269 29766 26345
rect 30138 26269 30246 26345
rect 30906 26269 31014 26345
rect 31386 26269 31494 26345
rect 32154 26269 32262 26345
rect 32634 26269 32742 26345
rect 33402 26269 33510 26345
rect 33882 26269 33990 26345
rect 34650 26269 34758 26345
rect 35130 26269 35238 26345
rect 35898 26269 36006 26345
rect 36378 26269 36486 26345
rect 37146 26269 37254 26345
rect 37626 26269 37734 26345
rect 38394 26269 38502 26345
rect 38874 26269 38982 26345
rect 39642 26269 39750 26345
rect 0 26173 39936 26221
rect 186 26015 294 26125
rect 954 26015 1062 26125
rect 1434 26015 1542 26125
rect 2202 26015 2310 26125
rect 2682 26015 2790 26125
rect 3450 26015 3558 26125
rect 3930 26015 4038 26125
rect 4698 26015 4806 26125
rect 5178 26015 5286 26125
rect 5946 26015 6054 26125
rect 6426 26015 6534 26125
rect 7194 26015 7302 26125
rect 7674 26015 7782 26125
rect 8442 26015 8550 26125
rect 8922 26015 9030 26125
rect 9690 26015 9798 26125
rect 10170 26015 10278 26125
rect 10938 26015 11046 26125
rect 11418 26015 11526 26125
rect 12186 26015 12294 26125
rect 12666 26015 12774 26125
rect 13434 26015 13542 26125
rect 13914 26015 14022 26125
rect 14682 26015 14790 26125
rect 15162 26015 15270 26125
rect 15930 26015 16038 26125
rect 16410 26015 16518 26125
rect 17178 26015 17286 26125
rect 17658 26015 17766 26125
rect 18426 26015 18534 26125
rect 18906 26015 19014 26125
rect 19674 26015 19782 26125
rect 20154 26015 20262 26125
rect 20922 26015 21030 26125
rect 21402 26015 21510 26125
rect 22170 26015 22278 26125
rect 22650 26015 22758 26125
rect 23418 26015 23526 26125
rect 23898 26015 24006 26125
rect 24666 26015 24774 26125
rect 25146 26015 25254 26125
rect 25914 26015 26022 26125
rect 26394 26015 26502 26125
rect 27162 26015 27270 26125
rect 27642 26015 27750 26125
rect 28410 26015 28518 26125
rect 28890 26015 28998 26125
rect 29658 26015 29766 26125
rect 30138 26015 30246 26125
rect 30906 26015 31014 26125
rect 31386 26015 31494 26125
rect 32154 26015 32262 26125
rect 32634 26015 32742 26125
rect 33402 26015 33510 26125
rect 33882 26015 33990 26125
rect 34650 26015 34758 26125
rect 35130 26015 35238 26125
rect 35898 26015 36006 26125
rect 36378 26015 36486 26125
rect 37146 26015 37254 26125
rect 37626 26015 37734 26125
rect 38394 26015 38502 26125
rect 38874 26015 38982 26125
rect 39642 26015 39750 26125
rect 0 25919 39936 25967
rect 186 25795 294 25871
rect 954 25795 1062 25871
rect 1434 25795 1542 25871
rect 2202 25795 2310 25871
rect 2682 25795 2790 25871
rect 3450 25795 3558 25871
rect 3930 25795 4038 25871
rect 4698 25795 4806 25871
rect 5178 25795 5286 25871
rect 5946 25795 6054 25871
rect 6426 25795 6534 25871
rect 7194 25795 7302 25871
rect 7674 25795 7782 25871
rect 8442 25795 8550 25871
rect 8922 25795 9030 25871
rect 9690 25795 9798 25871
rect 10170 25795 10278 25871
rect 10938 25795 11046 25871
rect 11418 25795 11526 25871
rect 12186 25795 12294 25871
rect 12666 25795 12774 25871
rect 13434 25795 13542 25871
rect 13914 25795 14022 25871
rect 14682 25795 14790 25871
rect 15162 25795 15270 25871
rect 15930 25795 16038 25871
rect 16410 25795 16518 25871
rect 17178 25795 17286 25871
rect 17658 25795 17766 25871
rect 18426 25795 18534 25871
rect 18906 25795 19014 25871
rect 19674 25795 19782 25871
rect 20154 25795 20262 25871
rect 20922 25795 21030 25871
rect 21402 25795 21510 25871
rect 22170 25795 22278 25871
rect 22650 25795 22758 25871
rect 23418 25795 23526 25871
rect 23898 25795 24006 25871
rect 24666 25795 24774 25871
rect 25146 25795 25254 25871
rect 25914 25795 26022 25871
rect 26394 25795 26502 25871
rect 27162 25795 27270 25871
rect 27642 25795 27750 25871
rect 28410 25795 28518 25871
rect 28890 25795 28998 25871
rect 29658 25795 29766 25871
rect 30138 25795 30246 25871
rect 30906 25795 31014 25871
rect 31386 25795 31494 25871
rect 32154 25795 32262 25871
rect 32634 25795 32742 25871
rect 33402 25795 33510 25871
rect 33882 25795 33990 25871
rect 34650 25795 34758 25871
rect 35130 25795 35238 25871
rect 35898 25795 36006 25871
rect 36378 25795 36486 25871
rect 37146 25795 37254 25871
rect 37626 25795 37734 25871
rect 38394 25795 38502 25871
rect 38874 25795 38982 25871
rect 39642 25795 39750 25871
rect 0 25699 39936 25747
rect 0 25603 39936 25651
rect 186 25479 294 25555
rect 954 25479 1062 25555
rect 1434 25479 1542 25555
rect 2202 25479 2310 25555
rect 2682 25479 2790 25555
rect 3450 25479 3558 25555
rect 3930 25479 4038 25555
rect 4698 25479 4806 25555
rect 5178 25479 5286 25555
rect 5946 25479 6054 25555
rect 6426 25479 6534 25555
rect 7194 25479 7302 25555
rect 7674 25479 7782 25555
rect 8442 25479 8550 25555
rect 8922 25479 9030 25555
rect 9690 25479 9798 25555
rect 10170 25479 10278 25555
rect 10938 25479 11046 25555
rect 11418 25479 11526 25555
rect 12186 25479 12294 25555
rect 12666 25479 12774 25555
rect 13434 25479 13542 25555
rect 13914 25479 14022 25555
rect 14682 25479 14790 25555
rect 15162 25479 15270 25555
rect 15930 25479 16038 25555
rect 16410 25479 16518 25555
rect 17178 25479 17286 25555
rect 17658 25479 17766 25555
rect 18426 25479 18534 25555
rect 18906 25479 19014 25555
rect 19674 25479 19782 25555
rect 20154 25479 20262 25555
rect 20922 25479 21030 25555
rect 21402 25479 21510 25555
rect 22170 25479 22278 25555
rect 22650 25479 22758 25555
rect 23418 25479 23526 25555
rect 23898 25479 24006 25555
rect 24666 25479 24774 25555
rect 25146 25479 25254 25555
rect 25914 25479 26022 25555
rect 26394 25479 26502 25555
rect 27162 25479 27270 25555
rect 27642 25479 27750 25555
rect 28410 25479 28518 25555
rect 28890 25479 28998 25555
rect 29658 25479 29766 25555
rect 30138 25479 30246 25555
rect 30906 25479 31014 25555
rect 31386 25479 31494 25555
rect 32154 25479 32262 25555
rect 32634 25479 32742 25555
rect 33402 25479 33510 25555
rect 33882 25479 33990 25555
rect 34650 25479 34758 25555
rect 35130 25479 35238 25555
rect 35898 25479 36006 25555
rect 36378 25479 36486 25555
rect 37146 25479 37254 25555
rect 37626 25479 37734 25555
rect 38394 25479 38502 25555
rect 38874 25479 38982 25555
rect 39642 25479 39750 25555
rect 0 25383 39936 25431
rect 186 25225 294 25335
rect 954 25225 1062 25335
rect 1434 25225 1542 25335
rect 2202 25225 2310 25335
rect 2682 25225 2790 25335
rect 3450 25225 3558 25335
rect 3930 25225 4038 25335
rect 4698 25225 4806 25335
rect 5178 25225 5286 25335
rect 5946 25225 6054 25335
rect 6426 25225 6534 25335
rect 7194 25225 7302 25335
rect 7674 25225 7782 25335
rect 8442 25225 8550 25335
rect 8922 25225 9030 25335
rect 9690 25225 9798 25335
rect 10170 25225 10278 25335
rect 10938 25225 11046 25335
rect 11418 25225 11526 25335
rect 12186 25225 12294 25335
rect 12666 25225 12774 25335
rect 13434 25225 13542 25335
rect 13914 25225 14022 25335
rect 14682 25225 14790 25335
rect 15162 25225 15270 25335
rect 15930 25225 16038 25335
rect 16410 25225 16518 25335
rect 17178 25225 17286 25335
rect 17658 25225 17766 25335
rect 18426 25225 18534 25335
rect 18906 25225 19014 25335
rect 19674 25225 19782 25335
rect 20154 25225 20262 25335
rect 20922 25225 21030 25335
rect 21402 25225 21510 25335
rect 22170 25225 22278 25335
rect 22650 25225 22758 25335
rect 23418 25225 23526 25335
rect 23898 25225 24006 25335
rect 24666 25225 24774 25335
rect 25146 25225 25254 25335
rect 25914 25225 26022 25335
rect 26394 25225 26502 25335
rect 27162 25225 27270 25335
rect 27642 25225 27750 25335
rect 28410 25225 28518 25335
rect 28890 25225 28998 25335
rect 29658 25225 29766 25335
rect 30138 25225 30246 25335
rect 30906 25225 31014 25335
rect 31386 25225 31494 25335
rect 32154 25225 32262 25335
rect 32634 25225 32742 25335
rect 33402 25225 33510 25335
rect 33882 25225 33990 25335
rect 34650 25225 34758 25335
rect 35130 25225 35238 25335
rect 35898 25225 36006 25335
rect 36378 25225 36486 25335
rect 37146 25225 37254 25335
rect 37626 25225 37734 25335
rect 38394 25225 38502 25335
rect 38874 25225 38982 25335
rect 39642 25225 39750 25335
rect 0 25129 39936 25177
rect 186 25005 294 25081
rect 954 25005 1062 25081
rect 1434 25005 1542 25081
rect 2202 25005 2310 25081
rect 2682 25005 2790 25081
rect 3450 25005 3558 25081
rect 3930 25005 4038 25081
rect 4698 25005 4806 25081
rect 5178 25005 5286 25081
rect 5946 25005 6054 25081
rect 6426 25005 6534 25081
rect 7194 25005 7302 25081
rect 7674 25005 7782 25081
rect 8442 25005 8550 25081
rect 8922 25005 9030 25081
rect 9690 25005 9798 25081
rect 10170 25005 10278 25081
rect 10938 25005 11046 25081
rect 11418 25005 11526 25081
rect 12186 25005 12294 25081
rect 12666 25005 12774 25081
rect 13434 25005 13542 25081
rect 13914 25005 14022 25081
rect 14682 25005 14790 25081
rect 15162 25005 15270 25081
rect 15930 25005 16038 25081
rect 16410 25005 16518 25081
rect 17178 25005 17286 25081
rect 17658 25005 17766 25081
rect 18426 25005 18534 25081
rect 18906 25005 19014 25081
rect 19674 25005 19782 25081
rect 20154 25005 20262 25081
rect 20922 25005 21030 25081
rect 21402 25005 21510 25081
rect 22170 25005 22278 25081
rect 22650 25005 22758 25081
rect 23418 25005 23526 25081
rect 23898 25005 24006 25081
rect 24666 25005 24774 25081
rect 25146 25005 25254 25081
rect 25914 25005 26022 25081
rect 26394 25005 26502 25081
rect 27162 25005 27270 25081
rect 27642 25005 27750 25081
rect 28410 25005 28518 25081
rect 28890 25005 28998 25081
rect 29658 25005 29766 25081
rect 30138 25005 30246 25081
rect 30906 25005 31014 25081
rect 31386 25005 31494 25081
rect 32154 25005 32262 25081
rect 32634 25005 32742 25081
rect 33402 25005 33510 25081
rect 33882 25005 33990 25081
rect 34650 25005 34758 25081
rect 35130 25005 35238 25081
rect 35898 25005 36006 25081
rect 36378 25005 36486 25081
rect 37146 25005 37254 25081
rect 37626 25005 37734 25081
rect 38394 25005 38502 25081
rect 38874 25005 38982 25081
rect 39642 25005 39750 25081
rect 0 24909 39936 24957
rect 0 24813 39936 24861
rect 186 24689 294 24765
rect 954 24689 1062 24765
rect 1434 24689 1542 24765
rect 2202 24689 2310 24765
rect 2682 24689 2790 24765
rect 3450 24689 3558 24765
rect 3930 24689 4038 24765
rect 4698 24689 4806 24765
rect 5178 24689 5286 24765
rect 5946 24689 6054 24765
rect 6426 24689 6534 24765
rect 7194 24689 7302 24765
rect 7674 24689 7782 24765
rect 8442 24689 8550 24765
rect 8922 24689 9030 24765
rect 9690 24689 9798 24765
rect 10170 24689 10278 24765
rect 10938 24689 11046 24765
rect 11418 24689 11526 24765
rect 12186 24689 12294 24765
rect 12666 24689 12774 24765
rect 13434 24689 13542 24765
rect 13914 24689 14022 24765
rect 14682 24689 14790 24765
rect 15162 24689 15270 24765
rect 15930 24689 16038 24765
rect 16410 24689 16518 24765
rect 17178 24689 17286 24765
rect 17658 24689 17766 24765
rect 18426 24689 18534 24765
rect 18906 24689 19014 24765
rect 19674 24689 19782 24765
rect 20154 24689 20262 24765
rect 20922 24689 21030 24765
rect 21402 24689 21510 24765
rect 22170 24689 22278 24765
rect 22650 24689 22758 24765
rect 23418 24689 23526 24765
rect 23898 24689 24006 24765
rect 24666 24689 24774 24765
rect 25146 24689 25254 24765
rect 25914 24689 26022 24765
rect 26394 24689 26502 24765
rect 27162 24689 27270 24765
rect 27642 24689 27750 24765
rect 28410 24689 28518 24765
rect 28890 24689 28998 24765
rect 29658 24689 29766 24765
rect 30138 24689 30246 24765
rect 30906 24689 31014 24765
rect 31386 24689 31494 24765
rect 32154 24689 32262 24765
rect 32634 24689 32742 24765
rect 33402 24689 33510 24765
rect 33882 24689 33990 24765
rect 34650 24689 34758 24765
rect 35130 24689 35238 24765
rect 35898 24689 36006 24765
rect 36378 24689 36486 24765
rect 37146 24689 37254 24765
rect 37626 24689 37734 24765
rect 38394 24689 38502 24765
rect 38874 24689 38982 24765
rect 39642 24689 39750 24765
rect 0 24593 39936 24641
rect 186 24435 294 24545
rect 954 24435 1062 24545
rect 1434 24435 1542 24545
rect 2202 24435 2310 24545
rect 2682 24435 2790 24545
rect 3450 24435 3558 24545
rect 3930 24435 4038 24545
rect 4698 24435 4806 24545
rect 5178 24435 5286 24545
rect 5946 24435 6054 24545
rect 6426 24435 6534 24545
rect 7194 24435 7302 24545
rect 7674 24435 7782 24545
rect 8442 24435 8550 24545
rect 8922 24435 9030 24545
rect 9690 24435 9798 24545
rect 10170 24435 10278 24545
rect 10938 24435 11046 24545
rect 11418 24435 11526 24545
rect 12186 24435 12294 24545
rect 12666 24435 12774 24545
rect 13434 24435 13542 24545
rect 13914 24435 14022 24545
rect 14682 24435 14790 24545
rect 15162 24435 15270 24545
rect 15930 24435 16038 24545
rect 16410 24435 16518 24545
rect 17178 24435 17286 24545
rect 17658 24435 17766 24545
rect 18426 24435 18534 24545
rect 18906 24435 19014 24545
rect 19674 24435 19782 24545
rect 20154 24435 20262 24545
rect 20922 24435 21030 24545
rect 21402 24435 21510 24545
rect 22170 24435 22278 24545
rect 22650 24435 22758 24545
rect 23418 24435 23526 24545
rect 23898 24435 24006 24545
rect 24666 24435 24774 24545
rect 25146 24435 25254 24545
rect 25914 24435 26022 24545
rect 26394 24435 26502 24545
rect 27162 24435 27270 24545
rect 27642 24435 27750 24545
rect 28410 24435 28518 24545
rect 28890 24435 28998 24545
rect 29658 24435 29766 24545
rect 30138 24435 30246 24545
rect 30906 24435 31014 24545
rect 31386 24435 31494 24545
rect 32154 24435 32262 24545
rect 32634 24435 32742 24545
rect 33402 24435 33510 24545
rect 33882 24435 33990 24545
rect 34650 24435 34758 24545
rect 35130 24435 35238 24545
rect 35898 24435 36006 24545
rect 36378 24435 36486 24545
rect 37146 24435 37254 24545
rect 37626 24435 37734 24545
rect 38394 24435 38502 24545
rect 38874 24435 38982 24545
rect 39642 24435 39750 24545
rect 0 24339 39936 24387
rect 186 24215 294 24291
rect 954 24215 1062 24291
rect 1434 24215 1542 24291
rect 2202 24215 2310 24291
rect 2682 24215 2790 24291
rect 3450 24215 3558 24291
rect 3930 24215 4038 24291
rect 4698 24215 4806 24291
rect 5178 24215 5286 24291
rect 5946 24215 6054 24291
rect 6426 24215 6534 24291
rect 7194 24215 7302 24291
rect 7674 24215 7782 24291
rect 8442 24215 8550 24291
rect 8922 24215 9030 24291
rect 9690 24215 9798 24291
rect 10170 24215 10278 24291
rect 10938 24215 11046 24291
rect 11418 24215 11526 24291
rect 12186 24215 12294 24291
rect 12666 24215 12774 24291
rect 13434 24215 13542 24291
rect 13914 24215 14022 24291
rect 14682 24215 14790 24291
rect 15162 24215 15270 24291
rect 15930 24215 16038 24291
rect 16410 24215 16518 24291
rect 17178 24215 17286 24291
rect 17658 24215 17766 24291
rect 18426 24215 18534 24291
rect 18906 24215 19014 24291
rect 19674 24215 19782 24291
rect 20154 24215 20262 24291
rect 20922 24215 21030 24291
rect 21402 24215 21510 24291
rect 22170 24215 22278 24291
rect 22650 24215 22758 24291
rect 23418 24215 23526 24291
rect 23898 24215 24006 24291
rect 24666 24215 24774 24291
rect 25146 24215 25254 24291
rect 25914 24215 26022 24291
rect 26394 24215 26502 24291
rect 27162 24215 27270 24291
rect 27642 24215 27750 24291
rect 28410 24215 28518 24291
rect 28890 24215 28998 24291
rect 29658 24215 29766 24291
rect 30138 24215 30246 24291
rect 30906 24215 31014 24291
rect 31386 24215 31494 24291
rect 32154 24215 32262 24291
rect 32634 24215 32742 24291
rect 33402 24215 33510 24291
rect 33882 24215 33990 24291
rect 34650 24215 34758 24291
rect 35130 24215 35238 24291
rect 35898 24215 36006 24291
rect 36378 24215 36486 24291
rect 37146 24215 37254 24291
rect 37626 24215 37734 24291
rect 38394 24215 38502 24291
rect 38874 24215 38982 24291
rect 39642 24215 39750 24291
rect 0 24119 39936 24167
rect 0 24023 39936 24071
rect 186 23899 294 23975
rect 954 23899 1062 23975
rect 1434 23899 1542 23975
rect 2202 23899 2310 23975
rect 2682 23899 2790 23975
rect 3450 23899 3558 23975
rect 3930 23899 4038 23975
rect 4698 23899 4806 23975
rect 5178 23899 5286 23975
rect 5946 23899 6054 23975
rect 6426 23899 6534 23975
rect 7194 23899 7302 23975
rect 7674 23899 7782 23975
rect 8442 23899 8550 23975
rect 8922 23899 9030 23975
rect 9690 23899 9798 23975
rect 10170 23899 10278 23975
rect 10938 23899 11046 23975
rect 11418 23899 11526 23975
rect 12186 23899 12294 23975
rect 12666 23899 12774 23975
rect 13434 23899 13542 23975
rect 13914 23899 14022 23975
rect 14682 23899 14790 23975
rect 15162 23899 15270 23975
rect 15930 23899 16038 23975
rect 16410 23899 16518 23975
rect 17178 23899 17286 23975
rect 17658 23899 17766 23975
rect 18426 23899 18534 23975
rect 18906 23899 19014 23975
rect 19674 23899 19782 23975
rect 20154 23899 20262 23975
rect 20922 23899 21030 23975
rect 21402 23899 21510 23975
rect 22170 23899 22278 23975
rect 22650 23899 22758 23975
rect 23418 23899 23526 23975
rect 23898 23899 24006 23975
rect 24666 23899 24774 23975
rect 25146 23899 25254 23975
rect 25914 23899 26022 23975
rect 26394 23899 26502 23975
rect 27162 23899 27270 23975
rect 27642 23899 27750 23975
rect 28410 23899 28518 23975
rect 28890 23899 28998 23975
rect 29658 23899 29766 23975
rect 30138 23899 30246 23975
rect 30906 23899 31014 23975
rect 31386 23899 31494 23975
rect 32154 23899 32262 23975
rect 32634 23899 32742 23975
rect 33402 23899 33510 23975
rect 33882 23899 33990 23975
rect 34650 23899 34758 23975
rect 35130 23899 35238 23975
rect 35898 23899 36006 23975
rect 36378 23899 36486 23975
rect 37146 23899 37254 23975
rect 37626 23899 37734 23975
rect 38394 23899 38502 23975
rect 38874 23899 38982 23975
rect 39642 23899 39750 23975
rect 0 23803 39936 23851
rect 186 23645 294 23755
rect 954 23645 1062 23755
rect 1434 23645 1542 23755
rect 2202 23645 2310 23755
rect 2682 23645 2790 23755
rect 3450 23645 3558 23755
rect 3930 23645 4038 23755
rect 4698 23645 4806 23755
rect 5178 23645 5286 23755
rect 5946 23645 6054 23755
rect 6426 23645 6534 23755
rect 7194 23645 7302 23755
rect 7674 23645 7782 23755
rect 8442 23645 8550 23755
rect 8922 23645 9030 23755
rect 9690 23645 9798 23755
rect 10170 23645 10278 23755
rect 10938 23645 11046 23755
rect 11418 23645 11526 23755
rect 12186 23645 12294 23755
rect 12666 23645 12774 23755
rect 13434 23645 13542 23755
rect 13914 23645 14022 23755
rect 14682 23645 14790 23755
rect 15162 23645 15270 23755
rect 15930 23645 16038 23755
rect 16410 23645 16518 23755
rect 17178 23645 17286 23755
rect 17658 23645 17766 23755
rect 18426 23645 18534 23755
rect 18906 23645 19014 23755
rect 19674 23645 19782 23755
rect 20154 23645 20262 23755
rect 20922 23645 21030 23755
rect 21402 23645 21510 23755
rect 22170 23645 22278 23755
rect 22650 23645 22758 23755
rect 23418 23645 23526 23755
rect 23898 23645 24006 23755
rect 24666 23645 24774 23755
rect 25146 23645 25254 23755
rect 25914 23645 26022 23755
rect 26394 23645 26502 23755
rect 27162 23645 27270 23755
rect 27642 23645 27750 23755
rect 28410 23645 28518 23755
rect 28890 23645 28998 23755
rect 29658 23645 29766 23755
rect 30138 23645 30246 23755
rect 30906 23645 31014 23755
rect 31386 23645 31494 23755
rect 32154 23645 32262 23755
rect 32634 23645 32742 23755
rect 33402 23645 33510 23755
rect 33882 23645 33990 23755
rect 34650 23645 34758 23755
rect 35130 23645 35238 23755
rect 35898 23645 36006 23755
rect 36378 23645 36486 23755
rect 37146 23645 37254 23755
rect 37626 23645 37734 23755
rect 38394 23645 38502 23755
rect 38874 23645 38982 23755
rect 39642 23645 39750 23755
rect 0 23549 39936 23597
rect 186 23425 294 23501
rect 954 23425 1062 23501
rect 1434 23425 1542 23501
rect 2202 23425 2310 23501
rect 2682 23425 2790 23501
rect 3450 23425 3558 23501
rect 3930 23425 4038 23501
rect 4698 23425 4806 23501
rect 5178 23425 5286 23501
rect 5946 23425 6054 23501
rect 6426 23425 6534 23501
rect 7194 23425 7302 23501
rect 7674 23425 7782 23501
rect 8442 23425 8550 23501
rect 8922 23425 9030 23501
rect 9690 23425 9798 23501
rect 10170 23425 10278 23501
rect 10938 23425 11046 23501
rect 11418 23425 11526 23501
rect 12186 23425 12294 23501
rect 12666 23425 12774 23501
rect 13434 23425 13542 23501
rect 13914 23425 14022 23501
rect 14682 23425 14790 23501
rect 15162 23425 15270 23501
rect 15930 23425 16038 23501
rect 16410 23425 16518 23501
rect 17178 23425 17286 23501
rect 17658 23425 17766 23501
rect 18426 23425 18534 23501
rect 18906 23425 19014 23501
rect 19674 23425 19782 23501
rect 20154 23425 20262 23501
rect 20922 23425 21030 23501
rect 21402 23425 21510 23501
rect 22170 23425 22278 23501
rect 22650 23425 22758 23501
rect 23418 23425 23526 23501
rect 23898 23425 24006 23501
rect 24666 23425 24774 23501
rect 25146 23425 25254 23501
rect 25914 23425 26022 23501
rect 26394 23425 26502 23501
rect 27162 23425 27270 23501
rect 27642 23425 27750 23501
rect 28410 23425 28518 23501
rect 28890 23425 28998 23501
rect 29658 23425 29766 23501
rect 30138 23425 30246 23501
rect 30906 23425 31014 23501
rect 31386 23425 31494 23501
rect 32154 23425 32262 23501
rect 32634 23425 32742 23501
rect 33402 23425 33510 23501
rect 33882 23425 33990 23501
rect 34650 23425 34758 23501
rect 35130 23425 35238 23501
rect 35898 23425 36006 23501
rect 36378 23425 36486 23501
rect 37146 23425 37254 23501
rect 37626 23425 37734 23501
rect 38394 23425 38502 23501
rect 38874 23425 38982 23501
rect 39642 23425 39750 23501
rect 0 23329 39936 23377
rect 0 23233 39936 23281
rect 186 23109 294 23185
rect 954 23109 1062 23185
rect 1434 23109 1542 23185
rect 2202 23109 2310 23185
rect 2682 23109 2790 23185
rect 3450 23109 3558 23185
rect 3930 23109 4038 23185
rect 4698 23109 4806 23185
rect 5178 23109 5286 23185
rect 5946 23109 6054 23185
rect 6426 23109 6534 23185
rect 7194 23109 7302 23185
rect 7674 23109 7782 23185
rect 8442 23109 8550 23185
rect 8922 23109 9030 23185
rect 9690 23109 9798 23185
rect 10170 23109 10278 23185
rect 10938 23109 11046 23185
rect 11418 23109 11526 23185
rect 12186 23109 12294 23185
rect 12666 23109 12774 23185
rect 13434 23109 13542 23185
rect 13914 23109 14022 23185
rect 14682 23109 14790 23185
rect 15162 23109 15270 23185
rect 15930 23109 16038 23185
rect 16410 23109 16518 23185
rect 17178 23109 17286 23185
rect 17658 23109 17766 23185
rect 18426 23109 18534 23185
rect 18906 23109 19014 23185
rect 19674 23109 19782 23185
rect 20154 23109 20262 23185
rect 20922 23109 21030 23185
rect 21402 23109 21510 23185
rect 22170 23109 22278 23185
rect 22650 23109 22758 23185
rect 23418 23109 23526 23185
rect 23898 23109 24006 23185
rect 24666 23109 24774 23185
rect 25146 23109 25254 23185
rect 25914 23109 26022 23185
rect 26394 23109 26502 23185
rect 27162 23109 27270 23185
rect 27642 23109 27750 23185
rect 28410 23109 28518 23185
rect 28890 23109 28998 23185
rect 29658 23109 29766 23185
rect 30138 23109 30246 23185
rect 30906 23109 31014 23185
rect 31386 23109 31494 23185
rect 32154 23109 32262 23185
rect 32634 23109 32742 23185
rect 33402 23109 33510 23185
rect 33882 23109 33990 23185
rect 34650 23109 34758 23185
rect 35130 23109 35238 23185
rect 35898 23109 36006 23185
rect 36378 23109 36486 23185
rect 37146 23109 37254 23185
rect 37626 23109 37734 23185
rect 38394 23109 38502 23185
rect 38874 23109 38982 23185
rect 39642 23109 39750 23185
rect 0 23013 39936 23061
rect 186 22855 294 22965
rect 954 22855 1062 22965
rect 1434 22855 1542 22965
rect 2202 22855 2310 22965
rect 2682 22855 2790 22965
rect 3450 22855 3558 22965
rect 3930 22855 4038 22965
rect 4698 22855 4806 22965
rect 5178 22855 5286 22965
rect 5946 22855 6054 22965
rect 6426 22855 6534 22965
rect 7194 22855 7302 22965
rect 7674 22855 7782 22965
rect 8442 22855 8550 22965
rect 8922 22855 9030 22965
rect 9690 22855 9798 22965
rect 10170 22855 10278 22965
rect 10938 22855 11046 22965
rect 11418 22855 11526 22965
rect 12186 22855 12294 22965
rect 12666 22855 12774 22965
rect 13434 22855 13542 22965
rect 13914 22855 14022 22965
rect 14682 22855 14790 22965
rect 15162 22855 15270 22965
rect 15930 22855 16038 22965
rect 16410 22855 16518 22965
rect 17178 22855 17286 22965
rect 17658 22855 17766 22965
rect 18426 22855 18534 22965
rect 18906 22855 19014 22965
rect 19674 22855 19782 22965
rect 20154 22855 20262 22965
rect 20922 22855 21030 22965
rect 21402 22855 21510 22965
rect 22170 22855 22278 22965
rect 22650 22855 22758 22965
rect 23418 22855 23526 22965
rect 23898 22855 24006 22965
rect 24666 22855 24774 22965
rect 25146 22855 25254 22965
rect 25914 22855 26022 22965
rect 26394 22855 26502 22965
rect 27162 22855 27270 22965
rect 27642 22855 27750 22965
rect 28410 22855 28518 22965
rect 28890 22855 28998 22965
rect 29658 22855 29766 22965
rect 30138 22855 30246 22965
rect 30906 22855 31014 22965
rect 31386 22855 31494 22965
rect 32154 22855 32262 22965
rect 32634 22855 32742 22965
rect 33402 22855 33510 22965
rect 33882 22855 33990 22965
rect 34650 22855 34758 22965
rect 35130 22855 35238 22965
rect 35898 22855 36006 22965
rect 36378 22855 36486 22965
rect 37146 22855 37254 22965
rect 37626 22855 37734 22965
rect 38394 22855 38502 22965
rect 38874 22855 38982 22965
rect 39642 22855 39750 22965
rect 0 22759 39936 22807
rect 186 22635 294 22711
rect 954 22635 1062 22711
rect 1434 22635 1542 22711
rect 2202 22635 2310 22711
rect 2682 22635 2790 22711
rect 3450 22635 3558 22711
rect 3930 22635 4038 22711
rect 4698 22635 4806 22711
rect 5178 22635 5286 22711
rect 5946 22635 6054 22711
rect 6426 22635 6534 22711
rect 7194 22635 7302 22711
rect 7674 22635 7782 22711
rect 8442 22635 8550 22711
rect 8922 22635 9030 22711
rect 9690 22635 9798 22711
rect 10170 22635 10278 22711
rect 10938 22635 11046 22711
rect 11418 22635 11526 22711
rect 12186 22635 12294 22711
rect 12666 22635 12774 22711
rect 13434 22635 13542 22711
rect 13914 22635 14022 22711
rect 14682 22635 14790 22711
rect 15162 22635 15270 22711
rect 15930 22635 16038 22711
rect 16410 22635 16518 22711
rect 17178 22635 17286 22711
rect 17658 22635 17766 22711
rect 18426 22635 18534 22711
rect 18906 22635 19014 22711
rect 19674 22635 19782 22711
rect 20154 22635 20262 22711
rect 20922 22635 21030 22711
rect 21402 22635 21510 22711
rect 22170 22635 22278 22711
rect 22650 22635 22758 22711
rect 23418 22635 23526 22711
rect 23898 22635 24006 22711
rect 24666 22635 24774 22711
rect 25146 22635 25254 22711
rect 25914 22635 26022 22711
rect 26394 22635 26502 22711
rect 27162 22635 27270 22711
rect 27642 22635 27750 22711
rect 28410 22635 28518 22711
rect 28890 22635 28998 22711
rect 29658 22635 29766 22711
rect 30138 22635 30246 22711
rect 30906 22635 31014 22711
rect 31386 22635 31494 22711
rect 32154 22635 32262 22711
rect 32634 22635 32742 22711
rect 33402 22635 33510 22711
rect 33882 22635 33990 22711
rect 34650 22635 34758 22711
rect 35130 22635 35238 22711
rect 35898 22635 36006 22711
rect 36378 22635 36486 22711
rect 37146 22635 37254 22711
rect 37626 22635 37734 22711
rect 38394 22635 38502 22711
rect 38874 22635 38982 22711
rect 39642 22635 39750 22711
rect 0 22539 39936 22587
rect 0 22443 39936 22491
rect 186 22319 294 22395
rect 954 22319 1062 22395
rect 1434 22319 1542 22395
rect 2202 22319 2310 22395
rect 2682 22319 2790 22395
rect 3450 22319 3558 22395
rect 3930 22319 4038 22395
rect 4698 22319 4806 22395
rect 5178 22319 5286 22395
rect 5946 22319 6054 22395
rect 6426 22319 6534 22395
rect 7194 22319 7302 22395
rect 7674 22319 7782 22395
rect 8442 22319 8550 22395
rect 8922 22319 9030 22395
rect 9690 22319 9798 22395
rect 10170 22319 10278 22395
rect 10938 22319 11046 22395
rect 11418 22319 11526 22395
rect 12186 22319 12294 22395
rect 12666 22319 12774 22395
rect 13434 22319 13542 22395
rect 13914 22319 14022 22395
rect 14682 22319 14790 22395
rect 15162 22319 15270 22395
rect 15930 22319 16038 22395
rect 16410 22319 16518 22395
rect 17178 22319 17286 22395
rect 17658 22319 17766 22395
rect 18426 22319 18534 22395
rect 18906 22319 19014 22395
rect 19674 22319 19782 22395
rect 20154 22319 20262 22395
rect 20922 22319 21030 22395
rect 21402 22319 21510 22395
rect 22170 22319 22278 22395
rect 22650 22319 22758 22395
rect 23418 22319 23526 22395
rect 23898 22319 24006 22395
rect 24666 22319 24774 22395
rect 25146 22319 25254 22395
rect 25914 22319 26022 22395
rect 26394 22319 26502 22395
rect 27162 22319 27270 22395
rect 27642 22319 27750 22395
rect 28410 22319 28518 22395
rect 28890 22319 28998 22395
rect 29658 22319 29766 22395
rect 30138 22319 30246 22395
rect 30906 22319 31014 22395
rect 31386 22319 31494 22395
rect 32154 22319 32262 22395
rect 32634 22319 32742 22395
rect 33402 22319 33510 22395
rect 33882 22319 33990 22395
rect 34650 22319 34758 22395
rect 35130 22319 35238 22395
rect 35898 22319 36006 22395
rect 36378 22319 36486 22395
rect 37146 22319 37254 22395
rect 37626 22319 37734 22395
rect 38394 22319 38502 22395
rect 38874 22319 38982 22395
rect 39642 22319 39750 22395
rect 0 22223 39936 22271
rect 186 22065 294 22175
rect 954 22065 1062 22175
rect 1434 22065 1542 22175
rect 2202 22065 2310 22175
rect 2682 22065 2790 22175
rect 3450 22065 3558 22175
rect 3930 22065 4038 22175
rect 4698 22065 4806 22175
rect 5178 22065 5286 22175
rect 5946 22065 6054 22175
rect 6426 22065 6534 22175
rect 7194 22065 7302 22175
rect 7674 22065 7782 22175
rect 8442 22065 8550 22175
rect 8922 22065 9030 22175
rect 9690 22065 9798 22175
rect 10170 22065 10278 22175
rect 10938 22065 11046 22175
rect 11418 22065 11526 22175
rect 12186 22065 12294 22175
rect 12666 22065 12774 22175
rect 13434 22065 13542 22175
rect 13914 22065 14022 22175
rect 14682 22065 14790 22175
rect 15162 22065 15270 22175
rect 15930 22065 16038 22175
rect 16410 22065 16518 22175
rect 17178 22065 17286 22175
rect 17658 22065 17766 22175
rect 18426 22065 18534 22175
rect 18906 22065 19014 22175
rect 19674 22065 19782 22175
rect 20154 22065 20262 22175
rect 20922 22065 21030 22175
rect 21402 22065 21510 22175
rect 22170 22065 22278 22175
rect 22650 22065 22758 22175
rect 23418 22065 23526 22175
rect 23898 22065 24006 22175
rect 24666 22065 24774 22175
rect 25146 22065 25254 22175
rect 25914 22065 26022 22175
rect 26394 22065 26502 22175
rect 27162 22065 27270 22175
rect 27642 22065 27750 22175
rect 28410 22065 28518 22175
rect 28890 22065 28998 22175
rect 29658 22065 29766 22175
rect 30138 22065 30246 22175
rect 30906 22065 31014 22175
rect 31386 22065 31494 22175
rect 32154 22065 32262 22175
rect 32634 22065 32742 22175
rect 33402 22065 33510 22175
rect 33882 22065 33990 22175
rect 34650 22065 34758 22175
rect 35130 22065 35238 22175
rect 35898 22065 36006 22175
rect 36378 22065 36486 22175
rect 37146 22065 37254 22175
rect 37626 22065 37734 22175
rect 38394 22065 38502 22175
rect 38874 22065 38982 22175
rect 39642 22065 39750 22175
rect 0 21969 39936 22017
rect 186 21845 294 21921
rect 954 21845 1062 21921
rect 1434 21845 1542 21921
rect 2202 21845 2310 21921
rect 2682 21845 2790 21921
rect 3450 21845 3558 21921
rect 3930 21845 4038 21921
rect 4698 21845 4806 21921
rect 5178 21845 5286 21921
rect 5946 21845 6054 21921
rect 6426 21845 6534 21921
rect 7194 21845 7302 21921
rect 7674 21845 7782 21921
rect 8442 21845 8550 21921
rect 8922 21845 9030 21921
rect 9690 21845 9798 21921
rect 10170 21845 10278 21921
rect 10938 21845 11046 21921
rect 11418 21845 11526 21921
rect 12186 21845 12294 21921
rect 12666 21845 12774 21921
rect 13434 21845 13542 21921
rect 13914 21845 14022 21921
rect 14682 21845 14790 21921
rect 15162 21845 15270 21921
rect 15930 21845 16038 21921
rect 16410 21845 16518 21921
rect 17178 21845 17286 21921
rect 17658 21845 17766 21921
rect 18426 21845 18534 21921
rect 18906 21845 19014 21921
rect 19674 21845 19782 21921
rect 20154 21845 20262 21921
rect 20922 21845 21030 21921
rect 21402 21845 21510 21921
rect 22170 21845 22278 21921
rect 22650 21845 22758 21921
rect 23418 21845 23526 21921
rect 23898 21845 24006 21921
rect 24666 21845 24774 21921
rect 25146 21845 25254 21921
rect 25914 21845 26022 21921
rect 26394 21845 26502 21921
rect 27162 21845 27270 21921
rect 27642 21845 27750 21921
rect 28410 21845 28518 21921
rect 28890 21845 28998 21921
rect 29658 21845 29766 21921
rect 30138 21845 30246 21921
rect 30906 21845 31014 21921
rect 31386 21845 31494 21921
rect 32154 21845 32262 21921
rect 32634 21845 32742 21921
rect 33402 21845 33510 21921
rect 33882 21845 33990 21921
rect 34650 21845 34758 21921
rect 35130 21845 35238 21921
rect 35898 21845 36006 21921
rect 36378 21845 36486 21921
rect 37146 21845 37254 21921
rect 37626 21845 37734 21921
rect 38394 21845 38502 21921
rect 38874 21845 38982 21921
rect 39642 21845 39750 21921
rect 0 21749 39936 21797
rect 0 21653 39936 21701
rect 186 21529 294 21605
rect 954 21529 1062 21605
rect 1434 21529 1542 21605
rect 2202 21529 2310 21605
rect 2682 21529 2790 21605
rect 3450 21529 3558 21605
rect 3930 21529 4038 21605
rect 4698 21529 4806 21605
rect 5178 21529 5286 21605
rect 5946 21529 6054 21605
rect 6426 21529 6534 21605
rect 7194 21529 7302 21605
rect 7674 21529 7782 21605
rect 8442 21529 8550 21605
rect 8922 21529 9030 21605
rect 9690 21529 9798 21605
rect 10170 21529 10278 21605
rect 10938 21529 11046 21605
rect 11418 21529 11526 21605
rect 12186 21529 12294 21605
rect 12666 21529 12774 21605
rect 13434 21529 13542 21605
rect 13914 21529 14022 21605
rect 14682 21529 14790 21605
rect 15162 21529 15270 21605
rect 15930 21529 16038 21605
rect 16410 21529 16518 21605
rect 17178 21529 17286 21605
rect 17658 21529 17766 21605
rect 18426 21529 18534 21605
rect 18906 21529 19014 21605
rect 19674 21529 19782 21605
rect 20154 21529 20262 21605
rect 20922 21529 21030 21605
rect 21402 21529 21510 21605
rect 22170 21529 22278 21605
rect 22650 21529 22758 21605
rect 23418 21529 23526 21605
rect 23898 21529 24006 21605
rect 24666 21529 24774 21605
rect 25146 21529 25254 21605
rect 25914 21529 26022 21605
rect 26394 21529 26502 21605
rect 27162 21529 27270 21605
rect 27642 21529 27750 21605
rect 28410 21529 28518 21605
rect 28890 21529 28998 21605
rect 29658 21529 29766 21605
rect 30138 21529 30246 21605
rect 30906 21529 31014 21605
rect 31386 21529 31494 21605
rect 32154 21529 32262 21605
rect 32634 21529 32742 21605
rect 33402 21529 33510 21605
rect 33882 21529 33990 21605
rect 34650 21529 34758 21605
rect 35130 21529 35238 21605
rect 35898 21529 36006 21605
rect 36378 21529 36486 21605
rect 37146 21529 37254 21605
rect 37626 21529 37734 21605
rect 38394 21529 38502 21605
rect 38874 21529 38982 21605
rect 39642 21529 39750 21605
rect 0 21433 39936 21481
rect 186 21275 294 21385
rect 954 21275 1062 21385
rect 1434 21275 1542 21385
rect 2202 21275 2310 21385
rect 2682 21275 2790 21385
rect 3450 21275 3558 21385
rect 3930 21275 4038 21385
rect 4698 21275 4806 21385
rect 5178 21275 5286 21385
rect 5946 21275 6054 21385
rect 6426 21275 6534 21385
rect 7194 21275 7302 21385
rect 7674 21275 7782 21385
rect 8442 21275 8550 21385
rect 8922 21275 9030 21385
rect 9690 21275 9798 21385
rect 10170 21275 10278 21385
rect 10938 21275 11046 21385
rect 11418 21275 11526 21385
rect 12186 21275 12294 21385
rect 12666 21275 12774 21385
rect 13434 21275 13542 21385
rect 13914 21275 14022 21385
rect 14682 21275 14790 21385
rect 15162 21275 15270 21385
rect 15930 21275 16038 21385
rect 16410 21275 16518 21385
rect 17178 21275 17286 21385
rect 17658 21275 17766 21385
rect 18426 21275 18534 21385
rect 18906 21275 19014 21385
rect 19674 21275 19782 21385
rect 20154 21275 20262 21385
rect 20922 21275 21030 21385
rect 21402 21275 21510 21385
rect 22170 21275 22278 21385
rect 22650 21275 22758 21385
rect 23418 21275 23526 21385
rect 23898 21275 24006 21385
rect 24666 21275 24774 21385
rect 25146 21275 25254 21385
rect 25914 21275 26022 21385
rect 26394 21275 26502 21385
rect 27162 21275 27270 21385
rect 27642 21275 27750 21385
rect 28410 21275 28518 21385
rect 28890 21275 28998 21385
rect 29658 21275 29766 21385
rect 30138 21275 30246 21385
rect 30906 21275 31014 21385
rect 31386 21275 31494 21385
rect 32154 21275 32262 21385
rect 32634 21275 32742 21385
rect 33402 21275 33510 21385
rect 33882 21275 33990 21385
rect 34650 21275 34758 21385
rect 35130 21275 35238 21385
rect 35898 21275 36006 21385
rect 36378 21275 36486 21385
rect 37146 21275 37254 21385
rect 37626 21275 37734 21385
rect 38394 21275 38502 21385
rect 38874 21275 38982 21385
rect 39642 21275 39750 21385
rect 0 21179 39936 21227
rect 186 21055 294 21131
rect 954 21055 1062 21131
rect 1434 21055 1542 21131
rect 2202 21055 2310 21131
rect 2682 21055 2790 21131
rect 3450 21055 3558 21131
rect 3930 21055 4038 21131
rect 4698 21055 4806 21131
rect 5178 21055 5286 21131
rect 5946 21055 6054 21131
rect 6426 21055 6534 21131
rect 7194 21055 7302 21131
rect 7674 21055 7782 21131
rect 8442 21055 8550 21131
rect 8922 21055 9030 21131
rect 9690 21055 9798 21131
rect 10170 21055 10278 21131
rect 10938 21055 11046 21131
rect 11418 21055 11526 21131
rect 12186 21055 12294 21131
rect 12666 21055 12774 21131
rect 13434 21055 13542 21131
rect 13914 21055 14022 21131
rect 14682 21055 14790 21131
rect 15162 21055 15270 21131
rect 15930 21055 16038 21131
rect 16410 21055 16518 21131
rect 17178 21055 17286 21131
rect 17658 21055 17766 21131
rect 18426 21055 18534 21131
rect 18906 21055 19014 21131
rect 19674 21055 19782 21131
rect 20154 21055 20262 21131
rect 20922 21055 21030 21131
rect 21402 21055 21510 21131
rect 22170 21055 22278 21131
rect 22650 21055 22758 21131
rect 23418 21055 23526 21131
rect 23898 21055 24006 21131
rect 24666 21055 24774 21131
rect 25146 21055 25254 21131
rect 25914 21055 26022 21131
rect 26394 21055 26502 21131
rect 27162 21055 27270 21131
rect 27642 21055 27750 21131
rect 28410 21055 28518 21131
rect 28890 21055 28998 21131
rect 29658 21055 29766 21131
rect 30138 21055 30246 21131
rect 30906 21055 31014 21131
rect 31386 21055 31494 21131
rect 32154 21055 32262 21131
rect 32634 21055 32742 21131
rect 33402 21055 33510 21131
rect 33882 21055 33990 21131
rect 34650 21055 34758 21131
rect 35130 21055 35238 21131
rect 35898 21055 36006 21131
rect 36378 21055 36486 21131
rect 37146 21055 37254 21131
rect 37626 21055 37734 21131
rect 38394 21055 38502 21131
rect 38874 21055 38982 21131
rect 39642 21055 39750 21131
rect 0 20959 39936 21007
rect 0 20863 39936 20911
rect 186 20739 294 20815
rect 954 20739 1062 20815
rect 1434 20739 1542 20815
rect 2202 20739 2310 20815
rect 2682 20739 2790 20815
rect 3450 20739 3558 20815
rect 3930 20739 4038 20815
rect 4698 20739 4806 20815
rect 5178 20739 5286 20815
rect 5946 20739 6054 20815
rect 6426 20739 6534 20815
rect 7194 20739 7302 20815
rect 7674 20739 7782 20815
rect 8442 20739 8550 20815
rect 8922 20739 9030 20815
rect 9690 20739 9798 20815
rect 10170 20739 10278 20815
rect 10938 20739 11046 20815
rect 11418 20739 11526 20815
rect 12186 20739 12294 20815
rect 12666 20739 12774 20815
rect 13434 20739 13542 20815
rect 13914 20739 14022 20815
rect 14682 20739 14790 20815
rect 15162 20739 15270 20815
rect 15930 20739 16038 20815
rect 16410 20739 16518 20815
rect 17178 20739 17286 20815
rect 17658 20739 17766 20815
rect 18426 20739 18534 20815
rect 18906 20739 19014 20815
rect 19674 20739 19782 20815
rect 20154 20739 20262 20815
rect 20922 20739 21030 20815
rect 21402 20739 21510 20815
rect 22170 20739 22278 20815
rect 22650 20739 22758 20815
rect 23418 20739 23526 20815
rect 23898 20739 24006 20815
rect 24666 20739 24774 20815
rect 25146 20739 25254 20815
rect 25914 20739 26022 20815
rect 26394 20739 26502 20815
rect 27162 20739 27270 20815
rect 27642 20739 27750 20815
rect 28410 20739 28518 20815
rect 28890 20739 28998 20815
rect 29658 20739 29766 20815
rect 30138 20739 30246 20815
rect 30906 20739 31014 20815
rect 31386 20739 31494 20815
rect 32154 20739 32262 20815
rect 32634 20739 32742 20815
rect 33402 20739 33510 20815
rect 33882 20739 33990 20815
rect 34650 20739 34758 20815
rect 35130 20739 35238 20815
rect 35898 20739 36006 20815
rect 36378 20739 36486 20815
rect 37146 20739 37254 20815
rect 37626 20739 37734 20815
rect 38394 20739 38502 20815
rect 38874 20739 38982 20815
rect 39642 20739 39750 20815
rect 0 20643 39936 20691
rect 186 20485 294 20595
rect 954 20485 1062 20595
rect 1434 20485 1542 20595
rect 2202 20485 2310 20595
rect 2682 20485 2790 20595
rect 3450 20485 3558 20595
rect 3930 20485 4038 20595
rect 4698 20485 4806 20595
rect 5178 20485 5286 20595
rect 5946 20485 6054 20595
rect 6426 20485 6534 20595
rect 7194 20485 7302 20595
rect 7674 20485 7782 20595
rect 8442 20485 8550 20595
rect 8922 20485 9030 20595
rect 9690 20485 9798 20595
rect 10170 20485 10278 20595
rect 10938 20485 11046 20595
rect 11418 20485 11526 20595
rect 12186 20485 12294 20595
rect 12666 20485 12774 20595
rect 13434 20485 13542 20595
rect 13914 20485 14022 20595
rect 14682 20485 14790 20595
rect 15162 20485 15270 20595
rect 15930 20485 16038 20595
rect 16410 20485 16518 20595
rect 17178 20485 17286 20595
rect 17658 20485 17766 20595
rect 18426 20485 18534 20595
rect 18906 20485 19014 20595
rect 19674 20485 19782 20595
rect 20154 20485 20262 20595
rect 20922 20485 21030 20595
rect 21402 20485 21510 20595
rect 22170 20485 22278 20595
rect 22650 20485 22758 20595
rect 23418 20485 23526 20595
rect 23898 20485 24006 20595
rect 24666 20485 24774 20595
rect 25146 20485 25254 20595
rect 25914 20485 26022 20595
rect 26394 20485 26502 20595
rect 27162 20485 27270 20595
rect 27642 20485 27750 20595
rect 28410 20485 28518 20595
rect 28890 20485 28998 20595
rect 29658 20485 29766 20595
rect 30138 20485 30246 20595
rect 30906 20485 31014 20595
rect 31386 20485 31494 20595
rect 32154 20485 32262 20595
rect 32634 20485 32742 20595
rect 33402 20485 33510 20595
rect 33882 20485 33990 20595
rect 34650 20485 34758 20595
rect 35130 20485 35238 20595
rect 35898 20485 36006 20595
rect 36378 20485 36486 20595
rect 37146 20485 37254 20595
rect 37626 20485 37734 20595
rect 38394 20485 38502 20595
rect 38874 20485 38982 20595
rect 39642 20485 39750 20595
rect 0 20389 39936 20437
rect 186 20265 294 20341
rect 954 20265 1062 20341
rect 1434 20265 1542 20341
rect 2202 20265 2310 20341
rect 2682 20265 2790 20341
rect 3450 20265 3558 20341
rect 3930 20265 4038 20341
rect 4698 20265 4806 20341
rect 5178 20265 5286 20341
rect 5946 20265 6054 20341
rect 6426 20265 6534 20341
rect 7194 20265 7302 20341
rect 7674 20265 7782 20341
rect 8442 20265 8550 20341
rect 8922 20265 9030 20341
rect 9690 20265 9798 20341
rect 10170 20265 10278 20341
rect 10938 20265 11046 20341
rect 11418 20265 11526 20341
rect 12186 20265 12294 20341
rect 12666 20265 12774 20341
rect 13434 20265 13542 20341
rect 13914 20265 14022 20341
rect 14682 20265 14790 20341
rect 15162 20265 15270 20341
rect 15930 20265 16038 20341
rect 16410 20265 16518 20341
rect 17178 20265 17286 20341
rect 17658 20265 17766 20341
rect 18426 20265 18534 20341
rect 18906 20265 19014 20341
rect 19674 20265 19782 20341
rect 20154 20265 20262 20341
rect 20922 20265 21030 20341
rect 21402 20265 21510 20341
rect 22170 20265 22278 20341
rect 22650 20265 22758 20341
rect 23418 20265 23526 20341
rect 23898 20265 24006 20341
rect 24666 20265 24774 20341
rect 25146 20265 25254 20341
rect 25914 20265 26022 20341
rect 26394 20265 26502 20341
rect 27162 20265 27270 20341
rect 27642 20265 27750 20341
rect 28410 20265 28518 20341
rect 28890 20265 28998 20341
rect 29658 20265 29766 20341
rect 30138 20265 30246 20341
rect 30906 20265 31014 20341
rect 31386 20265 31494 20341
rect 32154 20265 32262 20341
rect 32634 20265 32742 20341
rect 33402 20265 33510 20341
rect 33882 20265 33990 20341
rect 34650 20265 34758 20341
rect 35130 20265 35238 20341
rect 35898 20265 36006 20341
rect 36378 20265 36486 20341
rect 37146 20265 37254 20341
rect 37626 20265 37734 20341
rect 38394 20265 38502 20341
rect 38874 20265 38982 20341
rect 39642 20265 39750 20341
rect 0 20169 39936 20217
rect 0 20073 39936 20121
rect 186 19949 294 20025
rect 954 19949 1062 20025
rect 1434 19949 1542 20025
rect 2202 19949 2310 20025
rect 2682 19949 2790 20025
rect 3450 19949 3558 20025
rect 3930 19949 4038 20025
rect 4698 19949 4806 20025
rect 5178 19949 5286 20025
rect 5946 19949 6054 20025
rect 6426 19949 6534 20025
rect 7194 19949 7302 20025
rect 7674 19949 7782 20025
rect 8442 19949 8550 20025
rect 8922 19949 9030 20025
rect 9690 19949 9798 20025
rect 10170 19949 10278 20025
rect 10938 19949 11046 20025
rect 11418 19949 11526 20025
rect 12186 19949 12294 20025
rect 12666 19949 12774 20025
rect 13434 19949 13542 20025
rect 13914 19949 14022 20025
rect 14682 19949 14790 20025
rect 15162 19949 15270 20025
rect 15930 19949 16038 20025
rect 16410 19949 16518 20025
rect 17178 19949 17286 20025
rect 17658 19949 17766 20025
rect 18426 19949 18534 20025
rect 18906 19949 19014 20025
rect 19674 19949 19782 20025
rect 20154 19949 20262 20025
rect 20922 19949 21030 20025
rect 21402 19949 21510 20025
rect 22170 19949 22278 20025
rect 22650 19949 22758 20025
rect 23418 19949 23526 20025
rect 23898 19949 24006 20025
rect 24666 19949 24774 20025
rect 25146 19949 25254 20025
rect 25914 19949 26022 20025
rect 26394 19949 26502 20025
rect 27162 19949 27270 20025
rect 27642 19949 27750 20025
rect 28410 19949 28518 20025
rect 28890 19949 28998 20025
rect 29658 19949 29766 20025
rect 30138 19949 30246 20025
rect 30906 19949 31014 20025
rect 31386 19949 31494 20025
rect 32154 19949 32262 20025
rect 32634 19949 32742 20025
rect 33402 19949 33510 20025
rect 33882 19949 33990 20025
rect 34650 19949 34758 20025
rect 35130 19949 35238 20025
rect 35898 19949 36006 20025
rect 36378 19949 36486 20025
rect 37146 19949 37254 20025
rect 37626 19949 37734 20025
rect 38394 19949 38502 20025
rect 38874 19949 38982 20025
rect 39642 19949 39750 20025
rect 0 19853 39936 19901
rect 186 19695 294 19805
rect 954 19695 1062 19805
rect 1434 19695 1542 19805
rect 2202 19695 2310 19805
rect 2682 19695 2790 19805
rect 3450 19695 3558 19805
rect 3930 19695 4038 19805
rect 4698 19695 4806 19805
rect 5178 19695 5286 19805
rect 5946 19695 6054 19805
rect 6426 19695 6534 19805
rect 7194 19695 7302 19805
rect 7674 19695 7782 19805
rect 8442 19695 8550 19805
rect 8922 19695 9030 19805
rect 9690 19695 9798 19805
rect 10170 19695 10278 19805
rect 10938 19695 11046 19805
rect 11418 19695 11526 19805
rect 12186 19695 12294 19805
rect 12666 19695 12774 19805
rect 13434 19695 13542 19805
rect 13914 19695 14022 19805
rect 14682 19695 14790 19805
rect 15162 19695 15270 19805
rect 15930 19695 16038 19805
rect 16410 19695 16518 19805
rect 17178 19695 17286 19805
rect 17658 19695 17766 19805
rect 18426 19695 18534 19805
rect 18906 19695 19014 19805
rect 19674 19695 19782 19805
rect 20154 19695 20262 19805
rect 20922 19695 21030 19805
rect 21402 19695 21510 19805
rect 22170 19695 22278 19805
rect 22650 19695 22758 19805
rect 23418 19695 23526 19805
rect 23898 19695 24006 19805
rect 24666 19695 24774 19805
rect 25146 19695 25254 19805
rect 25914 19695 26022 19805
rect 26394 19695 26502 19805
rect 27162 19695 27270 19805
rect 27642 19695 27750 19805
rect 28410 19695 28518 19805
rect 28890 19695 28998 19805
rect 29658 19695 29766 19805
rect 30138 19695 30246 19805
rect 30906 19695 31014 19805
rect 31386 19695 31494 19805
rect 32154 19695 32262 19805
rect 32634 19695 32742 19805
rect 33402 19695 33510 19805
rect 33882 19695 33990 19805
rect 34650 19695 34758 19805
rect 35130 19695 35238 19805
rect 35898 19695 36006 19805
rect 36378 19695 36486 19805
rect 37146 19695 37254 19805
rect 37626 19695 37734 19805
rect 38394 19695 38502 19805
rect 38874 19695 38982 19805
rect 39642 19695 39750 19805
rect 0 19599 39936 19647
rect 186 19475 294 19551
rect 954 19475 1062 19551
rect 1434 19475 1542 19551
rect 2202 19475 2310 19551
rect 2682 19475 2790 19551
rect 3450 19475 3558 19551
rect 3930 19475 4038 19551
rect 4698 19475 4806 19551
rect 5178 19475 5286 19551
rect 5946 19475 6054 19551
rect 6426 19475 6534 19551
rect 7194 19475 7302 19551
rect 7674 19475 7782 19551
rect 8442 19475 8550 19551
rect 8922 19475 9030 19551
rect 9690 19475 9798 19551
rect 10170 19475 10278 19551
rect 10938 19475 11046 19551
rect 11418 19475 11526 19551
rect 12186 19475 12294 19551
rect 12666 19475 12774 19551
rect 13434 19475 13542 19551
rect 13914 19475 14022 19551
rect 14682 19475 14790 19551
rect 15162 19475 15270 19551
rect 15930 19475 16038 19551
rect 16410 19475 16518 19551
rect 17178 19475 17286 19551
rect 17658 19475 17766 19551
rect 18426 19475 18534 19551
rect 18906 19475 19014 19551
rect 19674 19475 19782 19551
rect 20154 19475 20262 19551
rect 20922 19475 21030 19551
rect 21402 19475 21510 19551
rect 22170 19475 22278 19551
rect 22650 19475 22758 19551
rect 23418 19475 23526 19551
rect 23898 19475 24006 19551
rect 24666 19475 24774 19551
rect 25146 19475 25254 19551
rect 25914 19475 26022 19551
rect 26394 19475 26502 19551
rect 27162 19475 27270 19551
rect 27642 19475 27750 19551
rect 28410 19475 28518 19551
rect 28890 19475 28998 19551
rect 29658 19475 29766 19551
rect 30138 19475 30246 19551
rect 30906 19475 31014 19551
rect 31386 19475 31494 19551
rect 32154 19475 32262 19551
rect 32634 19475 32742 19551
rect 33402 19475 33510 19551
rect 33882 19475 33990 19551
rect 34650 19475 34758 19551
rect 35130 19475 35238 19551
rect 35898 19475 36006 19551
rect 36378 19475 36486 19551
rect 37146 19475 37254 19551
rect 37626 19475 37734 19551
rect 38394 19475 38502 19551
rect 38874 19475 38982 19551
rect 39642 19475 39750 19551
rect 0 19379 39936 19427
rect 0 19283 39936 19331
rect 186 19159 294 19235
rect 954 19159 1062 19235
rect 1434 19159 1542 19235
rect 2202 19159 2310 19235
rect 2682 19159 2790 19235
rect 3450 19159 3558 19235
rect 3930 19159 4038 19235
rect 4698 19159 4806 19235
rect 5178 19159 5286 19235
rect 5946 19159 6054 19235
rect 6426 19159 6534 19235
rect 7194 19159 7302 19235
rect 7674 19159 7782 19235
rect 8442 19159 8550 19235
rect 8922 19159 9030 19235
rect 9690 19159 9798 19235
rect 10170 19159 10278 19235
rect 10938 19159 11046 19235
rect 11418 19159 11526 19235
rect 12186 19159 12294 19235
rect 12666 19159 12774 19235
rect 13434 19159 13542 19235
rect 13914 19159 14022 19235
rect 14682 19159 14790 19235
rect 15162 19159 15270 19235
rect 15930 19159 16038 19235
rect 16410 19159 16518 19235
rect 17178 19159 17286 19235
rect 17658 19159 17766 19235
rect 18426 19159 18534 19235
rect 18906 19159 19014 19235
rect 19674 19159 19782 19235
rect 20154 19159 20262 19235
rect 20922 19159 21030 19235
rect 21402 19159 21510 19235
rect 22170 19159 22278 19235
rect 22650 19159 22758 19235
rect 23418 19159 23526 19235
rect 23898 19159 24006 19235
rect 24666 19159 24774 19235
rect 25146 19159 25254 19235
rect 25914 19159 26022 19235
rect 26394 19159 26502 19235
rect 27162 19159 27270 19235
rect 27642 19159 27750 19235
rect 28410 19159 28518 19235
rect 28890 19159 28998 19235
rect 29658 19159 29766 19235
rect 30138 19159 30246 19235
rect 30906 19159 31014 19235
rect 31386 19159 31494 19235
rect 32154 19159 32262 19235
rect 32634 19159 32742 19235
rect 33402 19159 33510 19235
rect 33882 19159 33990 19235
rect 34650 19159 34758 19235
rect 35130 19159 35238 19235
rect 35898 19159 36006 19235
rect 36378 19159 36486 19235
rect 37146 19159 37254 19235
rect 37626 19159 37734 19235
rect 38394 19159 38502 19235
rect 38874 19159 38982 19235
rect 39642 19159 39750 19235
rect 0 19063 39936 19111
rect 186 18905 294 19015
rect 954 18905 1062 19015
rect 1434 18905 1542 19015
rect 2202 18905 2310 19015
rect 2682 18905 2790 19015
rect 3450 18905 3558 19015
rect 3930 18905 4038 19015
rect 4698 18905 4806 19015
rect 5178 18905 5286 19015
rect 5946 18905 6054 19015
rect 6426 18905 6534 19015
rect 7194 18905 7302 19015
rect 7674 18905 7782 19015
rect 8442 18905 8550 19015
rect 8922 18905 9030 19015
rect 9690 18905 9798 19015
rect 10170 18905 10278 19015
rect 10938 18905 11046 19015
rect 11418 18905 11526 19015
rect 12186 18905 12294 19015
rect 12666 18905 12774 19015
rect 13434 18905 13542 19015
rect 13914 18905 14022 19015
rect 14682 18905 14790 19015
rect 15162 18905 15270 19015
rect 15930 18905 16038 19015
rect 16410 18905 16518 19015
rect 17178 18905 17286 19015
rect 17658 18905 17766 19015
rect 18426 18905 18534 19015
rect 18906 18905 19014 19015
rect 19674 18905 19782 19015
rect 20154 18905 20262 19015
rect 20922 18905 21030 19015
rect 21402 18905 21510 19015
rect 22170 18905 22278 19015
rect 22650 18905 22758 19015
rect 23418 18905 23526 19015
rect 23898 18905 24006 19015
rect 24666 18905 24774 19015
rect 25146 18905 25254 19015
rect 25914 18905 26022 19015
rect 26394 18905 26502 19015
rect 27162 18905 27270 19015
rect 27642 18905 27750 19015
rect 28410 18905 28518 19015
rect 28890 18905 28998 19015
rect 29658 18905 29766 19015
rect 30138 18905 30246 19015
rect 30906 18905 31014 19015
rect 31386 18905 31494 19015
rect 32154 18905 32262 19015
rect 32634 18905 32742 19015
rect 33402 18905 33510 19015
rect 33882 18905 33990 19015
rect 34650 18905 34758 19015
rect 35130 18905 35238 19015
rect 35898 18905 36006 19015
rect 36378 18905 36486 19015
rect 37146 18905 37254 19015
rect 37626 18905 37734 19015
rect 38394 18905 38502 19015
rect 38874 18905 38982 19015
rect 39642 18905 39750 19015
rect 0 18809 39936 18857
rect 186 18685 294 18761
rect 954 18685 1062 18761
rect 1434 18685 1542 18761
rect 2202 18685 2310 18761
rect 2682 18685 2790 18761
rect 3450 18685 3558 18761
rect 3930 18685 4038 18761
rect 4698 18685 4806 18761
rect 5178 18685 5286 18761
rect 5946 18685 6054 18761
rect 6426 18685 6534 18761
rect 7194 18685 7302 18761
rect 7674 18685 7782 18761
rect 8442 18685 8550 18761
rect 8922 18685 9030 18761
rect 9690 18685 9798 18761
rect 10170 18685 10278 18761
rect 10938 18685 11046 18761
rect 11418 18685 11526 18761
rect 12186 18685 12294 18761
rect 12666 18685 12774 18761
rect 13434 18685 13542 18761
rect 13914 18685 14022 18761
rect 14682 18685 14790 18761
rect 15162 18685 15270 18761
rect 15930 18685 16038 18761
rect 16410 18685 16518 18761
rect 17178 18685 17286 18761
rect 17658 18685 17766 18761
rect 18426 18685 18534 18761
rect 18906 18685 19014 18761
rect 19674 18685 19782 18761
rect 20154 18685 20262 18761
rect 20922 18685 21030 18761
rect 21402 18685 21510 18761
rect 22170 18685 22278 18761
rect 22650 18685 22758 18761
rect 23418 18685 23526 18761
rect 23898 18685 24006 18761
rect 24666 18685 24774 18761
rect 25146 18685 25254 18761
rect 25914 18685 26022 18761
rect 26394 18685 26502 18761
rect 27162 18685 27270 18761
rect 27642 18685 27750 18761
rect 28410 18685 28518 18761
rect 28890 18685 28998 18761
rect 29658 18685 29766 18761
rect 30138 18685 30246 18761
rect 30906 18685 31014 18761
rect 31386 18685 31494 18761
rect 32154 18685 32262 18761
rect 32634 18685 32742 18761
rect 33402 18685 33510 18761
rect 33882 18685 33990 18761
rect 34650 18685 34758 18761
rect 35130 18685 35238 18761
rect 35898 18685 36006 18761
rect 36378 18685 36486 18761
rect 37146 18685 37254 18761
rect 37626 18685 37734 18761
rect 38394 18685 38502 18761
rect 38874 18685 38982 18761
rect 39642 18685 39750 18761
rect 0 18589 39936 18637
rect 0 18493 39936 18541
rect 186 18369 294 18445
rect 954 18369 1062 18445
rect 1434 18369 1542 18445
rect 2202 18369 2310 18445
rect 2682 18369 2790 18445
rect 3450 18369 3558 18445
rect 3930 18369 4038 18445
rect 4698 18369 4806 18445
rect 5178 18369 5286 18445
rect 5946 18369 6054 18445
rect 6426 18369 6534 18445
rect 7194 18369 7302 18445
rect 7674 18369 7782 18445
rect 8442 18369 8550 18445
rect 8922 18369 9030 18445
rect 9690 18369 9798 18445
rect 10170 18369 10278 18445
rect 10938 18369 11046 18445
rect 11418 18369 11526 18445
rect 12186 18369 12294 18445
rect 12666 18369 12774 18445
rect 13434 18369 13542 18445
rect 13914 18369 14022 18445
rect 14682 18369 14790 18445
rect 15162 18369 15270 18445
rect 15930 18369 16038 18445
rect 16410 18369 16518 18445
rect 17178 18369 17286 18445
rect 17658 18369 17766 18445
rect 18426 18369 18534 18445
rect 18906 18369 19014 18445
rect 19674 18369 19782 18445
rect 20154 18369 20262 18445
rect 20922 18369 21030 18445
rect 21402 18369 21510 18445
rect 22170 18369 22278 18445
rect 22650 18369 22758 18445
rect 23418 18369 23526 18445
rect 23898 18369 24006 18445
rect 24666 18369 24774 18445
rect 25146 18369 25254 18445
rect 25914 18369 26022 18445
rect 26394 18369 26502 18445
rect 27162 18369 27270 18445
rect 27642 18369 27750 18445
rect 28410 18369 28518 18445
rect 28890 18369 28998 18445
rect 29658 18369 29766 18445
rect 30138 18369 30246 18445
rect 30906 18369 31014 18445
rect 31386 18369 31494 18445
rect 32154 18369 32262 18445
rect 32634 18369 32742 18445
rect 33402 18369 33510 18445
rect 33882 18369 33990 18445
rect 34650 18369 34758 18445
rect 35130 18369 35238 18445
rect 35898 18369 36006 18445
rect 36378 18369 36486 18445
rect 37146 18369 37254 18445
rect 37626 18369 37734 18445
rect 38394 18369 38502 18445
rect 38874 18369 38982 18445
rect 39642 18369 39750 18445
rect 0 18273 39936 18321
rect 186 18115 294 18225
rect 954 18115 1062 18225
rect 1434 18115 1542 18225
rect 2202 18115 2310 18225
rect 2682 18115 2790 18225
rect 3450 18115 3558 18225
rect 3930 18115 4038 18225
rect 4698 18115 4806 18225
rect 5178 18115 5286 18225
rect 5946 18115 6054 18225
rect 6426 18115 6534 18225
rect 7194 18115 7302 18225
rect 7674 18115 7782 18225
rect 8442 18115 8550 18225
rect 8922 18115 9030 18225
rect 9690 18115 9798 18225
rect 10170 18115 10278 18225
rect 10938 18115 11046 18225
rect 11418 18115 11526 18225
rect 12186 18115 12294 18225
rect 12666 18115 12774 18225
rect 13434 18115 13542 18225
rect 13914 18115 14022 18225
rect 14682 18115 14790 18225
rect 15162 18115 15270 18225
rect 15930 18115 16038 18225
rect 16410 18115 16518 18225
rect 17178 18115 17286 18225
rect 17658 18115 17766 18225
rect 18426 18115 18534 18225
rect 18906 18115 19014 18225
rect 19674 18115 19782 18225
rect 20154 18115 20262 18225
rect 20922 18115 21030 18225
rect 21402 18115 21510 18225
rect 22170 18115 22278 18225
rect 22650 18115 22758 18225
rect 23418 18115 23526 18225
rect 23898 18115 24006 18225
rect 24666 18115 24774 18225
rect 25146 18115 25254 18225
rect 25914 18115 26022 18225
rect 26394 18115 26502 18225
rect 27162 18115 27270 18225
rect 27642 18115 27750 18225
rect 28410 18115 28518 18225
rect 28890 18115 28998 18225
rect 29658 18115 29766 18225
rect 30138 18115 30246 18225
rect 30906 18115 31014 18225
rect 31386 18115 31494 18225
rect 32154 18115 32262 18225
rect 32634 18115 32742 18225
rect 33402 18115 33510 18225
rect 33882 18115 33990 18225
rect 34650 18115 34758 18225
rect 35130 18115 35238 18225
rect 35898 18115 36006 18225
rect 36378 18115 36486 18225
rect 37146 18115 37254 18225
rect 37626 18115 37734 18225
rect 38394 18115 38502 18225
rect 38874 18115 38982 18225
rect 39642 18115 39750 18225
rect 0 18019 39936 18067
rect 186 17895 294 17971
rect 954 17895 1062 17971
rect 1434 17895 1542 17971
rect 2202 17895 2310 17971
rect 2682 17895 2790 17971
rect 3450 17895 3558 17971
rect 3930 17895 4038 17971
rect 4698 17895 4806 17971
rect 5178 17895 5286 17971
rect 5946 17895 6054 17971
rect 6426 17895 6534 17971
rect 7194 17895 7302 17971
rect 7674 17895 7782 17971
rect 8442 17895 8550 17971
rect 8922 17895 9030 17971
rect 9690 17895 9798 17971
rect 10170 17895 10278 17971
rect 10938 17895 11046 17971
rect 11418 17895 11526 17971
rect 12186 17895 12294 17971
rect 12666 17895 12774 17971
rect 13434 17895 13542 17971
rect 13914 17895 14022 17971
rect 14682 17895 14790 17971
rect 15162 17895 15270 17971
rect 15930 17895 16038 17971
rect 16410 17895 16518 17971
rect 17178 17895 17286 17971
rect 17658 17895 17766 17971
rect 18426 17895 18534 17971
rect 18906 17895 19014 17971
rect 19674 17895 19782 17971
rect 20154 17895 20262 17971
rect 20922 17895 21030 17971
rect 21402 17895 21510 17971
rect 22170 17895 22278 17971
rect 22650 17895 22758 17971
rect 23418 17895 23526 17971
rect 23898 17895 24006 17971
rect 24666 17895 24774 17971
rect 25146 17895 25254 17971
rect 25914 17895 26022 17971
rect 26394 17895 26502 17971
rect 27162 17895 27270 17971
rect 27642 17895 27750 17971
rect 28410 17895 28518 17971
rect 28890 17895 28998 17971
rect 29658 17895 29766 17971
rect 30138 17895 30246 17971
rect 30906 17895 31014 17971
rect 31386 17895 31494 17971
rect 32154 17895 32262 17971
rect 32634 17895 32742 17971
rect 33402 17895 33510 17971
rect 33882 17895 33990 17971
rect 34650 17895 34758 17971
rect 35130 17895 35238 17971
rect 35898 17895 36006 17971
rect 36378 17895 36486 17971
rect 37146 17895 37254 17971
rect 37626 17895 37734 17971
rect 38394 17895 38502 17971
rect 38874 17895 38982 17971
rect 39642 17895 39750 17971
rect 0 17799 39936 17847
rect 0 17703 39936 17751
rect 186 17579 294 17655
rect 954 17579 1062 17655
rect 1434 17579 1542 17655
rect 2202 17579 2310 17655
rect 2682 17579 2790 17655
rect 3450 17579 3558 17655
rect 3930 17579 4038 17655
rect 4698 17579 4806 17655
rect 5178 17579 5286 17655
rect 5946 17579 6054 17655
rect 6426 17579 6534 17655
rect 7194 17579 7302 17655
rect 7674 17579 7782 17655
rect 8442 17579 8550 17655
rect 8922 17579 9030 17655
rect 9690 17579 9798 17655
rect 10170 17579 10278 17655
rect 10938 17579 11046 17655
rect 11418 17579 11526 17655
rect 12186 17579 12294 17655
rect 12666 17579 12774 17655
rect 13434 17579 13542 17655
rect 13914 17579 14022 17655
rect 14682 17579 14790 17655
rect 15162 17579 15270 17655
rect 15930 17579 16038 17655
rect 16410 17579 16518 17655
rect 17178 17579 17286 17655
rect 17658 17579 17766 17655
rect 18426 17579 18534 17655
rect 18906 17579 19014 17655
rect 19674 17579 19782 17655
rect 20154 17579 20262 17655
rect 20922 17579 21030 17655
rect 21402 17579 21510 17655
rect 22170 17579 22278 17655
rect 22650 17579 22758 17655
rect 23418 17579 23526 17655
rect 23898 17579 24006 17655
rect 24666 17579 24774 17655
rect 25146 17579 25254 17655
rect 25914 17579 26022 17655
rect 26394 17579 26502 17655
rect 27162 17579 27270 17655
rect 27642 17579 27750 17655
rect 28410 17579 28518 17655
rect 28890 17579 28998 17655
rect 29658 17579 29766 17655
rect 30138 17579 30246 17655
rect 30906 17579 31014 17655
rect 31386 17579 31494 17655
rect 32154 17579 32262 17655
rect 32634 17579 32742 17655
rect 33402 17579 33510 17655
rect 33882 17579 33990 17655
rect 34650 17579 34758 17655
rect 35130 17579 35238 17655
rect 35898 17579 36006 17655
rect 36378 17579 36486 17655
rect 37146 17579 37254 17655
rect 37626 17579 37734 17655
rect 38394 17579 38502 17655
rect 38874 17579 38982 17655
rect 39642 17579 39750 17655
rect 0 17483 39936 17531
rect 186 17325 294 17435
rect 954 17325 1062 17435
rect 1434 17325 1542 17435
rect 2202 17325 2310 17435
rect 2682 17325 2790 17435
rect 3450 17325 3558 17435
rect 3930 17325 4038 17435
rect 4698 17325 4806 17435
rect 5178 17325 5286 17435
rect 5946 17325 6054 17435
rect 6426 17325 6534 17435
rect 7194 17325 7302 17435
rect 7674 17325 7782 17435
rect 8442 17325 8550 17435
rect 8922 17325 9030 17435
rect 9690 17325 9798 17435
rect 10170 17325 10278 17435
rect 10938 17325 11046 17435
rect 11418 17325 11526 17435
rect 12186 17325 12294 17435
rect 12666 17325 12774 17435
rect 13434 17325 13542 17435
rect 13914 17325 14022 17435
rect 14682 17325 14790 17435
rect 15162 17325 15270 17435
rect 15930 17325 16038 17435
rect 16410 17325 16518 17435
rect 17178 17325 17286 17435
rect 17658 17325 17766 17435
rect 18426 17325 18534 17435
rect 18906 17325 19014 17435
rect 19674 17325 19782 17435
rect 20154 17325 20262 17435
rect 20922 17325 21030 17435
rect 21402 17325 21510 17435
rect 22170 17325 22278 17435
rect 22650 17325 22758 17435
rect 23418 17325 23526 17435
rect 23898 17325 24006 17435
rect 24666 17325 24774 17435
rect 25146 17325 25254 17435
rect 25914 17325 26022 17435
rect 26394 17325 26502 17435
rect 27162 17325 27270 17435
rect 27642 17325 27750 17435
rect 28410 17325 28518 17435
rect 28890 17325 28998 17435
rect 29658 17325 29766 17435
rect 30138 17325 30246 17435
rect 30906 17325 31014 17435
rect 31386 17325 31494 17435
rect 32154 17325 32262 17435
rect 32634 17325 32742 17435
rect 33402 17325 33510 17435
rect 33882 17325 33990 17435
rect 34650 17325 34758 17435
rect 35130 17325 35238 17435
rect 35898 17325 36006 17435
rect 36378 17325 36486 17435
rect 37146 17325 37254 17435
rect 37626 17325 37734 17435
rect 38394 17325 38502 17435
rect 38874 17325 38982 17435
rect 39642 17325 39750 17435
rect 0 17229 39936 17277
rect 186 17105 294 17181
rect 954 17105 1062 17181
rect 1434 17105 1542 17181
rect 2202 17105 2310 17181
rect 2682 17105 2790 17181
rect 3450 17105 3558 17181
rect 3930 17105 4038 17181
rect 4698 17105 4806 17181
rect 5178 17105 5286 17181
rect 5946 17105 6054 17181
rect 6426 17105 6534 17181
rect 7194 17105 7302 17181
rect 7674 17105 7782 17181
rect 8442 17105 8550 17181
rect 8922 17105 9030 17181
rect 9690 17105 9798 17181
rect 10170 17105 10278 17181
rect 10938 17105 11046 17181
rect 11418 17105 11526 17181
rect 12186 17105 12294 17181
rect 12666 17105 12774 17181
rect 13434 17105 13542 17181
rect 13914 17105 14022 17181
rect 14682 17105 14790 17181
rect 15162 17105 15270 17181
rect 15930 17105 16038 17181
rect 16410 17105 16518 17181
rect 17178 17105 17286 17181
rect 17658 17105 17766 17181
rect 18426 17105 18534 17181
rect 18906 17105 19014 17181
rect 19674 17105 19782 17181
rect 20154 17105 20262 17181
rect 20922 17105 21030 17181
rect 21402 17105 21510 17181
rect 22170 17105 22278 17181
rect 22650 17105 22758 17181
rect 23418 17105 23526 17181
rect 23898 17105 24006 17181
rect 24666 17105 24774 17181
rect 25146 17105 25254 17181
rect 25914 17105 26022 17181
rect 26394 17105 26502 17181
rect 27162 17105 27270 17181
rect 27642 17105 27750 17181
rect 28410 17105 28518 17181
rect 28890 17105 28998 17181
rect 29658 17105 29766 17181
rect 30138 17105 30246 17181
rect 30906 17105 31014 17181
rect 31386 17105 31494 17181
rect 32154 17105 32262 17181
rect 32634 17105 32742 17181
rect 33402 17105 33510 17181
rect 33882 17105 33990 17181
rect 34650 17105 34758 17181
rect 35130 17105 35238 17181
rect 35898 17105 36006 17181
rect 36378 17105 36486 17181
rect 37146 17105 37254 17181
rect 37626 17105 37734 17181
rect 38394 17105 38502 17181
rect 38874 17105 38982 17181
rect 39642 17105 39750 17181
rect 0 17009 39936 17057
rect 0 16913 39936 16961
rect 186 16789 294 16865
rect 954 16789 1062 16865
rect 1434 16789 1542 16865
rect 2202 16789 2310 16865
rect 2682 16789 2790 16865
rect 3450 16789 3558 16865
rect 3930 16789 4038 16865
rect 4698 16789 4806 16865
rect 5178 16789 5286 16865
rect 5946 16789 6054 16865
rect 6426 16789 6534 16865
rect 7194 16789 7302 16865
rect 7674 16789 7782 16865
rect 8442 16789 8550 16865
rect 8922 16789 9030 16865
rect 9690 16789 9798 16865
rect 10170 16789 10278 16865
rect 10938 16789 11046 16865
rect 11418 16789 11526 16865
rect 12186 16789 12294 16865
rect 12666 16789 12774 16865
rect 13434 16789 13542 16865
rect 13914 16789 14022 16865
rect 14682 16789 14790 16865
rect 15162 16789 15270 16865
rect 15930 16789 16038 16865
rect 16410 16789 16518 16865
rect 17178 16789 17286 16865
rect 17658 16789 17766 16865
rect 18426 16789 18534 16865
rect 18906 16789 19014 16865
rect 19674 16789 19782 16865
rect 20154 16789 20262 16865
rect 20922 16789 21030 16865
rect 21402 16789 21510 16865
rect 22170 16789 22278 16865
rect 22650 16789 22758 16865
rect 23418 16789 23526 16865
rect 23898 16789 24006 16865
rect 24666 16789 24774 16865
rect 25146 16789 25254 16865
rect 25914 16789 26022 16865
rect 26394 16789 26502 16865
rect 27162 16789 27270 16865
rect 27642 16789 27750 16865
rect 28410 16789 28518 16865
rect 28890 16789 28998 16865
rect 29658 16789 29766 16865
rect 30138 16789 30246 16865
rect 30906 16789 31014 16865
rect 31386 16789 31494 16865
rect 32154 16789 32262 16865
rect 32634 16789 32742 16865
rect 33402 16789 33510 16865
rect 33882 16789 33990 16865
rect 34650 16789 34758 16865
rect 35130 16789 35238 16865
rect 35898 16789 36006 16865
rect 36378 16789 36486 16865
rect 37146 16789 37254 16865
rect 37626 16789 37734 16865
rect 38394 16789 38502 16865
rect 38874 16789 38982 16865
rect 39642 16789 39750 16865
rect 0 16693 39936 16741
rect 186 16535 294 16645
rect 954 16535 1062 16645
rect 1434 16535 1542 16645
rect 2202 16535 2310 16645
rect 2682 16535 2790 16645
rect 3450 16535 3558 16645
rect 3930 16535 4038 16645
rect 4698 16535 4806 16645
rect 5178 16535 5286 16645
rect 5946 16535 6054 16645
rect 6426 16535 6534 16645
rect 7194 16535 7302 16645
rect 7674 16535 7782 16645
rect 8442 16535 8550 16645
rect 8922 16535 9030 16645
rect 9690 16535 9798 16645
rect 10170 16535 10278 16645
rect 10938 16535 11046 16645
rect 11418 16535 11526 16645
rect 12186 16535 12294 16645
rect 12666 16535 12774 16645
rect 13434 16535 13542 16645
rect 13914 16535 14022 16645
rect 14682 16535 14790 16645
rect 15162 16535 15270 16645
rect 15930 16535 16038 16645
rect 16410 16535 16518 16645
rect 17178 16535 17286 16645
rect 17658 16535 17766 16645
rect 18426 16535 18534 16645
rect 18906 16535 19014 16645
rect 19674 16535 19782 16645
rect 20154 16535 20262 16645
rect 20922 16535 21030 16645
rect 21402 16535 21510 16645
rect 22170 16535 22278 16645
rect 22650 16535 22758 16645
rect 23418 16535 23526 16645
rect 23898 16535 24006 16645
rect 24666 16535 24774 16645
rect 25146 16535 25254 16645
rect 25914 16535 26022 16645
rect 26394 16535 26502 16645
rect 27162 16535 27270 16645
rect 27642 16535 27750 16645
rect 28410 16535 28518 16645
rect 28890 16535 28998 16645
rect 29658 16535 29766 16645
rect 30138 16535 30246 16645
rect 30906 16535 31014 16645
rect 31386 16535 31494 16645
rect 32154 16535 32262 16645
rect 32634 16535 32742 16645
rect 33402 16535 33510 16645
rect 33882 16535 33990 16645
rect 34650 16535 34758 16645
rect 35130 16535 35238 16645
rect 35898 16535 36006 16645
rect 36378 16535 36486 16645
rect 37146 16535 37254 16645
rect 37626 16535 37734 16645
rect 38394 16535 38502 16645
rect 38874 16535 38982 16645
rect 39642 16535 39750 16645
rect 0 16439 39936 16487
rect 186 16315 294 16391
rect 954 16315 1062 16391
rect 1434 16315 1542 16391
rect 2202 16315 2310 16391
rect 2682 16315 2790 16391
rect 3450 16315 3558 16391
rect 3930 16315 4038 16391
rect 4698 16315 4806 16391
rect 5178 16315 5286 16391
rect 5946 16315 6054 16391
rect 6426 16315 6534 16391
rect 7194 16315 7302 16391
rect 7674 16315 7782 16391
rect 8442 16315 8550 16391
rect 8922 16315 9030 16391
rect 9690 16315 9798 16391
rect 10170 16315 10278 16391
rect 10938 16315 11046 16391
rect 11418 16315 11526 16391
rect 12186 16315 12294 16391
rect 12666 16315 12774 16391
rect 13434 16315 13542 16391
rect 13914 16315 14022 16391
rect 14682 16315 14790 16391
rect 15162 16315 15270 16391
rect 15930 16315 16038 16391
rect 16410 16315 16518 16391
rect 17178 16315 17286 16391
rect 17658 16315 17766 16391
rect 18426 16315 18534 16391
rect 18906 16315 19014 16391
rect 19674 16315 19782 16391
rect 20154 16315 20262 16391
rect 20922 16315 21030 16391
rect 21402 16315 21510 16391
rect 22170 16315 22278 16391
rect 22650 16315 22758 16391
rect 23418 16315 23526 16391
rect 23898 16315 24006 16391
rect 24666 16315 24774 16391
rect 25146 16315 25254 16391
rect 25914 16315 26022 16391
rect 26394 16315 26502 16391
rect 27162 16315 27270 16391
rect 27642 16315 27750 16391
rect 28410 16315 28518 16391
rect 28890 16315 28998 16391
rect 29658 16315 29766 16391
rect 30138 16315 30246 16391
rect 30906 16315 31014 16391
rect 31386 16315 31494 16391
rect 32154 16315 32262 16391
rect 32634 16315 32742 16391
rect 33402 16315 33510 16391
rect 33882 16315 33990 16391
rect 34650 16315 34758 16391
rect 35130 16315 35238 16391
rect 35898 16315 36006 16391
rect 36378 16315 36486 16391
rect 37146 16315 37254 16391
rect 37626 16315 37734 16391
rect 38394 16315 38502 16391
rect 38874 16315 38982 16391
rect 39642 16315 39750 16391
rect 0 16219 39936 16267
rect 0 16123 39936 16171
rect 186 15999 294 16075
rect 954 15999 1062 16075
rect 1434 15999 1542 16075
rect 2202 15999 2310 16075
rect 2682 15999 2790 16075
rect 3450 15999 3558 16075
rect 3930 15999 4038 16075
rect 4698 15999 4806 16075
rect 5178 15999 5286 16075
rect 5946 15999 6054 16075
rect 6426 15999 6534 16075
rect 7194 15999 7302 16075
rect 7674 15999 7782 16075
rect 8442 15999 8550 16075
rect 8922 15999 9030 16075
rect 9690 15999 9798 16075
rect 10170 15999 10278 16075
rect 10938 15999 11046 16075
rect 11418 15999 11526 16075
rect 12186 15999 12294 16075
rect 12666 15999 12774 16075
rect 13434 15999 13542 16075
rect 13914 15999 14022 16075
rect 14682 15999 14790 16075
rect 15162 15999 15270 16075
rect 15930 15999 16038 16075
rect 16410 15999 16518 16075
rect 17178 15999 17286 16075
rect 17658 15999 17766 16075
rect 18426 15999 18534 16075
rect 18906 15999 19014 16075
rect 19674 15999 19782 16075
rect 20154 15999 20262 16075
rect 20922 15999 21030 16075
rect 21402 15999 21510 16075
rect 22170 15999 22278 16075
rect 22650 15999 22758 16075
rect 23418 15999 23526 16075
rect 23898 15999 24006 16075
rect 24666 15999 24774 16075
rect 25146 15999 25254 16075
rect 25914 15999 26022 16075
rect 26394 15999 26502 16075
rect 27162 15999 27270 16075
rect 27642 15999 27750 16075
rect 28410 15999 28518 16075
rect 28890 15999 28998 16075
rect 29658 15999 29766 16075
rect 30138 15999 30246 16075
rect 30906 15999 31014 16075
rect 31386 15999 31494 16075
rect 32154 15999 32262 16075
rect 32634 15999 32742 16075
rect 33402 15999 33510 16075
rect 33882 15999 33990 16075
rect 34650 15999 34758 16075
rect 35130 15999 35238 16075
rect 35898 15999 36006 16075
rect 36378 15999 36486 16075
rect 37146 15999 37254 16075
rect 37626 15999 37734 16075
rect 38394 15999 38502 16075
rect 38874 15999 38982 16075
rect 39642 15999 39750 16075
rect 0 15903 39936 15951
rect 186 15745 294 15855
rect 954 15745 1062 15855
rect 1434 15745 1542 15855
rect 2202 15745 2310 15855
rect 2682 15745 2790 15855
rect 3450 15745 3558 15855
rect 3930 15745 4038 15855
rect 4698 15745 4806 15855
rect 5178 15745 5286 15855
rect 5946 15745 6054 15855
rect 6426 15745 6534 15855
rect 7194 15745 7302 15855
rect 7674 15745 7782 15855
rect 8442 15745 8550 15855
rect 8922 15745 9030 15855
rect 9690 15745 9798 15855
rect 10170 15745 10278 15855
rect 10938 15745 11046 15855
rect 11418 15745 11526 15855
rect 12186 15745 12294 15855
rect 12666 15745 12774 15855
rect 13434 15745 13542 15855
rect 13914 15745 14022 15855
rect 14682 15745 14790 15855
rect 15162 15745 15270 15855
rect 15930 15745 16038 15855
rect 16410 15745 16518 15855
rect 17178 15745 17286 15855
rect 17658 15745 17766 15855
rect 18426 15745 18534 15855
rect 18906 15745 19014 15855
rect 19674 15745 19782 15855
rect 20154 15745 20262 15855
rect 20922 15745 21030 15855
rect 21402 15745 21510 15855
rect 22170 15745 22278 15855
rect 22650 15745 22758 15855
rect 23418 15745 23526 15855
rect 23898 15745 24006 15855
rect 24666 15745 24774 15855
rect 25146 15745 25254 15855
rect 25914 15745 26022 15855
rect 26394 15745 26502 15855
rect 27162 15745 27270 15855
rect 27642 15745 27750 15855
rect 28410 15745 28518 15855
rect 28890 15745 28998 15855
rect 29658 15745 29766 15855
rect 30138 15745 30246 15855
rect 30906 15745 31014 15855
rect 31386 15745 31494 15855
rect 32154 15745 32262 15855
rect 32634 15745 32742 15855
rect 33402 15745 33510 15855
rect 33882 15745 33990 15855
rect 34650 15745 34758 15855
rect 35130 15745 35238 15855
rect 35898 15745 36006 15855
rect 36378 15745 36486 15855
rect 37146 15745 37254 15855
rect 37626 15745 37734 15855
rect 38394 15745 38502 15855
rect 38874 15745 38982 15855
rect 39642 15745 39750 15855
rect 0 15649 39936 15697
rect 186 15525 294 15601
rect 954 15525 1062 15601
rect 1434 15525 1542 15601
rect 2202 15525 2310 15601
rect 2682 15525 2790 15601
rect 3450 15525 3558 15601
rect 3930 15525 4038 15601
rect 4698 15525 4806 15601
rect 5178 15525 5286 15601
rect 5946 15525 6054 15601
rect 6426 15525 6534 15601
rect 7194 15525 7302 15601
rect 7674 15525 7782 15601
rect 8442 15525 8550 15601
rect 8922 15525 9030 15601
rect 9690 15525 9798 15601
rect 10170 15525 10278 15601
rect 10938 15525 11046 15601
rect 11418 15525 11526 15601
rect 12186 15525 12294 15601
rect 12666 15525 12774 15601
rect 13434 15525 13542 15601
rect 13914 15525 14022 15601
rect 14682 15525 14790 15601
rect 15162 15525 15270 15601
rect 15930 15525 16038 15601
rect 16410 15525 16518 15601
rect 17178 15525 17286 15601
rect 17658 15525 17766 15601
rect 18426 15525 18534 15601
rect 18906 15525 19014 15601
rect 19674 15525 19782 15601
rect 20154 15525 20262 15601
rect 20922 15525 21030 15601
rect 21402 15525 21510 15601
rect 22170 15525 22278 15601
rect 22650 15525 22758 15601
rect 23418 15525 23526 15601
rect 23898 15525 24006 15601
rect 24666 15525 24774 15601
rect 25146 15525 25254 15601
rect 25914 15525 26022 15601
rect 26394 15525 26502 15601
rect 27162 15525 27270 15601
rect 27642 15525 27750 15601
rect 28410 15525 28518 15601
rect 28890 15525 28998 15601
rect 29658 15525 29766 15601
rect 30138 15525 30246 15601
rect 30906 15525 31014 15601
rect 31386 15525 31494 15601
rect 32154 15525 32262 15601
rect 32634 15525 32742 15601
rect 33402 15525 33510 15601
rect 33882 15525 33990 15601
rect 34650 15525 34758 15601
rect 35130 15525 35238 15601
rect 35898 15525 36006 15601
rect 36378 15525 36486 15601
rect 37146 15525 37254 15601
rect 37626 15525 37734 15601
rect 38394 15525 38502 15601
rect 38874 15525 38982 15601
rect 39642 15525 39750 15601
rect 0 15429 39936 15477
rect 0 15333 39936 15381
rect 186 15209 294 15285
rect 954 15209 1062 15285
rect 1434 15209 1542 15285
rect 2202 15209 2310 15285
rect 2682 15209 2790 15285
rect 3450 15209 3558 15285
rect 3930 15209 4038 15285
rect 4698 15209 4806 15285
rect 5178 15209 5286 15285
rect 5946 15209 6054 15285
rect 6426 15209 6534 15285
rect 7194 15209 7302 15285
rect 7674 15209 7782 15285
rect 8442 15209 8550 15285
rect 8922 15209 9030 15285
rect 9690 15209 9798 15285
rect 10170 15209 10278 15285
rect 10938 15209 11046 15285
rect 11418 15209 11526 15285
rect 12186 15209 12294 15285
rect 12666 15209 12774 15285
rect 13434 15209 13542 15285
rect 13914 15209 14022 15285
rect 14682 15209 14790 15285
rect 15162 15209 15270 15285
rect 15930 15209 16038 15285
rect 16410 15209 16518 15285
rect 17178 15209 17286 15285
rect 17658 15209 17766 15285
rect 18426 15209 18534 15285
rect 18906 15209 19014 15285
rect 19674 15209 19782 15285
rect 20154 15209 20262 15285
rect 20922 15209 21030 15285
rect 21402 15209 21510 15285
rect 22170 15209 22278 15285
rect 22650 15209 22758 15285
rect 23418 15209 23526 15285
rect 23898 15209 24006 15285
rect 24666 15209 24774 15285
rect 25146 15209 25254 15285
rect 25914 15209 26022 15285
rect 26394 15209 26502 15285
rect 27162 15209 27270 15285
rect 27642 15209 27750 15285
rect 28410 15209 28518 15285
rect 28890 15209 28998 15285
rect 29658 15209 29766 15285
rect 30138 15209 30246 15285
rect 30906 15209 31014 15285
rect 31386 15209 31494 15285
rect 32154 15209 32262 15285
rect 32634 15209 32742 15285
rect 33402 15209 33510 15285
rect 33882 15209 33990 15285
rect 34650 15209 34758 15285
rect 35130 15209 35238 15285
rect 35898 15209 36006 15285
rect 36378 15209 36486 15285
rect 37146 15209 37254 15285
rect 37626 15209 37734 15285
rect 38394 15209 38502 15285
rect 38874 15209 38982 15285
rect 39642 15209 39750 15285
rect 0 15113 39936 15161
rect 186 14955 294 15065
rect 954 14955 1062 15065
rect 1434 14955 1542 15065
rect 2202 14955 2310 15065
rect 2682 14955 2790 15065
rect 3450 14955 3558 15065
rect 3930 14955 4038 15065
rect 4698 14955 4806 15065
rect 5178 14955 5286 15065
rect 5946 14955 6054 15065
rect 6426 14955 6534 15065
rect 7194 14955 7302 15065
rect 7674 14955 7782 15065
rect 8442 14955 8550 15065
rect 8922 14955 9030 15065
rect 9690 14955 9798 15065
rect 10170 14955 10278 15065
rect 10938 14955 11046 15065
rect 11418 14955 11526 15065
rect 12186 14955 12294 15065
rect 12666 14955 12774 15065
rect 13434 14955 13542 15065
rect 13914 14955 14022 15065
rect 14682 14955 14790 15065
rect 15162 14955 15270 15065
rect 15930 14955 16038 15065
rect 16410 14955 16518 15065
rect 17178 14955 17286 15065
rect 17658 14955 17766 15065
rect 18426 14955 18534 15065
rect 18906 14955 19014 15065
rect 19674 14955 19782 15065
rect 20154 14955 20262 15065
rect 20922 14955 21030 15065
rect 21402 14955 21510 15065
rect 22170 14955 22278 15065
rect 22650 14955 22758 15065
rect 23418 14955 23526 15065
rect 23898 14955 24006 15065
rect 24666 14955 24774 15065
rect 25146 14955 25254 15065
rect 25914 14955 26022 15065
rect 26394 14955 26502 15065
rect 27162 14955 27270 15065
rect 27642 14955 27750 15065
rect 28410 14955 28518 15065
rect 28890 14955 28998 15065
rect 29658 14955 29766 15065
rect 30138 14955 30246 15065
rect 30906 14955 31014 15065
rect 31386 14955 31494 15065
rect 32154 14955 32262 15065
rect 32634 14955 32742 15065
rect 33402 14955 33510 15065
rect 33882 14955 33990 15065
rect 34650 14955 34758 15065
rect 35130 14955 35238 15065
rect 35898 14955 36006 15065
rect 36378 14955 36486 15065
rect 37146 14955 37254 15065
rect 37626 14955 37734 15065
rect 38394 14955 38502 15065
rect 38874 14955 38982 15065
rect 39642 14955 39750 15065
rect 0 14859 39936 14907
rect 186 14735 294 14811
rect 954 14735 1062 14811
rect 1434 14735 1542 14811
rect 2202 14735 2310 14811
rect 2682 14735 2790 14811
rect 3450 14735 3558 14811
rect 3930 14735 4038 14811
rect 4698 14735 4806 14811
rect 5178 14735 5286 14811
rect 5946 14735 6054 14811
rect 6426 14735 6534 14811
rect 7194 14735 7302 14811
rect 7674 14735 7782 14811
rect 8442 14735 8550 14811
rect 8922 14735 9030 14811
rect 9690 14735 9798 14811
rect 10170 14735 10278 14811
rect 10938 14735 11046 14811
rect 11418 14735 11526 14811
rect 12186 14735 12294 14811
rect 12666 14735 12774 14811
rect 13434 14735 13542 14811
rect 13914 14735 14022 14811
rect 14682 14735 14790 14811
rect 15162 14735 15270 14811
rect 15930 14735 16038 14811
rect 16410 14735 16518 14811
rect 17178 14735 17286 14811
rect 17658 14735 17766 14811
rect 18426 14735 18534 14811
rect 18906 14735 19014 14811
rect 19674 14735 19782 14811
rect 20154 14735 20262 14811
rect 20922 14735 21030 14811
rect 21402 14735 21510 14811
rect 22170 14735 22278 14811
rect 22650 14735 22758 14811
rect 23418 14735 23526 14811
rect 23898 14735 24006 14811
rect 24666 14735 24774 14811
rect 25146 14735 25254 14811
rect 25914 14735 26022 14811
rect 26394 14735 26502 14811
rect 27162 14735 27270 14811
rect 27642 14735 27750 14811
rect 28410 14735 28518 14811
rect 28890 14735 28998 14811
rect 29658 14735 29766 14811
rect 30138 14735 30246 14811
rect 30906 14735 31014 14811
rect 31386 14735 31494 14811
rect 32154 14735 32262 14811
rect 32634 14735 32742 14811
rect 33402 14735 33510 14811
rect 33882 14735 33990 14811
rect 34650 14735 34758 14811
rect 35130 14735 35238 14811
rect 35898 14735 36006 14811
rect 36378 14735 36486 14811
rect 37146 14735 37254 14811
rect 37626 14735 37734 14811
rect 38394 14735 38502 14811
rect 38874 14735 38982 14811
rect 39642 14735 39750 14811
rect 0 14639 39936 14687
rect 0 14543 39936 14591
rect 186 14419 294 14495
rect 954 14419 1062 14495
rect 1434 14419 1542 14495
rect 2202 14419 2310 14495
rect 2682 14419 2790 14495
rect 3450 14419 3558 14495
rect 3930 14419 4038 14495
rect 4698 14419 4806 14495
rect 5178 14419 5286 14495
rect 5946 14419 6054 14495
rect 6426 14419 6534 14495
rect 7194 14419 7302 14495
rect 7674 14419 7782 14495
rect 8442 14419 8550 14495
rect 8922 14419 9030 14495
rect 9690 14419 9798 14495
rect 10170 14419 10278 14495
rect 10938 14419 11046 14495
rect 11418 14419 11526 14495
rect 12186 14419 12294 14495
rect 12666 14419 12774 14495
rect 13434 14419 13542 14495
rect 13914 14419 14022 14495
rect 14682 14419 14790 14495
rect 15162 14419 15270 14495
rect 15930 14419 16038 14495
rect 16410 14419 16518 14495
rect 17178 14419 17286 14495
rect 17658 14419 17766 14495
rect 18426 14419 18534 14495
rect 18906 14419 19014 14495
rect 19674 14419 19782 14495
rect 20154 14419 20262 14495
rect 20922 14419 21030 14495
rect 21402 14419 21510 14495
rect 22170 14419 22278 14495
rect 22650 14419 22758 14495
rect 23418 14419 23526 14495
rect 23898 14419 24006 14495
rect 24666 14419 24774 14495
rect 25146 14419 25254 14495
rect 25914 14419 26022 14495
rect 26394 14419 26502 14495
rect 27162 14419 27270 14495
rect 27642 14419 27750 14495
rect 28410 14419 28518 14495
rect 28890 14419 28998 14495
rect 29658 14419 29766 14495
rect 30138 14419 30246 14495
rect 30906 14419 31014 14495
rect 31386 14419 31494 14495
rect 32154 14419 32262 14495
rect 32634 14419 32742 14495
rect 33402 14419 33510 14495
rect 33882 14419 33990 14495
rect 34650 14419 34758 14495
rect 35130 14419 35238 14495
rect 35898 14419 36006 14495
rect 36378 14419 36486 14495
rect 37146 14419 37254 14495
rect 37626 14419 37734 14495
rect 38394 14419 38502 14495
rect 38874 14419 38982 14495
rect 39642 14419 39750 14495
rect 0 14323 39936 14371
rect 186 14165 294 14275
rect 954 14165 1062 14275
rect 1434 14165 1542 14275
rect 2202 14165 2310 14275
rect 2682 14165 2790 14275
rect 3450 14165 3558 14275
rect 3930 14165 4038 14275
rect 4698 14165 4806 14275
rect 5178 14165 5286 14275
rect 5946 14165 6054 14275
rect 6426 14165 6534 14275
rect 7194 14165 7302 14275
rect 7674 14165 7782 14275
rect 8442 14165 8550 14275
rect 8922 14165 9030 14275
rect 9690 14165 9798 14275
rect 10170 14165 10278 14275
rect 10938 14165 11046 14275
rect 11418 14165 11526 14275
rect 12186 14165 12294 14275
rect 12666 14165 12774 14275
rect 13434 14165 13542 14275
rect 13914 14165 14022 14275
rect 14682 14165 14790 14275
rect 15162 14165 15270 14275
rect 15930 14165 16038 14275
rect 16410 14165 16518 14275
rect 17178 14165 17286 14275
rect 17658 14165 17766 14275
rect 18426 14165 18534 14275
rect 18906 14165 19014 14275
rect 19674 14165 19782 14275
rect 20154 14165 20262 14275
rect 20922 14165 21030 14275
rect 21402 14165 21510 14275
rect 22170 14165 22278 14275
rect 22650 14165 22758 14275
rect 23418 14165 23526 14275
rect 23898 14165 24006 14275
rect 24666 14165 24774 14275
rect 25146 14165 25254 14275
rect 25914 14165 26022 14275
rect 26394 14165 26502 14275
rect 27162 14165 27270 14275
rect 27642 14165 27750 14275
rect 28410 14165 28518 14275
rect 28890 14165 28998 14275
rect 29658 14165 29766 14275
rect 30138 14165 30246 14275
rect 30906 14165 31014 14275
rect 31386 14165 31494 14275
rect 32154 14165 32262 14275
rect 32634 14165 32742 14275
rect 33402 14165 33510 14275
rect 33882 14165 33990 14275
rect 34650 14165 34758 14275
rect 35130 14165 35238 14275
rect 35898 14165 36006 14275
rect 36378 14165 36486 14275
rect 37146 14165 37254 14275
rect 37626 14165 37734 14275
rect 38394 14165 38502 14275
rect 38874 14165 38982 14275
rect 39642 14165 39750 14275
rect 0 14069 39936 14117
rect 186 13945 294 14021
rect 954 13945 1062 14021
rect 1434 13945 1542 14021
rect 2202 13945 2310 14021
rect 2682 13945 2790 14021
rect 3450 13945 3558 14021
rect 3930 13945 4038 14021
rect 4698 13945 4806 14021
rect 5178 13945 5286 14021
rect 5946 13945 6054 14021
rect 6426 13945 6534 14021
rect 7194 13945 7302 14021
rect 7674 13945 7782 14021
rect 8442 13945 8550 14021
rect 8922 13945 9030 14021
rect 9690 13945 9798 14021
rect 10170 13945 10278 14021
rect 10938 13945 11046 14021
rect 11418 13945 11526 14021
rect 12186 13945 12294 14021
rect 12666 13945 12774 14021
rect 13434 13945 13542 14021
rect 13914 13945 14022 14021
rect 14682 13945 14790 14021
rect 15162 13945 15270 14021
rect 15930 13945 16038 14021
rect 16410 13945 16518 14021
rect 17178 13945 17286 14021
rect 17658 13945 17766 14021
rect 18426 13945 18534 14021
rect 18906 13945 19014 14021
rect 19674 13945 19782 14021
rect 20154 13945 20262 14021
rect 20922 13945 21030 14021
rect 21402 13945 21510 14021
rect 22170 13945 22278 14021
rect 22650 13945 22758 14021
rect 23418 13945 23526 14021
rect 23898 13945 24006 14021
rect 24666 13945 24774 14021
rect 25146 13945 25254 14021
rect 25914 13945 26022 14021
rect 26394 13945 26502 14021
rect 27162 13945 27270 14021
rect 27642 13945 27750 14021
rect 28410 13945 28518 14021
rect 28890 13945 28998 14021
rect 29658 13945 29766 14021
rect 30138 13945 30246 14021
rect 30906 13945 31014 14021
rect 31386 13945 31494 14021
rect 32154 13945 32262 14021
rect 32634 13945 32742 14021
rect 33402 13945 33510 14021
rect 33882 13945 33990 14021
rect 34650 13945 34758 14021
rect 35130 13945 35238 14021
rect 35898 13945 36006 14021
rect 36378 13945 36486 14021
rect 37146 13945 37254 14021
rect 37626 13945 37734 14021
rect 38394 13945 38502 14021
rect 38874 13945 38982 14021
rect 39642 13945 39750 14021
rect 0 13849 39936 13897
rect 0 13753 39936 13801
rect 186 13629 294 13705
rect 954 13629 1062 13705
rect 1434 13629 1542 13705
rect 2202 13629 2310 13705
rect 2682 13629 2790 13705
rect 3450 13629 3558 13705
rect 3930 13629 4038 13705
rect 4698 13629 4806 13705
rect 5178 13629 5286 13705
rect 5946 13629 6054 13705
rect 6426 13629 6534 13705
rect 7194 13629 7302 13705
rect 7674 13629 7782 13705
rect 8442 13629 8550 13705
rect 8922 13629 9030 13705
rect 9690 13629 9798 13705
rect 10170 13629 10278 13705
rect 10938 13629 11046 13705
rect 11418 13629 11526 13705
rect 12186 13629 12294 13705
rect 12666 13629 12774 13705
rect 13434 13629 13542 13705
rect 13914 13629 14022 13705
rect 14682 13629 14790 13705
rect 15162 13629 15270 13705
rect 15930 13629 16038 13705
rect 16410 13629 16518 13705
rect 17178 13629 17286 13705
rect 17658 13629 17766 13705
rect 18426 13629 18534 13705
rect 18906 13629 19014 13705
rect 19674 13629 19782 13705
rect 20154 13629 20262 13705
rect 20922 13629 21030 13705
rect 21402 13629 21510 13705
rect 22170 13629 22278 13705
rect 22650 13629 22758 13705
rect 23418 13629 23526 13705
rect 23898 13629 24006 13705
rect 24666 13629 24774 13705
rect 25146 13629 25254 13705
rect 25914 13629 26022 13705
rect 26394 13629 26502 13705
rect 27162 13629 27270 13705
rect 27642 13629 27750 13705
rect 28410 13629 28518 13705
rect 28890 13629 28998 13705
rect 29658 13629 29766 13705
rect 30138 13629 30246 13705
rect 30906 13629 31014 13705
rect 31386 13629 31494 13705
rect 32154 13629 32262 13705
rect 32634 13629 32742 13705
rect 33402 13629 33510 13705
rect 33882 13629 33990 13705
rect 34650 13629 34758 13705
rect 35130 13629 35238 13705
rect 35898 13629 36006 13705
rect 36378 13629 36486 13705
rect 37146 13629 37254 13705
rect 37626 13629 37734 13705
rect 38394 13629 38502 13705
rect 38874 13629 38982 13705
rect 39642 13629 39750 13705
rect 0 13533 39936 13581
rect 186 13375 294 13485
rect 954 13375 1062 13485
rect 1434 13375 1542 13485
rect 2202 13375 2310 13485
rect 2682 13375 2790 13485
rect 3450 13375 3558 13485
rect 3930 13375 4038 13485
rect 4698 13375 4806 13485
rect 5178 13375 5286 13485
rect 5946 13375 6054 13485
rect 6426 13375 6534 13485
rect 7194 13375 7302 13485
rect 7674 13375 7782 13485
rect 8442 13375 8550 13485
rect 8922 13375 9030 13485
rect 9690 13375 9798 13485
rect 10170 13375 10278 13485
rect 10938 13375 11046 13485
rect 11418 13375 11526 13485
rect 12186 13375 12294 13485
rect 12666 13375 12774 13485
rect 13434 13375 13542 13485
rect 13914 13375 14022 13485
rect 14682 13375 14790 13485
rect 15162 13375 15270 13485
rect 15930 13375 16038 13485
rect 16410 13375 16518 13485
rect 17178 13375 17286 13485
rect 17658 13375 17766 13485
rect 18426 13375 18534 13485
rect 18906 13375 19014 13485
rect 19674 13375 19782 13485
rect 20154 13375 20262 13485
rect 20922 13375 21030 13485
rect 21402 13375 21510 13485
rect 22170 13375 22278 13485
rect 22650 13375 22758 13485
rect 23418 13375 23526 13485
rect 23898 13375 24006 13485
rect 24666 13375 24774 13485
rect 25146 13375 25254 13485
rect 25914 13375 26022 13485
rect 26394 13375 26502 13485
rect 27162 13375 27270 13485
rect 27642 13375 27750 13485
rect 28410 13375 28518 13485
rect 28890 13375 28998 13485
rect 29658 13375 29766 13485
rect 30138 13375 30246 13485
rect 30906 13375 31014 13485
rect 31386 13375 31494 13485
rect 32154 13375 32262 13485
rect 32634 13375 32742 13485
rect 33402 13375 33510 13485
rect 33882 13375 33990 13485
rect 34650 13375 34758 13485
rect 35130 13375 35238 13485
rect 35898 13375 36006 13485
rect 36378 13375 36486 13485
rect 37146 13375 37254 13485
rect 37626 13375 37734 13485
rect 38394 13375 38502 13485
rect 38874 13375 38982 13485
rect 39642 13375 39750 13485
rect 0 13279 39936 13327
rect 186 13155 294 13231
rect 954 13155 1062 13231
rect 1434 13155 1542 13231
rect 2202 13155 2310 13231
rect 2682 13155 2790 13231
rect 3450 13155 3558 13231
rect 3930 13155 4038 13231
rect 4698 13155 4806 13231
rect 5178 13155 5286 13231
rect 5946 13155 6054 13231
rect 6426 13155 6534 13231
rect 7194 13155 7302 13231
rect 7674 13155 7782 13231
rect 8442 13155 8550 13231
rect 8922 13155 9030 13231
rect 9690 13155 9798 13231
rect 10170 13155 10278 13231
rect 10938 13155 11046 13231
rect 11418 13155 11526 13231
rect 12186 13155 12294 13231
rect 12666 13155 12774 13231
rect 13434 13155 13542 13231
rect 13914 13155 14022 13231
rect 14682 13155 14790 13231
rect 15162 13155 15270 13231
rect 15930 13155 16038 13231
rect 16410 13155 16518 13231
rect 17178 13155 17286 13231
rect 17658 13155 17766 13231
rect 18426 13155 18534 13231
rect 18906 13155 19014 13231
rect 19674 13155 19782 13231
rect 20154 13155 20262 13231
rect 20922 13155 21030 13231
rect 21402 13155 21510 13231
rect 22170 13155 22278 13231
rect 22650 13155 22758 13231
rect 23418 13155 23526 13231
rect 23898 13155 24006 13231
rect 24666 13155 24774 13231
rect 25146 13155 25254 13231
rect 25914 13155 26022 13231
rect 26394 13155 26502 13231
rect 27162 13155 27270 13231
rect 27642 13155 27750 13231
rect 28410 13155 28518 13231
rect 28890 13155 28998 13231
rect 29658 13155 29766 13231
rect 30138 13155 30246 13231
rect 30906 13155 31014 13231
rect 31386 13155 31494 13231
rect 32154 13155 32262 13231
rect 32634 13155 32742 13231
rect 33402 13155 33510 13231
rect 33882 13155 33990 13231
rect 34650 13155 34758 13231
rect 35130 13155 35238 13231
rect 35898 13155 36006 13231
rect 36378 13155 36486 13231
rect 37146 13155 37254 13231
rect 37626 13155 37734 13231
rect 38394 13155 38502 13231
rect 38874 13155 38982 13231
rect 39642 13155 39750 13231
rect 0 13059 39936 13107
rect 0 12963 39936 13011
rect 186 12839 294 12915
rect 954 12839 1062 12915
rect 1434 12839 1542 12915
rect 2202 12839 2310 12915
rect 2682 12839 2790 12915
rect 3450 12839 3558 12915
rect 3930 12839 4038 12915
rect 4698 12839 4806 12915
rect 5178 12839 5286 12915
rect 5946 12839 6054 12915
rect 6426 12839 6534 12915
rect 7194 12839 7302 12915
rect 7674 12839 7782 12915
rect 8442 12839 8550 12915
rect 8922 12839 9030 12915
rect 9690 12839 9798 12915
rect 10170 12839 10278 12915
rect 10938 12839 11046 12915
rect 11418 12839 11526 12915
rect 12186 12839 12294 12915
rect 12666 12839 12774 12915
rect 13434 12839 13542 12915
rect 13914 12839 14022 12915
rect 14682 12839 14790 12915
rect 15162 12839 15270 12915
rect 15930 12839 16038 12915
rect 16410 12839 16518 12915
rect 17178 12839 17286 12915
rect 17658 12839 17766 12915
rect 18426 12839 18534 12915
rect 18906 12839 19014 12915
rect 19674 12839 19782 12915
rect 20154 12839 20262 12915
rect 20922 12839 21030 12915
rect 21402 12839 21510 12915
rect 22170 12839 22278 12915
rect 22650 12839 22758 12915
rect 23418 12839 23526 12915
rect 23898 12839 24006 12915
rect 24666 12839 24774 12915
rect 25146 12839 25254 12915
rect 25914 12839 26022 12915
rect 26394 12839 26502 12915
rect 27162 12839 27270 12915
rect 27642 12839 27750 12915
rect 28410 12839 28518 12915
rect 28890 12839 28998 12915
rect 29658 12839 29766 12915
rect 30138 12839 30246 12915
rect 30906 12839 31014 12915
rect 31386 12839 31494 12915
rect 32154 12839 32262 12915
rect 32634 12839 32742 12915
rect 33402 12839 33510 12915
rect 33882 12839 33990 12915
rect 34650 12839 34758 12915
rect 35130 12839 35238 12915
rect 35898 12839 36006 12915
rect 36378 12839 36486 12915
rect 37146 12839 37254 12915
rect 37626 12839 37734 12915
rect 38394 12839 38502 12915
rect 38874 12839 38982 12915
rect 39642 12839 39750 12915
rect 0 12743 39936 12791
rect 186 12585 294 12695
rect 954 12585 1062 12695
rect 1434 12585 1542 12695
rect 2202 12585 2310 12695
rect 2682 12585 2790 12695
rect 3450 12585 3558 12695
rect 3930 12585 4038 12695
rect 4698 12585 4806 12695
rect 5178 12585 5286 12695
rect 5946 12585 6054 12695
rect 6426 12585 6534 12695
rect 7194 12585 7302 12695
rect 7674 12585 7782 12695
rect 8442 12585 8550 12695
rect 8922 12585 9030 12695
rect 9690 12585 9798 12695
rect 10170 12585 10278 12695
rect 10938 12585 11046 12695
rect 11418 12585 11526 12695
rect 12186 12585 12294 12695
rect 12666 12585 12774 12695
rect 13434 12585 13542 12695
rect 13914 12585 14022 12695
rect 14682 12585 14790 12695
rect 15162 12585 15270 12695
rect 15930 12585 16038 12695
rect 16410 12585 16518 12695
rect 17178 12585 17286 12695
rect 17658 12585 17766 12695
rect 18426 12585 18534 12695
rect 18906 12585 19014 12695
rect 19674 12585 19782 12695
rect 20154 12585 20262 12695
rect 20922 12585 21030 12695
rect 21402 12585 21510 12695
rect 22170 12585 22278 12695
rect 22650 12585 22758 12695
rect 23418 12585 23526 12695
rect 23898 12585 24006 12695
rect 24666 12585 24774 12695
rect 25146 12585 25254 12695
rect 25914 12585 26022 12695
rect 26394 12585 26502 12695
rect 27162 12585 27270 12695
rect 27642 12585 27750 12695
rect 28410 12585 28518 12695
rect 28890 12585 28998 12695
rect 29658 12585 29766 12695
rect 30138 12585 30246 12695
rect 30906 12585 31014 12695
rect 31386 12585 31494 12695
rect 32154 12585 32262 12695
rect 32634 12585 32742 12695
rect 33402 12585 33510 12695
rect 33882 12585 33990 12695
rect 34650 12585 34758 12695
rect 35130 12585 35238 12695
rect 35898 12585 36006 12695
rect 36378 12585 36486 12695
rect 37146 12585 37254 12695
rect 37626 12585 37734 12695
rect 38394 12585 38502 12695
rect 38874 12585 38982 12695
rect 39642 12585 39750 12695
rect 0 12489 39936 12537
rect 186 12365 294 12441
rect 954 12365 1062 12441
rect 1434 12365 1542 12441
rect 2202 12365 2310 12441
rect 2682 12365 2790 12441
rect 3450 12365 3558 12441
rect 3930 12365 4038 12441
rect 4698 12365 4806 12441
rect 5178 12365 5286 12441
rect 5946 12365 6054 12441
rect 6426 12365 6534 12441
rect 7194 12365 7302 12441
rect 7674 12365 7782 12441
rect 8442 12365 8550 12441
rect 8922 12365 9030 12441
rect 9690 12365 9798 12441
rect 10170 12365 10278 12441
rect 10938 12365 11046 12441
rect 11418 12365 11526 12441
rect 12186 12365 12294 12441
rect 12666 12365 12774 12441
rect 13434 12365 13542 12441
rect 13914 12365 14022 12441
rect 14682 12365 14790 12441
rect 15162 12365 15270 12441
rect 15930 12365 16038 12441
rect 16410 12365 16518 12441
rect 17178 12365 17286 12441
rect 17658 12365 17766 12441
rect 18426 12365 18534 12441
rect 18906 12365 19014 12441
rect 19674 12365 19782 12441
rect 20154 12365 20262 12441
rect 20922 12365 21030 12441
rect 21402 12365 21510 12441
rect 22170 12365 22278 12441
rect 22650 12365 22758 12441
rect 23418 12365 23526 12441
rect 23898 12365 24006 12441
rect 24666 12365 24774 12441
rect 25146 12365 25254 12441
rect 25914 12365 26022 12441
rect 26394 12365 26502 12441
rect 27162 12365 27270 12441
rect 27642 12365 27750 12441
rect 28410 12365 28518 12441
rect 28890 12365 28998 12441
rect 29658 12365 29766 12441
rect 30138 12365 30246 12441
rect 30906 12365 31014 12441
rect 31386 12365 31494 12441
rect 32154 12365 32262 12441
rect 32634 12365 32742 12441
rect 33402 12365 33510 12441
rect 33882 12365 33990 12441
rect 34650 12365 34758 12441
rect 35130 12365 35238 12441
rect 35898 12365 36006 12441
rect 36378 12365 36486 12441
rect 37146 12365 37254 12441
rect 37626 12365 37734 12441
rect 38394 12365 38502 12441
rect 38874 12365 38982 12441
rect 39642 12365 39750 12441
rect 0 12269 39936 12317
rect 0 12173 39936 12221
rect 186 12049 294 12125
rect 954 12049 1062 12125
rect 1434 12049 1542 12125
rect 2202 12049 2310 12125
rect 2682 12049 2790 12125
rect 3450 12049 3558 12125
rect 3930 12049 4038 12125
rect 4698 12049 4806 12125
rect 5178 12049 5286 12125
rect 5946 12049 6054 12125
rect 6426 12049 6534 12125
rect 7194 12049 7302 12125
rect 7674 12049 7782 12125
rect 8442 12049 8550 12125
rect 8922 12049 9030 12125
rect 9690 12049 9798 12125
rect 10170 12049 10278 12125
rect 10938 12049 11046 12125
rect 11418 12049 11526 12125
rect 12186 12049 12294 12125
rect 12666 12049 12774 12125
rect 13434 12049 13542 12125
rect 13914 12049 14022 12125
rect 14682 12049 14790 12125
rect 15162 12049 15270 12125
rect 15930 12049 16038 12125
rect 16410 12049 16518 12125
rect 17178 12049 17286 12125
rect 17658 12049 17766 12125
rect 18426 12049 18534 12125
rect 18906 12049 19014 12125
rect 19674 12049 19782 12125
rect 20154 12049 20262 12125
rect 20922 12049 21030 12125
rect 21402 12049 21510 12125
rect 22170 12049 22278 12125
rect 22650 12049 22758 12125
rect 23418 12049 23526 12125
rect 23898 12049 24006 12125
rect 24666 12049 24774 12125
rect 25146 12049 25254 12125
rect 25914 12049 26022 12125
rect 26394 12049 26502 12125
rect 27162 12049 27270 12125
rect 27642 12049 27750 12125
rect 28410 12049 28518 12125
rect 28890 12049 28998 12125
rect 29658 12049 29766 12125
rect 30138 12049 30246 12125
rect 30906 12049 31014 12125
rect 31386 12049 31494 12125
rect 32154 12049 32262 12125
rect 32634 12049 32742 12125
rect 33402 12049 33510 12125
rect 33882 12049 33990 12125
rect 34650 12049 34758 12125
rect 35130 12049 35238 12125
rect 35898 12049 36006 12125
rect 36378 12049 36486 12125
rect 37146 12049 37254 12125
rect 37626 12049 37734 12125
rect 38394 12049 38502 12125
rect 38874 12049 38982 12125
rect 39642 12049 39750 12125
rect 0 11953 39936 12001
rect 186 11795 294 11905
rect 954 11795 1062 11905
rect 1434 11795 1542 11905
rect 2202 11795 2310 11905
rect 2682 11795 2790 11905
rect 3450 11795 3558 11905
rect 3930 11795 4038 11905
rect 4698 11795 4806 11905
rect 5178 11795 5286 11905
rect 5946 11795 6054 11905
rect 6426 11795 6534 11905
rect 7194 11795 7302 11905
rect 7674 11795 7782 11905
rect 8442 11795 8550 11905
rect 8922 11795 9030 11905
rect 9690 11795 9798 11905
rect 10170 11795 10278 11905
rect 10938 11795 11046 11905
rect 11418 11795 11526 11905
rect 12186 11795 12294 11905
rect 12666 11795 12774 11905
rect 13434 11795 13542 11905
rect 13914 11795 14022 11905
rect 14682 11795 14790 11905
rect 15162 11795 15270 11905
rect 15930 11795 16038 11905
rect 16410 11795 16518 11905
rect 17178 11795 17286 11905
rect 17658 11795 17766 11905
rect 18426 11795 18534 11905
rect 18906 11795 19014 11905
rect 19674 11795 19782 11905
rect 20154 11795 20262 11905
rect 20922 11795 21030 11905
rect 21402 11795 21510 11905
rect 22170 11795 22278 11905
rect 22650 11795 22758 11905
rect 23418 11795 23526 11905
rect 23898 11795 24006 11905
rect 24666 11795 24774 11905
rect 25146 11795 25254 11905
rect 25914 11795 26022 11905
rect 26394 11795 26502 11905
rect 27162 11795 27270 11905
rect 27642 11795 27750 11905
rect 28410 11795 28518 11905
rect 28890 11795 28998 11905
rect 29658 11795 29766 11905
rect 30138 11795 30246 11905
rect 30906 11795 31014 11905
rect 31386 11795 31494 11905
rect 32154 11795 32262 11905
rect 32634 11795 32742 11905
rect 33402 11795 33510 11905
rect 33882 11795 33990 11905
rect 34650 11795 34758 11905
rect 35130 11795 35238 11905
rect 35898 11795 36006 11905
rect 36378 11795 36486 11905
rect 37146 11795 37254 11905
rect 37626 11795 37734 11905
rect 38394 11795 38502 11905
rect 38874 11795 38982 11905
rect 39642 11795 39750 11905
rect 0 11699 39936 11747
rect 186 11575 294 11651
rect 954 11575 1062 11651
rect 1434 11575 1542 11651
rect 2202 11575 2310 11651
rect 2682 11575 2790 11651
rect 3450 11575 3558 11651
rect 3930 11575 4038 11651
rect 4698 11575 4806 11651
rect 5178 11575 5286 11651
rect 5946 11575 6054 11651
rect 6426 11575 6534 11651
rect 7194 11575 7302 11651
rect 7674 11575 7782 11651
rect 8442 11575 8550 11651
rect 8922 11575 9030 11651
rect 9690 11575 9798 11651
rect 10170 11575 10278 11651
rect 10938 11575 11046 11651
rect 11418 11575 11526 11651
rect 12186 11575 12294 11651
rect 12666 11575 12774 11651
rect 13434 11575 13542 11651
rect 13914 11575 14022 11651
rect 14682 11575 14790 11651
rect 15162 11575 15270 11651
rect 15930 11575 16038 11651
rect 16410 11575 16518 11651
rect 17178 11575 17286 11651
rect 17658 11575 17766 11651
rect 18426 11575 18534 11651
rect 18906 11575 19014 11651
rect 19674 11575 19782 11651
rect 20154 11575 20262 11651
rect 20922 11575 21030 11651
rect 21402 11575 21510 11651
rect 22170 11575 22278 11651
rect 22650 11575 22758 11651
rect 23418 11575 23526 11651
rect 23898 11575 24006 11651
rect 24666 11575 24774 11651
rect 25146 11575 25254 11651
rect 25914 11575 26022 11651
rect 26394 11575 26502 11651
rect 27162 11575 27270 11651
rect 27642 11575 27750 11651
rect 28410 11575 28518 11651
rect 28890 11575 28998 11651
rect 29658 11575 29766 11651
rect 30138 11575 30246 11651
rect 30906 11575 31014 11651
rect 31386 11575 31494 11651
rect 32154 11575 32262 11651
rect 32634 11575 32742 11651
rect 33402 11575 33510 11651
rect 33882 11575 33990 11651
rect 34650 11575 34758 11651
rect 35130 11575 35238 11651
rect 35898 11575 36006 11651
rect 36378 11575 36486 11651
rect 37146 11575 37254 11651
rect 37626 11575 37734 11651
rect 38394 11575 38502 11651
rect 38874 11575 38982 11651
rect 39642 11575 39750 11651
rect 0 11479 39936 11527
rect 0 11383 39936 11431
rect 186 11259 294 11335
rect 954 11259 1062 11335
rect 1434 11259 1542 11335
rect 2202 11259 2310 11335
rect 2682 11259 2790 11335
rect 3450 11259 3558 11335
rect 3930 11259 4038 11335
rect 4698 11259 4806 11335
rect 5178 11259 5286 11335
rect 5946 11259 6054 11335
rect 6426 11259 6534 11335
rect 7194 11259 7302 11335
rect 7674 11259 7782 11335
rect 8442 11259 8550 11335
rect 8922 11259 9030 11335
rect 9690 11259 9798 11335
rect 10170 11259 10278 11335
rect 10938 11259 11046 11335
rect 11418 11259 11526 11335
rect 12186 11259 12294 11335
rect 12666 11259 12774 11335
rect 13434 11259 13542 11335
rect 13914 11259 14022 11335
rect 14682 11259 14790 11335
rect 15162 11259 15270 11335
rect 15930 11259 16038 11335
rect 16410 11259 16518 11335
rect 17178 11259 17286 11335
rect 17658 11259 17766 11335
rect 18426 11259 18534 11335
rect 18906 11259 19014 11335
rect 19674 11259 19782 11335
rect 20154 11259 20262 11335
rect 20922 11259 21030 11335
rect 21402 11259 21510 11335
rect 22170 11259 22278 11335
rect 22650 11259 22758 11335
rect 23418 11259 23526 11335
rect 23898 11259 24006 11335
rect 24666 11259 24774 11335
rect 25146 11259 25254 11335
rect 25914 11259 26022 11335
rect 26394 11259 26502 11335
rect 27162 11259 27270 11335
rect 27642 11259 27750 11335
rect 28410 11259 28518 11335
rect 28890 11259 28998 11335
rect 29658 11259 29766 11335
rect 30138 11259 30246 11335
rect 30906 11259 31014 11335
rect 31386 11259 31494 11335
rect 32154 11259 32262 11335
rect 32634 11259 32742 11335
rect 33402 11259 33510 11335
rect 33882 11259 33990 11335
rect 34650 11259 34758 11335
rect 35130 11259 35238 11335
rect 35898 11259 36006 11335
rect 36378 11259 36486 11335
rect 37146 11259 37254 11335
rect 37626 11259 37734 11335
rect 38394 11259 38502 11335
rect 38874 11259 38982 11335
rect 39642 11259 39750 11335
rect 0 11163 39936 11211
rect 186 11005 294 11115
rect 954 11005 1062 11115
rect 1434 11005 1542 11115
rect 2202 11005 2310 11115
rect 2682 11005 2790 11115
rect 3450 11005 3558 11115
rect 3930 11005 4038 11115
rect 4698 11005 4806 11115
rect 5178 11005 5286 11115
rect 5946 11005 6054 11115
rect 6426 11005 6534 11115
rect 7194 11005 7302 11115
rect 7674 11005 7782 11115
rect 8442 11005 8550 11115
rect 8922 11005 9030 11115
rect 9690 11005 9798 11115
rect 10170 11005 10278 11115
rect 10938 11005 11046 11115
rect 11418 11005 11526 11115
rect 12186 11005 12294 11115
rect 12666 11005 12774 11115
rect 13434 11005 13542 11115
rect 13914 11005 14022 11115
rect 14682 11005 14790 11115
rect 15162 11005 15270 11115
rect 15930 11005 16038 11115
rect 16410 11005 16518 11115
rect 17178 11005 17286 11115
rect 17658 11005 17766 11115
rect 18426 11005 18534 11115
rect 18906 11005 19014 11115
rect 19674 11005 19782 11115
rect 20154 11005 20262 11115
rect 20922 11005 21030 11115
rect 21402 11005 21510 11115
rect 22170 11005 22278 11115
rect 22650 11005 22758 11115
rect 23418 11005 23526 11115
rect 23898 11005 24006 11115
rect 24666 11005 24774 11115
rect 25146 11005 25254 11115
rect 25914 11005 26022 11115
rect 26394 11005 26502 11115
rect 27162 11005 27270 11115
rect 27642 11005 27750 11115
rect 28410 11005 28518 11115
rect 28890 11005 28998 11115
rect 29658 11005 29766 11115
rect 30138 11005 30246 11115
rect 30906 11005 31014 11115
rect 31386 11005 31494 11115
rect 32154 11005 32262 11115
rect 32634 11005 32742 11115
rect 33402 11005 33510 11115
rect 33882 11005 33990 11115
rect 34650 11005 34758 11115
rect 35130 11005 35238 11115
rect 35898 11005 36006 11115
rect 36378 11005 36486 11115
rect 37146 11005 37254 11115
rect 37626 11005 37734 11115
rect 38394 11005 38502 11115
rect 38874 11005 38982 11115
rect 39642 11005 39750 11115
rect 0 10909 39936 10957
rect 186 10785 294 10861
rect 954 10785 1062 10861
rect 1434 10785 1542 10861
rect 2202 10785 2310 10861
rect 2682 10785 2790 10861
rect 3450 10785 3558 10861
rect 3930 10785 4038 10861
rect 4698 10785 4806 10861
rect 5178 10785 5286 10861
rect 5946 10785 6054 10861
rect 6426 10785 6534 10861
rect 7194 10785 7302 10861
rect 7674 10785 7782 10861
rect 8442 10785 8550 10861
rect 8922 10785 9030 10861
rect 9690 10785 9798 10861
rect 10170 10785 10278 10861
rect 10938 10785 11046 10861
rect 11418 10785 11526 10861
rect 12186 10785 12294 10861
rect 12666 10785 12774 10861
rect 13434 10785 13542 10861
rect 13914 10785 14022 10861
rect 14682 10785 14790 10861
rect 15162 10785 15270 10861
rect 15930 10785 16038 10861
rect 16410 10785 16518 10861
rect 17178 10785 17286 10861
rect 17658 10785 17766 10861
rect 18426 10785 18534 10861
rect 18906 10785 19014 10861
rect 19674 10785 19782 10861
rect 20154 10785 20262 10861
rect 20922 10785 21030 10861
rect 21402 10785 21510 10861
rect 22170 10785 22278 10861
rect 22650 10785 22758 10861
rect 23418 10785 23526 10861
rect 23898 10785 24006 10861
rect 24666 10785 24774 10861
rect 25146 10785 25254 10861
rect 25914 10785 26022 10861
rect 26394 10785 26502 10861
rect 27162 10785 27270 10861
rect 27642 10785 27750 10861
rect 28410 10785 28518 10861
rect 28890 10785 28998 10861
rect 29658 10785 29766 10861
rect 30138 10785 30246 10861
rect 30906 10785 31014 10861
rect 31386 10785 31494 10861
rect 32154 10785 32262 10861
rect 32634 10785 32742 10861
rect 33402 10785 33510 10861
rect 33882 10785 33990 10861
rect 34650 10785 34758 10861
rect 35130 10785 35238 10861
rect 35898 10785 36006 10861
rect 36378 10785 36486 10861
rect 37146 10785 37254 10861
rect 37626 10785 37734 10861
rect 38394 10785 38502 10861
rect 38874 10785 38982 10861
rect 39642 10785 39750 10861
rect 0 10689 39936 10737
rect 0 10593 39936 10641
rect 186 10469 294 10545
rect 954 10469 1062 10545
rect 1434 10469 1542 10545
rect 2202 10469 2310 10545
rect 2682 10469 2790 10545
rect 3450 10469 3558 10545
rect 3930 10469 4038 10545
rect 4698 10469 4806 10545
rect 5178 10469 5286 10545
rect 5946 10469 6054 10545
rect 6426 10469 6534 10545
rect 7194 10469 7302 10545
rect 7674 10469 7782 10545
rect 8442 10469 8550 10545
rect 8922 10469 9030 10545
rect 9690 10469 9798 10545
rect 10170 10469 10278 10545
rect 10938 10469 11046 10545
rect 11418 10469 11526 10545
rect 12186 10469 12294 10545
rect 12666 10469 12774 10545
rect 13434 10469 13542 10545
rect 13914 10469 14022 10545
rect 14682 10469 14790 10545
rect 15162 10469 15270 10545
rect 15930 10469 16038 10545
rect 16410 10469 16518 10545
rect 17178 10469 17286 10545
rect 17658 10469 17766 10545
rect 18426 10469 18534 10545
rect 18906 10469 19014 10545
rect 19674 10469 19782 10545
rect 20154 10469 20262 10545
rect 20922 10469 21030 10545
rect 21402 10469 21510 10545
rect 22170 10469 22278 10545
rect 22650 10469 22758 10545
rect 23418 10469 23526 10545
rect 23898 10469 24006 10545
rect 24666 10469 24774 10545
rect 25146 10469 25254 10545
rect 25914 10469 26022 10545
rect 26394 10469 26502 10545
rect 27162 10469 27270 10545
rect 27642 10469 27750 10545
rect 28410 10469 28518 10545
rect 28890 10469 28998 10545
rect 29658 10469 29766 10545
rect 30138 10469 30246 10545
rect 30906 10469 31014 10545
rect 31386 10469 31494 10545
rect 32154 10469 32262 10545
rect 32634 10469 32742 10545
rect 33402 10469 33510 10545
rect 33882 10469 33990 10545
rect 34650 10469 34758 10545
rect 35130 10469 35238 10545
rect 35898 10469 36006 10545
rect 36378 10469 36486 10545
rect 37146 10469 37254 10545
rect 37626 10469 37734 10545
rect 38394 10469 38502 10545
rect 38874 10469 38982 10545
rect 39642 10469 39750 10545
rect 0 10373 39936 10421
rect 186 10215 294 10325
rect 954 10215 1062 10325
rect 1434 10215 1542 10325
rect 2202 10215 2310 10325
rect 2682 10215 2790 10325
rect 3450 10215 3558 10325
rect 3930 10215 4038 10325
rect 4698 10215 4806 10325
rect 5178 10215 5286 10325
rect 5946 10215 6054 10325
rect 6426 10215 6534 10325
rect 7194 10215 7302 10325
rect 7674 10215 7782 10325
rect 8442 10215 8550 10325
rect 8922 10215 9030 10325
rect 9690 10215 9798 10325
rect 10170 10215 10278 10325
rect 10938 10215 11046 10325
rect 11418 10215 11526 10325
rect 12186 10215 12294 10325
rect 12666 10215 12774 10325
rect 13434 10215 13542 10325
rect 13914 10215 14022 10325
rect 14682 10215 14790 10325
rect 15162 10215 15270 10325
rect 15930 10215 16038 10325
rect 16410 10215 16518 10325
rect 17178 10215 17286 10325
rect 17658 10215 17766 10325
rect 18426 10215 18534 10325
rect 18906 10215 19014 10325
rect 19674 10215 19782 10325
rect 20154 10215 20262 10325
rect 20922 10215 21030 10325
rect 21402 10215 21510 10325
rect 22170 10215 22278 10325
rect 22650 10215 22758 10325
rect 23418 10215 23526 10325
rect 23898 10215 24006 10325
rect 24666 10215 24774 10325
rect 25146 10215 25254 10325
rect 25914 10215 26022 10325
rect 26394 10215 26502 10325
rect 27162 10215 27270 10325
rect 27642 10215 27750 10325
rect 28410 10215 28518 10325
rect 28890 10215 28998 10325
rect 29658 10215 29766 10325
rect 30138 10215 30246 10325
rect 30906 10215 31014 10325
rect 31386 10215 31494 10325
rect 32154 10215 32262 10325
rect 32634 10215 32742 10325
rect 33402 10215 33510 10325
rect 33882 10215 33990 10325
rect 34650 10215 34758 10325
rect 35130 10215 35238 10325
rect 35898 10215 36006 10325
rect 36378 10215 36486 10325
rect 37146 10215 37254 10325
rect 37626 10215 37734 10325
rect 38394 10215 38502 10325
rect 38874 10215 38982 10325
rect 39642 10215 39750 10325
rect 0 10119 39936 10167
rect 186 9995 294 10071
rect 954 9995 1062 10071
rect 1434 9995 1542 10071
rect 2202 9995 2310 10071
rect 2682 9995 2790 10071
rect 3450 9995 3558 10071
rect 3930 9995 4038 10071
rect 4698 9995 4806 10071
rect 5178 9995 5286 10071
rect 5946 9995 6054 10071
rect 6426 9995 6534 10071
rect 7194 9995 7302 10071
rect 7674 9995 7782 10071
rect 8442 9995 8550 10071
rect 8922 9995 9030 10071
rect 9690 9995 9798 10071
rect 10170 9995 10278 10071
rect 10938 9995 11046 10071
rect 11418 9995 11526 10071
rect 12186 9995 12294 10071
rect 12666 9995 12774 10071
rect 13434 9995 13542 10071
rect 13914 9995 14022 10071
rect 14682 9995 14790 10071
rect 15162 9995 15270 10071
rect 15930 9995 16038 10071
rect 16410 9995 16518 10071
rect 17178 9995 17286 10071
rect 17658 9995 17766 10071
rect 18426 9995 18534 10071
rect 18906 9995 19014 10071
rect 19674 9995 19782 10071
rect 20154 9995 20262 10071
rect 20922 9995 21030 10071
rect 21402 9995 21510 10071
rect 22170 9995 22278 10071
rect 22650 9995 22758 10071
rect 23418 9995 23526 10071
rect 23898 9995 24006 10071
rect 24666 9995 24774 10071
rect 25146 9995 25254 10071
rect 25914 9995 26022 10071
rect 26394 9995 26502 10071
rect 27162 9995 27270 10071
rect 27642 9995 27750 10071
rect 28410 9995 28518 10071
rect 28890 9995 28998 10071
rect 29658 9995 29766 10071
rect 30138 9995 30246 10071
rect 30906 9995 31014 10071
rect 31386 9995 31494 10071
rect 32154 9995 32262 10071
rect 32634 9995 32742 10071
rect 33402 9995 33510 10071
rect 33882 9995 33990 10071
rect 34650 9995 34758 10071
rect 35130 9995 35238 10071
rect 35898 9995 36006 10071
rect 36378 9995 36486 10071
rect 37146 9995 37254 10071
rect 37626 9995 37734 10071
rect 38394 9995 38502 10071
rect 38874 9995 38982 10071
rect 39642 9995 39750 10071
rect 0 9899 39936 9947
rect 0 9803 39936 9851
rect 186 9679 294 9755
rect 954 9679 1062 9755
rect 1434 9679 1542 9755
rect 2202 9679 2310 9755
rect 2682 9679 2790 9755
rect 3450 9679 3558 9755
rect 3930 9679 4038 9755
rect 4698 9679 4806 9755
rect 5178 9679 5286 9755
rect 5946 9679 6054 9755
rect 6426 9679 6534 9755
rect 7194 9679 7302 9755
rect 7674 9679 7782 9755
rect 8442 9679 8550 9755
rect 8922 9679 9030 9755
rect 9690 9679 9798 9755
rect 10170 9679 10278 9755
rect 10938 9679 11046 9755
rect 11418 9679 11526 9755
rect 12186 9679 12294 9755
rect 12666 9679 12774 9755
rect 13434 9679 13542 9755
rect 13914 9679 14022 9755
rect 14682 9679 14790 9755
rect 15162 9679 15270 9755
rect 15930 9679 16038 9755
rect 16410 9679 16518 9755
rect 17178 9679 17286 9755
rect 17658 9679 17766 9755
rect 18426 9679 18534 9755
rect 18906 9679 19014 9755
rect 19674 9679 19782 9755
rect 20154 9679 20262 9755
rect 20922 9679 21030 9755
rect 21402 9679 21510 9755
rect 22170 9679 22278 9755
rect 22650 9679 22758 9755
rect 23418 9679 23526 9755
rect 23898 9679 24006 9755
rect 24666 9679 24774 9755
rect 25146 9679 25254 9755
rect 25914 9679 26022 9755
rect 26394 9679 26502 9755
rect 27162 9679 27270 9755
rect 27642 9679 27750 9755
rect 28410 9679 28518 9755
rect 28890 9679 28998 9755
rect 29658 9679 29766 9755
rect 30138 9679 30246 9755
rect 30906 9679 31014 9755
rect 31386 9679 31494 9755
rect 32154 9679 32262 9755
rect 32634 9679 32742 9755
rect 33402 9679 33510 9755
rect 33882 9679 33990 9755
rect 34650 9679 34758 9755
rect 35130 9679 35238 9755
rect 35898 9679 36006 9755
rect 36378 9679 36486 9755
rect 37146 9679 37254 9755
rect 37626 9679 37734 9755
rect 38394 9679 38502 9755
rect 38874 9679 38982 9755
rect 39642 9679 39750 9755
rect 0 9583 39936 9631
rect 186 9425 294 9535
rect 954 9425 1062 9535
rect 1434 9425 1542 9535
rect 2202 9425 2310 9535
rect 2682 9425 2790 9535
rect 3450 9425 3558 9535
rect 3930 9425 4038 9535
rect 4698 9425 4806 9535
rect 5178 9425 5286 9535
rect 5946 9425 6054 9535
rect 6426 9425 6534 9535
rect 7194 9425 7302 9535
rect 7674 9425 7782 9535
rect 8442 9425 8550 9535
rect 8922 9425 9030 9535
rect 9690 9425 9798 9535
rect 10170 9425 10278 9535
rect 10938 9425 11046 9535
rect 11418 9425 11526 9535
rect 12186 9425 12294 9535
rect 12666 9425 12774 9535
rect 13434 9425 13542 9535
rect 13914 9425 14022 9535
rect 14682 9425 14790 9535
rect 15162 9425 15270 9535
rect 15930 9425 16038 9535
rect 16410 9425 16518 9535
rect 17178 9425 17286 9535
rect 17658 9425 17766 9535
rect 18426 9425 18534 9535
rect 18906 9425 19014 9535
rect 19674 9425 19782 9535
rect 20154 9425 20262 9535
rect 20922 9425 21030 9535
rect 21402 9425 21510 9535
rect 22170 9425 22278 9535
rect 22650 9425 22758 9535
rect 23418 9425 23526 9535
rect 23898 9425 24006 9535
rect 24666 9425 24774 9535
rect 25146 9425 25254 9535
rect 25914 9425 26022 9535
rect 26394 9425 26502 9535
rect 27162 9425 27270 9535
rect 27642 9425 27750 9535
rect 28410 9425 28518 9535
rect 28890 9425 28998 9535
rect 29658 9425 29766 9535
rect 30138 9425 30246 9535
rect 30906 9425 31014 9535
rect 31386 9425 31494 9535
rect 32154 9425 32262 9535
rect 32634 9425 32742 9535
rect 33402 9425 33510 9535
rect 33882 9425 33990 9535
rect 34650 9425 34758 9535
rect 35130 9425 35238 9535
rect 35898 9425 36006 9535
rect 36378 9425 36486 9535
rect 37146 9425 37254 9535
rect 37626 9425 37734 9535
rect 38394 9425 38502 9535
rect 38874 9425 38982 9535
rect 39642 9425 39750 9535
rect 0 9329 39936 9377
rect 186 9205 294 9281
rect 954 9205 1062 9281
rect 1434 9205 1542 9281
rect 2202 9205 2310 9281
rect 2682 9205 2790 9281
rect 3450 9205 3558 9281
rect 3930 9205 4038 9281
rect 4698 9205 4806 9281
rect 5178 9205 5286 9281
rect 5946 9205 6054 9281
rect 6426 9205 6534 9281
rect 7194 9205 7302 9281
rect 7674 9205 7782 9281
rect 8442 9205 8550 9281
rect 8922 9205 9030 9281
rect 9690 9205 9798 9281
rect 10170 9205 10278 9281
rect 10938 9205 11046 9281
rect 11418 9205 11526 9281
rect 12186 9205 12294 9281
rect 12666 9205 12774 9281
rect 13434 9205 13542 9281
rect 13914 9205 14022 9281
rect 14682 9205 14790 9281
rect 15162 9205 15270 9281
rect 15930 9205 16038 9281
rect 16410 9205 16518 9281
rect 17178 9205 17286 9281
rect 17658 9205 17766 9281
rect 18426 9205 18534 9281
rect 18906 9205 19014 9281
rect 19674 9205 19782 9281
rect 20154 9205 20262 9281
rect 20922 9205 21030 9281
rect 21402 9205 21510 9281
rect 22170 9205 22278 9281
rect 22650 9205 22758 9281
rect 23418 9205 23526 9281
rect 23898 9205 24006 9281
rect 24666 9205 24774 9281
rect 25146 9205 25254 9281
rect 25914 9205 26022 9281
rect 26394 9205 26502 9281
rect 27162 9205 27270 9281
rect 27642 9205 27750 9281
rect 28410 9205 28518 9281
rect 28890 9205 28998 9281
rect 29658 9205 29766 9281
rect 30138 9205 30246 9281
rect 30906 9205 31014 9281
rect 31386 9205 31494 9281
rect 32154 9205 32262 9281
rect 32634 9205 32742 9281
rect 33402 9205 33510 9281
rect 33882 9205 33990 9281
rect 34650 9205 34758 9281
rect 35130 9205 35238 9281
rect 35898 9205 36006 9281
rect 36378 9205 36486 9281
rect 37146 9205 37254 9281
rect 37626 9205 37734 9281
rect 38394 9205 38502 9281
rect 38874 9205 38982 9281
rect 39642 9205 39750 9281
rect 0 9109 39936 9157
rect 0 9013 39936 9061
rect 186 8889 294 8965
rect 954 8889 1062 8965
rect 1434 8889 1542 8965
rect 2202 8889 2310 8965
rect 2682 8889 2790 8965
rect 3450 8889 3558 8965
rect 3930 8889 4038 8965
rect 4698 8889 4806 8965
rect 5178 8889 5286 8965
rect 5946 8889 6054 8965
rect 6426 8889 6534 8965
rect 7194 8889 7302 8965
rect 7674 8889 7782 8965
rect 8442 8889 8550 8965
rect 8922 8889 9030 8965
rect 9690 8889 9798 8965
rect 10170 8889 10278 8965
rect 10938 8889 11046 8965
rect 11418 8889 11526 8965
rect 12186 8889 12294 8965
rect 12666 8889 12774 8965
rect 13434 8889 13542 8965
rect 13914 8889 14022 8965
rect 14682 8889 14790 8965
rect 15162 8889 15270 8965
rect 15930 8889 16038 8965
rect 16410 8889 16518 8965
rect 17178 8889 17286 8965
rect 17658 8889 17766 8965
rect 18426 8889 18534 8965
rect 18906 8889 19014 8965
rect 19674 8889 19782 8965
rect 20154 8889 20262 8965
rect 20922 8889 21030 8965
rect 21402 8889 21510 8965
rect 22170 8889 22278 8965
rect 22650 8889 22758 8965
rect 23418 8889 23526 8965
rect 23898 8889 24006 8965
rect 24666 8889 24774 8965
rect 25146 8889 25254 8965
rect 25914 8889 26022 8965
rect 26394 8889 26502 8965
rect 27162 8889 27270 8965
rect 27642 8889 27750 8965
rect 28410 8889 28518 8965
rect 28890 8889 28998 8965
rect 29658 8889 29766 8965
rect 30138 8889 30246 8965
rect 30906 8889 31014 8965
rect 31386 8889 31494 8965
rect 32154 8889 32262 8965
rect 32634 8889 32742 8965
rect 33402 8889 33510 8965
rect 33882 8889 33990 8965
rect 34650 8889 34758 8965
rect 35130 8889 35238 8965
rect 35898 8889 36006 8965
rect 36378 8889 36486 8965
rect 37146 8889 37254 8965
rect 37626 8889 37734 8965
rect 38394 8889 38502 8965
rect 38874 8889 38982 8965
rect 39642 8889 39750 8965
rect 0 8793 39936 8841
rect 186 8635 294 8745
rect 954 8635 1062 8745
rect 1434 8635 1542 8745
rect 2202 8635 2310 8745
rect 2682 8635 2790 8745
rect 3450 8635 3558 8745
rect 3930 8635 4038 8745
rect 4698 8635 4806 8745
rect 5178 8635 5286 8745
rect 5946 8635 6054 8745
rect 6426 8635 6534 8745
rect 7194 8635 7302 8745
rect 7674 8635 7782 8745
rect 8442 8635 8550 8745
rect 8922 8635 9030 8745
rect 9690 8635 9798 8745
rect 10170 8635 10278 8745
rect 10938 8635 11046 8745
rect 11418 8635 11526 8745
rect 12186 8635 12294 8745
rect 12666 8635 12774 8745
rect 13434 8635 13542 8745
rect 13914 8635 14022 8745
rect 14682 8635 14790 8745
rect 15162 8635 15270 8745
rect 15930 8635 16038 8745
rect 16410 8635 16518 8745
rect 17178 8635 17286 8745
rect 17658 8635 17766 8745
rect 18426 8635 18534 8745
rect 18906 8635 19014 8745
rect 19674 8635 19782 8745
rect 20154 8635 20262 8745
rect 20922 8635 21030 8745
rect 21402 8635 21510 8745
rect 22170 8635 22278 8745
rect 22650 8635 22758 8745
rect 23418 8635 23526 8745
rect 23898 8635 24006 8745
rect 24666 8635 24774 8745
rect 25146 8635 25254 8745
rect 25914 8635 26022 8745
rect 26394 8635 26502 8745
rect 27162 8635 27270 8745
rect 27642 8635 27750 8745
rect 28410 8635 28518 8745
rect 28890 8635 28998 8745
rect 29658 8635 29766 8745
rect 30138 8635 30246 8745
rect 30906 8635 31014 8745
rect 31386 8635 31494 8745
rect 32154 8635 32262 8745
rect 32634 8635 32742 8745
rect 33402 8635 33510 8745
rect 33882 8635 33990 8745
rect 34650 8635 34758 8745
rect 35130 8635 35238 8745
rect 35898 8635 36006 8745
rect 36378 8635 36486 8745
rect 37146 8635 37254 8745
rect 37626 8635 37734 8745
rect 38394 8635 38502 8745
rect 38874 8635 38982 8745
rect 39642 8635 39750 8745
rect 0 8539 39936 8587
rect 186 8415 294 8491
rect 954 8415 1062 8491
rect 1434 8415 1542 8491
rect 2202 8415 2310 8491
rect 2682 8415 2790 8491
rect 3450 8415 3558 8491
rect 3930 8415 4038 8491
rect 4698 8415 4806 8491
rect 5178 8415 5286 8491
rect 5946 8415 6054 8491
rect 6426 8415 6534 8491
rect 7194 8415 7302 8491
rect 7674 8415 7782 8491
rect 8442 8415 8550 8491
rect 8922 8415 9030 8491
rect 9690 8415 9798 8491
rect 10170 8415 10278 8491
rect 10938 8415 11046 8491
rect 11418 8415 11526 8491
rect 12186 8415 12294 8491
rect 12666 8415 12774 8491
rect 13434 8415 13542 8491
rect 13914 8415 14022 8491
rect 14682 8415 14790 8491
rect 15162 8415 15270 8491
rect 15930 8415 16038 8491
rect 16410 8415 16518 8491
rect 17178 8415 17286 8491
rect 17658 8415 17766 8491
rect 18426 8415 18534 8491
rect 18906 8415 19014 8491
rect 19674 8415 19782 8491
rect 20154 8415 20262 8491
rect 20922 8415 21030 8491
rect 21402 8415 21510 8491
rect 22170 8415 22278 8491
rect 22650 8415 22758 8491
rect 23418 8415 23526 8491
rect 23898 8415 24006 8491
rect 24666 8415 24774 8491
rect 25146 8415 25254 8491
rect 25914 8415 26022 8491
rect 26394 8415 26502 8491
rect 27162 8415 27270 8491
rect 27642 8415 27750 8491
rect 28410 8415 28518 8491
rect 28890 8415 28998 8491
rect 29658 8415 29766 8491
rect 30138 8415 30246 8491
rect 30906 8415 31014 8491
rect 31386 8415 31494 8491
rect 32154 8415 32262 8491
rect 32634 8415 32742 8491
rect 33402 8415 33510 8491
rect 33882 8415 33990 8491
rect 34650 8415 34758 8491
rect 35130 8415 35238 8491
rect 35898 8415 36006 8491
rect 36378 8415 36486 8491
rect 37146 8415 37254 8491
rect 37626 8415 37734 8491
rect 38394 8415 38502 8491
rect 38874 8415 38982 8491
rect 39642 8415 39750 8491
rect 0 8319 39936 8367
rect 0 8223 39936 8271
rect 186 8099 294 8175
rect 954 8099 1062 8175
rect 1434 8099 1542 8175
rect 2202 8099 2310 8175
rect 2682 8099 2790 8175
rect 3450 8099 3558 8175
rect 3930 8099 4038 8175
rect 4698 8099 4806 8175
rect 5178 8099 5286 8175
rect 5946 8099 6054 8175
rect 6426 8099 6534 8175
rect 7194 8099 7302 8175
rect 7674 8099 7782 8175
rect 8442 8099 8550 8175
rect 8922 8099 9030 8175
rect 9690 8099 9798 8175
rect 10170 8099 10278 8175
rect 10938 8099 11046 8175
rect 11418 8099 11526 8175
rect 12186 8099 12294 8175
rect 12666 8099 12774 8175
rect 13434 8099 13542 8175
rect 13914 8099 14022 8175
rect 14682 8099 14790 8175
rect 15162 8099 15270 8175
rect 15930 8099 16038 8175
rect 16410 8099 16518 8175
rect 17178 8099 17286 8175
rect 17658 8099 17766 8175
rect 18426 8099 18534 8175
rect 18906 8099 19014 8175
rect 19674 8099 19782 8175
rect 20154 8099 20262 8175
rect 20922 8099 21030 8175
rect 21402 8099 21510 8175
rect 22170 8099 22278 8175
rect 22650 8099 22758 8175
rect 23418 8099 23526 8175
rect 23898 8099 24006 8175
rect 24666 8099 24774 8175
rect 25146 8099 25254 8175
rect 25914 8099 26022 8175
rect 26394 8099 26502 8175
rect 27162 8099 27270 8175
rect 27642 8099 27750 8175
rect 28410 8099 28518 8175
rect 28890 8099 28998 8175
rect 29658 8099 29766 8175
rect 30138 8099 30246 8175
rect 30906 8099 31014 8175
rect 31386 8099 31494 8175
rect 32154 8099 32262 8175
rect 32634 8099 32742 8175
rect 33402 8099 33510 8175
rect 33882 8099 33990 8175
rect 34650 8099 34758 8175
rect 35130 8099 35238 8175
rect 35898 8099 36006 8175
rect 36378 8099 36486 8175
rect 37146 8099 37254 8175
rect 37626 8099 37734 8175
rect 38394 8099 38502 8175
rect 38874 8099 38982 8175
rect 39642 8099 39750 8175
rect 0 8003 39936 8051
rect 186 7845 294 7955
rect 954 7845 1062 7955
rect 1434 7845 1542 7955
rect 2202 7845 2310 7955
rect 2682 7845 2790 7955
rect 3450 7845 3558 7955
rect 3930 7845 4038 7955
rect 4698 7845 4806 7955
rect 5178 7845 5286 7955
rect 5946 7845 6054 7955
rect 6426 7845 6534 7955
rect 7194 7845 7302 7955
rect 7674 7845 7782 7955
rect 8442 7845 8550 7955
rect 8922 7845 9030 7955
rect 9690 7845 9798 7955
rect 10170 7845 10278 7955
rect 10938 7845 11046 7955
rect 11418 7845 11526 7955
rect 12186 7845 12294 7955
rect 12666 7845 12774 7955
rect 13434 7845 13542 7955
rect 13914 7845 14022 7955
rect 14682 7845 14790 7955
rect 15162 7845 15270 7955
rect 15930 7845 16038 7955
rect 16410 7845 16518 7955
rect 17178 7845 17286 7955
rect 17658 7845 17766 7955
rect 18426 7845 18534 7955
rect 18906 7845 19014 7955
rect 19674 7845 19782 7955
rect 20154 7845 20262 7955
rect 20922 7845 21030 7955
rect 21402 7845 21510 7955
rect 22170 7845 22278 7955
rect 22650 7845 22758 7955
rect 23418 7845 23526 7955
rect 23898 7845 24006 7955
rect 24666 7845 24774 7955
rect 25146 7845 25254 7955
rect 25914 7845 26022 7955
rect 26394 7845 26502 7955
rect 27162 7845 27270 7955
rect 27642 7845 27750 7955
rect 28410 7845 28518 7955
rect 28890 7845 28998 7955
rect 29658 7845 29766 7955
rect 30138 7845 30246 7955
rect 30906 7845 31014 7955
rect 31386 7845 31494 7955
rect 32154 7845 32262 7955
rect 32634 7845 32742 7955
rect 33402 7845 33510 7955
rect 33882 7845 33990 7955
rect 34650 7845 34758 7955
rect 35130 7845 35238 7955
rect 35898 7845 36006 7955
rect 36378 7845 36486 7955
rect 37146 7845 37254 7955
rect 37626 7845 37734 7955
rect 38394 7845 38502 7955
rect 38874 7845 38982 7955
rect 39642 7845 39750 7955
rect 0 7749 39936 7797
rect 186 7625 294 7701
rect 954 7625 1062 7701
rect 1434 7625 1542 7701
rect 2202 7625 2310 7701
rect 2682 7625 2790 7701
rect 3450 7625 3558 7701
rect 3930 7625 4038 7701
rect 4698 7625 4806 7701
rect 5178 7625 5286 7701
rect 5946 7625 6054 7701
rect 6426 7625 6534 7701
rect 7194 7625 7302 7701
rect 7674 7625 7782 7701
rect 8442 7625 8550 7701
rect 8922 7625 9030 7701
rect 9690 7625 9798 7701
rect 10170 7625 10278 7701
rect 10938 7625 11046 7701
rect 11418 7625 11526 7701
rect 12186 7625 12294 7701
rect 12666 7625 12774 7701
rect 13434 7625 13542 7701
rect 13914 7625 14022 7701
rect 14682 7625 14790 7701
rect 15162 7625 15270 7701
rect 15930 7625 16038 7701
rect 16410 7625 16518 7701
rect 17178 7625 17286 7701
rect 17658 7625 17766 7701
rect 18426 7625 18534 7701
rect 18906 7625 19014 7701
rect 19674 7625 19782 7701
rect 20154 7625 20262 7701
rect 20922 7625 21030 7701
rect 21402 7625 21510 7701
rect 22170 7625 22278 7701
rect 22650 7625 22758 7701
rect 23418 7625 23526 7701
rect 23898 7625 24006 7701
rect 24666 7625 24774 7701
rect 25146 7625 25254 7701
rect 25914 7625 26022 7701
rect 26394 7625 26502 7701
rect 27162 7625 27270 7701
rect 27642 7625 27750 7701
rect 28410 7625 28518 7701
rect 28890 7625 28998 7701
rect 29658 7625 29766 7701
rect 30138 7625 30246 7701
rect 30906 7625 31014 7701
rect 31386 7625 31494 7701
rect 32154 7625 32262 7701
rect 32634 7625 32742 7701
rect 33402 7625 33510 7701
rect 33882 7625 33990 7701
rect 34650 7625 34758 7701
rect 35130 7625 35238 7701
rect 35898 7625 36006 7701
rect 36378 7625 36486 7701
rect 37146 7625 37254 7701
rect 37626 7625 37734 7701
rect 38394 7625 38502 7701
rect 38874 7625 38982 7701
rect 39642 7625 39750 7701
rect 0 7529 39936 7577
rect 0 7433 39936 7481
rect 186 7309 294 7385
rect 954 7309 1062 7385
rect 1434 7309 1542 7385
rect 2202 7309 2310 7385
rect 2682 7309 2790 7385
rect 3450 7309 3558 7385
rect 3930 7309 4038 7385
rect 4698 7309 4806 7385
rect 5178 7309 5286 7385
rect 5946 7309 6054 7385
rect 6426 7309 6534 7385
rect 7194 7309 7302 7385
rect 7674 7309 7782 7385
rect 8442 7309 8550 7385
rect 8922 7309 9030 7385
rect 9690 7309 9798 7385
rect 10170 7309 10278 7385
rect 10938 7309 11046 7385
rect 11418 7309 11526 7385
rect 12186 7309 12294 7385
rect 12666 7309 12774 7385
rect 13434 7309 13542 7385
rect 13914 7309 14022 7385
rect 14682 7309 14790 7385
rect 15162 7309 15270 7385
rect 15930 7309 16038 7385
rect 16410 7309 16518 7385
rect 17178 7309 17286 7385
rect 17658 7309 17766 7385
rect 18426 7309 18534 7385
rect 18906 7309 19014 7385
rect 19674 7309 19782 7385
rect 20154 7309 20262 7385
rect 20922 7309 21030 7385
rect 21402 7309 21510 7385
rect 22170 7309 22278 7385
rect 22650 7309 22758 7385
rect 23418 7309 23526 7385
rect 23898 7309 24006 7385
rect 24666 7309 24774 7385
rect 25146 7309 25254 7385
rect 25914 7309 26022 7385
rect 26394 7309 26502 7385
rect 27162 7309 27270 7385
rect 27642 7309 27750 7385
rect 28410 7309 28518 7385
rect 28890 7309 28998 7385
rect 29658 7309 29766 7385
rect 30138 7309 30246 7385
rect 30906 7309 31014 7385
rect 31386 7309 31494 7385
rect 32154 7309 32262 7385
rect 32634 7309 32742 7385
rect 33402 7309 33510 7385
rect 33882 7309 33990 7385
rect 34650 7309 34758 7385
rect 35130 7309 35238 7385
rect 35898 7309 36006 7385
rect 36378 7309 36486 7385
rect 37146 7309 37254 7385
rect 37626 7309 37734 7385
rect 38394 7309 38502 7385
rect 38874 7309 38982 7385
rect 39642 7309 39750 7385
rect 0 7213 39936 7261
rect 186 7055 294 7165
rect 954 7055 1062 7165
rect 1434 7055 1542 7165
rect 2202 7055 2310 7165
rect 2682 7055 2790 7165
rect 3450 7055 3558 7165
rect 3930 7055 4038 7165
rect 4698 7055 4806 7165
rect 5178 7055 5286 7165
rect 5946 7055 6054 7165
rect 6426 7055 6534 7165
rect 7194 7055 7302 7165
rect 7674 7055 7782 7165
rect 8442 7055 8550 7165
rect 8922 7055 9030 7165
rect 9690 7055 9798 7165
rect 10170 7055 10278 7165
rect 10938 7055 11046 7165
rect 11418 7055 11526 7165
rect 12186 7055 12294 7165
rect 12666 7055 12774 7165
rect 13434 7055 13542 7165
rect 13914 7055 14022 7165
rect 14682 7055 14790 7165
rect 15162 7055 15270 7165
rect 15930 7055 16038 7165
rect 16410 7055 16518 7165
rect 17178 7055 17286 7165
rect 17658 7055 17766 7165
rect 18426 7055 18534 7165
rect 18906 7055 19014 7165
rect 19674 7055 19782 7165
rect 20154 7055 20262 7165
rect 20922 7055 21030 7165
rect 21402 7055 21510 7165
rect 22170 7055 22278 7165
rect 22650 7055 22758 7165
rect 23418 7055 23526 7165
rect 23898 7055 24006 7165
rect 24666 7055 24774 7165
rect 25146 7055 25254 7165
rect 25914 7055 26022 7165
rect 26394 7055 26502 7165
rect 27162 7055 27270 7165
rect 27642 7055 27750 7165
rect 28410 7055 28518 7165
rect 28890 7055 28998 7165
rect 29658 7055 29766 7165
rect 30138 7055 30246 7165
rect 30906 7055 31014 7165
rect 31386 7055 31494 7165
rect 32154 7055 32262 7165
rect 32634 7055 32742 7165
rect 33402 7055 33510 7165
rect 33882 7055 33990 7165
rect 34650 7055 34758 7165
rect 35130 7055 35238 7165
rect 35898 7055 36006 7165
rect 36378 7055 36486 7165
rect 37146 7055 37254 7165
rect 37626 7055 37734 7165
rect 38394 7055 38502 7165
rect 38874 7055 38982 7165
rect 39642 7055 39750 7165
rect 0 6959 39936 7007
rect 186 6835 294 6911
rect 954 6835 1062 6911
rect 1434 6835 1542 6911
rect 2202 6835 2310 6911
rect 2682 6835 2790 6911
rect 3450 6835 3558 6911
rect 3930 6835 4038 6911
rect 4698 6835 4806 6911
rect 5178 6835 5286 6911
rect 5946 6835 6054 6911
rect 6426 6835 6534 6911
rect 7194 6835 7302 6911
rect 7674 6835 7782 6911
rect 8442 6835 8550 6911
rect 8922 6835 9030 6911
rect 9690 6835 9798 6911
rect 10170 6835 10278 6911
rect 10938 6835 11046 6911
rect 11418 6835 11526 6911
rect 12186 6835 12294 6911
rect 12666 6835 12774 6911
rect 13434 6835 13542 6911
rect 13914 6835 14022 6911
rect 14682 6835 14790 6911
rect 15162 6835 15270 6911
rect 15930 6835 16038 6911
rect 16410 6835 16518 6911
rect 17178 6835 17286 6911
rect 17658 6835 17766 6911
rect 18426 6835 18534 6911
rect 18906 6835 19014 6911
rect 19674 6835 19782 6911
rect 20154 6835 20262 6911
rect 20922 6835 21030 6911
rect 21402 6835 21510 6911
rect 22170 6835 22278 6911
rect 22650 6835 22758 6911
rect 23418 6835 23526 6911
rect 23898 6835 24006 6911
rect 24666 6835 24774 6911
rect 25146 6835 25254 6911
rect 25914 6835 26022 6911
rect 26394 6835 26502 6911
rect 27162 6835 27270 6911
rect 27642 6835 27750 6911
rect 28410 6835 28518 6911
rect 28890 6835 28998 6911
rect 29658 6835 29766 6911
rect 30138 6835 30246 6911
rect 30906 6835 31014 6911
rect 31386 6835 31494 6911
rect 32154 6835 32262 6911
rect 32634 6835 32742 6911
rect 33402 6835 33510 6911
rect 33882 6835 33990 6911
rect 34650 6835 34758 6911
rect 35130 6835 35238 6911
rect 35898 6835 36006 6911
rect 36378 6835 36486 6911
rect 37146 6835 37254 6911
rect 37626 6835 37734 6911
rect 38394 6835 38502 6911
rect 38874 6835 38982 6911
rect 39642 6835 39750 6911
rect 0 6739 39936 6787
rect 0 6643 39936 6691
rect 186 6519 294 6595
rect 954 6519 1062 6595
rect 1434 6519 1542 6595
rect 2202 6519 2310 6595
rect 2682 6519 2790 6595
rect 3450 6519 3558 6595
rect 3930 6519 4038 6595
rect 4698 6519 4806 6595
rect 5178 6519 5286 6595
rect 5946 6519 6054 6595
rect 6426 6519 6534 6595
rect 7194 6519 7302 6595
rect 7674 6519 7782 6595
rect 8442 6519 8550 6595
rect 8922 6519 9030 6595
rect 9690 6519 9798 6595
rect 10170 6519 10278 6595
rect 10938 6519 11046 6595
rect 11418 6519 11526 6595
rect 12186 6519 12294 6595
rect 12666 6519 12774 6595
rect 13434 6519 13542 6595
rect 13914 6519 14022 6595
rect 14682 6519 14790 6595
rect 15162 6519 15270 6595
rect 15930 6519 16038 6595
rect 16410 6519 16518 6595
rect 17178 6519 17286 6595
rect 17658 6519 17766 6595
rect 18426 6519 18534 6595
rect 18906 6519 19014 6595
rect 19674 6519 19782 6595
rect 20154 6519 20262 6595
rect 20922 6519 21030 6595
rect 21402 6519 21510 6595
rect 22170 6519 22278 6595
rect 22650 6519 22758 6595
rect 23418 6519 23526 6595
rect 23898 6519 24006 6595
rect 24666 6519 24774 6595
rect 25146 6519 25254 6595
rect 25914 6519 26022 6595
rect 26394 6519 26502 6595
rect 27162 6519 27270 6595
rect 27642 6519 27750 6595
rect 28410 6519 28518 6595
rect 28890 6519 28998 6595
rect 29658 6519 29766 6595
rect 30138 6519 30246 6595
rect 30906 6519 31014 6595
rect 31386 6519 31494 6595
rect 32154 6519 32262 6595
rect 32634 6519 32742 6595
rect 33402 6519 33510 6595
rect 33882 6519 33990 6595
rect 34650 6519 34758 6595
rect 35130 6519 35238 6595
rect 35898 6519 36006 6595
rect 36378 6519 36486 6595
rect 37146 6519 37254 6595
rect 37626 6519 37734 6595
rect 38394 6519 38502 6595
rect 38874 6519 38982 6595
rect 39642 6519 39750 6595
rect 0 6423 39936 6471
rect 186 6265 294 6375
rect 954 6265 1062 6375
rect 1434 6265 1542 6375
rect 2202 6265 2310 6375
rect 2682 6265 2790 6375
rect 3450 6265 3558 6375
rect 3930 6265 4038 6375
rect 4698 6265 4806 6375
rect 5178 6265 5286 6375
rect 5946 6265 6054 6375
rect 6426 6265 6534 6375
rect 7194 6265 7302 6375
rect 7674 6265 7782 6375
rect 8442 6265 8550 6375
rect 8922 6265 9030 6375
rect 9690 6265 9798 6375
rect 10170 6265 10278 6375
rect 10938 6265 11046 6375
rect 11418 6265 11526 6375
rect 12186 6265 12294 6375
rect 12666 6265 12774 6375
rect 13434 6265 13542 6375
rect 13914 6265 14022 6375
rect 14682 6265 14790 6375
rect 15162 6265 15270 6375
rect 15930 6265 16038 6375
rect 16410 6265 16518 6375
rect 17178 6265 17286 6375
rect 17658 6265 17766 6375
rect 18426 6265 18534 6375
rect 18906 6265 19014 6375
rect 19674 6265 19782 6375
rect 20154 6265 20262 6375
rect 20922 6265 21030 6375
rect 21402 6265 21510 6375
rect 22170 6265 22278 6375
rect 22650 6265 22758 6375
rect 23418 6265 23526 6375
rect 23898 6265 24006 6375
rect 24666 6265 24774 6375
rect 25146 6265 25254 6375
rect 25914 6265 26022 6375
rect 26394 6265 26502 6375
rect 27162 6265 27270 6375
rect 27642 6265 27750 6375
rect 28410 6265 28518 6375
rect 28890 6265 28998 6375
rect 29658 6265 29766 6375
rect 30138 6265 30246 6375
rect 30906 6265 31014 6375
rect 31386 6265 31494 6375
rect 32154 6265 32262 6375
rect 32634 6265 32742 6375
rect 33402 6265 33510 6375
rect 33882 6265 33990 6375
rect 34650 6265 34758 6375
rect 35130 6265 35238 6375
rect 35898 6265 36006 6375
rect 36378 6265 36486 6375
rect 37146 6265 37254 6375
rect 37626 6265 37734 6375
rect 38394 6265 38502 6375
rect 38874 6265 38982 6375
rect 39642 6265 39750 6375
rect 0 6169 39936 6217
rect 186 6045 294 6121
rect 954 6045 1062 6121
rect 1434 6045 1542 6121
rect 2202 6045 2310 6121
rect 2682 6045 2790 6121
rect 3450 6045 3558 6121
rect 3930 6045 4038 6121
rect 4698 6045 4806 6121
rect 5178 6045 5286 6121
rect 5946 6045 6054 6121
rect 6426 6045 6534 6121
rect 7194 6045 7302 6121
rect 7674 6045 7782 6121
rect 8442 6045 8550 6121
rect 8922 6045 9030 6121
rect 9690 6045 9798 6121
rect 10170 6045 10278 6121
rect 10938 6045 11046 6121
rect 11418 6045 11526 6121
rect 12186 6045 12294 6121
rect 12666 6045 12774 6121
rect 13434 6045 13542 6121
rect 13914 6045 14022 6121
rect 14682 6045 14790 6121
rect 15162 6045 15270 6121
rect 15930 6045 16038 6121
rect 16410 6045 16518 6121
rect 17178 6045 17286 6121
rect 17658 6045 17766 6121
rect 18426 6045 18534 6121
rect 18906 6045 19014 6121
rect 19674 6045 19782 6121
rect 20154 6045 20262 6121
rect 20922 6045 21030 6121
rect 21402 6045 21510 6121
rect 22170 6045 22278 6121
rect 22650 6045 22758 6121
rect 23418 6045 23526 6121
rect 23898 6045 24006 6121
rect 24666 6045 24774 6121
rect 25146 6045 25254 6121
rect 25914 6045 26022 6121
rect 26394 6045 26502 6121
rect 27162 6045 27270 6121
rect 27642 6045 27750 6121
rect 28410 6045 28518 6121
rect 28890 6045 28998 6121
rect 29658 6045 29766 6121
rect 30138 6045 30246 6121
rect 30906 6045 31014 6121
rect 31386 6045 31494 6121
rect 32154 6045 32262 6121
rect 32634 6045 32742 6121
rect 33402 6045 33510 6121
rect 33882 6045 33990 6121
rect 34650 6045 34758 6121
rect 35130 6045 35238 6121
rect 35898 6045 36006 6121
rect 36378 6045 36486 6121
rect 37146 6045 37254 6121
rect 37626 6045 37734 6121
rect 38394 6045 38502 6121
rect 38874 6045 38982 6121
rect 39642 6045 39750 6121
rect 0 5949 39936 5997
rect 0 5853 39936 5901
rect 186 5729 294 5805
rect 954 5729 1062 5805
rect 1434 5729 1542 5805
rect 2202 5729 2310 5805
rect 2682 5729 2790 5805
rect 3450 5729 3558 5805
rect 3930 5729 4038 5805
rect 4698 5729 4806 5805
rect 5178 5729 5286 5805
rect 5946 5729 6054 5805
rect 6426 5729 6534 5805
rect 7194 5729 7302 5805
rect 7674 5729 7782 5805
rect 8442 5729 8550 5805
rect 8922 5729 9030 5805
rect 9690 5729 9798 5805
rect 10170 5729 10278 5805
rect 10938 5729 11046 5805
rect 11418 5729 11526 5805
rect 12186 5729 12294 5805
rect 12666 5729 12774 5805
rect 13434 5729 13542 5805
rect 13914 5729 14022 5805
rect 14682 5729 14790 5805
rect 15162 5729 15270 5805
rect 15930 5729 16038 5805
rect 16410 5729 16518 5805
rect 17178 5729 17286 5805
rect 17658 5729 17766 5805
rect 18426 5729 18534 5805
rect 18906 5729 19014 5805
rect 19674 5729 19782 5805
rect 20154 5729 20262 5805
rect 20922 5729 21030 5805
rect 21402 5729 21510 5805
rect 22170 5729 22278 5805
rect 22650 5729 22758 5805
rect 23418 5729 23526 5805
rect 23898 5729 24006 5805
rect 24666 5729 24774 5805
rect 25146 5729 25254 5805
rect 25914 5729 26022 5805
rect 26394 5729 26502 5805
rect 27162 5729 27270 5805
rect 27642 5729 27750 5805
rect 28410 5729 28518 5805
rect 28890 5729 28998 5805
rect 29658 5729 29766 5805
rect 30138 5729 30246 5805
rect 30906 5729 31014 5805
rect 31386 5729 31494 5805
rect 32154 5729 32262 5805
rect 32634 5729 32742 5805
rect 33402 5729 33510 5805
rect 33882 5729 33990 5805
rect 34650 5729 34758 5805
rect 35130 5729 35238 5805
rect 35898 5729 36006 5805
rect 36378 5729 36486 5805
rect 37146 5729 37254 5805
rect 37626 5729 37734 5805
rect 38394 5729 38502 5805
rect 38874 5729 38982 5805
rect 39642 5729 39750 5805
rect 0 5633 39936 5681
rect 186 5475 294 5585
rect 954 5475 1062 5585
rect 1434 5475 1542 5585
rect 2202 5475 2310 5585
rect 2682 5475 2790 5585
rect 3450 5475 3558 5585
rect 3930 5475 4038 5585
rect 4698 5475 4806 5585
rect 5178 5475 5286 5585
rect 5946 5475 6054 5585
rect 6426 5475 6534 5585
rect 7194 5475 7302 5585
rect 7674 5475 7782 5585
rect 8442 5475 8550 5585
rect 8922 5475 9030 5585
rect 9690 5475 9798 5585
rect 10170 5475 10278 5585
rect 10938 5475 11046 5585
rect 11418 5475 11526 5585
rect 12186 5475 12294 5585
rect 12666 5475 12774 5585
rect 13434 5475 13542 5585
rect 13914 5475 14022 5585
rect 14682 5475 14790 5585
rect 15162 5475 15270 5585
rect 15930 5475 16038 5585
rect 16410 5475 16518 5585
rect 17178 5475 17286 5585
rect 17658 5475 17766 5585
rect 18426 5475 18534 5585
rect 18906 5475 19014 5585
rect 19674 5475 19782 5585
rect 20154 5475 20262 5585
rect 20922 5475 21030 5585
rect 21402 5475 21510 5585
rect 22170 5475 22278 5585
rect 22650 5475 22758 5585
rect 23418 5475 23526 5585
rect 23898 5475 24006 5585
rect 24666 5475 24774 5585
rect 25146 5475 25254 5585
rect 25914 5475 26022 5585
rect 26394 5475 26502 5585
rect 27162 5475 27270 5585
rect 27642 5475 27750 5585
rect 28410 5475 28518 5585
rect 28890 5475 28998 5585
rect 29658 5475 29766 5585
rect 30138 5475 30246 5585
rect 30906 5475 31014 5585
rect 31386 5475 31494 5585
rect 32154 5475 32262 5585
rect 32634 5475 32742 5585
rect 33402 5475 33510 5585
rect 33882 5475 33990 5585
rect 34650 5475 34758 5585
rect 35130 5475 35238 5585
rect 35898 5475 36006 5585
rect 36378 5475 36486 5585
rect 37146 5475 37254 5585
rect 37626 5475 37734 5585
rect 38394 5475 38502 5585
rect 38874 5475 38982 5585
rect 39642 5475 39750 5585
rect 0 5379 39936 5427
rect 186 5255 294 5331
rect 954 5255 1062 5331
rect 1434 5255 1542 5331
rect 2202 5255 2310 5331
rect 2682 5255 2790 5331
rect 3450 5255 3558 5331
rect 3930 5255 4038 5331
rect 4698 5255 4806 5331
rect 5178 5255 5286 5331
rect 5946 5255 6054 5331
rect 6426 5255 6534 5331
rect 7194 5255 7302 5331
rect 7674 5255 7782 5331
rect 8442 5255 8550 5331
rect 8922 5255 9030 5331
rect 9690 5255 9798 5331
rect 10170 5255 10278 5331
rect 10938 5255 11046 5331
rect 11418 5255 11526 5331
rect 12186 5255 12294 5331
rect 12666 5255 12774 5331
rect 13434 5255 13542 5331
rect 13914 5255 14022 5331
rect 14682 5255 14790 5331
rect 15162 5255 15270 5331
rect 15930 5255 16038 5331
rect 16410 5255 16518 5331
rect 17178 5255 17286 5331
rect 17658 5255 17766 5331
rect 18426 5255 18534 5331
rect 18906 5255 19014 5331
rect 19674 5255 19782 5331
rect 20154 5255 20262 5331
rect 20922 5255 21030 5331
rect 21402 5255 21510 5331
rect 22170 5255 22278 5331
rect 22650 5255 22758 5331
rect 23418 5255 23526 5331
rect 23898 5255 24006 5331
rect 24666 5255 24774 5331
rect 25146 5255 25254 5331
rect 25914 5255 26022 5331
rect 26394 5255 26502 5331
rect 27162 5255 27270 5331
rect 27642 5255 27750 5331
rect 28410 5255 28518 5331
rect 28890 5255 28998 5331
rect 29658 5255 29766 5331
rect 30138 5255 30246 5331
rect 30906 5255 31014 5331
rect 31386 5255 31494 5331
rect 32154 5255 32262 5331
rect 32634 5255 32742 5331
rect 33402 5255 33510 5331
rect 33882 5255 33990 5331
rect 34650 5255 34758 5331
rect 35130 5255 35238 5331
rect 35898 5255 36006 5331
rect 36378 5255 36486 5331
rect 37146 5255 37254 5331
rect 37626 5255 37734 5331
rect 38394 5255 38502 5331
rect 38874 5255 38982 5331
rect 39642 5255 39750 5331
rect 0 5159 39936 5207
rect 0 5063 39936 5111
rect 186 4939 294 5015
rect 954 4939 1062 5015
rect 1434 4939 1542 5015
rect 2202 4939 2310 5015
rect 2682 4939 2790 5015
rect 3450 4939 3558 5015
rect 3930 4939 4038 5015
rect 4698 4939 4806 5015
rect 5178 4939 5286 5015
rect 5946 4939 6054 5015
rect 6426 4939 6534 5015
rect 7194 4939 7302 5015
rect 7674 4939 7782 5015
rect 8442 4939 8550 5015
rect 8922 4939 9030 5015
rect 9690 4939 9798 5015
rect 10170 4939 10278 5015
rect 10938 4939 11046 5015
rect 11418 4939 11526 5015
rect 12186 4939 12294 5015
rect 12666 4939 12774 5015
rect 13434 4939 13542 5015
rect 13914 4939 14022 5015
rect 14682 4939 14790 5015
rect 15162 4939 15270 5015
rect 15930 4939 16038 5015
rect 16410 4939 16518 5015
rect 17178 4939 17286 5015
rect 17658 4939 17766 5015
rect 18426 4939 18534 5015
rect 18906 4939 19014 5015
rect 19674 4939 19782 5015
rect 20154 4939 20262 5015
rect 20922 4939 21030 5015
rect 21402 4939 21510 5015
rect 22170 4939 22278 5015
rect 22650 4939 22758 5015
rect 23418 4939 23526 5015
rect 23898 4939 24006 5015
rect 24666 4939 24774 5015
rect 25146 4939 25254 5015
rect 25914 4939 26022 5015
rect 26394 4939 26502 5015
rect 27162 4939 27270 5015
rect 27642 4939 27750 5015
rect 28410 4939 28518 5015
rect 28890 4939 28998 5015
rect 29658 4939 29766 5015
rect 30138 4939 30246 5015
rect 30906 4939 31014 5015
rect 31386 4939 31494 5015
rect 32154 4939 32262 5015
rect 32634 4939 32742 5015
rect 33402 4939 33510 5015
rect 33882 4939 33990 5015
rect 34650 4939 34758 5015
rect 35130 4939 35238 5015
rect 35898 4939 36006 5015
rect 36378 4939 36486 5015
rect 37146 4939 37254 5015
rect 37626 4939 37734 5015
rect 38394 4939 38502 5015
rect 38874 4939 38982 5015
rect 39642 4939 39750 5015
rect 0 4843 39936 4891
rect 186 4685 294 4795
rect 954 4685 1062 4795
rect 1434 4685 1542 4795
rect 2202 4685 2310 4795
rect 2682 4685 2790 4795
rect 3450 4685 3558 4795
rect 3930 4685 4038 4795
rect 4698 4685 4806 4795
rect 5178 4685 5286 4795
rect 5946 4685 6054 4795
rect 6426 4685 6534 4795
rect 7194 4685 7302 4795
rect 7674 4685 7782 4795
rect 8442 4685 8550 4795
rect 8922 4685 9030 4795
rect 9690 4685 9798 4795
rect 10170 4685 10278 4795
rect 10938 4685 11046 4795
rect 11418 4685 11526 4795
rect 12186 4685 12294 4795
rect 12666 4685 12774 4795
rect 13434 4685 13542 4795
rect 13914 4685 14022 4795
rect 14682 4685 14790 4795
rect 15162 4685 15270 4795
rect 15930 4685 16038 4795
rect 16410 4685 16518 4795
rect 17178 4685 17286 4795
rect 17658 4685 17766 4795
rect 18426 4685 18534 4795
rect 18906 4685 19014 4795
rect 19674 4685 19782 4795
rect 20154 4685 20262 4795
rect 20922 4685 21030 4795
rect 21402 4685 21510 4795
rect 22170 4685 22278 4795
rect 22650 4685 22758 4795
rect 23418 4685 23526 4795
rect 23898 4685 24006 4795
rect 24666 4685 24774 4795
rect 25146 4685 25254 4795
rect 25914 4685 26022 4795
rect 26394 4685 26502 4795
rect 27162 4685 27270 4795
rect 27642 4685 27750 4795
rect 28410 4685 28518 4795
rect 28890 4685 28998 4795
rect 29658 4685 29766 4795
rect 30138 4685 30246 4795
rect 30906 4685 31014 4795
rect 31386 4685 31494 4795
rect 32154 4685 32262 4795
rect 32634 4685 32742 4795
rect 33402 4685 33510 4795
rect 33882 4685 33990 4795
rect 34650 4685 34758 4795
rect 35130 4685 35238 4795
rect 35898 4685 36006 4795
rect 36378 4685 36486 4795
rect 37146 4685 37254 4795
rect 37626 4685 37734 4795
rect 38394 4685 38502 4795
rect 38874 4685 38982 4795
rect 39642 4685 39750 4795
rect 0 4589 39936 4637
rect 186 4465 294 4541
rect 954 4465 1062 4541
rect 1434 4465 1542 4541
rect 2202 4465 2310 4541
rect 2682 4465 2790 4541
rect 3450 4465 3558 4541
rect 3930 4465 4038 4541
rect 4698 4465 4806 4541
rect 5178 4465 5286 4541
rect 5946 4465 6054 4541
rect 6426 4465 6534 4541
rect 7194 4465 7302 4541
rect 7674 4465 7782 4541
rect 8442 4465 8550 4541
rect 8922 4465 9030 4541
rect 9690 4465 9798 4541
rect 10170 4465 10278 4541
rect 10938 4465 11046 4541
rect 11418 4465 11526 4541
rect 12186 4465 12294 4541
rect 12666 4465 12774 4541
rect 13434 4465 13542 4541
rect 13914 4465 14022 4541
rect 14682 4465 14790 4541
rect 15162 4465 15270 4541
rect 15930 4465 16038 4541
rect 16410 4465 16518 4541
rect 17178 4465 17286 4541
rect 17658 4465 17766 4541
rect 18426 4465 18534 4541
rect 18906 4465 19014 4541
rect 19674 4465 19782 4541
rect 20154 4465 20262 4541
rect 20922 4465 21030 4541
rect 21402 4465 21510 4541
rect 22170 4465 22278 4541
rect 22650 4465 22758 4541
rect 23418 4465 23526 4541
rect 23898 4465 24006 4541
rect 24666 4465 24774 4541
rect 25146 4465 25254 4541
rect 25914 4465 26022 4541
rect 26394 4465 26502 4541
rect 27162 4465 27270 4541
rect 27642 4465 27750 4541
rect 28410 4465 28518 4541
rect 28890 4465 28998 4541
rect 29658 4465 29766 4541
rect 30138 4465 30246 4541
rect 30906 4465 31014 4541
rect 31386 4465 31494 4541
rect 32154 4465 32262 4541
rect 32634 4465 32742 4541
rect 33402 4465 33510 4541
rect 33882 4465 33990 4541
rect 34650 4465 34758 4541
rect 35130 4465 35238 4541
rect 35898 4465 36006 4541
rect 36378 4465 36486 4541
rect 37146 4465 37254 4541
rect 37626 4465 37734 4541
rect 38394 4465 38502 4541
rect 38874 4465 38982 4541
rect 39642 4465 39750 4541
rect 0 4369 39936 4417
rect 0 4273 39936 4321
rect 186 4149 294 4225
rect 954 4149 1062 4225
rect 1434 4149 1542 4225
rect 2202 4149 2310 4225
rect 2682 4149 2790 4225
rect 3450 4149 3558 4225
rect 3930 4149 4038 4225
rect 4698 4149 4806 4225
rect 5178 4149 5286 4225
rect 5946 4149 6054 4225
rect 6426 4149 6534 4225
rect 7194 4149 7302 4225
rect 7674 4149 7782 4225
rect 8442 4149 8550 4225
rect 8922 4149 9030 4225
rect 9690 4149 9798 4225
rect 10170 4149 10278 4225
rect 10938 4149 11046 4225
rect 11418 4149 11526 4225
rect 12186 4149 12294 4225
rect 12666 4149 12774 4225
rect 13434 4149 13542 4225
rect 13914 4149 14022 4225
rect 14682 4149 14790 4225
rect 15162 4149 15270 4225
rect 15930 4149 16038 4225
rect 16410 4149 16518 4225
rect 17178 4149 17286 4225
rect 17658 4149 17766 4225
rect 18426 4149 18534 4225
rect 18906 4149 19014 4225
rect 19674 4149 19782 4225
rect 20154 4149 20262 4225
rect 20922 4149 21030 4225
rect 21402 4149 21510 4225
rect 22170 4149 22278 4225
rect 22650 4149 22758 4225
rect 23418 4149 23526 4225
rect 23898 4149 24006 4225
rect 24666 4149 24774 4225
rect 25146 4149 25254 4225
rect 25914 4149 26022 4225
rect 26394 4149 26502 4225
rect 27162 4149 27270 4225
rect 27642 4149 27750 4225
rect 28410 4149 28518 4225
rect 28890 4149 28998 4225
rect 29658 4149 29766 4225
rect 30138 4149 30246 4225
rect 30906 4149 31014 4225
rect 31386 4149 31494 4225
rect 32154 4149 32262 4225
rect 32634 4149 32742 4225
rect 33402 4149 33510 4225
rect 33882 4149 33990 4225
rect 34650 4149 34758 4225
rect 35130 4149 35238 4225
rect 35898 4149 36006 4225
rect 36378 4149 36486 4225
rect 37146 4149 37254 4225
rect 37626 4149 37734 4225
rect 38394 4149 38502 4225
rect 38874 4149 38982 4225
rect 39642 4149 39750 4225
rect 0 4053 39936 4101
rect 186 3895 294 4005
rect 954 3895 1062 4005
rect 1434 3895 1542 4005
rect 2202 3895 2310 4005
rect 2682 3895 2790 4005
rect 3450 3895 3558 4005
rect 3930 3895 4038 4005
rect 4698 3895 4806 4005
rect 5178 3895 5286 4005
rect 5946 3895 6054 4005
rect 6426 3895 6534 4005
rect 7194 3895 7302 4005
rect 7674 3895 7782 4005
rect 8442 3895 8550 4005
rect 8922 3895 9030 4005
rect 9690 3895 9798 4005
rect 10170 3895 10278 4005
rect 10938 3895 11046 4005
rect 11418 3895 11526 4005
rect 12186 3895 12294 4005
rect 12666 3895 12774 4005
rect 13434 3895 13542 4005
rect 13914 3895 14022 4005
rect 14682 3895 14790 4005
rect 15162 3895 15270 4005
rect 15930 3895 16038 4005
rect 16410 3895 16518 4005
rect 17178 3895 17286 4005
rect 17658 3895 17766 4005
rect 18426 3895 18534 4005
rect 18906 3895 19014 4005
rect 19674 3895 19782 4005
rect 20154 3895 20262 4005
rect 20922 3895 21030 4005
rect 21402 3895 21510 4005
rect 22170 3895 22278 4005
rect 22650 3895 22758 4005
rect 23418 3895 23526 4005
rect 23898 3895 24006 4005
rect 24666 3895 24774 4005
rect 25146 3895 25254 4005
rect 25914 3895 26022 4005
rect 26394 3895 26502 4005
rect 27162 3895 27270 4005
rect 27642 3895 27750 4005
rect 28410 3895 28518 4005
rect 28890 3895 28998 4005
rect 29658 3895 29766 4005
rect 30138 3895 30246 4005
rect 30906 3895 31014 4005
rect 31386 3895 31494 4005
rect 32154 3895 32262 4005
rect 32634 3895 32742 4005
rect 33402 3895 33510 4005
rect 33882 3895 33990 4005
rect 34650 3895 34758 4005
rect 35130 3895 35238 4005
rect 35898 3895 36006 4005
rect 36378 3895 36486 4005
rect 37146 3895 37254 4005
rect 37626 3895 37734 4005
rect 38394 3895 38502 4005
rect 38874 3895 38982 4005
rect 39642 3895 39750 4005
rect 0 3799 39936 3847
rect 186 3675 294 3751
rect 954 3675 1062 3751
rect 1434 3675 1542 3751
rect 2202 3675 2310 3751
rect 2682 3675 2790 3751
rect 3450 3675 3558 3751
rect 3930 3675 4038 3751
rect 4698 3675 4806 3751
rect 5178 3675 5286 3751
rect 5946 3675 6054 3751
rect 6426 3675 6534 3751
rect 7194 3675 7302 3751
rect 7674 3675 7782 3751
rect 8442 3675 8550 3751
rect 8922 3675 9030 3751
rect 9690 3675 9798 3751
rect 10170 3675 10278 3751
rect 10938 3675 11046 3751
rect 11418 3675 11526 3751
rect 12186 3675 12294 3751
rect 12666 3675 12774 3751
rect 13434 3675 13542 3751
rect 13914 3675 14022 3751
rect 14682 3675 14790 3751
rect 15162 3675 15270 3751
rect 15930 3675 16038 3751
rect 16410 3675 16518 3751
rect 17178 3675 17286 3751
rect 17658 3675 17766 3751
rect 18426 3675 18534 3751
rect 18906 3675 19014 3751
rect 19674 3675 19782 3751
rect 20154 3675 20262 3751
rect 20922 3675 21030 3751
rect 21402 3675 21510 3751
rect 22170 3675 22278 3751
rect 22650 3675 22758 3751
rect 23418 3675 23526 3751
rect 23898 3675 24006 3751
rect 24666 3675 24774 3751
rect 25146 3675 25254 3751
rect 25914 3675 26022 3751
rect 26394 3675 26502 3751
rect 27162 3675 27270 3751
rect 27642 3675 27750 3751
rect 28410 3675 28518 3751
rect 28890 3675 28998 3751
rect 29658 3675 29766 3751
rect 30138 3675 30246 3751
rect 30906 3675 31014 3751
rect 31386 3675 31494 3751
rect 32154 3675 32262 3751
rect 32634 3675 32742 3751
rect 33402 3675 33510 3751
rect 33882 3675 33990 3751
rect 34650 3675 34758 3751
rect 35130 3675 35238 3751
rect 35898 3675 36006 3751
rect 36378 3675 36486 3751
rect 37146 3675 37254 3751
rect 37626 3675 37734 3751
rect 38394 3675 38502 3751
rect 38874 3675 38982 3751
rect 39642 3675 39750 3751
rect 0 3579 39936 3627
rect 0 3483 39936 3531
rect 186 3359 294 3435
rect 954 3359 1062 3435
rect 1434 3359 1542 3435
rect 2202 3359 2310 3435
rect 2682 3359 2790 3435
rect 3450 3359 3558 3435
rect 3930 3359 4038 3435
rect 4698 3359 4806 3435
rect 5178 3359 5286 3435
rect 5946 3359 6054 3435
rect 6426 3359 6534 3435
rect 7194 3359 7302 3435
rect 7674 3359 7782 3435
rect 8442 3359 8550 3435
rect 8922 3359 9030 3435
rect 9690 3359 9798 3435
rect 10170 3359 10278 3435
rect 10938 3359 11046 3435
rect 11418 3359 11526 3435
rect 12186 3359 12294 3435
rect 12666 3359 12774 3435
rect 13434 3359 13542 3435
rect 13914 3359 14022 3435
rect 14682 3359 14790 3435
rect 15162 3359 15270 3435
rect 15930 3359 16038 3435
rect 16410 3359 16518 3435
rect 17178 3359 17286 3435
rect 17658 3359 17766 3435
rect 18426 3359 18534 3435
rect 18906 3359 19014 3435
rect 19674 3359 19782 3435
rect 20154 3359 20262 3435
rect 20922 3359 21030 3435
rect 21402 3359 21510 3435
rect 22170 3359 22278 3435
rect 22650 3359 22758 3435
rect 23418 3359 23526 3435
rect 23898 3359 24006 3435
rect 24666 3359 24774 3435
rect 25146 3359 25254 3435
rect 25914 3359 26022 3435
rect 26394 3359 26502 3435
rect 27162 3359 27270 3435
rect 27642 3359 27750 3435
rect 28410 3359 28518 3435
rect 28890 3359 28998 3435
rect 29658 3359 29766 3435
rect 30138 3359 30246 3435
rect 30906 3359 31014 3435
rect 31386 3359 31494 3435
rect 32154 3359 32262 3435
rect 32634 3359 32742 3435
rect 33402 3359 33510 3435
rect 33882 3359 33990 3435
rect 34650 3359 34758 3435
rect 35130 3359 35238 3435
rect 35898 3359 36006 3435
rect 36378 3359 36486 3435
rect 37146 3359 37254 3435
rect 37626 3359 37734 3435
rect 38394 3359 38502 3435
rect 38874 3359 38982 3435
rect 39642 3359 39750 3435
rect 0 3263 39936 3311
rect 186 3105 294 3215
rect 954 3105 1062 3215
rect 1434 3105 1542 3215
rect 2202 3105 2310 3215
rect 2682 3105 2790 3215
rect 3450 3105 3558 3215
rect 3930 3105 4038 3215
rect 4698 3105 4806 3215
rect 5178 3105 5286 3215
rect 5946 3105 6054 3215
rect 6426 3105 6534 3215
rect 7194 3105 7302 3215
rect 7674 3105 7782 3215
rect 8442 3105 8550 3215
rect 8922 3105 9030 3215
rect 9690 3105 9798 3215
rect 10170 3105 10278 3215
rect 10938 3105 11046 3215
rect 11418 3105 11526 3215
rect 12186 3105 12294 3215
rect 12666 3105 12774 3215
rect 13434 3105 13542 3215
rect 13914 3105 14022 3215
rect 14682 3105 14790 3215
rect 15162 3105 15270 3215
rect 15930 3105 16038 3215
rect 16410 3105 16518 3215
rect 17178 3105 17286 3215
rect 17658 3105 17766 3215
rect 18426 3105 18534 3215
rect 18906 3105 19014 3215
rect 19674 3105 19782 3215
rect 20154 3105 20262 3215
rect 20922 3105 21030 3215
rect 21402 3105 21510 3215
rect 22170 3105 22278 3215
rect 22650 3105 22758 3215
rect 23418 3105 23526 3215
rect 23898 3105 24006 3215
rect 24666 3105 24774 3215
rect 25146 3105 25254 3215
rect 25914 3105 26022 3215
rect 26394 3105 26502 3215
rect 27162 3105 27270 3215
rect 27642 3105 27750 3215
rect 28410 3105 28518 3215
rect 28890 3105 28998 3215
rect 29658 3105 29766 3215
rect 30138 3105 30246 3215
rect 30906 3105 31014 3215
rect 31386 3105 31494 3215
rect 32154 3105 32262 3215
rect 32634 3105 32742 3215
rect 33402 3105 33510 3215
rect 33882 3105 33990 3215
rect 34650 3105 34758 3215
rect 35130 3105 35238 3215
rect 35898 3105 36006 3215
rect 36378 3105 36486 3215
rect 37146 3105 37254 3215
rect 37626 3105 37734 3215
rect 38394 3105 38502 3215
rect 38874 3105 38982 3215
rect 39642 3105 39750 3215
rect 0 3009 39936 3057
rect 186 2885 294 2961
rect 954 2885 1062 2961
rect 1434 2885 1542 2961
rect 2202 2885 2310 2961
rect 2682 2885 2790 2961
rect 3450 2885 3558 2961
rect 3930 2885 4038 2961
rect 4698 2885 4806 2961
rect 5178 2885 5286 2961
rect 5946 2885 6054 2961
rect 6426 2885 6534 2961
rect 7194 2885 7302 2961
rect 7674 2885 7782 2961
rect 8442 2885 8550 2961
rect 8922 2885 9030 2961
rect 9690 2885 9798 2961
rect 10170 2885 10278 2961
rect 10938 2885 11046 2961
rect 11418 2885 11526 2961
rect 12186 2885 12294 2961
rect 12666 2885 12774 2961
rect 13434 2885 13542 2961
rect 13914 2885 14022 2961
rect 14682 2885 14790 2961
rect 15162 2885 15270 2961
rect 15930 2885 16038 2961
rect 16410 2885 16518 2961
rect 17178 2885 17286 2961
rect 17658 2885 17766 2961
rect 18426 2885 18534 2961
rect 18906 2885 19014 2961
rect 19674 2885 19782 2961
rect 20154 2885 20262 2961
rect 20922 2885 21030 2961
rect 21402 2885 21510 2961
rect 22170 2885 22278 2961
rect 22650 2885 22758 2961
rect 23418 2885 23526 2961
rect 23898 2885 24006 2961
rect 24666 2885 24774 2961
rect 25146 2885 25254 2961
rect 25914 2885 26022 2961
rect 26394 2885 26502 2961
rect 27162 2885 27270 2961
rect 27642 2885 27750 2961
rect 28410 2885 28518 2961
rect 28890 2885 28998 2961
rect 29658 2885 29766 2961
rect 30138 2885 30246 2961
rect 30906 2885 31014 2961
rect 31386 2885 31494 2961
rect 32154 2885 32262 2961
rect 32634 2885 32742 2961
rect 33402 2885 33510 2961
rect 33882 2885 33990 2961
rect 34650 2885 34758 2961
rect 35130 2885 35238 2961
rect 35898 2885 36006 2961
rect 36378 2885 36486 2961
rect 37146 2885 37254 2961
rect 37626 2885 37734 2961
rect 38394 2885 38502 2961
rect 38874 2885 38982 2961
rect 39642 2885 39750 2961
rect 0 2789 39936 2837
rect 0 2693 39936 2741
rect 186 2569 294 2645
rect 954 2569 1062 2645
rect 1434 2569 1542 2645
rect 2202 2569 2310 2645
rect 2682 2569 2790 2645
rect 3450 2569 3558 2645
rect 3930 2569 4038 2645
rect 4698 2569 4806 2645
rect 5178 2569 5286 2645
rect 5946 2569 6054 2645
rect 6426 2569 6534 2645
rect 7194 2569 7302 2645
rect 7674 2569 7782 2645
rect 8442 2569 8550 2645
rect 8922 2569 9030 2645
rect 9690 2569 9798 2645
rect 10170 2569 10278 2645
rect 10938 2569 11046 2645
rect 11418 2569 11526 2645
rect 12186 2569 12294 2645
rect 12666 2569 12774 2645
rect 13434 2569 13542 2645
rect 13914 2569 14022 2645
rect 14682 2569 14790 2645
rect 15162 2569 15270 2645
rect 15930 2569 16038 2645
rect 16410 2569 16518 2645
rect 17178 2569 17286 2645
rect 17658 2569 17766 2645
rect 18426 2569 18534 2645
rect 18906 2569 19014 2645
rect 19674 2569 19782 2645
rect 20154 2569 20262 2645
rect 20922 2569 21030 2645
rect 21402 2569 21510 2645
rect 22170 2569 22278 2645
rect 22650 2569 22758 2645
rect 23418 2569 23526 2645
rect 23898 2569 24006 2645
rect 24666 2569 24774 2645
rect 25146 2569 25254 2645
rect 25914 2569 26022 2645
rect 26394 2569 26502 2645
rect 27162 2569 27270 2645
rect 27642 2569 27750 2645
rect 28410 2569 28518 2645
rect 28890 2569 28998 2645
rect 29658 2569 29766 2645
rect 30138 2569 30246 2645
rect 30906 2569 31014 2645
rect 31386 2569 31494 2645
rect 32154 2569 32262 2645
rect 32634 2569 32742 2645
rect 33402 2569 33510 2645
rect 33882 2569 33990 2645
rect 34650 2569 34758 2645
rect 35130 2569 35238 2645
rect 35898 2569 36006 2645
rect 36378 2569 36486 2645
rect 37146 2569 37254 2645
rect 37626 2569 37734 2645
rect 38394 2569 38502 2645
rect 38874 2569 38982 2645
rect 39642 2569 39750 2645
rect 0 2473 39936 2521
rect 186 2315 294 2425
rect 954 2315 1062 2425
rect 1434 2315 1542 2425
rect 2202 2315 2310 2425
rect 2682 2315 2790 2425
rect 3450 2315 3558 2425
rect 3930 2315 4038 2425
rect 4698 2315 4806 2425
rect 5178 2315 5286 2425
rect 5946 2315 6054 2425
rect 6426 2315 6534 2425
rect 7194 2315 7302 2425
rect 7674 2315 7782 2425
rect 8442 2315 8550 2425
rect 8922 2315 9030 2425
rect 9690 2315 9798 2425
rect 10170 2315 10278 2425
rect 10938 2315 11046 2425
rect 11418 2315 11526 2425
rect 12186 2315 12294 2425
rect 12666 2315 12774 2425
rect 13434 2315 13542 2425
rect 13914 2315 14022 2425
rect 14682 2315 14790 2425
rect 15162 2315 15270 2425
rect 15930 2315 16038 2425
rect 16410 2315 16518 2425
rect 17178 2315 17286 2425
rect 17658 2315 17766 2425
rect 18426 2315 18534 2425
rect 18906 2315 19014 2425
rect 19674 2315 19782 2425
rect 20154 2315 20262 2425
rect 20922 2315 21030 2425
rect 21402 2315 21510 2425
rect 22170 2315 22278 2425
rect 22650 2315 22758 2425
rect 23418 2315 23526 2425
rect 23898 2315 24006 2425
rect 24666 2315 24774 2425
rect 25146 2315 25254 2425
rect 25914 2315 26022 2425
rect 26394 2315 26502 2425
rect 27162 2315 27270 2425
rect 27642 2315 27750 2425
rect 28410 2315 28518 2425
rect 28890 2315 28998 2425
rect 29658 2315 29766 2425
rect 30138 2315 30246 2425
rect 30906 2315 31014 2425
rect 31386 2315 31494 2425
rect 32154 2315 32262 2425
rect 32634 2315 32742 2425
rect 33402 2315 33510 2425
rect 33882 2315 33990 2425
rect 34650 2315 34758 2425
rect 35130 2315 35238 2425
rect 35898 2315 36006 2425
rect 36378 2315 36486 2425
rect 37146 2315 37254 2425
rect 37626 2315 37734 2425
rect 38394 2315 38502 2425
rect 38874 2315 38982 2425
rect 39642 2315 39750 2425
rect 0 2219 39936 2267
rect 186 2095 294 2171
rect 954 2095 1062 2171
rect 1434 2095 1542 2171
rect 2202 2095 2310 2171
rect 2682 2095 2790 2171
rect 3450 2095 3558 2171
rect 3930 2095 4038 2171
rect 4698 2095 4806 2171
rect 5178 2095 5286 2171
rect 5946 2095 6054 2171
rect 6426 2095 6534 2171
rect 7194 2095 7302 2171
rect 7674 2095 7782 2171
rect 8442 2095 8550 2171
rect 8922 2095 9030 2171
rect 9690 2095 9798 2171
rect 10170 2095 10278 2171
rect 10938 2095 11046 2171
rect 11418 2095 11526 2171
rect 12186 2095 12294 2171
rect 12666 2095 12774 2171
rect 13434 2095 13542 2171
rect 13914 2095 14022 2171
rect 14682 2095 14790 2171
rect 15162 2095 15270 2171
rect 15930 2095 16038 2171
rect 16410 2095 16518 2171
rect 17178 2095 17286 2171
rect 17658 2095 17766 2171
rect 18426 2095 18534 2171
rect 18906 2095 19014 2171
rect 19674 2095 19782 2171
rect 20154 2095 20262 2171
rect 20922 2095 21030 2171
rect 21402 2095 21510 2171
rect 22170 2095 22278 2171
rect 22650 2095 22758 2171
rect 23418 2095 23526 2171
rect 23898 2095 24006 2171
rect 24666 2095 24774 2171
rect 25146 2095 25254 2171
rect 25914 2095 26022 2171
rect 26394 2095 26502 2171
rect 27162 2095 27270 2171
rect 27642 2095 27750 2171
rect 28410 2095 28518 2171
rect 28890 2095 28998 2171
rect 29658 2095 29766 2171
rect 30138 2095 30246 2171
rect 30906 2095 31014 2171
rect 31386 2095 31494 2171
rect 32154 2095 32262 2171
rect 32634 2095 32742 2171
rect 33402 2095 33510 2171
rect 33882 2095 33990 2171
rect 34650 2095 34758 2171
rect 35130 2095 35238 2171
rect 35898 2095 36006 2171
rect 36378 2095 36486 2171
rect 37146 2095 37254 2171
rect 37626 2095 37734 2171
rect 38394 2095 38502 2171
rect 38874 2095 38982 2171
rect 39642 2095 39750 2171
rect 0 1999 39936 2047
rect 0 1903 39936 1951
rect 186 1779 294 1855
rect 954 1779 1062 1855
rect 1434 1779 1542 1855
rect 2202 1779 2310 1855
rect 2682 1779 2790 1855
rect 3450 1779 3558 1855
rect 3930 1779 4038 1855
rect 4698 1779 4806 1855
rect 5178 1779 5286 1855
rect 5946 1779 6054 1855
rect 6426 1779 6534 1855
rect 7194 1779 7302 1855
rect 7674 1779 7782 1855
rect 8442 1779 8550 1855
rect 8922 1779 9030 1855
rect 9690 1779 9798 1855
rect 10170 1779 10278 1855
rect 10938 1779 11046 1855
rect 11418 1779 11526 1855
rect 12186 1779 12294 1855
rect 12666 1779 12774 1855
rect 13434 1779 13542 1855
rect 13914 1779 14022 1855
rect 14682 1779 14790 1855
rect 15162 1779 15270 1855
rect 15930 1779 16038 1855
rect 16410 1779 16518 1855
rect 17178 1779 17286 1855
rect 17658 1779 17766 1855
rect 18426 1779 18534 1855
rect 18906 1779 19014 1855
rect 19674 1779 19782 1855
rect 20154 1779 20262 1855
rect 20922 1779 21030 1855
rect 21402 1779 21510 1855
rect 22170 1779 22278 1855
rect 22650 1779 22758 1855
rect 23418 1779 23526 1855
rect 23898 1779 24006 1855
rect 24666 1779 24774 1855
rect 25146 1779 25254 1855
rect 25914 1779 26022 1855
rect 26394 1779 26502 1855
rect 27162 1779 27270 1855
rect 27642 1779 27750 1855
rect 28410 1779 28518 1855
rect 28890 1779 28998 1855
rect 29658 1779 29766 1855
rect 30138 1779 30246 1855
rect 30906 1779 31014 1855
rect 31386 1779 31494 1855
rect 32154 1779 32262 1855
rect 32634 1779 32742 1855
rect 33402 1779 33510 1855
rect 33882 1779 33990 1855
rect 34650 1779 34758 1855
rect 35130 1779 35238 1855
rect 35898 1779 36006 1855
rect 36378 1779 36486 1855
rect 37146 1779 37254 1855
rect 37626 1779 37734 1855
rect 38394 1779 38502 1855
rect 38874 1779 38982 1855
rect 39642 1779 39750 1855
rect 0 1683 39936 1731
rect 186 1525 294 1635
rect 954 1525 1062 1635
rect 1434 1525 1542 1635
rect 2202 1525 2310 1635
rect 2682 1525 2790 1635
rect 3450 1525 3558 1635
rect 3930 1525 4038 1635
rect 4698 1525 4806 1635
rect 5178 1525 5286 1635
rect 5946 1525 6054 1635
rect 6426 1525 6534 1635
rect 7194 1525 7302 1635
rect 7674 1525 7782 1635
rect 8442 1525 8550 1635
rect 8922 1525 9030 1635
rect 9690 1525 9798 1635
rect 10170 1525 10278 1635
rect 10938 1525 11046 1635
rect 11418 1525 11526 1635
rect 12186 1525 12294 1635
rect 12666 1525 12774 1635
rect 13434 1525 13542 1635
rect 13914 1525 14022 1635
rect 14682 1525 14790 1635
rect 15162 1525 15270 1635
rect 15930 1525 16038 1635
rect 16410 1525 16518 1635
rect 17178 1525 17286 1635
rect 17658 1525 17766 1635
rect 18426 1525 18534 1635
rect 18906 1525 19014 1635
rect 19674 1525 19782 1635
rect 20154 1525 20262 1635
rect 20922 1525 21030 1635
rect 21402 1525 21510 1635
rect 22170 1525 22278 1635
rect 22650 1525 22758 1635
rect 23418 1525 23526 1635
rect 23898 1525 24006 1635
rect 24666 1525 24774 1635
rect 25146 1525 25254 1635
rect 25914 1525 26022 1635
rect 26394 1525 26502 1635
rect 27162 1525 27270 1635
rect 27642 1525 27750 1635
rect 28410 1525 28518 1635
rect 28890 1525 28998 1635
rect 29658 1525 29766 1635
rect 30138 1525 30246 1635
rect 30906 1525 31014 1635
rect 31386 1525 31494 1635
rect 32154 1525 32262 1635
rect 32634 1525 32742 1635
rect 33402 1525 33510 1635
rect 33882 1525 33990 1635
rect 34650 1525 34758 1635
rect 35130 1525 35238 1635
rect 35898 1525 36006 1635
rect 36378 1525 36486 1635
rect 37146 1525 37254 1635
rect 37626 1525 37734 1635
rect 38394 1525 38502 1635
rect 38874 1525 38982 1635
rect 39642 1525 39750 1635
rect 0 1429 39936 1477
rect 186 1305 294 1381
rect 954 1305 1062 1381
rect 1434 1305 1542 1381
rect 2202 1305 2310 1381
rect 2682 1305 2790 1381
rect 3450 1305 3558 1381
rect 3930 1305 4038 1381
rect 4698 1305 4806 1381
rect 5178 1305 5286 1381
rect 5946 1305 6054 1381
rect 6426 1305 6534 1381
rect 7194 1305 7302 1381
rect 7674 1305 7782 1381
rect 8442 1305 8550 1381
rect 8922 1305 9030 1381
rect 9690 1305 9798 1381
rect 10170 1305 10278 1381
rect 10938 1305 11046 1381
rect 11418 1305 11526 1381
rect 12186 1305 12294 1381
rect 12666 1305 12774 1381
rect 13434 1305 13542 1381
rect 13914 1305 14022 1381
rect 14682 1305 14790 1381
rect 15162 1305 15270 1381
rect 15930 1305 16038 1381
rect 16410 1305 16518 1381
rect 17178 1305 17286 1381
rect 17658 1305 17766 1381
rect 18426 1305 18534 1381
rect 18906 1305 19014 1381
rect 19674 1305 19782 1381
rect 20154 1305 20262 1381
rect 20922 1305 21030 1381
rect 21402 1305 21510 1381
rect 22170 1305 22278 1381
rect 22650 1305 22758 1381
rect 23418 1305 23526 1381
rect 23898 1305 24006 1381
rect 24666 1305 24774 1381
rect 25146 1305 25254 1381
rect 25914 1305 26022 1381
rect 26394 1305 26502 1381
rect 27162 1305 27270 1381
rect 27642 1305 27750 1381
rect 28410 1305 28518 1381
rect 28890 1305 28998 1381
rect 29658 1305 29766 1381
rect 30138 1305 30246 1381
rect 30906 1305 31014 1381
rect 31386 1305 31494 1381
rect 32154 1305 32262 1381
rect 32634 1305 32742 1381
rect 33402 1305 33510 1381
rect 33882 1305 33990 1381
rect 34650 1305 34758 1381
rect 35130 1305 35238 1381
rect 35898 1305 36006 1381
rect 36378 1305 36486 1381
rect 37146 1305 37254 1381
rect 37626 1305 37734 1381
rect 38394 1305 38502 1381
rect 38874 1305 38982 1381
rect 39642 1305 39750 1381
rect 0 1209 39936 1257
rect 0 1113 39936 1161
rect 186 989 294 1065
rect 954 989 1062 1065
rect 1434 989 1542 1065
rect 2202 989 2310 1065
rect 2682 989 2790 1065
rect 3450 989 3558 1065
rect 3930 989 4038 1065
rect 4698 989 4806 1065
rect 5178 989 5286 1065
rect 5946 989 6054 1065
rect 6426 989 6534 1065
rect 7194 989 7302 1065
rect 7674 989 7782 1065
rect 8442 989 8550 1065
rect 8922 989 9030 1065
rect 9690 989 9798 1065
rect 10170 989 10278 1065
rect 10938 989 11046 1065
rect 11418 989 11526 1065
rect 12186 989 12294 1065
rect 12666 989 12774 1065
rect 13434 989 13542 1065
rect 13914 989 14022 1065
rect 14682 989 14790 1065
rect 15162 989 15270 1065
rect 15930 989 16038 1065
rect 16410 989 16518 1065
rect 17178 989 17286 1065
rect 17658 989 17766 1065
rect 18426 989 18534 1065
rect 18906 989 19014 1065
rect 19674 989 19782 1065
rect 20154 989 20262 1065
rect 20922 989 21030 1065
rect 21402 989 21510 1065
rect 22170 989 22278 1065
rect 22650 989 22758 1065
rect 23418 989 23526 1065
rect 23898 989 24006 1065
rect 24666 989 24774 1065
rect 25146 989 25254 1065
rect 25914 989 26022 1065
rect 26394 989 26502 1065
rect 27162 989 27270 1065
rect 27642 989 27750 1065
rect 28410 989 28518 1065
rect 28890 989 28998 1065
rect 29658 989 29766 1065
rect 30138 989 30246 1065
rect 30906 989 31014 1065
rect 31386 989 31494 1065
rect 32154 989 32262 1065
rect 32634 989 32742 1065
rect 33402 989 33510 1065
rect 33882 989 33990 1065
rect 34650 989 34758 1065
rect 35130 989 35238 1065
rect 35898 989 36006 1065
rect 36378 989 36486 1065
rect 37146 989 37254 1065
rect 37626 989 37734 1065
rect 38394 989 38502 1065
rect 38874 989 38982 1065
rect 39642 989 39750 1065
rect 0 893 39936 941
rect 186 735 294 845
rect 954 735 1062 845
rect 1434 735 1542 845
rect 2202 735 2310 845
rect 2682 735 2790 845
rect 3450 735 3558 845
rect 3930 735 4038 845
rect 4698 735 4806 845
rect 5178 735 5286 845
rect 5946 735 6054 845
rect 6426 735 6534 845
rect 7194 735 7302 845
rect 7674 735 7782 845
rect 8442 735 8550 845
rect 8922 735 9030 845
rect 9690 735 9798 845
rect 10170 735 10278 845
rect 10938 735 11046 845
rect 11418 735 11526 845
rect 12186 735 12294 845
rect 12666 735 12774 845
rect 13434 735 13542 845
rect 13914 735 14022 845
rect 14682 735 14790 845
rect 15162 735 15270 845
rect 15930 735 16038 845
rect 16410 735 16518 845
rect 17178 735 17286 845
rect 17658 735 17766 845
rect 18426 735 18534 845
rect 18906 735 19014 845
rect 19674 735 19782 845
rect 20154 735 20262 845
rect 20922 735 21030 845
rect 21402 735 21510 845
rect 22170 735 22278 845
rect 22650 735 22758 845
rect 23418 735 23526 845
rect 23898 735 24006 845
rect 24666 735 24774 845
rect 25146 735 25254 845
rect 25914 735 26022 845
rect 26394 735 26502 845
rect 27162 735 27270 845
rect 27642 735 27750 845
rect 28410 735 28518 845
rect 28890 735 28998 845
rect 29658 735 29766 845
rect 30138 735 30246 845
rect 30906 735 31014 845
rect 31386 735 31494 845
rect 32154 735 32262 845
rect 32634 735 32742 845
rect 33402 735 33510 845
rect 33882 735 33990 845
rect 34650 735 34758 845
rect 35130 735 35238 845
rect 35898 735 36006 845
rect 36378 735 36486 845
rect 37146 735 37254 845
rect 37626 735 37734 845
rect 38394 735 38502 845
rect 38874 735 38982 845
rect 39642 735 39750 845
rect 0 639 39936 687
rect 186 515 294 591
rect 954 515 1062 591
rect 1434 515 1542 591
rect 2202 515 2310 591
rect 2682 515 2790 591
rect 3450 515 3558 591
rect 3930 515 4038 591
rect 4698 515 4806 591
rect 5178 515 5286 591
rect 5946 515 6054 591
rect 6426 515 6534 591
rect 7194 515 7302 591
rect 7674 515 7782 591
rect 8442 515 8550 591
rect 8922 515 9030 591
rect 9690 515 9798 591
rect 10170 515 10278 591
rect 10938 515 11046 591
rect 11418 515 11526 591
rect 12186 515 12294 591
rect 12666 515 12774 591
rect 13434 515 13542 591
rect 13914 515 14022 591
rect 14682 515 14790 591
rect 15162 515 15270 591
rect 15930 515 16038 591
rect 16410 515 16518 591
rect 17178 515 17286 591
rect 17658 515 17766 591
rect 18426 515 18534 591
rect 18906 515 19014 591
rect 19674 515 19782 591
rect 20154 515 20262 591
rect 20922 515 21030 591
rect 21402 515 21510 591
rect 22170 515 22278 591
rect 22650 515 22758 591
rect 23418 515 23526 591
rect 23898 515 24006 591
rect 24666 515 24774 591
rect 25146 515 25254 591
rect 25914 515 26022 591
rect 26394 515 26502 591
rect 27162 515 27270 591
rect 27642 515 27750 591
rect 28410 515 28518 591
rect 28890 515 28998 591
rect 29658 515 29766 591
rect 30138 515 30246 591
rect 30906 515 31014 591
rect 31386 515 31494 591
rect 32154 515 32262 591
rect 32634 515 32742 591
rect 33402 515 33510 591
rect 33882 515 33990 591
rect 34650 515 34758 591
rect 35130 515 35238 591
rect 35898 515 36006 591
rect 36378 515 36486 591
rect 37146 515 37254 591
rect 37626 515 37734 591
rect 38394 515 38502 591
rect 38874 515 38982 591
rect 39642 515 39750 591
rect 0 419 39936 467
rect 0 323 39936 371
rect 186 199 294 275
rect 954 199 1062 275
rect 1434 199 1542 275
rect 2202 199 2310 275
rect 2682 199 2790 275
rect 3450 199 3558 275
rect 3930 199 4038 275
rect 4698 199 4806 275
rect 5178 199 5286 275
rect 5946 199 6054 275
rect 6426 199 6534 275
rect 7194 199 7302 275
rect 7674 199 7782 275
rect 8442 199 8550 275
rect 8922 199 9030 275
rect 9690 199 9798 275
rect 10170 199 10278 275
rect 10938 199 11046 275
rect 11418 199 11526 275
rect 12186 199 12294 275
rect 12666 199 12774 275
rect 13434 199 13542 275
rect 13914 199 14022 275
rect 14682 199 14790 275
rect 15162 199 15270 275
rect 15930 199 16038 275
rect 16410 199 16518 275
rect 17178 199 17286 275
rect 17658 199 17766 275
rect 18426 199 18534 275
rect 18906 199 19014 275
rect 19674 199 19782 275
rect 20154 199 20262 275
rect 20922 199 21030 275
rect 21402 199 21510 275
rect 22170 199 22278 275
rect 22650 199 22758 275
rect 23418 199 23526 275
rect 23898 199 24006 275
rect 24666 199 24774 275
rect 25146 199 25254 275
rect 25914 199 26022 275
rect 26394 199 26502 275
rect 27162 199 27270 275
rect 27642 199 27750 275
rect 28410 199 28518 275
rect 28890 199 28998 275
rect 29658 199 29766 275
rect 30138 199 30246 275
rect 30906 199 31014 275
rect 31386 199 31494 275
rect 32154 199 32262 275
rect 32634 199 32742 275
rect 33402 199 33510 275
rect 33882 199 33990 275
rect 34650 199 34758 275
rect 35130 199 35238 275
rect 35898 199 36006 275
rect 36378 199 36486 275
rect 37146 199 37254 275
rect 37626 199 37734 275
rect 38394 199 38502 275
rect 38874 199 38982 275
rect 39642 199 39750 275
rect 0 103 39936 151
rect 186 -55 294 55
rect 954 -55 1062 55
rect 1434 -55 1542 55
rect 2202 -55 2310 55
rect 2682 -55 2790 55
rect 3450 -55 3558 55
rect 3930 -55 4038 55
rect 4698 -55 4806 55
rect 5178 -55 5286 55
rect 5946 -55 6054 55
rect 6426 -55 6534 55
rect 7194 -55 7302 55
rect 7674 -55 7782 55
rect 8442 -55 8550 55
rect 8922 -55 9030 55
rect 9690 -55 9798 55
rect 10170 -55 10278 55
rect 10938 -55 11046 55
rect 11418 -55 11526 55
rect 12186 -55 12294 55
rect 12666 -55 12774 55
rect 13434 -55 13542 55
rect 13914 -55 14022 55
rect 14682 -55 14790 55
rect 15162 -55 15270 55
rect 15930 -55 16038 55
rect 16410 -55 16518 55
rect 17178 -55 17286 55
rect 17658 -55 17766 55
rect 18426 -55 18534 55
rect 18906 -55 19014 55
rect 19674 -55 19782 55
rect 20154 -55 20262 55
rect 20922 -55 21030 55
rect 21402 -55 21510 55
rect 22170 -55 22278 55
rect 22650 -55 22758 55
rect 23418 -55 23526 55
rect 23898 -55 24006 55
rect 24666 -55 24774 55
rect 25146 -55 25254 55
rect 25914 -55 26022 55
rect 26394 -55 26502 55
rect 27162 -55 27270 55
rect 27642 -55 27750 55
rect 28410 -55 28518 55
rect 28890 -55 28998 55
rect 29658 -55 29766 55
rect 30138 -55 30246 55
rect 30906 -55 31014 55
rect 31386 -55 31494 55
rect 32154 -55 32262 55
rect 32634 -55 32742 55
rect 33402 -55 33510 55
rect 33882 -55 33990 55
rect 34650 -55 34758 55
rect 35130 -55 35238 55
rect 35898 -55 36006 55
rect 36378 -55 36486 55
rect 37146 -55 37254 55
rect 37626 -55 37734 55
rect 38394 -55 38502 55
rect 38874 -55 38982 55
rect 39642 -55 39750 55
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_0
timestamp 1666464484
transform -1 0 39936 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1
timestamp 1666464484
transform -1 0 39936 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2
timestamp 1666464484
transform -1 0 38688 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3
timestamp 1666464484
transform 1 0 38688 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4
timestamp 1666464484
transform 1 0 38688 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5
timestamp 1666464484
transform -1 0 38688 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6
timestamp 1666464484
transform -1 0 38688 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7
timestamp 1666464484
transform -1 0 38688 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8
timestamp 1666464484
transform -1 0 38688 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_9
timestamp 1666464484
transform -1 0 38688 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_10
timestamp 1666464484
transform -1 0 38688 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_11
timestamp 1666464484
transform 1 0 38688 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_12
timestamp 1666464484
transform 1 0 38688 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_13
timestamp 1666464484
transform 1 0 38688 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_14
timestamp 1666464484
transform 1 0 38688 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_15
timestamp 1666464484
transform 1 0 38688 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_16
timestamp 1666464484
transform -1 0 39936 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_17
timestamp 1666464484
transform -1 0 39936 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_18
timestamp 1666464484
transform -1 0 39936 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_19
timestamp 1666464484
transform -1 0 39936 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_20
timestamp 1666464484
transform -1 0 39936 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_21
timestamp 1666464484
transform 1 0 36192 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_22
timestamp 1666464484
transform 1 0 36192 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_23
timestamp 1666464484
transform 1 0 36192 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_24
timestamp 1666464484
transform 1 0 36192 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_25
timestamp 1666464484
transform 1 0 36192 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_26
timestamp 1666464484
transform 1 0 36192 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_27
timestamp 1666464484
transform -1 0 36192 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_28
timestamp 1666464484
transform -1 0 36192 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_29
timestamp 1666464484
transform -1 0 36192 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_30
timestamp 1666464484
transform -1 0 36192 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_31
timestamp 1666464484
transform -1 0 36192 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_32
timestamp 1666464484
transform -1 0 36192 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_33
timestamp 1666464484
transform -1 0 36192 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_34
timestamp 1666464484
transform 1 0 36192 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_35
timestamp 1666464484
transform 1 0 36192 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_36
timestamp 1666464484
transform 1 0 36192 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_37
timestamp 1666464484
transform 1 0 36192 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_38
timestamp 1666464484
transform 1 0 36192 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_39
timestamp 1666464484
transform 1 0 36192 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_40
timestamp 1666464484
transform 1 0 36192 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_41
timestamp 1666464484
transform -1 0 36192 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_42
timestamp 1666464484
transform -1 0 36192 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_43
timestamp 1666464484
transform -1 0 36192 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_44
timestamp 1666464484
transform -1 0 36192 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_45
timestamp 1666464484
transform -1 0 36192 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_46
timestamp 1666464484
transform -1 0 36192 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_47
timestamp 1666464484
transform -1 0 38688 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_48
timestamp 1666464484
transform 1 0 38688 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_49
timestamp 1666464484
transform 1 0 38688 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_50
timestamp 1666464484
transform 1 0 38688 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_51
timestamp 1666464484
transform 1 0 38688 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_52
timestamp 1666464484
transform 1 0 38688 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_53
timestamp 1666464484
transform 1 0 38688 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_54
timestamp 1666464484
transform -1 0 38688 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_55
timestamp 1666464484
transform -1 0 39936 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_56
timestamp 1666464484
transform -1 0 39936 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_57
timestamp 1666464484
transform -1 0 39936 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_58
timestamp 1666464484
transform -1 0 39936 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_59
timestamp 1666464484
transform -1 0 39936 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_60
timestamp 1666464484
transform -1 0 39936 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_61
timestamp 1666464484
transform -1 0 38688 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_62
timestamp 1666464484
transform -1 0 38688 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_63
timestamp 1666464484
transform -1 0 38688 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_64
timestamp 1666464484
transform -1 0 38688 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_65
timestamp 1666464484
transform -1 0 38688 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_66
timestamp 1666464484
transform 1 0 38688 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_67
timestamp 1666464484
transform -1 0 39936 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_68
timestamp 1666464484
transform -1 0 39936 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_69
timestamp 1666464484
transform 1 0 38688 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_70
timestamp 1666464484
transform -1 0 37440 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_71
timestamp 1666464484
transform -1 0 37440 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_72
timestamp 1666464484
transform -1 0 37440 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_73
timestamp 1666464484
transform -1 0 37440 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_74
timestamp 1666464484
transform -1 0 37440 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_75
timestamp 1666464484
transform -1 0 37440 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_76
timestamp 1666464484
transform 1 0 37440 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_77
timestamp 1666464484
transform 1 0 37440 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_78
timestamp 1666464484
transform 1 0 37440 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_79
timestamp 1666464484
transform 1 0 37440 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_80
timestamp 1666464484
transform 1 0 37440 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_81
timestamp 1666464484
transform 1 0 37440 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_82
timestamp 1666464484
transform 1 0 37440 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_83
timestamp 1666464484
transform 1 0 37440 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_84
timestamp 1666464484
transform 1 0 37440 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_85
timestamp 1666464484
transform 1 0 37440 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_86
timestamp 1666464484
transform 1 0 37440 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_87
timestamp 1666464484
transform 1 0 37440 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_88
timestamp 1666464484
transform 1 0 37440 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_89
timestamp 1666464484
transform 1 0 37440 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_90
timestamp 1666464484
transform 1 0 37440 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_91
timestamp 1666464484
transform -1 0 37440 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_92
timestamp 1666464484
transform -1 0 37440 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_93
timestamp 1666464484
transform -1 0 37440 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_94
timestamp 1666464484
transform -1 0 37440 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_95
timestamp 1666464484
transform -1 0 37440 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_96
timestamp 1666464484
transform -1 0 37440 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_97
timestamp 1666464484
transform -1 0 37440 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_98
timestamp 1666464484
transform -1 0 37440 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_99
timestamp 1666464484
transform -1 0 37440 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_100
timestamp 1666464484
transform -1 0 38688 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_101
timestamp 1666464484
transform -1 0 36192 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_102
timestamp 1666464484
transform -1 0 36192 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_103
timestamp 1666464484
transform 1 0 36192 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_104
timestamp 1666464484
transform 1 0 36192 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_105
timestamp 1666464484
transform 1 0 31200 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_106
timestamp 1666464484
transform 1 0 31200 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_107
timestamp 1666464484
transform 1 0 31200 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_108
timestamp 1666464484
transform 1 0 31200 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_109
timestamp 1666464484
transform 1 0 31200 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_110
timestamp 1666464484
transform 1 0 31200 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_111
timestamp 1666464484
transform -1 0 32448 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_112
timestamp 1666464484
transform -1 0 32448 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_113
timestamp 1666464484
transform -1 0 33696 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_114
timestamp 1666464484
transform -1 0 33696 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_115
timestamp 1666464484
transform -1 0 33696 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_116
timestamp 1666464484
transform -1 0 33696 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_117
timestamp 1666464484
transform -1 0 33696 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_118
timestamp 1666464484
transform 1 0 32448 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_119
timestamp 1666464484
transform 1 0 32448 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_120
timestamp 1666464484
transform 1 0 32448 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_121
timestamp 1666464484
transform 1 0 32448 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_122
timestamp 1666464484
transform 1 0 31200 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_123
timestamp 1666464484
transform 1 0 31200 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_124
timestamp 1666464484
transform 1 0 31200 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_125
timestamp 1666464484
transform 1 0 31200 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_126
timestamp 1666464484
transform -1 0 32448 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_127
timestamp 1666464484
transform 1 0 32448 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_128
timestamp 1666464484
transform 1 0 32448 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_129
timestamp 1666464484
transform 1 0 32448 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_130
timestamp 1666464484
transform 1 0 32448 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_131
timestamp 1666464484
transform 1 0 32448 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_132
timestamp 1666464484
transform 1 0 32448 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_133
timestamp 1666464484
transform 1 0 32448 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_134
timestamp 1666464484
transform 1 0 32448 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_135
timestamp 1666464484
transform 1 0 32448 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_136
timestamp 1666464484
transform 1 0 32448 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_137
timestamp 1666464484
transform 1 0 32448 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_138
timestamp 1666464484
transform -1 0 31200 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_139
timestamp 1666464484
transform -1 0 31200 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_140
timestamp 1666464484
transform 1 0 33696 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_141
timestamp 1666464484
transform 1 0 33696 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_142
timestamp 1666464484
transform 1 0 33696 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_143
timestamp 1666464484
transform 1 0 33696 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_144
timestamp 1666464484
transform 1 0 33696 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_145
timestamp 1666464484
transform 1 0 33696 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_146
timestamp 1666464484
transform 1 0 33696 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_147
timestamp 1666464484
transform 1 0 33696 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_148
timestamp 1666464484
transform 1 0 33696 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_149
timestamp 1666464484
transform 1 0 33696 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_150
timestamp 1666464484
transform 1 0 33696 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_151
timestamp 1666464484
transform 1 0 33696 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_152
timestamp 1666464484
transform 1 0 33696 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_153
timestamp 1666464484
transform 1 0 33696 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_154
timestamp 1666464484
transform 1 0 33696 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_155
timestamp 1666464484
transform -1 0 32448 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_156
timestamp 1666464484
transform -1 0 32448 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_157
timestamp 1666464484
transform -1 0 32448 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_158
timestamp 1666464484
transform -1 0 32448 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_159
timestamp 1666464484
transform -1 0 32448 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_160
timestamp 1666464484
transform -1 0 32448 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_161
timestamp 1666464484
transform -1 0 32448 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_162
timestamp 1666464484
transform -1 0 32448 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_163
timestamp 1666464484
transform -1 0 32448 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_164
timestamp 1666464484
transform -1 0 32448 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_165
timestamp 1666464484
transform -1 0 32448 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_166
timestamp 1666464484
transform -1 0 32448 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_167
timestamp 1666464484
transform 1 0 31200 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_168
timestamp 1666464484
transform 1 0 31200 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_169
timestamp 1666464484
transform 1 0 31200 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_170
timestamp 1666464484
transform -1 0 33696 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_171
timestamp 1666464484
transform -1 0 33696 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_172
timestamp 1666464484
transform -1 0 33696 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_173
timestamp 1666464484
transform -1 0 33696 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_174
timestamp 1666464484
transform -1 0 33696 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_175
timestamp 1666464484
transform -1 0 33696 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_176
timestamp 1666464484
transform -1 0 33696 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_177
timestamp 1666464484
transform -1 0 33696 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_178
timestamp 1666464484
transform -1 0 33696 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_179
timestamp 1666464484
transform -1 0 33696 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_180
timestamp 1666464484
transform 1 0 31200 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_181
timestamp 1666464484
transform -1 0 31200 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_182
timestamp 1666464484
transform -1 0 31200 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_183
timestamp 1666464484
transform -1 0 31200 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_184
timestamp 1666464484
transform -1 0 31200 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_185
timestamp 1666464484
transform -1 0 31200 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_186
timestamp 1666464484
transform -1 0 31200 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_187
timestamp 1666464484
transform -1 0 31200 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_188
timestamp 1666464484
transform -1 0 31200 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_189
timestamp 1666464484
transform -1 0 31200 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_190
timestamp 1666464484
transform -1 0 31200 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_191
timestamp 1666464484
transform -1 0 31200 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_192
timestamp 1666464484
transform -1 0 31200 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_193
timestamp 1666464484
transform -1 0 31200 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_194
timestamp 1666464484
transform 1 0 31200 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_195
timestamp 1666464484
transform 1 0 31200 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_196
timestamp 1666464484
transform 1 0 31200 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_197
timestamp 1666464484
transform 1 0 31200 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_198
timestamp 1666464484
transform 1 0 31200 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_199
timestamp 1666464484
transform 1 0 31200 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_200
timestamp 1666464484
transform 1 0 31200 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_201
timestamp 1666464484
transform 1 0 31200 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_202
timestamp 1666464484
transform 1 0 31200 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_203
timestamp 1666464484
transform -1 0 32448 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_204
timestamp 1666464484
transform 1 0 33696 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_205
timestamp 1666464484
transform 1 0 32448 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_206
timestamp 1666464484
transform 1 0 32448 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_207
timestamp 1666464484
transform 1 0 32448 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_208
timestamp 1666464484
transform 1 0 32448 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_209
timestamp 1666464484
transform 1 0 32448 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_210
timestamp 1666464484
transform 1 0 32448 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_211
timestamp 1666464484
transform 1 0 32448 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_212
timestamp 1666464484
transform 1 0 32448 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_213
timestamp 1666464484
transform 1 0 32448 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_214
timestamp 1666464484
transform 1 0 32448 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_215
timestamp 1666464484
transform 1 0 32448 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_216
timestamp 1666464484
transform 1 0 32448 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_217
timestamp 1666464484
transform 1 0 32448 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_218
timestamp 1666464484
transform 1 0 32448 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_219
timestamp 1666464484
transform 1 0 33696 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_220
timestamp 1666464484
transform 1 0 33696 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_221
timestamp 1666464484
transform -1 0 33696 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_222
timestamp 1666464484
transform -1 0 33696 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_223
timestamp 1666464484
transform -1 0 33696 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_224
timestamp 1666464484
transform -1 0 33696 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_225
timestamp 1666464484
transform -1 0 33696 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_226
timestamp 1666464484
transform -1 0 33696 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_227
timestamp 1666464484
transform -1 0 33696 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_228
timestamp 1666464484
transform 1 0 33696 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_229
timestamp 1666464484
transform 1 0 33696 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_230
timestamp 1666464484
transform 1 0 33696 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_231
timestamp 1666464484
transform 1 0 33696 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_232
timestamp 1666464484
transform 1 0 33696 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_233
timestamp 1666464484
transform 1 0 33696 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_234
timestamp 1666464484
transform 1 0 33696 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_235
timestamp 1666464484
transform 1 0 33696 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_236
timestamp 1666464484
transform 1 0 33696 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_237
timestamp 1666464484
transform 1 0 33696 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_238
timestamp 1666464484
transform -1 0 31200 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_239
timestamp 1666464484
transform -1 0 31200 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_240
timestamp 1666464484
transform -1 0 31200 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_241
timestamp 1666464484
transform -1 0 31200 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_242
timestamp 1666464484
transform -1 0 31200 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_243
timestamp 1666464484
transform -1 0 31200 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_244
timestamp 1666464484
transform -1 0 33696 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_245
timestamp 1666464484
transform -1 0 33696 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_246
timestamp 1666464484
transform -1 0 33696 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_247
timestamp 1666464484
transform -1 0 33696 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_248
timestamp 1666464484
transform -1 0 33696 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_249
timestamp 1666464484
transform -1 0 33696 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_250
timestamp 1666464484
transform -1 0 33696 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_251
timestamp 1666464484
transform -1 0 31200 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_252
timestamp 1666464484
transform -1 0 31200 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_253
timestamp 1666464484
transform 1 0 31200 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_254
timestamp 1666464484
transform 1 0 31200 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_255
timestamp 1666464484
transform 1 0 31200 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_256
timestamp 1666464484
transform 1 0 31200 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_257
timestamp 1666464484
transform 1 0 31200 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_258
timestamp 1666464484
transform 1 0 31200 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_259
timestamp 1666464484
transform -1 0 31200 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_260
timestamp 1666464484
transform -1 0 31200 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_261
timestamp 1666464484
transform -1 0 31200 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_262
timestamp 1666464484
transform -1 0 31200 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_263
timestamp 1666464484
transform -1 0 32448 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_264
timestamp 1666464484
transform -1 0 32448 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_265
timestamp 1666464484
transform -1 0 32448 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_266
timestamp 1666464484
transform -1 0 31200 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_267
timestamp 1666464484
transform -1 0 31200 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_268
timestamp 1666464484
transform 1 0 33696 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_269
timestamp 1666464484
transform -1 0 32448 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_270
timestamp 1666464484
transform -1 0 32448 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_271
timestamp 1666464484
transform -1 0 32448 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_272
timestamp 1666464484
transform -1 0 32448 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_273
timestamp 1666464484
transform -1 0 32448 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_274
timestamp 1666464484
transform -1 0 32448 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_275
timestamp 1666464484
transform -1 0 32448 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_276
timestamp 1666464484
transform -1 0 32448 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_277
timestamp 1666464484
transform -1 0 32448 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_278
timestamp 1666464484
transform -1 0 32448 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_279
timestamp 1666464484
transform -1 0 38688 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_280
timestamp 1666464484
transform -1 0 38688 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_281
timestamp 1666464484
transform -1 0 38688 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_282
timestamp 1666464484
transform 1 0 38688 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_283
timestamp 1666464484
transform 1 0 38688 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_284
timestamp 1666464484
transform 1 0 38688 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_285
timestamp 1666464484
transform 1 0 38688 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_286
timestamp 1666464484
transform 1 0 38688 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_287
timestamp 1666464484
transform 1 0 38688 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_288
timestamp 1666464484
transform 1 0 38688 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_289
timestamp 1666464484
transform 1 0 38688 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_290
timestamp 1666464484
transform 1 0 37440 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_291
timestamp 1666464484
transform 1 0 37440 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_292
timestamp 1666464484
transform 1 0 37440 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_293
timestamp 1666464484
transform 1 0 37440 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_294
timestamp 1666464484
transform 1 0 37440 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_295
timestamp 1666464484
transform 1 0 37440 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_296
timestamp 1666464484
transform 1 0 37440 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_297
timestamp 1666464484
transform 1 0 37440 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_298
timestamp 1666464484
transform 1 0 37440 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_299
timestamp 1666464484
transform 1 0 37440 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_300
timestamp 1666464484
transform 1 0 37440 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_301
timestamp 1666464484
transform 1 0 37440 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_302
timestamp 1666464484
transform 1 0 37440 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_303
timestamp 1666464484
transform 1 0 37440 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_304
timestamp 1666464484
transform 1 0 38688 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_305
timestamp 1666464484
transform 1 0 38688 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_306
timestamp 1666464484
transform 1 0 38688 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_307
timestamp 1666464484
transform 1 0 38688 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_308
timestamp 1666464484
transform 1 0 38688 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_309
timestamp 1666464484
transform 1 0 38688 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_310
timestamp 1666464484
transform -1 0 38688 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_311
timestamp 1666464484
transform -1 0 38688 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_312
timestamp 1666464484
transform -1 0 38688 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_313
timestamp 1666464484
transform -1 0 38688 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_314
timestamp 1666464484
transform -1 0 38688 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_315
timestamp 1666464484
transform -1 0 38688 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_316
timestamp 1666464484
transform -1 0 38688 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_317
timestamp 1666464484
transform -1 0 38688 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_318
timestamp 1666464484
transform -1 0 36192 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_319
timestamp 1666464484
transform -1 0 36192 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_320
timestamp 1666464484
transform -1 0 36192 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_321
timestamp 1666464484
transform -1 0 36192 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_322
timestamp 1666464484
transform -1 0 36192 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_323
timestamp 1666464484
transform -1 0 36192 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_324
timestamp 1666464484
transform -1 0 36192 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_325
timestamp 1666464484
transform -1 0 36192 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_326
timestamp 1666464484
transform -1 0 36192 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_327
timestamp 1666464484
transform -1 0 36192 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_328
timestamp 1666464484
transform -1 0 36192 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_329
timestamp 1666464484
transform -1 0 36192 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_330
timestamp 1666464484
transform -1 0 36192 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_331
timestamp 1666464484
transform -1 0 36192 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_332
timestamp 1666464484
transform 1 0 36192 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_333
timestamp 1666464484
transform 1 0 36192 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_334
timestamp 1666464484
transform 1 0 36192 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_335
timestamp 1666464484
transform 1 0 36192 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_336
timestamp 1666464484
transform 1 0 36192 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_337
timestamp 1666464484
transform 1 0 36192 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_338
timestamp 1666464484
transform 1 0 36192 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_339
timestamp 1666464484
transform 1 0 36192 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_340
timestamp 1666464484
transform 1 0 36192 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_341
timestamp 1666464484
transform -1 0 39936 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_342
timestamp 1666464484
transform -1 0 39936 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_343
timestamp 1666464484
transform -1 0 39936 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_344
timestamp 1666464484
transform -1 0 39936 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_345
timestamp 1666464484
transform -1 0 39936 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_346
timestamp 1666464484
transform -1 0 39936 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_347
timestamp 1666464484
transform -1 0 39936 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_348
timestamp 1666464484
transform -1 0 39936 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_349
timestamp 1666464484
transform -1 0 39936 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_350
timestamp 1666464484
transform -1 0 39936 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_351
timestamp 1666464484
transform -1 0 39936 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_352
timestamp 1666464484
transform -1 0 39936 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_353
timestamp 1666464484
transform -1 0 39936 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_354
timestamp 1666464484
transform -1 0 39936 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_355
timestamp 1666464484
transform 1 0 36192 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_356
timestamp 1666464484
transform 1 0 36192 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_357
timestamp 1666464484
transform 1 0 36192 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_358
timestamp 1666464484
transform 1 0 36192 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_359
timestamp 1666464484
transform 1 0 36192 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_360
timestamp 1666464484
transform -1 0 38688 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_361
timestamp 1666464484
transform -1 0 38688 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_362
timestamp 1666464484
transform -1 0 37440 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_363
timestamp 1666464484
transform -1 0 37440 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_364
timestamp 1666464484
transform -1 0 37440 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_365
timestamp 1666464484
transform -1 0 37440 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_366
timestamp 1666464484
transform -1 0 37440 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_367
timestamp 1666464484
transform -1 0 37440 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_368
timestamp 1666464484
transform -1 0 37440 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_369
timestamp 1666464484
transform -1 0 37440 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_370
timestamp 1666464484
transform -1 0 37440 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_371
timestamp 1666464484
transform -1 0 37440 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_372
timestamp 1666464484
transform -1 0 37440 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_373
timestamp 1666464484
transform -1 0 37440 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_374
timestamp 1666464484
transform -1 0 37440 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_375
timestamp 1666464484
transform -1 0 37440 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_376
timestamp 1666464484
transform -1 0 38688 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_377
timestamp 1666464484
transform -1 0 34944 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_378
timestamp 1666464484
transform -1 0 34944 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_379
timestamp 1666464484
transform -1 0 34944 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_380
timestamp 1666464484
transform -1 0 34944 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_381
timestamp 1666464484
transform -1 0 34944 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_382
timestamp 1666464484
transform -1 0 34944 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_383
timestamp 1666464484
transform -1 0 34944 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_384
timestamp 1666464484
transform -1 0 34944 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_385
timestamp 1666464484
transform -1 0 34944 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_386
timestamp 1666464484
transform -1 0 34944 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_387
timestamp 1666464484
transform -1 0 34944 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_388
timestamp 1666464484
transform 1 0 37440 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_389
timestamp 1666464484
transform 1 0 37440 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_390
timestamp 1666464484
transform -1 0 34944 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_391
timestamp 1666464484
transform -1 0 34944 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_392
timestamp 1666464484
transform -1 0 34944 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_393
timestamp 1666464484
transform -1 0 34944 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_394
timestamp 1666464484
transform -1 0 34944 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_395
timestamp 1666464484
transform -1 0 34944 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_396
timestamp 1666464484
transform -1 0 34944 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_397
timestamp 1666464484
transform -1 0 34944 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_398
timestamp 1666464484
transform -1 0 34944 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_399
timestamp 1666464484
transform -1 0 34944 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_400
timestamp 1666464484
transform -1 0 34944 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_401
timestamp 1666464484
transform -1 0 34944 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_402
timestamp 1666464484
transform -1 0 36192 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_403
timestamp 1666464484
transform -1 0 36192 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_404
timestamp 1666464484
transform -1 0 34944 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_405
timestamp 1666464484
transform -1 0 34944 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_406
timestamp 1666464484
transform -1 0 34944 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_407
timestamp 1666464484
transform -1 0 34944 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_408
timestamp 1666464484
transform -1 0 34944 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_409
timestamp 1666464484
transform -1 0 34944 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_410
timestamp 1666464484
transform -1 0 34944 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_411
timestamp 1666464484
transform -1 0 39936 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_412
timestamp 1666464484
transform -1 0 39936 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_413
timestamp 1666464484
transform -1 0 34944 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_414
timestamp 1666464484
transform 1 0 31200 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_415
timestamp 1666464484
transform 1 0 31200 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_416
timestamp 1666464484
transform 1 0 32448 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_417
timestamp 1666464484
transform 1 0 32448 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_418
timestamp 1666464484
transform -1 0 37440 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_419
timestamp 1666464484
transform -1 0 37440 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_420
timestamp 1666464484
transform -1 0 33696 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_421
timestamp 1666464484
transform -1 0 33696 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_422
timestamp 1666464484
transform 1 0 38688 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_423
timestamp 1666464484
transform 1 0 38688 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_424
timestamp 1666464484
transform 1 0 34944 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_425
timestamp 1666464484
transform 1 0 34944 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_426
timestamp 1666464484
transform 1 0 34944 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_427
timestamp 1666464484
transform 1 0 34944 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_428
timestamp 1666464484
transform 1 0 34944 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_429
timestamp 1666464484
transform 1 0 34944 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_430
timestamp 1666464484
transform 1 0 34944 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_431
timestamp 1666464484
transform 1 0 34944 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_432
timestamp 1666464484
transform 1 0 34944 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_433
timestamp 1666464484
transform 1 0 34944 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_434
timestamp 1666464484
transform 1 0 34944 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_435
timestamp 1666464484
transform 1 0 34944 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_436
timestamp 1666464484
transform 1 0 34944 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_437
timestamp 1666464484
transform 1 0 34944 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_438
timestamp 1666464484
transform 1 0 34944 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_439
timestamp 1666464484
transform 1 0 34944 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_440
timestamp 1666464484
transform 1 0 34944 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_441
timestamp 1666464484
transform 1 0 34944 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_442
timestamp 1666464484
transform 1 0 34944 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_443
timestamp 1666464484
transform 1 0 34944 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_444
timestamp 1666464484
transform 1 0 34944 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_445
timestamp 1666464484
transform 1 0 34944 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_446
timestamp 1666464484
transform 1 0 34944 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_447
timestamp 1666464484
transform 1 0 34944 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_448
timestamp 1666464484
transform 1 0 34944 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_449
timestamp 1666464484
transform 1 0 34944 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_450
timestamp 1666464484
transform 1 0 34944 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_451
timestamp 1666464484
transform 1 0 34944 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_452
timestamp 1666464484
transform 1 0 34944 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_453
timestamp 1666464484
transform 1 0 34944 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_454
timestamp 1666464484
transform 1 0 34944 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_455
timestamp 1666464484
transform -1 0 32448 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_456
timestamp 1666464484
transform -1 0 32448 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_457
timestamp 1666464484
transform 1 0 33696 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_458
timestamp 1666464484
transform 1 0 36192 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_459
timestamp 1666464484
transform 1 0 36192 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_460
timestamp 1666464484
transform -1 0 38688 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_461
timestamp 1666464484
transform -1 0 38688 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_462
timestamp 1666464484
transform 1 0 33696 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_463
timestamp 1666464484
transform -1 0 31200 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_464
timestamp 1666464484
transform -1 0 31200 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_465
timestamp 1666464484
transform -1 0 26208 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_466
timestamp 1666464484
transform -1 0 26208 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_467
timestamp 1666464484
transform -1 0 26208 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_468
timestamp 1666464484
transform -1 0 26208 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_469
timestamp 1666464484
transform -1 0 26208 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_470
timestamp 1666464484
transform -1 0 26208 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_471
timestamp 1666464484
transform 1 0 27456 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_472
timestamp 1666464484
transform 1 0 27456 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_473
timestamp 1666464484
transform -1 0 27456 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_474
timestamp 1666464484
transform -1 0 27456 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_475
timestamp 1666464484
transform -1 0 27456 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_476
timestamp 1666464484
transform -1 0 26208 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_477
timestamp 1666464484
transform -1 0 27456 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_478
timestamp 1666464484
transform -1 0 27456 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_479
timestamp 1666464484
transform -1 0 27456 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_480
timestamp 1666464484
transform -1 0 27456 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_481
timestamp 1666464484
transform -1 0 27456 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_482
timestamp 1666464484
transform -1 0 27456 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_483
timestamp 1666464484
transform -1 0 27456 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_484
timestamp 1666464484
transform 1 0 27456 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_485
timestamp 1666464484
transform -1 0 28704 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_486
timestamp 1666464484
transform -1 0 28704 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_487
timestamp 1666464484
transform -1 0 28704 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_488
timestamp 1666464484
transform -1 0 28704 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_489
timestamp 1666464484
transform -1 0 28704 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_490
timestamp 1666464484
transform 1 0 26208 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_491
timestamp 1666464484
transform 1 0 26208 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_492
timestamp 1666464484
transform 1 0 26208 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_493
timestamp 1666464484
transform -1 0 28704 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_494
timestamp 1666464484
transform -1 0 28704 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_495
timestamp 1666464484
transform -1 0 28704 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_496
timestamp 1666464484
transform -1 0 28704 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_497
timestamp 1666464484
transform -1 0 28704 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_498
timestamp 1666464484
transform -1 0 26208 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_499
timestamp 1666464484
transform -1 0 26208 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_500
timestamp 1666464484
transform 1 0 26208 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_501
timestamp 1666464484
transform 1 0 26208 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_502
timestamp 1666464484
transform 1 0 26208 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_503
timestamp 1666464484
transform 1 0 26208 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_504
timestamp 1666464484
transform 1 0 26208 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_505
timestamp 1666464484
transform 1 0 26208 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_506
timestamp 1666464484
transform 1 0 26208 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_507
timestamp 1666464484
transform 1 0 27456 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_508
timestamp 1666464484
transform 1 0 27456 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_509
timestamp 1666464484
transform 1 0 26208 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_510
timestamp 1666464484
transform 1 0 26208 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_511
timestamp 1666464484
transform 1 0 26208 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_512
timestamp 1666464484
transform -1 0 27456 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_513
timestamp 1666464484
transform -1 0 27456 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_514
timestamp 1666464484
transform -1 0 27456 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_515
timestamp 1666464484
transform -1 0 27456 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_516
timestamp 1666464484
transform -1 0 27456 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_517
timestamp 1666464484
transform 1 0 26208 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_518
timestamp 1666464484
transform 1 0 26208 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_519
timestamp 1666464484
transform -1 0 26208 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_520
timestamp 1666464484
transform -1 0 26208 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_521
timestamp 1666464484
transform -1 0 26208 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_522
timestamp 1666464484
transform -1 0 26208 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_523
timestamp 1666464484
transform -1 0 26208 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_524
timestamp 1666464484
transform -1 0 26208 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_525
timestamp 1666464484
transform -1 0 28704 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_526
timestamp 1666464484
transform -1 0 28704 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_527
timestamp 1666464484
transform -1 0 28704 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_528
timestamp 1666464484
transform 1 0 28704 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_529
timestamp 1666464484
transform 1 0 28704 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_530
timestamp 1666464484
transform 1 0 28704 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_531
timestamp 1666464484
transform 1 0 28704 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_532
timestamp 1666464484
transform 1 0 28704 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_533
timestamp 1666464484
transform 1 0 28704 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_534
timestamp 1666464484
transform 1 0 28704 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_535
timestamp 1666464484
transform 1 0 28704 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_536
timestamp 1666464484
transform 1 0 28704 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_537
timestamp 1666464484
transform 1 0 28704 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_538
timestamp 1666464484
transform 1 0 28704 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_539
timestamp 1666464484
transform 1 0 28704 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_540
timestamp 1666464484
transform 1 0 28704 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_541
timestamp 1666464484
transform 1 0 28704 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_542
timestamp 1666464484
transform 1 0 28704 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_543
timestamp 1666464484
transform -1 0 28704 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_544
timestamp 1666464484
transform -1 0 28704 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_545
timestamp 1666464484
transform 1 0 27456 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_546
timestamp 1666464484
transform 1 0 27456 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_547
timestamp 1666464484
transform 1 0 27456 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_548
timestamp 1666464484
transform 1 0 27456 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_549
timestamp 1666464484
transform 1 0 27456 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_550
timestamp 1666464484
transform 1 0 27456 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_551
timestamp 1666464484
transform 1 0 27456 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_552
timestamp 1666464484
transform 1 0 27456 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_553
timestamp 1666464484
transform 1 0 27456 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_554
timestamp 1666464484
transform 1 0 27456 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_555
timestamp 1666464484
transform -1 0 22464 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_556
timestamp 1666464484
transform -1 0 22464 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_557
timestamp 1666464484
transform -1 0 22464 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_558
timestamp 1666464484
transform -1 0 22464 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_559
timestamp 1666464484
transform -1 0 22464 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_560
timestamp 1666464484
transform -1 0 22464 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_561
timestamp 1666464484
transform -1 0 22464 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_562
timestamp 1666464484
transform -1 0 22464 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_563
timestamp 1666464484
transform 1 0 22464 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_564
timestamp 1666464484
transform 1 0 22464 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_565
timestamp 1666464484
transform 1 0 22464 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_566
timestamp 1666464484
transform 1 0 22464 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_567
timestamp 1666464484
transform -1 0 21216 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_568
timestamp 1666464484
transform -1 0 21216 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_569
timestamp 1666464484
transform 1 0 23712 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_570
timestamp 1666464484
transform 1 0 23712 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_571
timestamp 1666464484
transform 1 0 23712 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_572
timestamp 1666464484
transform 1 0 23712 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_573
timestamp 1666464484
transform -1 0 22464 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_574
timestamp 1666464484
transform 1 0 21216 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_575
timestamp 1666464484
transform 1 0 21216 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_576
timestamp 1666464484
transform 1 0 21216 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_577
timestamp 1666464484
transform 1 0 21216 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_578
timestamp 1666464484
transform -1 0 23712 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_579
timestamp 1666464484
transform 1 0 21216 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_580
timestamp 1666464484
transform -1 0 23712 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_581
timestamp 1666464484
transform 1 0 21216 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_582
timestamp 1666464484
transform 1 0 21216 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_583
timestamp 1666464484
transform -1 0 23712 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_584
timestamp 1666464484
transform -1 0 23712 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_585
timestamp 1666464484
transform -1 0 23712 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_586
timestamp 1666464484
transform -1 0 23712 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_587
timestamp 1666464484
transform -1 0 23712 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_588
timestamp 1666464484
transform -1 0 23712 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_589
timestamp 1666464484
transform -1 0 23712 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_590
timestamp 1666464484
transform -1 0 23712 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_591
timestamp 1666464484
transform -1 0 23712 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_592
timestamp 1666464484
transform -1 0 23712 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_593
timestamp 1666464484
transform -1 0 23712 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_594
timestamp 1666464484
transform 1 0 23712 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_595
timestamp 1666464484
transform -1 0 21216 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_596
timestamp 1666464484
transform -1 0 21216 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_597
timestamp 1666464484
transform -1 0 21216 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_598
timestamp 1666464484
transform -1 0 21216 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_599
timestamp 1666464484
transform -1 0 21216 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_600
timestamp 1666464484
transform -1 0 21216 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_601
timestamp 1666464484
transform -1 0 21216 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_602
timestamp 1666464484
transform -1 0 21216 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_603
timestamp 1666464484
transform 1 0 22464 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_604
timestamp 1666464484
transform 1 0 22464 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_605
timestamp 1666464484
transform -1 0 21216 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_606
timestamp 1666464484
transform -1 0 23712 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_607
timestamp 1666464484
transform -1 0 23712 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_608
timestamp 1666464484
transform -1 0 22464 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_609
timestamp 1666464484
transform -1 0 22464 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_610
timestamp 1666464484
transform -1 0 22464 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_611
timestamp 1666464484
transform 1 0 22464 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_612
timestamp 1666464484
transform 1 0 22464 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_613
timestamp 1666464484
transform 1 0 22464 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_614
timestamp 1666464484
transform 1 0 22464 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_615
timestamp 1666464484
transform 1 0 22464 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_616
timestamp 1666464484
transform 1 0 22464 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_617
timestamp 1666464484
transform 1 0 22464 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_618
timestamp 1666464484
transform 1 0 22464 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_619
timestamp 1666464484
transform 1 0 22464 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_620
timestamp 1666464484
transform 1 0 23712 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_621
timestamp 1666464484
transform 1 0 23712 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_622
timestamp 1666464484
transform 1 0 23712 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_623
timestamp 1666464484
transform 1 0 23712 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_624
timestamp 1666464484
transform 1 0 23712 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_625
timestamp 1666464484
transform 1 0 23712 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_626
timestamp 1666464484
transform 1 0 23712 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_627
timestamp 1666464484
transform 1 0 23712 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_628
timestamp 1666464484
transform 1 0 23712 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_629
timestamp 1666464484
transform 1 0 23712 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_630
timestamp 1666464484
transform 1 0 21216 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_631
timestamp 1666464484
transform 1 0 21216 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_632
timestamp 1666464484
transform 1 0 21216 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_633
timestamp 1666464484
transform 1 0 21216 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_634
timestamp 1666464484
transform 1 0 21216 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_635
timestamp 1666464484
transform 1 0 21216 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_636
timestamp 1666464484
transform -1 0 22464 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_637
timestamp 1666464484
transform 1 0 21216 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_638
timestamp 1666464484
transform 1 0 21216 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_639
timestamp 1666464484
transform -1 0 21216 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_640
timestamp 1666464484
transform -1 0 21216 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_641
timestamp 1666464484
transform -1 0 21216 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_642
timestamp 1666464484
transform -1 0 21216 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_643
timestamp 1666464484
transform -1 0 22464 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_644
timestamp 1666464484
transform -1 0 22464 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_645
timestamp 1666464484
transform -1 0 23712 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_646
timestamp 1666464484
transform -1 0 23712 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_647
timestamp 1666464484
transform -1 0 23712 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_648
timestamp 1666464484
transform -1 0 23712 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_649
timestamp 1666464484
transform -1 0 23712 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_650
timestamp 1666464484
transform -1 0 23712 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_651
timestamp 1666464484
transform -1 0 23712 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_652
timestamp 1666464484
transform -1 0 23712 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_653
timestamp 1666464484
transform -1 0 23712 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_654
timestamp 1666464484
transform -1 0 23712 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_655
timestamp 1666464484
transform -1 0 23712 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_656
timestamp 1666464484
transform 1 0 23712 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_657
timestamp 1666464484
transform 1 0 23712 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_658
timestamp 1666464484
transform 1 0 23712 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_659
timestamp 1666464484
transform 1 0 23712 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_660
timestamp 1666464484
transform -1 0 22464 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_661
timestamp 1666464484
transform -1 0 22464 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_662
timestamp 1666464484
transform -1 0 22464 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_663
timestamp 1666464484
transform -1 0 22464 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_664
timestamp 1666464484
transform -1 0 22464 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_665
timestamp 1666464484
transform -1 0 22464 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_666
timestamp 1666464484
transform -1 0 22464 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_667
timestamp 1666464484
transform -1 0 22464 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_668
timestamp 1666464484
transform -1 0 21216 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_669
timestamp 1666464484
transform -1 0 22464 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_670
timestamp 1666464484
transform -1 0 22464 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_671
timestamp 1666464484
transform -1 0 22464 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_672
timestamp 1666464484
transform -1 0 22464 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_673
timestamp 1666464484
transform -1 0 22464 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_674
timestamp 1666464484
transform 1 0 22464 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_675
timestamp 1666464484
transform 1 0 22464 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_676
timestamp 1666464484
transform -1 0 23712 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_677
timestamp 1666464484
transform -1 0 23712 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_678
timestamp 1666464484
transform 1 0 22464 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_679
timestamp 1666464484
transform 1 0 21216 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_680
timestamp 1666464484
transform 1 0 21216 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_681
timestamp 1666464484
transform 1 0 21216 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_682
timestamp 1666464484
transform 1 0 21216 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_683
timestamp 1666464484
transform 1 0 21216 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_684
timestamp 1666464484
transform 1 0 21216 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_685
timestamp 1666464484
transform 1 0 21216 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_686
timestamp 1666464484
transform 1 0 21216 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_687
timestamp 1666464484
transform 1 0 21216 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_688
timestamp 1666464484
transform 1 0 21216 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_689
timestamp 1666464484
transform 1 0 21216 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_690
timestamp 1666464484
transform 1 0 22464 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_691
timestamp 1666464484
transform 1 0 22464 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_692
timestamp 1666464484
transform 1 0 22464 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_693
timestamp 1666464484
transform 1 0 22464 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_694
timestamp 1666464484
transform 1 0 22464 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_695
timestamp 1666464484
transform 1 0 22464 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_696
timestamp 1666464484
transform 1 0 22464 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_697
timestamp 1666464484
transform 1 0 22464 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_698
timestamp 1666464484
transform 1 0 22464 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_699
timestamp 1666464484
transform 1 0 23712 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_700
timestamp 1666464484
transform 1 0 23712 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_701
timestamp 1666464484
transform 1 0 23712 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_702
timestamp 1666464484
transform -1 0 23712 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_703
timestamp 1666464484
transform 1 0 23712 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_704
timestamp 1666464484
transform 1 0 23712 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_705
timestamp 1666464484
transform 1 0 23712 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_706
timestamp 1666464484
transform -1 0 21216 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_707
timestamp 1666464484
transform -1 0 21216 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_708
timestamp 1666464484
transform -1 0 21216 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_709
timestamp 1666464484
transform -1 0 21216 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_710
timestamp 1666464484
transform -1 0 21216 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_711
timestamp 1666464484
transform -1 0 21216 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_712
timestamp 1666464484
transform -1 0 21216 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_713
timestamp 1666464484
transform -1 0 21216 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_714
timestamp 1666464484
transform -1 0 21216 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_715
timestamp 1666464484
transform -1 0 21216 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_716
timestamp 1666464484
transform -1 0 21216 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_717
timestamp 1666464484
transform -1 0 21216 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_718
timestamp 1666464484
transform -1 0 21216 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_719
timestamp 1666464484
transform 1 0 23712 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_720
timestamp 1666464484
transform 1 0 23712 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_721
timestamp 1666464484
transform 1 0 21216 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_722
timestamp 1666464484
transform 1 0 21216 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_723
timestamp 1666464484
transform 1 0 21216 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_724
timestamp 1666464484
transform 1 0 23712 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_725
timestamp 1666464484
transform 1 0 23712 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_726
timestamp 1666464484
transform 1 0 22464 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_727
timestamp 1666464484
transform 1 0 22464 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_728
timestamp 1666464484
transform -1 0 22464 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_729
timestamp 1666464484
transform 1 0 26208 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_730
timestamp 1666464484
transform 1 0 26208 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_731
timestamp 1666464484
transform 1 0 28704 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_732
timestamp 1666464484
transform 1 0 28704 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_733
timestamp 1666464484
transform 1 0 28704 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_734
timestamp 1666464484
transform 1 0 28704 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_735
timestamp 1666464484
transform 1 0 28704 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_736
timestamp 1666464484
transform 1 0 26208 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_737
timestamp 1666464484
transform 1 0 26208 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_738
timestamp 1666464484
transform 1 0 26208 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_739
timestamp 1666464484
transform 1 0 26208 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_740
timestamp 1666464484
transform 1 0 26208 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_741
timestamp 1666464484
transform 1 0 26208 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_742
timestamp 1666464484
transform 1 0 26208 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_743
timestamp 1666464484
transform 1 0 26208 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_744
timestamp 1666464484
transform 1 0 26208 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_745
timestamp 1666464484
transform 1 0 26208 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_746
timestamp 1666464484
transform 1 0 26208 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_747
timestamp 1666464484
transform -1 0 27456 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_748
timestamp 1666464484
transform -1 0 27456 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_749
timestamp 1666464484
transform -1 0 27456 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_750
timestamp 1666464484
transform -1 0 28704 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_751
timestamp 1666464484
transform 1 0 27456 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_752
timestamp 1666464484
transform 1 0 27456 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_753
timestamp 1666464484
transform 1 0 27456 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_754
timestamp 1666464484
transform 1 0 27456 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_755
timestamp 1666464484
transform 1 0 27456 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_756
timestamp 1666464484
transform 1 0 27456 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_757
timestamp 1666464484
transform 1 0 27456 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_758
timestamp 1666464484
transform 1 0 27456 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_759
timestamp 1666464484
transform 1 0 27456 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_760
timestamp 1666464484
transform -1 0 28704 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_761
timestamp 1666464484
transform 1 0 28704 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_762
timestamp 1666464484
transform 1 0 28704 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_763
timestamp 1666464484
transform 1 0 28704 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_764
timestamp 1666464484
transform 1 0 28704 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_765
timestamp 1666464484
transform 1 0 28704 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_766
timestamp 1666464484
transform 1 0 28704 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_767
timestamp 1666464484
transform 1 0 28704 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_768
timestamp 1666464484
transform 1 0 28704 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_769
timestamp 1666464484
transform 1 0 28704 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_770
timestamp 1666464484
transform -1 0 28704 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_771
timestamp 1666464484
transform -1 0 28704 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_772
timestamp 1666464484
transform -1 0 28704 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_773
timestamp 1666464484
transform -1 0 28704 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_774
timestamp 1666464484
transform 1 0 27456 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_775
timestamp 1666464484
transform 1 0 27456 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_776
timestamp 1666464484
transform 1 0 27456 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_777
timestamp 1666464484
transform 1 0 27456 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_778
timestamp 1666464484
transform 1 0 27456 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_779
timestamp 1666464484
transform -1 0 27456 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_780
timestamp 1666464484
transform -1 0 27456 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_781
timestamp 1666464484
transform -1 0 27456 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_782
timestamp 1666464484
transform -1 0 27456 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_783
timestamp 1666464484
transform -1 0 27456 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_784
timestamp 1666464484
transform -1 0 27456 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_785
timestamp 1666464484
transform -1 0 27456 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_786
timestamp 1666464484
transform -1 0 27456 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_787
timestamp 1666464484
transform -1 0 26208 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_788
timestamp 1666464484
transform -1 0 26208 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_789
timestamp 1666464484
transform -1 0 26208 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_790
timestamp 1666464484
transform -1 0 26208 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_791
timestamp 1666464484
transform -1 0 26208 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_792
timestamp 1666464484
transform -1 0 26208 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_793
timestamp 1666464484
transform -1 0 26208 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_794
timestamp 1666464484
transform -1 0 26208 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_795
timestamp 1666464484
transform -1 0 27456 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_796
timestamp 1666464484
transform 1 0 26208 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_797
timestamp 1666464484
transform -1 0 27456 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_798
timestamp 1666464484
transform -1 0 27456 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_799
timestamp 1666464484
transform -1 0 28704 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_800
timestamp 1666464484
transform -1 0 28704 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_801
timestamp 1666464484
transform -1 0 28704 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_802
timestamp 1666464484
transform -1 0 28704 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_803
timestamp 1666464484
transform -1 0 28704 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_804
timestamp 1666464484
transform -1 0 26208 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_805
timestamp 1666464484
transform -1 0 26208 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_806
timestamp 1666464484
transform -1 0 26208 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_807
timestamp 1666464484
transform -1 0 26208 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_808
timestamp 1666464484
transform -1 0 26208 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_809
timestamp 1666464484
transform -1 0 26208 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_810
timestamp 1666464484
transform -1 0 28704 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_811
timestamp 1666464484
transform -1 0 28704 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_812
timestamp 1666464484
transform -1 0 28704 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_813
timestamp 1666464484
transform -1 0 27456 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_814
timestamp 1666464484
transform -1 0 27456 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_815
timestamp 1666464484
transform 1 0 28704 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_816
timestamp 1666464484
transform 1 0 28704 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_817
timestamp 1666464484
transform 1 0 22464 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_818
timestamp 1666464484
transform 1 0 22464 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_819
timestamp 1666464484
transform 1 0 27456 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_820
timestamp 1666464484
transform 1 0 27456 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_821
timestamp 1666464484
transform -1 0 21216 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_822
timestamp 1666464484
transform -1 0 21216 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_823
timestamp 1666464484
transform 1 0 21216 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_824
timestamp 1666464484
transform 1 0 21216 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_825
timestamp 1666464484
transform -1 0 24960 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_826
timestamp 1666464484
transform -1 0 24960 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_827
timestamp 1666464484
transform -1 0 24960 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_828
timestamp 1666464484
transform -1 0 24960 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_829
timestamp 1666464484
transform -1 0 24960 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_830
timestamp 1666464484
transform -1 0 24960 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_831
timestamp 1666464484
transform -1 0 24960 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_832
timestamp 1666464484
transform -1 0 24960 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_833
timestamp 1666464484
transform -1 0 24960 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_834
timestamp 1666464484
transform -1 0 24960 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_835
timestamp 1666464484
transform -1 0 24960 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_836
timestamp 1666464484
transform -1 0 24960 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_837
timestamp 1666464484
transform -1 0 24960 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_838
timestamp 1666464484
transform -1 0 24960 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_839
timestamp 1666464484
transform -1 0 24960 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_840
timestamp 1666464484
transform -1 0 24960 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_841
timestamp 1666464484
transform -1 0 24960 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_842
timestamp 1666464484
transform -1 0 24960 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_843
timestamp 1666464484
transform -1 0 24960 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_844
timestamp 1666464484
transform 1 0 24960 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_845
timestamp 1666464484
transform 1 0 24960 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_846
timestamp 1666464484
transform 1 0 24960 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_847
timestamp 1666464484
transform 1 0 24960 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_848
timestamp 1666464484
transform 1 0 24960 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_849
timestamp 1666464484
transform 1 0 24960 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_850
timestamp 1666464484
transform 1 0 24960 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_851
timestamp 1666464484
transform 1 0 24960 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_852
timestamp 1666464484
transform 1 0 24960 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_853
timestamp 1666464484
transform 1 0 24960 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_854
timestamp 1666464484
transform 1 0 24960 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_855
timestamp 1666464484
transform 1 0 24960 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_856
timestamp 1666464484
transform 1 0 24960 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_857
timestamp 1666464484
transform 1 0 24960 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_858
timestamp 1666464484
transform 1 0 24960 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_859
timestamp 1666464484
transform 1 0 24960 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_860
timestamp 1666464484
transform 1 0 24960 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_861
timestamp 1666464484
transform -1 0 26208 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_862
timestamp 1666464484
transform 1 0 26208 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_863
timestamp 1666464484
transform 1 0 26208 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_864
timestamp 1666464484
transform -1 0 28704 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_865
timestamp 1666464484
transform -1 0 28704 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_866
timestamp 1666464484
transform -1 0 24960 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_867
timestamp 1666464484
transform -1 0 24960 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_868
timestamp 1666464484
transform -1 0 24960 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_869
timestamp 1666464484
transform -1 0 24960 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_870
timestamp 1666464484
transform -1 0 24960 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_871
timestamp 1666464484
transform -1 0 24960 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_872
timestamp 1666464484
transform -1 0 24960 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_873
timestamp 1666464484
transform -1 0 24960 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_874
timestamp 1666464484
transform -1 0 24960 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_875
timestamp 1666464484
transform -1 0 24960 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_876
timestamp 1666464484
transform -1 0 24960 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_877
timestamp 1666464484
transform -1 0 24960 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_878
timestamp 1666464484
transform 1 0 24960 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_879
timestamp 1666464484
transform 1 0 24960 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_880
timestamp 1666464484
transform 1 0 24960 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_881
timestamp 1666464484
transform 1 0 24960 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_882
timestamp 1666464484
transform 1 0 24960 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_883
timestamp 1666464484
transform 1 0 24960 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_884
timestamp 1666464484
transform 1 0 24960 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_885
timestamp 1666464484
transform 1 0 24960 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_886
timestamp 1666464484
transform 1 0 24960 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_887
timestamp 1666464484
transform 1 0 24960 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_888
timestamp 1666464484
transform 1 0 24960 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_889
timestamp 1666464484
transform 1 0 24960 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_890
timestamp 1666464484
transform 1 0 24960 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_891
timestamp 1666464484
transform 1 0 24960 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_892
timestamp 1666464484
transform 1 0 23712 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_893
timestamp 1666464484
transform 1 0 23712 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_894
timestamp 1666464484
transform -1 0 22464 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_895
timestamp 1666464484
transform -1 0 22464 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_896
timestamp 1666464484
transform -1 0 23712 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_897
timestamp 1666464484
transform -1 0 23712 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_898
timestamp 1666464484
transform -1 0 26208 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_899
timestamp 1666464484
transform -1 0 26208 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_900
timestamp 1666464484
transform 1 0 28704 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_901
timestamp 1666464484
transform 1 0 28704 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_902
timestamp 1666464484
transform -1 0 26208 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_903
timestamp 1666464484
transform -1 0 26208 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_904
timestamp 1666464484
transform -1 0 26208 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_905
timestamp 1666464484
transform -1 0 26208 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_906
timestamp 1666464484
transform -1 0 26208 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_907
timestamp 1666464484
transform -1 0 26208 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_908
timestamp 1666464484
transform -1 0 26208 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_909
timestamp 1666464484
transform -1 0 26208 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_910
timestamp 1666464484
transform -1 0 26208 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_911
timestamp 1666464484
transform -1 0 26208 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_912
timestamp 1666464484
transform -1 0 26208 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_913
timestamp 1666464484
transform -1 0 26208 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_914
timestamp 1666464484
transform 1 0 28704 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_915
timestamp 1666464484
transform 1 0 28704 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_916
timestamp 1666464484
transform 1 0 28704 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_917
timestamp 1666464484
transform -1 0 28704 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_918
timestamp 1666464484
transform -1 0 28704 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_919
timestamp 1666464484
transform -1 0 28704 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_920
timestamp 1666464484
transform -1 0 28704 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_921
timestamp 1666464484
transform -1 0 28704 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_922
timestamp 1666464484
transform -1 0 28704 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_923
timestamp 1666464484
transform -1 0 28704 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_924
timestamp 1666464484
transform -1 0 28704 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_925
timestamp 1666464484
transform -1 0 28704 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_926
timestamp 1666464484
transform -1 0 28704 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_927
timestamp 1666464484
transform -1 0 28704 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_928
timestamp 1666464484
transform -1 0 28704 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_929
timestamp 1666464484
transform -1 0 28704 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_930
timestamp 1666464484
transform -1 0 28704 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_931
timestamp 1666464484
transform 1 0 28704 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_932
timestamp 1666464484
transform -1 0 27456 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_933
timestamp 1666464484
transform -1 0 27456 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_934
timestamp 1666464484
transform -1 0 27456 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_935
timestamp 1666464484
transform -1 0 27456 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_936
timestamp 1666464484
transform -1 0 27456 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_937
timestamp 1666464484
transform -1 0 27456 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_938
timestamp 1666464484
transform -1 0 27456 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_939
timestamp 1666464484
transform -1 0 27456 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_940
timestamp 1666464484
transform -1 0 27456 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_941
timestamp 1666464484
transform 1 0 28704 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_942
timestamp 1666464484
transform 1 0 28704 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_943
timestamp 1666464484
transform 1 0 28704 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_944
timestamp 1666464484
transform 1 0 28704 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_945
timestamp 1666464484
transform 1 0 28704 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_946
timestamp 1666464484
transform 1 0 27456 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_947
timestamp 1666464484
transform 1 0 27456 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_948
timestamp 1666464484
transform 1 0 27456 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_949
timestamp 1666464484
transform 1 0 27456 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_950
timestamp 1666464484
transform 1 0 27456 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_951
timestamp 1666464484
transform 1 0 27456 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_952
timestamp 1666464484
transform 1 0 27456 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_953
timestamp 1666464484
transform 1 0 27456 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_954
timestamp 1666464484
transform 1 0 27456 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_955
timestamp 1666464484
transform 1 0 27456 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_956
timestamp 1666464484
transform 1 0 27456 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_957
timestamp 1666464484
transform 1 0 27456 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_958
timestamp 1666464484
transform 1 0 26208 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_959
timestamp 1666464484
transform 1 0 26208 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_960
timestamp 1666464484
transform 1 0 26208 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_961
timestamp 1666464484
transform 1 0 26208 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_962
timestamp 1666464484
transform 1 0 26208 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_963
timestamp 1666464484
transform 1 0 26208 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_964
timestamp 1666464484
transform 1 0 26208 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_965
timestamp 1666464484
transform 1 0 27456 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_966
timestamp 1666464484
transform 1 0 27456 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_967
timestamp 1666464484
transform -1 0 27456 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_968
timestamp 1666464484
transform -1 0 27456 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_969
timestamp 1666464484
transform -1 0 27456 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_970
timestamp 1666464484
transform -1 0 27456 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_971
timestamp 1666464484
transform -1 0 27456 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_972
timestamp 1666464484
transform 1 0 26208 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_973
timestamp 1666464484
transform 1 0 26208 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_974
timestamp 1666464484
transform 1 0 26208 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_975
timestamp 1666464484
transform 1 0 26208 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_976
timestamp 1666464484
transform 1 0 26208 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_977
timestamp 1666464484
transform 1 0 26208 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_978
timestamp 1666464484
transform 1 0 26208 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_979
timestamp 1666464484
transform 1 0 28704 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_980
timestamp 1666464484
transform 1 0 28704 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_981
timestamp 1666464484
transform 1 0 28704 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_982
timestamp 1666464484
transform -1 0 26208 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_983
timestamp 1666464484
transform 1 0 21216 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_984
timestamp 1666464484
transform -1 0 22464 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_985
timestamp 1666464484
transform -1 0 22464 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_986
timestamp 1666464484
transform 1 0 23712 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_987
timestamp 1666464484
transform 1 0 23712 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_988
timestamp 1666464484
transform 1 0 22464 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_989
timestamp 1666464484
transform 1 0 22464 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_990
timestamp 1666464484
transform 1 0 22464 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_991
timestamp 1666464484
transform 1 0 22464 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_992
timestamp 1666464484
transform 1 0 22464 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_993
timestamp 1666464484
transform 1 0 22464 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_994
timestamp 1666464484
transform 1 0 22464 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_995
timestamp 1666464484
transform 1 0 22464 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_996
timestamp 1666464484
transform 1 0 22464 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_997
timestamp 1666464484
transform 1 0 22464 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_998
timestamp 1666464484
transform -1 0 21216 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_999
timestamp 1666464484
transform -1 0 21216 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1000
timestamp 1666464484
transform -1 0 21216 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1001
timestamp 1666464484
transform -1 0 21216 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1002
timestamp 1666464484
transform -1 0 21216 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1003
timestamp 1666464484
transform -1 0 21216 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1004
timestamp 1666464484
transform -1 0 21216 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1005
timestamp 1666464484
transform -1 0 21216 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1006
timestamp 1666464484
transform -1 0 21216 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1007
timestamp 1666464484
transform -1 0 21216 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1008
timestamp 1666464484
transform -1 0 21216 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1009
timestamp 1666464484
transform -1 0 21216 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1010
timestamp 1666464484
transform -1 0 21216 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1011
timestamp 1666464484
transform -1 0 21216 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1012
timestamp 1666464484
transform 1 0 22464 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1013
timestamp 1666464484
transform 1 0 22464 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1014
timestamp 1666464484
transform 1 0 22464 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1015
timestamp 1666464484
transform 1 0 22464 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1016
timestamp 1666464484
transform 1 0 23712 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1017
timestamp 1666464484
transform 1 0 23712 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1018
timestamp 1666464484
transform 1 0 23712 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1019
timestamp 1666464484
transform 1 0 23712 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1020
timestamp 1666464484
transform 1 0 23712 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1021
timestamp 1666464484
transform 1 0 23712 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1022
timestamp 1666464484
transform 1 0 23712 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1023
timestamp 1666464484
transform 1 0 23712 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1024
timestamp 1666464484
transform -1 0 22464 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1025
timestamp 1666464484
transform 1 0 21216 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1026
timestamp 1666464484
transform 1 0 21216 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1027
timestamp 1666464484
transform 1 0 21216 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1028
timestamp 1666464484
transform -1 0 23712 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1029
timestamp 1666464484
transform -1 0 23712 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1030
timestamp 1666464484
transform -1 0 23712 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1031
timestamp 1666464484
transform 1 0 21216 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1032
timestamp 1666464484
transform 1 0 21216 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1033
timestamp 1666464484
transform 1 0 21216 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1034
timestamp 1666464484
transform 1 0 21216 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1035
timestamp 1666464484
transform 1 0 21216 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1036
timestamp 1666464484
transform 1 0 21216 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1037
timestamp 1666464484
transform 1 0 21216 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1038
timestamp 1666464484
transform 1 0 21216 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1039
timestamp 1666464484
transform -1 0 22464 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1040
timestamp 1666464484
transform -1 0 22464 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1041
timestamp 1666464484
transform 1 0 23712 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1042
timestamp 1666464484
transform 1 0 23712 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1043
timestamp 1666464484
transform 1 0 23712 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1044
timestamp 1666464484
transform 1 0 23712 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1045
timestamp 1666464484
transform -1 0 23712 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1046
timestamp 1666464484
transform -1 0 23712 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1047
timestamp 1666464484
transform -1 0 23712 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1048
timestamp 1666464484
transform -1 0 23712 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1049
timestamp 1666464484
transform -1 0 23712 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1050
timestamp 1666464484
transform -1 0 23712 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1051
timestamp 1666464484
transform -1 0 23712 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1052
timestamp 1666464484
transform -1 0 23712 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1053
timestamp 1666464484
transform -1 0 23712 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1054
timestamp 1666464484
transform -1 0 22464 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1055
timestamp 1666464484
transform -1 0 23712 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1056
timestamp 1666464484
transform -1 0 23712 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1057
timestamp 1666464484
transform -1 0 22464 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1058
timestamp 1666464484
transform -1 0 22464 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1059
timestamp 1666464484
transform -1 0 22464 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1060
timestamp 1666464484
transform -1 0 22464 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1061
timestamp 1666464484
transform -1 0 22464 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1062
timestamp 1666464484
transform -1 0 22464 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1063
timestamp 1666464484
transform -1 0 22464 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1064
timestamp 1666464484
transform -1 0 22464 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1065
timestamp 1666464484
transform 1 0 21216 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1066
timestamp 1666464484
transform 1 0 21216 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1067
timestamp 1666464484
transform -1 0 21216 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1068
timestamp 1666464484
transform -1 0 21216 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1069
timestamp 1666464484
transform -1 0 21216 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1070
timestamp 1666464484
transform -1 0 21216 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1071
timestamp 1666464484
transform -1 0 21216 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1072
timestamp 1666464484
transform -1 0 21216 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1073
timestamp 1666464484
transform -1 0 21216 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1074
timestamp 1666464484
transform -1 0 21216 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1075
timestamp 1666464484
transform -1 0 21216 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1076
timestamp 1666464484
transform -1 0 21216 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1077
timestamp 1666464484
transform -1 0 21216 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1078
timestamp 1666464484
transform -1 0 21216 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1079
timestamp 1666464484
transform -1 0 21216 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1080
timestamp 1666464484
transform -1 0 22464 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1081
timestamp 1666464484
transform -1 0 22464 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1082
timestamp 1666464484
transform -1 0 22464 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1083
timestamp 1666464484
transform -1 0 22464 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1084
timestamp 1666464484
transform -1 0 23712 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1085
timestamp 1666464484
transform -1 0 23712 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1086
timestamp 1666464484
transform -1 0 23712 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1087
timestamp 1666464484
transform -1 0 23712 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1088
timestamp 1666464484
transform -1 0 23712 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1089
timestamp 1666464484
transform 1 0 23712 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1090
timestamp 1666464484
transform 1 0 23712 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1091
timestamp 1666464484
transform 1 0 23712 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1092
timestamp 1666464484
transform 1 0 23712 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1093
timestamp 1666464484
transform 1 0 23712 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1094
timestamp 1666464484
transform 1 0 23712 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1095
timestamp 1666464484
transform 1 0 23712 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1096
timestamp 1666464484
transform 1 0 23712 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1097
timestamp 1666464484
transform -1 0 21216 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1098
timestamp 1666464484
transform 1 0 23712 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1099
timestamp 1666464484
transform 1 0 23712 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1100
timestamp 1666464484
transform 1 0 23712 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1101
timestamp 1666464484
transform 1 0 23712 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1102
timestamp 1666464484
transform 1 0 23712 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1103
timestamp 1666464484
transform 1 0 22464 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1104
timestamp 1666464484
transform 1 0 21216 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1105
timestamp 1666464484
transform 1 0 21216 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1106
timestamp 1666464484
transform 1 0 21216 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1107
timestamp 1666464484
transform 1 0 21216 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1108
timestamp 1666464484
transform 1 0 21216 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1109
timestamp 1666464484
transform 1 0 21216 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1110
timestamp 1666464484
transform 1 0 21216 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1111
timestamp 1666464484
transform 1 0 21216 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1112
timestamp 1666464484
transform 1 0 22464 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1113
timestamp 1666464484
transform 1 0 22464 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1114
timestamp 1666464484
transform 1 0 22464 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1115
timestamp 1666464484
transform 1 0 22464 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1116
timestamp 1666464484
transform 1 0 22464 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1117
timestamp 1666464484
transform 1 0 22464 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1118
timestamp 1666464484
transform 1 0 22464 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1119
timestamp 1666464484
transform 1 0 22464 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1120
timestamp 1666464484
transform 1 0 22464 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1121
timestamp 1666464484
transform 1 0 22464 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1122
timestamp 1666464484
transform 1 0 22464 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1123
timestamp 1666464484
transform 1 0 21216 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1124
timestamp 1666464484
transform 1 0 21216 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1125
timestamp 1666464484
transform 1 0 21216 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1126
timestamp 1666464484
transform 1 0 21216 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1127
timestamp 1666464484
transform 1 0 21216 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1128
timestamp 1666464484
transform 1 0 21216 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1129
timestamp 1666464484
transform 1 0 22464 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1130
timestamp 1666464484
transform 1 0 22464 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1131
timestamp 1666464484
transform 1 0 23712 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1132
timestamp 1666464484
transform -1 0 23712 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1133
timestamp 1666464484
transform -1 0 23712 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1134
timestamp 1666464484
transform -1 0 23712 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1135
timestamp 1666464484
transform -1 0 23712 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1136
timestamp 1666464484
transform -1 0 23712 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1137
timestamp 1666464484
transform -1 0 23712 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1138
timestamp 1666464484
transform -1 0 23712 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1139
timestamp 1666464484
transform -1 0 23712 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1140
timestamp 1666464484
transform -1 0 23712 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1141
timestamp 1666464484
transform -1 0 22464 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1142
timestamp 1666464484
transform -1 0 22464 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1143
timestamp 1666464484
transform -1 0 22464 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1144
timestamp 1666464484
transform -1 0 22464 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1145
timestamp 1666464484
transform -1 0 22464 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1146
timestamp 1666464484
transform -1 0 22464 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1147
timestamp 1666464484
transform -1 0 22464 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1148
timestamp 1666464484
transform -1 0 22464 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1149
timestamp 1666464484
transform -1 0 22464 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1150
timestamp 1666464484
transform -1 0 22464 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1151
timestamp 1666464484
transform 1 0 27456 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1152
timestamp 1666464484
transform 1 0 27456 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1153
timestamp 1666464484
transform 1 0 27456 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1154
timestamp 1666464484
transform 1 0 28704 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1155
timestamp 1666464484
transform -1 0 26208 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1156
timestamp 1666464484
transform -1 0 26208 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1157
timestamp 1666464484
transform -1 0 26208 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1158
timestamp 1666464484
transform -1 0 26208 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1159
timestamp 1666464484
transform -1 0 26208 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1160
timestamp 1666464484
transform -1 0 26208 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1161
timestamp 1666464484
transform 1 0 28704 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1162
timestamp 1666464484
transform 1 0 26208 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1163
timestamp 1666464484
transform 1 0 26208 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1164
timestamp 1666464484
transform 1 0 26208 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1165
timestamp 1666464484
transform 1 0 26208 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1166
timestamp 1666464484
transform 1 0 28704 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1167
timestamp 1666464484
transform 1 0 28704 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1168
timestamp 1666464484
transform 1 0 28704 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1169
timestamp 1666464484
transform 1 0 28704 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1170
timestamp 1666464484
transform 1 0 28704 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1171
timestamp 1666464484
transform 1 0 26208 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1172
timestamp 1666464484
transform 1 0 26208 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1173
timestamp 1666464484
transform 1 0 26208 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1174
timestamp 1666464484
transform 1 0 26208 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1175
timestamp 1666464484
transform 1 0 26208 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1176
timestamp 1666464484
transform 1 0 26208 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1177
timestamp 1666464484
transform 1 0 26208 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1178
timestamp 1666464484
transform 1 0 26208 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1179
timestamp 1666464484
transform 1 0 26208 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1180
timestamp 1666464484
transform 1 0 26208 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1181
timestamp 1666464484
transform 1 0 28704 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1182
timestamp 1666464484
transform 1 0 28704 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1183
timestamp 1666464484
transform -1 0 27456 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1184
timestamp 1666464484
transform -1 0 27456 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1185
timestamp 1666464484
transform -1 0 27456 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1186
timestamp 1666464484
transform -1 0 27456 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1187
timestamp 1666464484
transform -1 0 27456 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1188
timestamp 1666464484
transform -1 0 27456 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1189
timestamp 1666464484
transform -1 0 27456 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1190
timestamp 1666464484
transform -1 0 27456 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1191
timestamp 1666464484
transform -1 0 27456 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1192
timestamp 1666464484
transform -1 0 27456 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1193
timestamp 1666464484
transform -1 0 27456 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1194
timestamp 1666464484
transform -1 0 27456 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1195
timestamp 1666464484
transform -1 0 27456 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1196
timestamp 1666464484
transform 1 0 28704 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1197
timestamp 1666464484
transform -1 0 26208 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1198
timestamp 1666464484
transform -1 0 26208 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1199
timestamp 1666464484
transform -1 0 26208 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1200
timestamp 1666464484
transform -1 0 26208 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1201
timestamp 1666464484
transform -1 0 27456 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1202
timestamp 1666464484
transform -1 0 26208 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1203
timestamp 1666464484
transform -1 0 28704 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1204
timestamp 1666464484
transform -1 0 28704 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1205
timestamp 1666464484
transform -1 0 28704 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1206
timestamp 1666464484
transform -1 0 28704 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1207
timestamp 1666464484
transform -1 0 28704 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1208
timestamp 1666464484
transform -1 0 28704 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1209
timestamp 1666464484
transform -1 0 28704 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1210
timestamp 1666464484
transform -1 0 28704 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1211
timestamp 1666464484
transform -1 0 28704 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1212
timestamp 1666464484
transform -1 0 28704 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1213
timestamp 1666464484
transform -1 0 28704 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1214
timestamp 1666464484
transform -1 0 28704 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1215
timestamp 1666464484
transform -1 0 28704 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1216
timestamp 1666464484
transform -1 0 28704 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1217
timestamp 1666464484
transform -1 0 26208 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1218
timestamp 1666464484
transform -1 0 26208 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1219
timestamp 1666464484
transform -1 0 26208 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1220
timestamp 1666464484
transform 1 0 28704 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1221
timestamp 1666464484
transform 1 0 28704 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1222
timestamp 1666464484
transform 1 0 28704 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1223
timestamp 1666464484
transform 1 0 28704 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1224
timestamp 1666464484
transform 1 0 27456 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1225
timestamp 1666464484
transform 1 0 27456 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1226
timestamp 1666464484
transform 1 0 27456 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1227
timestamp 1666464484
transform 1 0 27456 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1228
timestamp 1666464484
transform 1 0 27456 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1229
timestamp 1666464484
transform 1 0 27456 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1230
timestamp 1666464484
transform 1 0 27456 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1231
timestamp 1666464484
transform 1 0 27456 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1232
timestamp 1666464484
transform 1 0 27456 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1233
timestamp 1666464484
transform 1 0 27456 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1234
timestamp 1666464484
transform 1 0 27456 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1235
timestamp 1666464484
transform -1 0 21216 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1236
timestamp 1666464484
transform -1 0 21216 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1237
timestamp 1666464484
transform -1 0 24960 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1238
timestamp 1666464484
transform -1 0 24960 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1239
timestamp 1666464484
transform -1 0 24960 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1240
timestamp 1666464484
transform -1 0 24960 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1241
timestamp 1666464484
transform -1 0 24960 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1242
timestamp 1666464484
transform -1 0 24960 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1243
timestamp 1666464484
transform -1 0 24960 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1244
timestamp 1666464484
transform -1 0 24960 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1245
timestamp 1666464484
transform -1 0 24960 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1246
timestamp 1666464484
transform -1 0 24960 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1247
timestamp 1666464484
transform -1 0 24960 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1248
timestamp 1666464484
transform -1 0 24960 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1249
timestamp 1666464484
transform -1 0 24960 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1250
timestamp 1666464484
transform -1 0 24960 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1251
timestamp 1666464484
transform -1 0 24960 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1252
timestamp 1666464484
transform -1 0 24960 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1253
timestamp 1666464484
transform -1 0 24960 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1254
timestamp 1666464484
transform -1 0 24960 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1255
timestamp 1666464484
transform 1 0 26208 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1256
timestamp 1666464484
transform 1 0 26208 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1257
timestamp 1666464484
transform -1 0 24960 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1258
timestamp 1666464484
transform -1 0 24960 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1259
timestamp 1666464484
transform -1 0 24960 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1260
timestamp 1666464484
transform -1 0 24960 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1261
timestamp 1666464484
transform -1 0 24960 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1262
timestamp 1666464484
transform -1 0 27456 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1263
timestamp 1666464484
transform -1 0 28704 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1264
timestamp 1666464484
transform -1 0 28704 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1265
timestamp 1666464484
transform -1 0 27456 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1266
timestamp 1666464484
transform 1 0 24960 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1267
timestamp 1666464484
transform 1 0 24960 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1268
timestamp 1666464484
transform 1 0 24960 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1269
timestamp 1666464484
transform 1 0 24960 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1270
timestamp 1666464484
transform 1 0 24960 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1271
timestamp 1666464484
transform 1 0 24960 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1272
timestamp 1666464484
transform 1 0 24960 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1273
timestamp 1666464484
transform 1 0 24960 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1274
timestamp 1666464484
transform 1 0 24960 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1275
timestamp 1666464484
transform 1 0 24960 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1276
timestamp 1666464484
transform 1 0 24960 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1277
timestamp 1666464484
transform 1 0 24960 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1278
timestamp 1666464484
transform 1 0 24960 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1279
timestamp 1666464484
transform 1 0 24960 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1280
timestamp 1666464484
transform 1 0 24960 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1281
timestamp 1666464484
transform 1 0 24960 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1282
timestamp 1666464484
transform 1 0 24960 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1283
timestamp 1666464484
transform 1 0 24960 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1284
timestamp 1666464484
transform 1 0 24960 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1285
timestamp 1666464484
transform 1 0 24960 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1286
timestamp 1666464484
transform 1 0 24960 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1287
timestamp 1666464484
transform 1 0 24960 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1288
timestamp 1666464484
transform 1 0 24960 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1289
timestamp 1666464484
transform 1 0 24960 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1290
timestamp 1666464484
transform 1 0 24960 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1291
timestamp 1666464484
transform 1 0 24960 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1292
timestamp 1666464484
transform 1 0 24960 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1293
timestamp 1666464484
transform 1 0 24960 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1294
timestamp 1666464484
transform 1 0 24960 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1295
timestamp 1666464484
transform 1 0 24960 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1296
timestamp 1666464484
transform 1 0 21216 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1297
timestamp 1666464484
transform 1 0 21216 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1298
timestamp 1666464484
transform -1 0 26208 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1299
timestamp 1666464484
transform -1 0 26208 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1300
timestamp 1666464484
transform -1 0 22464 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1301
timestamp 1666464484
transform -1 0 22464 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1302
timestamp 1666464484
transform 1 0 27456 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1303
timestamp 1666464484
transform 1 0 27456 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1304
timestamp 1666464484
transform 1 0 22464 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1305
timestamp 1666464484
transform -1 0 23712 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1306
timestamp 1666464484
transform -1 0 23712 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1307
timestamp 1666464484
transform 1 0 22464 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1308
timestamp 1666464484
transform 1 0 28704 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1309
timestamp 1666464484
transform 1 0 28704 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1310
timestamp 1666464484
transform 1 0 23712 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1311
timestamp 1666464484
transform 1 0 23712 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1312
timestamp 1666464484
transform -1 0 24960 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1313
timestamp 1666464484
transform -1 0 24960 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1314
timestamp 1666464484
transform -1 0 24960 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1315
timestamp 1666464484
transform -1 0 24960 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1316
timestamp 1666464484
transform -1 0 24960 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1317
timestamp 1666464484
transform -1 0 24960 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1318
timestamp 1666464484
transform -1 0 24960 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1319
timestamp 1666464484
transform -1 0 38688 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1320
timestamp 1666464484
transform -1 0 38688 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1321
timestamp 1666464484
transform -1 0 38688 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1322
timestamp 1666464484
transform -1 0 38688 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1323
timestamp 1666464484
transform -1 0 38688 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1324
timestamp 1666464484
transform -1 0 38688 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1325
timestamp 1666464484
transform -1 0 38688 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1326
timestamp 1666464484
transform -1 0 38688 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1327
timestamp 1666464484
transform -1 0 38688 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1328
timestamp 1666464484
transform -1 0 38688 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1329
timestamp 1666464484
transform -1 0 38688 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1330
timestamp 1666464484
transform -1 0 38688 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1331
timestamp 1666464484
transform -1 0 38688 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1332
timestamp 1666464484
transform -1 0 38688 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1333
timestamp 1666464484
transform 1 0 37440 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1334
timestamp 1666464484
transform 1 0 38688 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1335
timestamp 1666464484
transform 1 0 38688 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1336
timestamp 1666464484
transform 1 0 38688 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1337
timestamp 1666464484
transform 1 0 38688 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1338
timestamp 1666464484
transform 1 0 38688 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1339
timestamp 1666464484
transform 1 0 38688 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1340
timestamp 1666464484
transform 1 0 38688 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1341
timestamp 1666464484
transform 1 0 38688 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1342
timestamp 1666464484
transform 1 0 38688 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1343
timestamp 1666464484
transform 1 0 38688 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1344
timestamp 1666464484
transform 1 0 38688 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1345
timestamp 1666464484
transform 1 0 38688 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1346
timestamp 1666464484
transform 1 0 38688 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1347
timestamp 1666464484
transform 1 0 38688 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1348
timestamp 1666464484
transform 1 0 37440 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1349
timestamp 1666464484
transform 1 0 37440 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1350
timestamp 1666464484
transform 1 0 37440 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1351
timestamp 1666464484
transform -1 0 36192 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1352
timestamp 1666464484
transform -1 0 36192 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1353
timestamp 1666464484
transform -1 0 36192 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1354
timestamp 1666464484
transform -1 0 36192 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1355
timestamp 1666464484
transform -1 0 36192 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1356
timestamp 1666464484
transform -1 0 36192 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1357
timestamp 1666464484
transform -1 0 36192 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1358
timestamp 1666464484
transform -1 0 36192 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1359
timestamp 1666464484
transform -1 0 36192 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1360
timestamp 1666464484
transform -1 0 36192 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1361
timestamp 1666464484
transform -1 0 36192 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1362
timestamp 1666464484
transform -1 0 36192 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1363
timestamp 1666464484
transform 1 0 36192 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1364
timestamp 1666464484
transform 1 0 36192 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1365
timestamp 1666464484
transform 1 0 36192 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1366
timestamp 1666464484
transform 1 0 36192 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1367
timestamp 1666464484
transform 1 0 36192 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1368
timestamp 1666464484
transform 1 0 36192 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1369
timestamp 1666464484
transform 1 0 36192 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1370
timestamp 1666464484
transform -1 0 39936 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1371
timestamp 1666464484
transform -1 0 39936 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1372
timestamp 1666464484
transform -1 0 39936 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1373
timestamp 1666464484
transform -1 0 39936 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1374
timestamp 1666464484
transform -1 0 39936 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1375
timestamp 1666464484
transform -1 0 39936 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1376
timestamp 1666464484
transform -1 0 39936 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1377
timestamp 1666464484
transform -1 0 39936 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1378
timestamp 1666464484
transform -1 0 39936 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1379
timestamp 1666464484
transform -1 0 39936 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1380
timestamp 1666464484
transform -1 0 39936 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1381
timestamp 1666464484
transform -1 0 39936 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1382
timestamp 1666464484
transform -1 0 39936 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1383
timestamp 1666464484
transform -1 0 39936 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1384
timestamp 1666464484
transform 1 0 36192 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1385
timestamp 1666464484
transform 1 0 36192 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1386
timestamp 1666464484
transform 1 0 36192 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1387
timestamp 1666464484
transform -1 0 37440 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1388
timestamp 1666464484
transform -1 0 37440 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1389
timestamp 1666464484
transform -1 0 37440 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1390
timestamp 1666464484
transform -1 0 37440 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1391
timestamp 1666464484
transform -1 0 37440 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1392
timestamp 1666464484
transform -1 0 37440 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1393
timestamp 1666464484
transform -1 0 37440 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1394
timestamp 1666464484
transform -1 0 37440 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1395
timestamp 1666464484
transform -1 0 37440 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1396
timestamp 1666464484
transform -1 0 37440 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1397
timestamp 1666464484
transform -1 0 37440 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1398
timestamp 1666464484
transform -1 0 37440 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1399
timestamp 1666464484
transform -1 0 37440 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1400
timestamp 1666464484
transform -1 0 37440 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1401
timestamp 1666464484
transform 1 0 36192 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1402
timestamp 1666464484
transform 1 0 36192 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1403
timestamp 1666464484
transform 1 0 36192 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1404
timestamp 1666464484
transform 1 0 36192 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1405
timestamp 1666464484
transform -1 0 36192 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1406
timestamp 1666464484
transform -1 0 36192 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1407
timestamp 1666464484
transform 1 0 37440 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1408
timestamp 1666464484
transform 1 0 37440 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1409
timestamp 1666464484
transform 1 0 37440 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1410
timestamp 1666464484
transform 1 0 37440 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1411
timestamp 1666464484
transform 1 0 37440 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1412
timestamp 1666464484
transform 1 0 37440 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1413
timestamp 1666464484
transform 1 0 37440 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1414
timestamp 1666464484
transform 1 0 37440 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1415
timestamp 1666464484
transform 1 0 37440 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1416
timestamp 1666464484
transform 1 0 37440 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1417
timestamp 1666464484
transform 1 0 33696 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1418
timestamp 1666464484
transform 1 0 33696 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1419
timestamp 1666464484
transform 1 0 33696 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1420
timestamp 1666464484
transform 1 0 33696 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1421
timestamp 1666464484
transform 1 0 33696 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1422
timestamp 1666464484
transform 1 0 33696 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1423
timestamp 1666464484
transform 1 0 33696 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1424
timestamp 1666464484
transform 1 0 33696 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1425
timestamp 1666464484
transform 1 0 33696 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1426
timestamp 1666464484
transform 1 0 33696 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1427
timestamp 1666464484
transform 1 0 33696 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1428
timestamp 1666464484
transform -1 0 31200 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1429
timestamp 1666464484
transform 1 0 33696 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1430
timestamp 1666464484
transform 1 0 33696 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1431
timestamp 1666464484
transform 1 0 31200 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1432
timestamp 1666464484
transform 1 0 31200 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1433
timestamp 1666464484
transform 1 0 31200 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1434
timestamp 1666464484
transform 1 0 31200 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1435
timestamp 1666464484
transform 1 0 31200 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1436
timestamp 1666464484
transform 1 0 31200 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1437
timestamp 1666464484
transform 1 0 31200 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1438
timestamp 1666464484
transform 1 0 31200 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1439
timestamp 1666464484
transform 1 0 31200 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1440
timestamp 1666464484
transform 1 0 31200 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1441
timestamp 1666464484
transform 1 0 31200 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1442
timestamp 1666464484
transform -1 0 32448 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1443
timestamp 1666464484
transform 1 0 32448 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1444
timestamp 1666464484
transform 1 0 32448 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1445
timestamp 1666464484
transform 1 0 32448 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1446
timestamp 1666464484
transform 1 0 32448 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1447
timestamp 1666464484
transform 1 0 32448 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1448
timestamp 1666464484
transform 1 0 32448 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1449
timestamp 1666464484
transform -1 0 33696 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1450
timestamp 1666464484
transform -1 0 33696 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1451
timestamp 1666464484
transform -1 0 33696 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1452
timestamp 1666464484
transform 1 0 32448 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1453
timestamp 1666464484
transform 1 0 32448 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1454
timestamp 1666464484
transform 1 0 32448 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1455
timestamp 1666464484
transform 1 0 32448 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1456
timestamp 1666464484
transform 1 0 32448 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1457
timestamp 1666464484
transform -1 0 31200 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1458
timestamp 1666464484
transform -1 0 31200 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1459
timestamp 1666464484
transform -1 0 31200 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1460
timestamp 1666464484
transform -1 0 31200 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1461
timestamp 1666464484
transform -1 0 31200 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1462
timestamp 1666464484
transform -1 0 31200 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1463
timestamp 1666464484
transform -1 0 32448 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1464
timestamp 1666464484
transform -1 0 32448 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1465
timestamp 1666464484
transform -1 0 32448 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1466
timestamp 1666464484
transform -1 0 32448 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1467
timestamp 1666464484
transform -1 0 32448 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1468
timestamp 1666464484
transform -1 0 33696 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1469
timestamp 1666464484
transform -1 0 33696 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1470
timestamp 1666464484
transform -1 0 33696 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1471
timestamp 1666464484
transform -1 0 33696 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1472
timestamp 1666464484
transform -1 0 33696 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1473
timestamp 1666464484
transform -1 0 33696 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1474
timestamp 1666464484
transform -1 0 33696 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1475
timestamp 1666464484
transform -1 0 33696 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1476
timestamp 1666464484
transform -1 0 33696 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1477
timestamp 1666464484
transform -1 0 33696 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1478
timestamp 1666464484
transform -1 0 33696 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1479
timestamp 1666464484
transform -1 0 32448 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1480
timestamp 1666464484
transform -1 0 32448 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1481
timestamp 1666464484
transform -1 0 31200 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1482
timestamp 1666464484
transform -1 0 31200 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1483
timestamp 1666464484
transform -1 0 31200 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1484
timestamp 1666464484
transform -1 0 31200 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1485
timestamp 1666464484
transform 1 0 31200 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1486
timestamp 1666464484
transform -1 0 31200 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1487
timestamp 1666464484
transform -1 0 31200 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1488
timestamp 1666464484
transform 1 0 31200 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1489
timestamp 1666464484
transform 1 0 31200 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1490
timestamp 1666464484
transform -1 0 32448 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1491
timestamp 1666464484
transform -1 0 32448 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1492
timestamp 1666464484
transform -1 0 32448 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1493
timestamp 1666464484
transform -1 0 32448 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1494
timestamp 1666464484
transform -1 0 32448 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1495
timestamp 1666464484
transform -1 0 32448 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1496
timestamp 1666464484
transform 1 0 33696 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1497
timestamp 1666464484
transform 1 0 32448 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1498
timestamp 1666464484
transform 1 0 32448 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1499
timestamp 1666464484
transform 1 0 32448 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1500
timestamp 1666464484
transform -1 0 31200 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1501
timestamp 1666464484
transform -1 0 31200 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1502
timestamp 1666464484
transform -1 0 31200 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1503
timestamp 1666464484
transform -1 0 31200 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1504
timestamp 1666464484
transform -1 0 31200 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1505
timestamp 1666464484
transform -1 0 31200 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1506
timestamp 1666464484
transform -1 0 33696 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1507
timestamp 1666464484
transform -1 0 33696 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1508
timestamp 1666464484
transform -1 0 33696 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1509
timestamp 1666464484
transform -1 0 33696 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1510
timestamp 1666464484
transform -1 0 33696 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1511
timestamp 1666464484
transform -1 0 33696 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1512
timestamp 1666464484
transform -1 0 33696 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1513
timestamp 1666464484
transform -1 0 33696 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1514
timestamp 1666464484
transform -1 0 33696 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1515
timestamp 1666464484
transform -1 0 33696 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1516
timestamp 1666464484
transform -1 0 33696 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1517
timestamp 1666464484
transform -1 0 33696 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1518
timestamp 1666464484
transform -1 0 33696 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1519
timestamp 1666464484
transform -1 0 33696 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1520
timestamp 1666464484
transform -1 0 32448 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1521
timestamp 1666464484
transform -1 0 31200 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1522
timestamp 1666464484
transform -1 0 31200 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1523
timestamp 1666464484
transform -1 0 31200 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1524
timestamp 1666464484
transform -1 0 31200 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1525
timestamp 1666464484
transform -1 0 31200 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1526
timestamp 1666464484
transform 1 0 33696 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1527
timestamp 1666464484
transform 1 0 33696 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1528
timestamp 1666464484
transform 1 0 33696 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1529
timestamp 1666464484
transform 1 0 33696 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1530
timestamp 1666464484
transform 1 0 33696 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1531
timestamp 1666464484
transform 1 0 33696 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1532
timestamp 1666464484
transform 1 0 33696 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1533
timestamp 1666464484
transform 1 0 33696 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1534
timestamp 1666464484
transform 1 0 33696 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1535
timestamp 1666464484
transform 1 0 33696 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1536
timestamp 1666464484
transform 1 0 33696 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1537
timestamp 1666464484
transform 1 0 33696 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1538
timestamp 1666464484
transform 1 0 33696 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1539
timestamp 1666464484
transform 1 0 31200 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1540
timestamp 1666464484
transform 1 0 32448 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1541
timestamp 1666464484
transform 1 0 32448 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1542
timestamp 1666464484
transform 1 0 32448 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1543
timestamp 1666464484
transform 1 0 32448 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1544
timestamp 1666464484
transform 1 0 32448 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1545
timestamp 1666464484
transform 1 0 32448 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1546
timestamp 1666464484
transform 1 0 32448 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1547
timestamp 1666464484
transform 1 0 32448 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1548
timestamp 1666464484
transform 1 0 32448 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1549
timestamp 1666464484
transform 1 0 32448 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1550
timestamp 1666464484
transform 1 0 32448 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1551
timestamp 1666464484
transform 1 0 32448 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1552
timestamp 1666464484
transform 1 0 32448 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1553
timestamp 1666464484
transform 1 0 32448 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1554
timestamp 1666464484
transform 1 0 31200 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1555
timestamp 1666464484
transform 1 0 31200 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1556
timestamp 1666464484
transform 1 0 31200 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1557
timestamp 1666464484
transform 1 0 31200 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1558
timestamp 1666464484
transform 1 0 31200 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1559
timestamp 1666464484
transform 1 0 31200 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1560
timestamp 1666464484
transform 1 0 31200 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1561
timestamp 1666464484
transform 1 0 31200 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1562
timestamp 1666464484
transform 1 0 31200 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1563
timestamp 1666464484
transform 1 0 31200 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1564
timestamp 1666464484
transform 1 0 31200 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1565
timestamp 1666464484
transform 1 0 31200 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1566
timestamp 1666464484
transform 1 0 31200 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1567
timestamp 1666464484
transform -1 0 31200 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1568
timestamp 1666464484
transform -1 0 31200 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1569
timestamp 1666464484
transform -1 0 31200 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1570
timestamp 1666464484
transform 1 0 33696 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1571
timestamp 1666464484
transform -1 0 31200 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1572
timestamp 1666464484
transform -1 0 32448 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1573
timestamp 1666464484
transform -1 0 32448 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1574
timestamp 1666464484
transform -1 0 32448 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1575
timestamp 1666464484
transform -1 0 32448 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1576
timestamp 1666464484
transform -1 0 32448 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1577
timestamp 1666464484
transform -1 0 32448 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1578
timestamp 1666464484
transform -1 0 32448 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1579
timestamp 1666464484
transform -1 0 32448 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1580
timestamp 1666464484
transform -1 0 32448 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1581
timestamp 1666464484
transform -1 0 32448 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1582
timestamp 1666464484
transform -1 0 32448 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1583
timestamp 1666464484
transform -1 0 32448 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1584
timestamp 1666464484
transform -1 0 32448 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1585
timestamp 1666464484
transform 1 0 36192 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1586
timestamp 1666464484
transform 1 0 36192 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1587
timestamp 1666464484
transform -1 0 39936 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1588
timestamp 1666464484
transform -1 0 39936 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1589
timestamp 1666464484
transform -1 0 39936 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1590
timestamp 1666464484
transform -1 0 39936 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1591
timestamp 1666464484
transform -1 0 39936 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1592
timestamp 1666464484
transform -1 0 39936 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1593
timestamp 1666464484
transform -1 0 39936 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1594
timestamp 1666464484
transform -1 0 39936 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1595
timestamp 1666464484
transform -1 0 39936 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1596
timestamp 1666464484
transform -1 0 39936 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1597
timestamp 1666464484
transform -1 0 39936 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1598
timestamp 1666464484
transform -1 0 39936 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1599
timestamp 1666464484
transform -1 0 39936 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1600
timestamp 1666464484
transform -1 0 39936 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1601
timestamp 1666464484
transform 1 0 36192 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1602
timestamp 1666464484
transform 1 0 36192 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1603
timestamp 1666464484
transform 1 0 36192 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1604
timestamp 1666464484
transform 1 0 36192 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1605
timestamp 1666464484
transform -1 0 36192 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1606
timestamp 1666464484
transform -1 0 36192 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1607
timestamp 1666464484
transform 1 0 38688 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1608
timestamp 1666464484
transform 1 0 38688 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1609
timestamp 1666464484
transform 1 0 38688 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1610
timestamp 1666464484
transform 1 0 38688 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1611
timestamp 1666464484
transform 1 0 38688 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1612
timestamp 1666464484
transform 1 0 38688 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1613
timestamp 1666464484
transform 1 0 38688 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1614
timestamp 1666464484
transform 1 0 38688 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1615
timestamp 1666464484
transform 1 0 38688 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1616
timestamp 1666464484
transform 1 0 38688 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1617
timestamp 1666464484
transform 1 0 38688 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1618
timestamp 1666464484
transform 1 0 38688 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1619
timestamp 1666464484
transform 1 0 38688 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1620
timestamp 1666464484
transform 1 0 38688 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1621
timestamp 1666464484
transform -1 0 36192 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1622
timestamp 1666464484
transform -1 0 36192 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1623
timestamp 1666464484
transform -1 0 36192 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1624
timestamp 1666464484
transform -1 0 36192 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1625
timestamp 1666464484
transform -1 0 38688 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1626
timestamp 1666464484
transform -1 0 38688 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1627
timestamp 1666464484
transform -1 0 38688 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1628
timestamp 1666464484
transform -1 0 38688 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1629
timestamp 1666464484
transform -1 0 38688 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1630
timestamp 1666464484
transform -1 0 38688 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1631
timestamp 1666464484
transform -1 0 38688 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1632
timestamp 1666464484
transform -1 0 38688 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1633
timestamp 1666464484
transform -1 0 38688 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1634
timestamp 1666464484
transform -1 0 38688 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1635
timestamp 1666464484
transform -1 0 38688 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1636
timestamp 1666464484
transform -1 0 38688 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1637
timestamp 1666464484
transform -1 0 38688 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1638
timestamp 1666464484
transform -1 0 38688 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1639
timestamp 1666464484
transform -1 0 36192 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1640
timestamp 1666464484
transform -1 0 36192 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1641
timestamp 1666464484
transform -1 0 36192 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1642
timestamp 1666464484
transform -1 0 36192 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1643
timestamp 1666464484
transform 1 0 37440 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1644
timestamp 1666464484
transform 1 0 37440 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1645
timestamp 1666464484
transform 1 0 37440 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1646
timestamp 1666464484
transform 1 0 37440 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1647
timestamp 1666464484
transform 1 0 37440 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1648
timestamp 1666464484
transform 1 0 37440 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1649
timestamp 1666464484
transform 1 0 37440 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1650
timestamp 1666464484
transform 1 0 37440 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1651
timestamp 1666464484
transform 1 0 37440 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1652
timestamp 1666464484
transform 1 0 37440 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1653
timestamp 1666464484
transform 1 0 37440 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1654
timestamp 1666464484
transform 1 0 37440 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1655
timestamp 1666464484
transform 1 0 37440 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1656
timestamp 1666464484
transform 1 0 37440 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1657
timestamp 1666464484
transform -1 0 36192 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1658
timestamp 1666464484
transform -1 0 36192 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1659
timestamp 1666464484
transform -1 0 37440 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1660
timestamp 1666464484
transform -1 0 37440 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1661
timestamp 1666464484
transform -1 0 37440 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1662
timestamp 1666464484
transform -1 0 37440 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1663
timestamp 1666464484
transform -1 0 37440 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1664
timestamp 1666464484
transform -1 0 37440 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1665
timestamp 1666464484
transform -1 0 37440 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1666
timestamp 1666464484
transform -1 0 37440 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1667
timestamp 1666464484
transform -1 0 37440 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1668
timestamp 1666464484
transform -1 0 37440 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1669
timestamp 1666464484
transform -1 0 37440 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1670
timestamp 1666464484
transform -1 0 37440 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1671
timestamp 1666464484
transform -1 0 37440 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1672
timestamp 1666464484
transform -1 0 37440 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1673
timestamp 1666464484
transform -1 0 36192 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1674
timestamp 1666464484
transform -1 0 36192 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1675
timestamp 1666464484
transform 1 0 36192 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1676
timestamp 1666464484
transform 1 0 36192 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1677
timestamp 1666464484
transform 1 0 36192 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1678
timestamp 1666464484
transform 1 0 36192 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1679
timestamp 1666464484
transform 1 0 36192 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1680
timestamp 1666464484
transform 1 0 36192 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1681
timestamp 1666464484
transform 1 0 36192 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1682
timestamp 1666464484
transform 1 0 36192 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1683
timestamp 1666464484
transform -1 0 33696 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1684
timestamp 1666464484
transform -1 0 33696 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1685
timestamp 1666464484
transform -1 0 39936 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1686
timestamp 1666464484
transform -1 0 39936 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1687
timestamp 1666464484
transform -1 0 31200 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1688
timestamp 1666464484
transform -1 0 31200 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1689
timestamp 1666464484
transform 1 0 32448 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1690
timestamp 1666464484
transform 1 0 32448 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1691
timestamp 1666464484
transform 1 0 38688 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1692
timestamp 1666464484
transform 1 0 38688 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1693
timestamp 1666464484
transform -1 0 32448 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1694
timestamp 1666464484
transform -1 0 32448 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1695
timestamp 1666464484
transform -1 0 38688 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1696
timestamp 1666464484
transform -1 0 38688 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1697
timestamp 1666464484
transform 1 0 31200 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1698
timestamp 1666464484
transform 1 0 31200 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1699
timestamp 1666464484
transform 1 0 37440 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1700
timestamp 1666464484
transform 1 0 37440 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1701
timestamp 1666464484
transform -1 0 37440 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1702
timestamp 1666464484
transform -1 0 37440 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1703
timestamp 1666464484
transform 1 0 36192 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1704
timestamp 1666464484
transform 1 0 36192 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1705
timestamp 1666464484
transform -1 0 36192 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1706
timestamp 1666464484
transform -1 0 36192 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1707
timestamp 1666464484
transform 1 0 34944 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1708
timestamp 1666464484
transform 1 0 34944 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1709
timestamp 1666464484
transform 1 0 34944 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1710
timestamp 1666464484
transform 1 0 34944 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1711
timestamp 1666464484
transform 1 0 34944 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1712
timestamp 1666464484
transform 1 0 34944 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1713
timestamp 1666464484
transform 1 0 34944 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1714
timestamp 1666464484
transform 1 0 34944 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1715
timestamp 1666464484
transform 1 0 34944 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1716
timestamp 1666464484
transform 1 0 34944 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1717
timestamp 1666464484
transform 1 0 34944 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1718
timestamp 1666464484
transform 1 0 34944 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1719
timestamp 1666464484
transform 1 0 34944 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1720
timestamp 1666464484
transform 1 0 34944 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1721
timestamp 1666464484
transform 1 0 34944 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1722
timestamp 1666464484
transform 1 0 34944 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1723
timestamp 1666464484
transform 1 0 34944 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1724
timestamp 1666464484
transform 1 0 34944 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1725
timestamp 1666464484
transform 1 0 34944 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1726
timestamp 1666464484
transform 1 0 34944 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1727
timestamp 1666464484
transform 1 0 34944 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1728
timestamp 1666464484
transform 1 0 34944 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1729
timestamp 1666464484
transform 1 0 34944 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1730
timestamp 1666464484
transform 1 0 34944 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1731
timestamp 1666464484
transform 1 0 34944 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1732
timestamp 1666464484
transform 1 0 34944 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1733
timestamp 1666464484
transform 1 0 34944 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1734
timestamp 1666464484
transform 1 0 34944 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1735
timestamp 1666464484
transform 1 0 34944 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1736
timestamp 1666464484
transform 1 0 34944 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1737
timestamp 1666464484
transform -1 0 34944 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1738
timestamp 1666464484
transform -1 0 34944 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1739
timestamp 1666464484
transform -1 0 34944 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1740
timestamp 1666464484
transform -1 0 34944 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1741
timestamp 1666464484
transform -1 0 34944 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1742
timestamp 1666464484
transform -1 0 34944 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1743
timestamp 1666464484
transform -1 0 34944 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1744
timestamp 1666464484
transform -1 0 34944 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1745
timestamp 1666464484
transform -1 0 34944 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1746
timestamp 1666464484
transform -1 0 34944 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1747
timestamp 1666464484
transform -1 0 34944 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1748
timestamp 1666464484
transform -1 0 34944 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1749
timestamp 1666464484
transform -1 0 34944 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1750
timestamp 1666464484
transform -1 0 34944 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1751
timestamp 1666464484
transform -1 0 34944 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1752
timestamp 1666464484
transform -1 0 34944 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1753
timestamp 1666464484
transform -1 0 34944 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1754
timestamp 1666464484
transform -1 0 34944 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1755
timestamp 1666464484
transform -1 0 34944 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1756
timestamp 1666464484
transform -1 0 34944 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1757
timestamp 1666464484
transform -1 0 34944 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1758
timestamp 1666464484
transform -1 0 34944 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1759
timestamp 1666464484
transform -1 0 34944 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1760
timestamp 1666464484
transform -1 0 34944 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1761
timestamp 1666464484
transform -1 0 34944 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1762
timestamp 1666464484
transform -1 0 34944 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1763
timestamp 1666464484
transform -1 0 34944 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1764
timestamp 1666464484
transform -1 0 34944 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1765
timestamp 1666464484
transform -1 0 34944 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1766
timestamp 1666464484
transform -1 0 34944 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1767
timestamp 1666464484
transform 1 0 33696 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1768
timestamp 1666464484
transform 1 0 33696 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1769
timestamp 1666464484
transform -1 0 21216 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1770
timestamp 1666464484
transform -1 0 21216 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1771
timestamp 1666464484
transform 1 0 29952 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1772
timestamp 1666464484
transform 1 0 29952 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1773
timestamp 1666464484
transform 1 0 29952 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1774
timestamp 1666464484
transform 1 0 29952 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1775
timestamp 1666464484
transform 1 0 29952 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1776
timestamp 1666464484
transform 1 0 29952 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1777
timestamp 1666464484
transform 1 0 29952 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1778
timestamp 1666464484
transform 1 0 29952 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1779
timestamp 1666464484
transform 1 0 29952 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1780
timestamp 1666464484
transform 1 0 29952 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1781
timestamp 1666464484
transform 1 0 29952 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1782
timestamp 1666464484
transform 1 0 29952 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1783
timestamp 1666464484
transform 1 0 29952 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1784
timestamp 1666464484
transform 1 0 29952 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1785
timestamp 1666464484
transform 1 0 29952 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1786
timestamp 1666464484
transform 1 0 29952 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1787
timestamp 1666464484
transform 1 0 29952 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1788
timestamp 1666464484
transform 1 0 29952 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1789
timestamp 1666464484
transform 1 0 29952 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1790
timestamp 1666464484
transform 1 0 29952 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1791
timestamp 1666464484
transform 1 0 29952 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1792
timestamp 1666464484
transform 1 0 29952 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1793
timestamp 1666464484
transform 1 0 29952 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1794
timestamp 1666464484
transform 1 0 29952 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1795
timestamp 1666464484
transform 1 0 29952 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1796
timestamp 1666464484
transform 1 0 29952 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1797
timestamp 1666464484
transform 1 0 29952 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1798
timestamp 1666464484
transform 1 0 29952 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1799
timestamp 1666464484
transform 1 0 29952 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1800
timestamp 1666464484
transform 1 0 29952 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1801
timestamp 1666464484
transform 1 0 29952 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1802
timestamp 1666464484
transform 1 0 29952 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1803
timestamp 1666464484
transform 1 0 29952 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1804
timestamp 1666464484
transform -1 0 39936 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1805
timestamp 1666464484
transform -1 0 39936 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1806
timestamp 1666464484
transform 1 0 29952 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1807
timestamp 1666464484
transform 1 0 29952 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1808
timestamp 1666464484
transform 1 0 29952 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1809
timestamp 1666464484
transform 1 0 29952 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1810
timestamp 1666464484
transform 1 0 29952 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1811
timestamp 1666464484
transform 1 0 29952 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1812
timestamp 1666464484
transform 1 0 29952 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1813
timestamp 1666464484
transform 1 0 29952 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1814
timestamp 1666464484
transform 1 0 29952 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1815
timestamp 1666464484
transform 1 0 29952 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1816
timestamp 1666464484
transform 1 0 29952 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1817
timestamp 1666464484
transform 1 0 29952 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1818
timestamp 1666464484
transform 1 0 29952 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1819
timestamp 1666464484
transform 1 0 29952 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1820
timestamp 1666464484
transform 1 0 29952 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1821
timestamp 1666464484
transform 1 0 29952 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1822
timestamp 1666464484
transform 1 0 29952 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1823
timestamp 1666464484
transform 1 0 29952 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1824
timestamp 1666464484
transform 1 0 29952 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1825
timestamp 1666464484
transform 1 0 29952 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1826
timestamp 1666464484
transform 1 0 29952 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1827
timestamp 1666464484
transform 1 0 29952 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1828
timestamp 1666464484
transform 1 0 29952 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1829
timestamp 1666464484
transform 1 0 29952 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1830
timestamp 1666464484
transform 1 0 29952 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1831
timestamp 1666464484
transform 1 0 29952 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1832
timestamp 1666464484
transform 1 0 29952 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1833
timestamp 1666464484
transform 1 0 29952 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1834
timestamp 1666464484
transform 1 0 29952 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1835
timestamp 1666464484
transform 1 0 29952 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1836
timestamp 1666464484
transform 1 0 38688 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1837
timestamp 1666464484
transform 1 0 38688 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1838
timestamp 1666464484
transform 1 0 24960 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1839
timestamp 1666464484
transform 1 0 24960 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1840
timestamp 1666464484
transform -1 0 29952 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1841
timestamp 1666464484
transform -1 0 29952 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1842
timestamp 1666464484
transform -1 0 29952 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1843
timestamp 1666464484
transform -1 0 29952 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1844
timestamp 1666464484
transform -1 0 29952 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1845
timestamp 1666464484
transform -1 0 29952 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1846
timestamp 1666464484
transform -1 0 29952 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1847
timestamp 1666464484
transform -1 0 29952 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1848
timestamp 1666464484
transform -1 0 29952 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1849
timestamp 1666464484
transform -1 0 29952 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1850
timestamp 1666464484
transform -1 0 29952 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1851
timestamp 1666464484
transform -1 0 29952 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1852
timestamp 1666464484
transform -1 0 29952 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1853
timestamp 1666464484
transform -1 0 29952 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1854
timestamp 1666464484
transform -1 0 29952 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1855
timestamp 1666464484
transform -1 0 29952 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1856
timestamp 1666464484
transform -1 0 29952 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1857
timestamp 1666464484
transform -1 0 29952 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1858
timestamp 1666464484
transform -1 0 29952 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1859
timestamp 1666464484
transform -1 0 29952 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1860
timestamp 1666464484
transform -1 0 29952 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1861
timestamp 1666464484
transform -1 0 29952 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1862
timestamp 1666464484
transform -1 0 29952 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1863
timestamp 1666464484
transform -1 0 29952 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1864
timestamp 1666464484
transform -1 0 29952 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1865
timestamp 1666464484
transform -1 0 29952 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1866
timestamp 1666464484
transform -1 0 29952 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1867
timestamp 1666464484
transform -1 0 29952 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1868
timestamp 1666464484
transform -1 0 29952 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1869
timestamp 1666464484
transform -1 0 29952 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1870
timestamp 1666464484
transform -1 0 29952 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1871
timestamp 1666464484
transform -1 0 29952 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1872
timestamp 1666464484
transform -1 0 29952 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1873
timestamp 1666464484
transform -1 0 29952 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1874
timestamp 1666464484
transform -1 0 29952 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1875
timestamp 1666464484
transform -1 0 38688 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1876
timestamp 1666464484
transform -1 0 38688 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1877
timestamp 1666464484
transform -1 0 29952 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1878
timestamp 1666464484
transform -1 0 29952 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1879
timestamp 1666464484
transform -1 0 29952 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1880
timestamp 1666464484
transform -1 0 29952 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1881
timestamp 1666464484
transform -1 0 29952 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1882
timestamp 1666464484
transform -1 0 29952 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1883
timestamp 1666464484
transform -1 0 29952 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1884
timestamp 1666464484
transform -1 0 29952 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1885
timestamp 1666464484
transform -1 0 29952 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1886
timestamp 1666464484
transform -1 0 29952 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1887
timestamp 1666464484
transform -1 0 29952 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1888
timestamp 1666464484
transform -1 0 29952 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1889
timestamp 1666464484
transform -1 0 29952 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1890
timestamp 1666464484
transform -1 0 29952 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1891
timestamp 1666464484
transform -1 0 29952 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1892
timestamp 1666464484
transform -1 0 29952 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1893
timestamp 1666464484
transform -1 0 29952 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1894
timestamp 1666464484
transform -1 0 29952 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1895
timestamp 1666464484
transform -1 0 29952 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1896
timestamp 1666464484
transform -1 0 29952 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1897
timestamp 1666464484
transform -1 0 29952 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1898
timestamp 1666464484
transform -1 0 29952 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1899
timestamp 1666464484
transform -1 0 29952 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1900
timestamp 1666464484
transform -1 0 29952 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1901
timestamp 1666464484
transform -1 0 29952 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1902
timestamp 1666464484
transform -1 0 29952 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1903
timestamp 1666464484
transform -1 0 29952 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1904
timestamp 1666464484
transform -1 0 29952 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1905
timestamp 1666464484
transform 1 0 37440 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1906
timestamp 1666464484
transform 1 0 37440 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1907
timestamp 1666464484
transform 1 0 22464 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1908
timestamp 1666464484
transform 1 0 22464 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1909
timestamp 1666464484
transform 1 0 28704 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1910
timestamp 1666464484
transform 1 0 28704 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1911
timestamp 1666464484
transform -1 0 37440 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1912
timestamp 1666464484
transform -1 0 37440 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1913
timestamp 1666464484
transform 1 0 36192 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1914
timestamp 1666464484
transform 1 0 36192 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1915
timestamp 1666464484
transform -1 0 24960 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1916
timestamp 1666464484
transform -1 0 24960 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1917
timestamp 1666464484
transform -1 0 28704 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1918
timestamp 1666464484
transform -1 0 28704 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1919
timestamp 1666464484
transform -1 0 36192 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1920
timestamp 1666464484
transform -1 0 36192 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1921
timestamp 1666464484
transform 1 0 34944 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1922
timestamp 1666464484
transform 1 0 34944 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1923
timestamp 1666464484
transform 1 0 21216 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1924
timestamp 1666464484
transform 1 0 21216 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1925
timestamp 1666464484
transform 1 0 27456 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1926
timestamp 1666464484
transform 1 0 27456 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1927
timestamp 1666464484
transform -1 0 34944 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1928
timestamp 1666464484
transform -1 0 34944 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1929
timestamp 1666464484
transform 1 0 23712 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1930
timestamp 1666464484
transform 1 0 33696 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1931
timestamp 1666464484
transform 1 0 33696 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1932
timestamp 1666464484
transform 1 0 23712 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1933
timestamp 1666464484
transform -1 0 27456 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1934
timestamp 1666464484
transform -1 0 27456 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1935
timestamp 1666464484
transform -1 0 33696 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1936
timestamp 1666464484
transform -1 0 33696 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1937
timestamp 1666464484
transform 1 0 32448 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1938
timestamp 1666464484
transform 1 0 32448 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1939
timestamp 1666464484
transform -1 0 22464 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1940
timestamp 1666464484
transform -1 0 22464 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1941
timestamp 1666464484
transform 1 0 26208 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1942
timestamp 1666464484
transform 1 0 26208 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1943
timestamp 1666464484
transform -1 0 32448 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1944
timestamp 1666464484
transform -1 0 32448 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1945
timestamp 1666464484
transform -1 0 23712 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1946
timestamp 1666464484
transform -1 0 23712 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1947
timestamp 1666464484
transform 1 0 31200 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1948
timestamp 1666464484
transform 1 0 31200 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1949
timestamp 1666464484
transform -1 0 26208 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1950
timestamp 1666464484
transform -1 0 26208 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1951
timestamp 1666464484
transform -1 0 31200 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1952
timestamp 1666464484
transform -1 0 31200 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1953
timestamp 1666464484
transform -1 0 18720 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1954
timestamp 1666464484
transform -1 0 18720 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1955
timestamp 1666464484
transform -1 0 18720 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1956
timestamp 1666464484
transform -1 0 18720 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1957
timestamp 1666464484
transform -1 0 18720 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1958
timestamp 1666464484
transform -1 0 18720 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1959
timestamp 1666464484
transform -1 0 18720 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1960
timestamp 1666464484
transform -1 0 18720 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1961
timestamp 1666464484
transform -1 0 18720 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1962
timestamp 1666464484
transform -1 0 18720 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1963
timestamp 1666464484
transform -1 0 18720 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1964
timestamp 1666464484
transform -1 0 18720 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1965
timestamp 1666464484
transform -1 0 18720 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1966
timestamp 1666464484
transform -1 0 18720 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1967
timestamp 1666464484
transform 1 0 16224 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1968
timestamp 1666464484
transform 1 0 16224 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1969
timestamp 1666464484
transform 1 0 16224 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1970
timestamp 1666464484
transform 1 0 16224 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1971
timestamp 1666464484
transform 1 0 16224 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1972
timestamp 1666464484
transform 1 0 16224 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1973
timestamp 1666464484
transform 1 0 17472 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1974
timestamp 1666464484
transform 1 0 17472 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1975
timestamp 1666464484
transform 1 0 18720 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1976
timestamp 1666464484
transform 1 0 18720 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1977
timestamp 1666464484
transform 1 0 18720 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1978
timestamp 1666464484
transform 1 0 17472 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1979
timestamp 1666464484
transform 1 0 17472 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1980
timestamp 1666464484
transform 1 0 17472 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1981
timestamp 1666464484
transform 1 0 17472 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1982
timestamp 1666464484
transform 1 0 18720 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1983
timestamp 1666464484
transform 1 0 18720 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1984
timestamp 1666464484
transform 1 0 18720 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1985
timestamp 1666464484
transform 1 0 18720 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1986
timestamp 1666464484
transform 1 0 18720 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1987
timestamp 1666464484
transform 1 0 18720 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1988
timestamp 1666464484
transform 1 0 18720 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1989
timestamp 1666464484
transform 1 0 18720 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1990
timestamp 1666464484
transform 1 0 18720 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1991
timestamp 1666464484
transform 1 0 18720 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1992
timestamp 1666464484
transform 1 0 18720 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1993
timestamp 1666464484
transform 1 0 18720 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1994
timestamp 1666464484
transform 1 0 17472 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1995
timestamp 1666464484
transform -1 0 16224 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1996
timestamp 1666464484
transform -1 0 16224 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1997
timestamp 1666464484
transform -1 0 16224 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1998
timestamp 1666464484
transform -1 0 16224 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_1999
timestamp 1666464484
transform -1 0 16224 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2000
timestamp 1666464484
transform -1 0 16224 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2001
timestamp 1666464484
transform -1 0 16224 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2002
timestamp 1666464484
transform -1 0 16224 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2003
timestamp 1666464484
transform -1 0 16224 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2004
timestamp 1666464484
transform 1 0 17472 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2005
timestamp 1666464484
transform 1 0 17472 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2006
timestamp 1666464484
transform 1 0 17472 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2007
timestamp 1666464484
transform 1 0 17472 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2008
timestamp 1666464484
transform 1 0 17472 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2009
timestamp 1666464484
transform 1 0 17472 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2010
timestamp 1666464484
transform 1 0 17472 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2011
timestamp 1666464484
transform 1 0 17472 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2012
timestamp 1666464484
transform 1 0 16224 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2013
timestamp 1666464484
transform 1 0 16224 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2014
timestamp 1666464484
transform 1 0 16224 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2015
timestamp 1666464484
transform 1 0 16224 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2016
timestamp 1666464484
transform 1 0 16224 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2017
timestamp 1666464484
transform 1 0 16224 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2018
timestamp 1666464484
transform 1 0 16224 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2019
timestamp 1666464484
transform 1 0 16224 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2020
timestamp 1666464484
transform -1 0 17472 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2021
timestamp 1666464484
transform -1 0 17472 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2022
timestamp 1666464484
transform -1 0 17472 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2023
timestamp 1666464484
transform -1 0 17472 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2024
timestamp 1666464484
transform -1 0 17472 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2025
timestamp 1666464484
transform -1 0 17472 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2026
timestamp 1666464484
transform -1 0 17472 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2027
timestamp 1666464484
transform -1 0 17472 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2028
timestamp 1666464484
transform -1 0 17472 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2029
timestamp 1666464484
transform -1 0 17472 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2030
timestamp 1666464484
transform -1 0 17472 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2031
timestamp 1666464484
transform -1 0 17472 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2032
timestamp 1666464484
transform -1 0 17472 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2033
timestamp 1666464484
transform -1 0 17472 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2034
timestamp 1666464484
transform -1 0 17472 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2035
timestamp 1666464484
transform -1 0 16224 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2036
timestamp 1666464484
transform -1 0 16224 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2037
timestamp 1666464484
transform -1 0 16224 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2038
timestamp 1666464484
transform -1 0 16224 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2039
timestamp 1666464484
transform -1 0 16224 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2040
timestamp 1666464484
transform -1 0 16224 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2041
timestamp 1666464484
transform 1 0 16224 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2042
timestamp 1666464484
transform -1 0 18720 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2043
timestamp 1666464484
transform -1 0 13728 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2044
timestamp 1666464484
transform 1 0 12480 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2045
timestamp 1666464484
transform 1 0 12480 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2046
timestamp 1666464484
transform 1 0 12480 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2047
timestamp 1666464484
transform 1 0 12480 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2048
timestamp 1666464484
transform 1 0 12480 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2049
timestamp 1666464484
transform -1 0 12480 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2050
timestamp 1666464484
transform -1 0 12480 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2051
timestamp 1666464484
transform -1 0 12480 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2052
timestamp 1666464484
transform -1 0 12480 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2053
timestamp 1666464484
transform -1 0 11232 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2054
timestamp 1666464484
transform -1 0 11232 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2055
timestamp 1666464484
transform -1 0 11232 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2056
timestamp 1666464484
transform -1 0 11232 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2057
timestamp 1666464484
transform 1 0 11232 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2058
timestamp 1666464484
transform 1 0 11232 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2059
timestamp 1666464484
transform 1 0 11232 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2060
timestamp 1666464484
transform 1 0 11232 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2061
timestamp 1666464484
transform 1 0 11232 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2062
timestamp 1666464484
transform 1 0 11232 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2063
timestamp 1666464484
transform 1 0 11232 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2064
timestamp 1666464484
transform 1 0 11232 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2065
timestamp 1666464484
transform 1 0 11232 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2066
timestamp 1666464484
transform 1 0 11232 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2067
timestamp 1666464484
transform 1 0 11232 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2068
timestamp 1666464484
transform 1 0 11232 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2069
timestamp 1666464484
transform 1 0 11232 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2070
timestamp 1666464484
transform 1 0 11232 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2071
timestamp 1666464484
transform 1 0 11232 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2072
timestamp 1666464484
transform -1 0 11232 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2073
timestamp 1666464484
transform -1 0 11232 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2074
timestamp 1666464484
transform -1 0 11232 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2075
timestamp 1666464484
transform -1 0 11232 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2076
timestamp 1666464484
transform -1 0 11232 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2077
timestamp 1666464484
transform -1 0 11232 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2078
timestamp 1666464484
transform -1 0 11232 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2079
timestamp 1666464484
transform -1 0 11232 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2080
timestamp 1666464484
transform -1 0 11232 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2081
timestamp 1666464484
transform -1 0 11232 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2082
timestamp 1666464484
transform -1 0 11232 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2083
timestamp 1666464484
transform -1 0 12480 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2084
timestamp 1666464484
transform -1 0 12480 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2085
timestamp 1666464484
transform -1 0 13728 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2086
timestamp 1666464484
transform -1 0 13728 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2087
timestamp 1666464484
transform -1 0 13728 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2088
timestamp 1666464484
transform -1 0 13728 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2089
timestamp 1666464484
transform 1 0 12480 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2090
timestamp 1666464484
transform 1 0 12480 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2091
timestamp 1666464484
transform 1 0 12480 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2092
timestamp 1666464484
transform 1 0 12480 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2093
timestamp 1666464484
transform 1 0 12480 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2094
timestamp 1666464484
transform 1 0 12480 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2095
timestamp 1666464484
transform 1 0 12480 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2096
timestamp 1666464484
transform 1 0 12480 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2097
timestamp 1666464484
transform -1 0 13728 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2098
timestamp 1666464484
transform 1 0 13728 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2099
timestamp 1666464484
transform 1 0 13728 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2100
timestamp 1666464484
transform 1 0 12480 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2101
timestamp 1666464484
transform 1 0 12480 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2102
timestamp 1666464484
transform -1 0 13728 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2103
timestamp 1666464484
transform -1 0 13728 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2104
timestamp 1666464484
transform -1 0 13728 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2105
timestamp 1666464484
transform -1 0 13728 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2106
timestamp 1666464484
transform -1 0 13728 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2107
timestamp 1666464484
transform -1 0 13728 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2108
timestamp 1666464484
transform -1 0 13728 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2109
timestamp 1666464484
transform -1 0 12480 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2110
timestamp 1666464484
transform -1 0 12480 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2111
timestamp 1666464484
transform -1 0 12480 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2112
timestamp 1666464484
transform -1 0 12480 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2113
timestamp 1666464484
transform 1 0 13728 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2114
timestamp 1666464484
transform 1 0 13728 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2115
timestamp 1666464484
transform 1 0 13728 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2116
timestamp 1666464484
transform 1 0 13728 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2117
timestamp 1666464484
transform 1 0 13728 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2118
timestamp 1666464484
transform 1 0 13728 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2119
timestamp 1666464484
transform 1 0 13728 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2120
timestamp 1666464484
transform 1 0 13728 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2121
timestamp 1666464484
transform 1 0 13728 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2122
timestamp 1666464484
transform 1 0 13728 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2123
timestamp 1666464484
transform 1 0 13728 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2124
timestamp 1666464484
transform 1 0 13728 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2125
timestamp 1666464484
transform 1 0 13728 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2126
timestamp 1666464484
transform -1 0 12480 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2127
timestamp 1666464484
transform -1 0 12480 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2128
timestamp 1666464484
transform -1 0 12480 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2129
timestamp 1666464484
transform -1 0 12480 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2130
timestamp 1666464484
transform -1 0 12480 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2131
timestamp 1666464484
transform -1 0 13728 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2132
timestamp 1666464484
transform -1 0 13728 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2133
timestamp 1666464484
transform 1 0 11232 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2134
timestamp 1666464484
transform 1 0 11232 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2135
timestamp 1666464484
transform 1 0 11232 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2136
timestamp 1666464484
transform 1 0 11232 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2137
timestamp 1666464484
transform 1 0 11232 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2138
timestamp 1666464484
transform 1 0 11232 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2139
timestamp 1666464484
transform 1 0 11232 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2140
timestamp 1666464484
transform 1 0 11232 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2141
timestamp 1666464484
transform 1 0 11232 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2142
timestamp 1666464484
transform 1 0 11232 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2143
timestamp 1666464484
transform 1 0 11232 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2144
timestamp 1666464484
transform 1 0 11232 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2145
timestamp 1666464484
transform 1 0 12480 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2146
timestamp 1666464484
transform -1 0 12480 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2147
timestamp 1666464484
transform -1 0 12480 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2148
timestamp 1666464484
transform -1 0 12480 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2149
timestamp 1666464484
transform -1 0 12480 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2150
timestamp 1666464484
transform -1 0 12480 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2151
timestamp 1666464484
transform -1 0 12480 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2152
timestamp 1666464484
transform -1 0 12480 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2153
timestamp 1666464484
transform -1 0 12480 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2154
timestamp 1666464484
transform -1 0 12480 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2155
timestamp 1666464484
transform -1 0 12480 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2156
timestamp 1666464484
transform -1 0 12480 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2157
timestamp 1666464484
transform -1 0 12480 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2158
timestamp 1666464484
transform 1 0 12480 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2159
timestamp 1666464484
transform 1 0 12480 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2160
timestamp 1666464484
transform 1 0 11232 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2161
timestamp 1666464484
transform 1 0 11232 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2162
timestamp 1666464484
transform -1 0 12480 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2163
timestamp 1666464484
transform -1 0 12480 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2164
timestamp 1666464484
transform 1 0 13728 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2165
timestamp 1666464484
transform 1 0 13728 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2166
timestamp 1666464484
transform 1 0 13728 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2167
timestamp 1666464484
transform 1 0 13728 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2168
timestamp 1666464484
transform 1 0 13728 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2169
timestamp 1666464484
transform 1 0 13728 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2170
timestamp 1666464484
transform 1 0 13728 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2171
timestamp 1666464484
transform 1 0 13728 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2172
timestamp 1666464484
transform 1 0 13728 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2173
timestamp 1666464484
transform 1 0 13728 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2174
timestamp 1666464484
transform 1 0 13728 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2175
timestamp 1666464484
transform 1 0 13728 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2176
timestamp 1666464484
transform 1 0 13728 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2177
timestamp 1666464484
transform 1 0 13728 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2178
timestamp 1666464484
transform 1 0 12480 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2179
timestamp 1666464484
transform 1 0 12480 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2180
timestamp 1666464484
transform 1 0 12480 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2181
timestamp 1666464484
transform -1 0 11232 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2182
timestamp 1666464484
transform -1 0 11232 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2183
timestamp 1666464484
transform -1 0 11232 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2184
timestamp 1666464484
transform -1 0 11232 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2185
timestamp 1666464484
transform -1 0 11232 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2186
timestamp 1666464484
transform -1 0 11232 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2187
timestamp 1666464484
transform -1 0 11232 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2188
timestamp 1666464484
transform -1 0 11232 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2189
timestamp 1666464484
transform -1 0 11232 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2190
timestamp 1666464484
transform -1 0 11232 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2191
timestamp 1666464484
transform -1 0 11232 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2192
timestamp 1666464484
transform -1 0 11232 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2193
timestamp 1666464484
transform -1 0 11232 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2194
timestamp 1666464484
transform -1 0 11232 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2195
timestamp 1666464484
transform 1 0 12480 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2196
timestamp 1666464484
transform 1 0 12480 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2197
timestamp 1666464484
transform 1 0 12480 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2198
timestamp 1666464484
transform 1 0 12480 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2199
timestamp 1666464484
transform -1 0 13728 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2200
timestamp 1666464484
transform -1 0 13728 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2201
timestamp 1666464484
transform -1 0 13728 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2202
timestamp 1666464484
transform -1 0 13728 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2203
timestamp 1666464484
transform -1 0 13728 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2204
timestamp 1666464484
transform -1 0 13728 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2205
timestamp 1666464484
transform -1 0 13728 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2206
timestamp 1666464484
transform -1 0 13728 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2207
timestamp 1666464484
transform -1 0 13728 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2208
timestamp 1666464484
transform -1 0 13728 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2209
timestamp 1666464484
transform -1 0 13728 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2210
timestamp 1666464484
transform -1 0 13728 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2211
timestamp 1666464484
transform -1 0 13728 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2212
timestamp 1666464484
transform -1 0 13728 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2213
timestamp 1666464484
transform 1 0 12480 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2214
timestamp 1666464484
transform 1 0 12480 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2215
timestamp 1666464484
transform 1 0 12480 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2216
timestamp 1666464484
transform 1 0 12480 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2217
timestamp 1666464484
transform 1 0 16224 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2218
timestamp 1666464484
transform 1 0 16224 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2219
timestamp 1666464484
transform 1 0 18720 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2220
timestamp 1666464484
transform -1 0 17472 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2221
timestamp 1666464484
transform -1 0 17472 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2222
timestamp 1666464484
transform -1 0 17472 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2223
timestamp 1666464484
transform -1 0 17472 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2224
timestamp 1666464484
transform -1 0 17472 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2225
timestamp 1666464484
transform -1 0 17472 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2226
timestamp 1666464484
transform -1 0 17472 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2227
timestamp 1666464484
transform -1 0 17472 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2228
timestamp 1666464484
transform -1 0 17472 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2229
timestamp 1666464484
transform -1 0 17472 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2230
timestamp 1666464484
transform -1 0 17472 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2231
timestamp 1666464484
transform -1 0 17472 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2232
timestamp 1666464484
transform -1 0 17472 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2233
timestamp 1666464484
transform -1 0 17472 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2234
timestamp 1666464484
transform 1 0 18720 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2235
timestamp 1666464484
transform 1 0 18720 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2236
timestamp 1666464484
transform 1 0 18720 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2237
timestamp 1666464484
transform 1 0 18720 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2238
timestamp 1666464484
transform 1 0 18720 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2239
timestamp 1666464484
transform 1 0 18720 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2240
timestamp 1666464484
transform 1 0 18720 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2241
timestamp 1666464484
transform 1 0 18720 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2242
timestamp 1666464484
transform 1 0 18720 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2243
timestamp 1666464484
transform 1 0 18720 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2244
timestamp 1666464484
transform -1 0 16224 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2245
timestamp 1666464484
transform -1 0 16224 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2246
timestamp 1666464484
transform -1 0 16224 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2247
timestamp 1666464484
transform -1 0 16224 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2248
timestamp 1666464484
transform -1 0 16224 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2249
timestamp 1666464484
transform -1 0 16224 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2250
timestamp 1666464484
transform -1 0 16224 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2251
timestamp 1666464484
transform -1 0 16224 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2252
timestamp 1666464484
transform -1 0 16224 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2253
timestamp 1666464484
transform -1 0 18720 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2254
timestamp 1666464484
transform -1 0 18720 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2255
timestamp 1666464484
transform -1 0 18720 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2256
timestamp 1666464484
transform -1 0 18720 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2257
timestamp 1666464484
transform -1 0 18720 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2258
timestamp 1666464484
transform -1 0 18720 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2259
timestamp 1666464484
transform -1 0 18720 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2260
timestamp 1666464484
transform -1 0 18720 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2261
timestamp 1666464484
transform -1 0 18720 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2262
timestamp 1666464484
transform -1 0 18720 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2263
timestamp 1666464484
transform -1 0 18720 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2264
timestamp 1666464484
transform -1 0 18720 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2265
timestamp 1666464484
transform -1 0 18720 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2266
timestamp 1666464484
transform -1 0 18720 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2267
timestamp 1666464484
transform -1 0 16224 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2268
timestamp 1666464484
transform 1 0 17472 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2269
timestamp 1666464484
transform 1 0 17472 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2270
timestamp 1666464484
transform 1 0 17472 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2271
timestamp 1666464484
transform 1 0 17472 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2272
timestamp 1666464484
transform 1 0 17472 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2273
timestamp 1666464484
transform 1 0 17472 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2274
timestamp 1666464484
transform 1 0 17472 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2275
timestamp 1666464484
transform 1 0 17472 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2276
timestamp 1666464484
transform 1 0 17472 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2277
timestamp 1666464484
transform 1 0 17472 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2278
timestamp 1666464484
transform 1 0 17472 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2279
timestamp 1666464484
transform 1 0 17472 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2280
timestamp 1666464484
transform 1 0 17472 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2281
timestamp 1666464484
transform 1 0 17472 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2282
timestamp 1666464484
transform -1 0 16224 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2283
timestamp 1666464484
transform -1 0 16224 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2284
timestamp 1666464484
transform -1 0 16224 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2285
timestamp 1666464484
transform -1 0 16224 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2286
timestamp 1666464484
transform 1 0 18720 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2287
timestamp 1666464484
transform 1 0 18720 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2288
timestamp 1666464484
transform 1 0 18720 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2289
timestamp 1666464484
transform 1 0 16224 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2290
timestamp 1666464484
transform 1 0 16224 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2291
timestamp 1666464484
transform 1 0 16224 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2292
timestamp 1666464484
transform 1 0 16224 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2293
timestamp 1666464484
transform 1 0 16224 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2294
timestamp 1666464484
transform 1 0 16224 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2295
timestamp 1666464484
transform 1 0 16224 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2296
timestamp 1666464484
transform 1 0 16224 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2297
timestamp 1666464484
transform 1 0 16224 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2298
timestamp 1666464484
transform 1 0 16224 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2299
timestamp 1666464484
transform 1 0 16224 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2300
timestamp 1666464484
transform 1 0 16224 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2301
timestamp 1666464484
transform 1 0 11232 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2302
timestamp 1666464484
transform 1 0 11232 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2303
timestamp 1666464484
transform -1 0 16224 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2304
timestamp 1666464484
transform -1 0 17472 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2305
timestamp 1666464484
transform -1 0 17472 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2306
timestamp 1666464484
transform 1 0 13728 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2307
timestamp 1666464484
transform 1 0 13728 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2308
timestamp 1666464484
transform -1 0 14976 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2309
timestamp 1666464484
transform -1 0 11232 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2310
timestamp 1666464484
transform -1 0 11232 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2311
timestamp 1666464484
transform -1 0 14976 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2312
timestamp 1666464484
transform -1 0 14976 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2313
timestamp 1666464484
transform -1 0 14976 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2314
timestamp 1666464484
transform -1 0 14976 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2315
timestamp 1666464484
transform -1 0 14976 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2316
timestamp 1666464484
transform -1 0 14976 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2317
timestamp 1666464484
transform -1 0 14976 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2318
timestamp 1666464484
transform -1 0 14976 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2319
timestamp 1666464484
transform -1 0 14976 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2320
timestamp 1666464484
transform -1 0 14976 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2321
timestamp 1666464484
transform -1 0 14976 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2322
timestamp 1666464484
transform -1 0 14976 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2323
timestamp 1666464484
transform -1 0 18720 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2324
timestamp 1666464484
transform -1 0 18720 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2325
timestamp 1666464484
transform -1 0 14976 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2326
timestamp 1666464484
transform -1 0 14976 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2327
timestamp 1666464484
transform -1 0 14976 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2328
timestamp 1666464484
transform -1 0 14976 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2329
timestamp 1666464484
transform -1 0 14976 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2330
timestamp 1666464484
transform -1 0 14976 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2331
timestamp 1666464484
transform -1 0 14976 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2332
timestamp 1666464484
transform -1 0 14976 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2333
timestamp 1666464484
transform -1 0 14976 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2334
timestamp 1666464484
transform -1 0 14976 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2335
timestamp 1666464484
transform -1 0 14976 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2336
timestamp 1666464484
transform -1 0 14976 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2337
timestamp 1666464484
transform -1 0 14976 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2338
timestamp 1666464484
transform -1 0 14976 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2339
timestamp 1666464484
transform -1 0 14976 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2340
timestamp 1666464484
transform -1 0 14976 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2341
timestamp 1666464484
transform -1 0 14976 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2342
timestamp 1666464484
transform -1 0 14976 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2343
timestamp 1666464484
transform -1 0 13728 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2344
timestamp 1666464484
transform -1 0 13728 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2345
timestamp 1666464484
transform 1 0 16224 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2346
timestamp 1666464484
transform 1 0 16224 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2347
timestamp 1666464484
transform 1 0 14976 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2348
timestamp 1666464484
transform 1 0 14976 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2349
timestamp 1666464484
transform 1 0 14976 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2350
timestamp 1666464484
transform 1 0 14976 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2351
timestamp 1666464484
transform 1 0 14976 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2352
timestamp 1666464484
transform 1 0 14976 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2353
timestamp 1666464484
transform 1 0 14976 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2354
timestamp 1666464484
transform 1 0 14976 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2355
timestamp 1666464484
transform 1 0 14976 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2356
timestamp 1666464484
transform 1 0 14976 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2357
timestamp 1666464484
transform 1 0 14976 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2358
timestamp 1666464484
transform 1 0 14976 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2359
timestamp 1666464484
transform 1 0 14976 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2360
timestamp 1666464484
transform 1 0 14976 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2361
timestamp 1666464484
transform 1 0 14976 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2362
timestamp 1666464484
transform 1 0 14976 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2363
timestamp 1666464484
transform 1 0 14976 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2364
timestamp 1666464484
transform 1 0 14976 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2365
timestamp 1666464484
transform 1 0 14976 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2366
timestamp 1666464484
transform 1 0 17472 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2367
timestamp 1666464484
transform 1 0 17472 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2368
timestamp 1666464484
transform 1 0 14976 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2369
timestamp 1666464484
transform 1 0 14976 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2370
timestamp 1666464484
transform 1 0 14976 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2371
timestamp 1666464484
transform 1 0 14976 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2372
timestamp 1666464484
transform 1 0 14976 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2373
timestamp 1666464484
transform 1 0 14976 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2374
timestamp 1666464484
transform 1 0 14976 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2375
timestamp 1666464484
transform 1 0 14976 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2376
timestamp 1666464484
transform 1 0 14976 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2377
timestamp 1666464484
transform 1 0 14976 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2378
timestamp 1666464484
transform 1 0 14976 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2379
timestamp 1666464484
transform 1 0 14976 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2380
timestamp 1666464484
transform -1 0 12480 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2381
timestamp 1666464484
transform -1 0 12480 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2382
timestamp 1666464484
transform 1 0 12480 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2383
timestamp 1666464484
transform 1 0 12480 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2384
timestamp 1666464484
transform -1 0 16224 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2385
timestamp 1666464484
transform 1 0 18720 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2386
timestamp 1666464484
transform 1 0 18720 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2387
timestamp 1666464484
transform 1 0 8736 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2388
timestamp 1666464484
transform 1 0 8736 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2389
timestamp 1666464484
transform 1 0 8736 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2390
timestamp 1666464484
transform -1 0 6240 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2391
timestamp 1666464484
transform -1 0 6240 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2392
timestamp 1666464484
transform -1 0 6240 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2393
timestamp 1666464484
transform -1 0 6240 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2394
timestamp 1666464484
transform -1 0 6240 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2395
timestamp 1666464484
transform -1 0 6240 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2396
timestamp 1666464484
transform -1 0 6240 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2397
timestamp 1666464484
transform -1 0 6240 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2398
timestamp 1666464484
transform -1 0 6240 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2399
timestamp 1666464484
transform -1 0 6240 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2400
timestamp 1666464484
transform -1 0 6240 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2401
timestamp 1666464484
transform -1 0 6240 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2402
timestamp 1666464484
transform -1 0 6240 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2403
timestamp 1666464484
transform -1 0 6240 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2404
timestamp 1666464484
transform -1 0 6240 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2405
timestamp 1666464484
transform 1 0 8736 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2406
timestamp 1666464484
transform 1 0 8736 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2407
timestamp 1666464484
transform 1 0 8736 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2408
timestamp 1666464484
transform 1 0 8736 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2409
timestamp 1666464484
transform 1 0 8736 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2410
timestamp 1666464484
transform 1 0 8736 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2411
timestamp 1666464484
transform 1 0 8736 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2412
timestamp 1666464484
transform 1 0 8736 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2413
timestamp 1666464484
transform 1 0 8736 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2414
timestamp 1666464484
transform 1 0 8736 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2415
timestamp 1666464484
transform 1 0 6240 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2416
timestamp 1666464484
transform -1 0 8736 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2417
timestamp 1666464484
transform -1 0 8736 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2418
timestamp 1666464484
transform -1 0 8736 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2419
timestamp 1666464484
transform -1 0 8736 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2420
timestamp 1666464484
transform -1 0 8736 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2421
timestamp 1666464484
transform -1 0 8736 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2422
timestamp 1666464484
transform -1 0 8736 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2423
timestamp 1666464484
transform -1 0 7488 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2424
timestamp 1666464484
transform -1 0 7488 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2425
timestamp 1666464484
transform -1 0 7488 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2426
timestamp 1666464484
transform -1 0 7488 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2427
timestamp 1666464484
transform -1 0 7488 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2428
timestamp 1666464484
transform 1 0 7488 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2429
timestamp 1666464484
transform 1 0 7488 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2430
timestamp 1666464484
transform 1 0 7488 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2431
timestamp 1666464484
transform 1 0 7488 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2432
timestamp 1666464484
transform 1 0 7488 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2433
timestamp 1666464484
transform 1 0 7488 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2434
timestamp 1666464484
transform 1 0 7488 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2435
timestamp 1666464484
transform 1 0 7488 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2436
timestamp 1666464484
transform 1 0 7488 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2437
timestamp 1666464484
transform 1 0 7488 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2438
timestamp 1666464484
transform 1 0 7488 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2439
timestamp 1666464484
transform 1 0 7488 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2440
timestamp 1666464484
transform 1 0 7488 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2441
timestamp 1666464484
transform 1 0 7488 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2442
timestamp 1666464484
transform 1 0 7488 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2443
timestamp 1666464484
transform -1 0 7488 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2444
timestamp 1666464484
transform -1 0 7488 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2445
timestamp 1666464484
transform -1 0 7488 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2446
timestamp 1666464484
transform -1 0 7488 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2447
timestamp 1666464484
transform -1 0 7488 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2448
timestamp 1666464484
transform -1 0 7488 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2449
timestamp 1666464484
transform -1 0 7488 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2450
timestamp 1666464484
transform -1 0 7488 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2451
timestamp 1666464484
transform -1 0 7488 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2452
timestamp 1666464484
transform -1 0 7488 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2453
timestamp 1666464484
transform 1 0 6240 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2454
timestamp 1666464484
transform 1 0 6240 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2455
timestamp 1666464484
transform 1 0 6240 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2456
timestamp 1666464484
transform 1 0 6240 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2457
timestamp 1666464484
transform 1 0 6240 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2458
timestamp 1666464484
transform 1 0 6240 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2459
timestamp 1666464484
transform 1 0 6240 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2460
timestamp 1666464484
transform 1 0 6240 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2461
timestamp 1666464484
transform 1 0 6240 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2462
timestamp 1666464484
transform 1 0 6240 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2463
timestamp 1666464484
transform -1 0 8736 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2464
timestamp 1666464484
transform -1 0 8736 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2465
timestamp 1666464484
transform -1 0 8736 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2466
timestamp 1666464484
transform -1 0 8736 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2467
timestamp 1666464484
transform -1 0 8736 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2468
timestamp 1666464484
transform -1 0 8736 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2469
timestamp 1666464484
transform -1 0 8736 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2470
timestamp 1666464484
transform -1 0 8736 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2471
timestamp 1666464484
transform 1 0 6240 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2472
timestamp 1666464484
transform 1 0 6240 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2473
timestamp 1666464484
transform 1 0 6240 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2474
timestamp 1666464484
transform 1 0 6240 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2475
timestamp 1666464484
transform 1 0 8736 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2476
timestamp 1666464484
transform 1 0 8736 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2477
timestamp 1666464484
transform 1 0 3744 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2478
timestamp 1666464484
transform 1 0 3744 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2479
timestamp 1666464484
transform 1 0 3744 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2480
timestamp 1666464484
transform 1 0 3744 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2481
timestamp 1666464484
transform -1 0 3744 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2482
timestamp 1666464484
transform -1 0 3744 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2483
timestamp 1666464484
transform -1 0 3744 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2484
timestamp 1666464484
transform -1 0 3744 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2485
timestamp 1666464484
transform -1 0 3744 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2486
timestamp 1666464484
transform -1 0 3744 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2487
timestamp 1666464484
transform -1 0 3744 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2488
timestamp 1666464484
transform 1 0 3744 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2489
timestamp 1666464484
transform 1 0 3744 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2490
timestamp 1666464484
transform 1 0 3744 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2491
timestamp 1666464484
transform 1 0 1248 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2492
timestamp 1666464484
transform 1 0 1248 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2493
timestamp 1666464484
transform -1 0 1248 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2494
timestamp 1666464484
transform -1 0 1248 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2495
timestamp 1666464484
transform 1 0 0 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2496
timestamp 1666464484
transform 1 0 0 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2497
timestamp 1666464484
transform -1 0 1248 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2498
timestamp 1666464484
transform -1 0 1248 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2499
timestamp 1666464484
transform 1 0 0 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2500
timestamp 1666464484
transform -1 0 1248 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2501
timestamp 1666464484
transform 1 0 1248 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2502
timestamp 1666464484
transform 1 0 1248 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2503
timestamp 1666464484
transform 1 0 1248 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2504
timestamp 1666464484
transform -1 0 1248 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2505
timestamp 1666464484
transform 1 0 0 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2506
timestamp 1666464484
transform 1 0 0 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2507
timestamp 1666464484
transform -1 0 1248 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2508
timestamp 1666464484
transform 1 0 0 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2509
timestamp 1666464484
transform 1 0 0 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2510
timestamp 1666464484
transform 1 0 1248 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2511
timestamp 1666464484
transform 1 0 1248 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2512
timestamp 1666464484
transform 1 0 0 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2513
timestamp 1666464484
transform 1 0 0 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2514
timestamp 1666464484
transform 1 0 0 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2515
timestamp 1666464484
transform 1 0 1248 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2516
timestamp 1666464484
transform 1 0 1248 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2517
timestamp 1666464484
transform 1 0 1248 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2518
timestamp 1666464484
transform 1 0 1248 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2519
timestamp 1666464484
transform 1 0 1248 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2520
timestamp 1666464484
transform 1 0 0 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2521
timestamp 1666464484
transform -1 0 1248 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2522
timestamp 1666464484
transform -1 0 1248 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2523
timestamp 1666464484
transform -1 0 1248 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2524
timestamp 1666464484
transform -1 0 1248 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2525
timestamp 1666464484
transform -1 0 1248 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2526
timestamp 1666464484
transform 1 0 1248 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2527
timestamp 1666464484
transform -1 0 1248 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2528
timestamp 1666464484
transform 1 0 0 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2529
timestamp 1666464484
transform 1 0 0 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2530
timestamp 1666464484
transform 1 0 3744 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2531
timestamp 1666464484
transform 1 0 3744 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2532
timestamp 1666464484
transform -1 0 3744 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2533
timestamp 1666464484
transform 1 0 3744 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2534
timestamp 1666464484
transform -1 0 3744 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2535
timestamp 1666464484
transform -1 0 3744 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2536
timestamp 1666464484
transform 1 0 3744 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2537
timestamp 1666464484
transform 1 0 3744 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2538
timestamp 1666464484
transform 1 0 3744 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2539
timestamp 1666464484
transform -1 0 3744 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2540
timestamp 1666464484
transform -1 0 3744 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2541
timestamp 1666464484
transform -1 0 3744 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2542
timestamp 1666464484
transform -1 0 2496 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2543
timestamp 1666464484
transform 1 0 1248 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2544
timestamp 1666464484
transform 1 0 1248 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2545
timestamp 1666464484
transform -1 0 1248 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2546
timestamp 1666464484
transform 1 0 3744 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2547
timestamp 1666464484
transform 1 0 3744 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2548
timestamp 1666464484
transform -1 0 2496 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2549
timestamp 1666464484
transform -1 0 2496 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2550
timestamp 1666464484
transform 1 0 2496 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2551
timestamp 1666464484
transform 1 0 2496 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2552
timestamp 1666464484
transform 1 0 2496 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2553
timestamp 1666464484
transform 1 0 2496 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2554
timestamp 1666464484
transform 1 0 2496 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2555
timestamp 1666464484
transform 1 0 2496 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2556
timestamp 1666464484
transform 1 0 2496 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2557
timestamp 1666464484
transform 1 0 2496 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2558
timestamp 1666464484
transform -1 0 3744 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2559
timestamp 1666464484
transform -1 0 3744 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2560
timestamp 1666464484
transform -1 0 2496 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2561
timestamp 1666464484
transform -1 0 2496 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2562
timestamp 1666464484
transform -1 0 2496 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2563
timestamp 1666464484
transform -1 0 2496 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2564
timestamp 1666464484
transform 1 0 0 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2565
timestamp 1666464484
transform 1 0 0 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2566
timestamp 1666464484
transform -1 0 1248 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2567
timestamp 1666464484
transform -1 0 2496 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2568
timestamp 1666464484
transform -1 0 2496 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2569
timestamp 1666464484
transform -1 0 2496 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2570
timestamp 1666464484
transform -1 0 2496 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2571
timestamp 1666464484
transform 1 0 2496 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2572
timestamp 1666464484
transform 1 0 2496 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2573
timestamp 1666464484
transform 1 0 2496 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2574
timestamp 1666464484
transform 1 0 2496 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2575
timestamp 1666464484
transform 1 0 2496 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2576
timestamp 1666464484
transform 1 0 2496 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2577
timestamp 1666464484
transform 1 0 2496 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2578
timestamp 1666464484
transform -1 0 2496 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2579
timestamp 1666464484
transform -1 0 2496 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2580
timestamp 1666464484
transform -1 0 2496 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2581
timestamp 1666464484
transform -1 0 2496 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2582
timestamp 1666464484
transform -1 0 3744 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2583
timestamp 1666464484
transform -1 0 3744 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2584
timestamp 1666464484
transform -1 0 3744 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2585
timestamp 1666464484
transform -1 0 2496 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2586
timestamp 1666464484
transform 1 0 0 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2587
timestamp 1666464484
transform 1 0 0 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2588
timestamp 1666464484
transform 1 0 0 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2589
timestamp 1666464484
transform 1 0 0 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2590
timestamp 1666464484
transform 1 0 0 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2591
timestamp 1666464484
transform 1 0 0 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2592
timestamp 1666464484
transform -1 0 1248 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2593
timestamp 1666464484
transform -1 0 3744 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2594
timestamp 1666464484
transform -1 0 3744 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2595
timestamp 1666464484
transform -1 0 3744 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2596
timestamp 1666464484
transform -1 0 3744 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2597
timestamp 1666464484
transform 1 0 0 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2598
timestamp 1666464484
transform -1 0 1248 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2599
timestamp 1666464484
transform -1 0 1248 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2600
timestamp 1666464484
transform 1 0 0 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2601
timestamp 1666464484
transform 1 0 0 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2602
timestamp 1666464484
transform 1 0 0 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2603
timestamp 1666464484
transform 1 0 0 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2604
timestamp 1666464484
transform 1 0 0 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2605
timestamp 1666464484
transform -1 0 2496 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2606
timestamp 1666464484
transform -1 0 2496 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2607
timestamp 1666464484
transform -1 0 2496 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2608
timestamp 1666464484
transform -1 0 1248 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2609
timestamp 1666464484
transform -1 0 1248 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2610
timestamp 1666464484
transform -1 0 1248 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2611
timestamp 1666464484
transform -1 0 1248 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2612
timestamp 1666464484
transform -1 0 1248 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2613
timestamp 1666464484
transform -1 0 1248 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2614
timestamp 1666464484
transform -1 0 1248 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2615
timestamp 1666464484
transform 1 0 2496 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2616
timestamp 1666464484
transform 1 0 2496 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2617
timestamp 1666464484
transform 1 0 2496 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2618
timestamp 1666464484
transform 1 0 2496 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2619
timestamp 1666464484
transform 1 0 2496 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2620
timestamp 1666464484
transform -1 0 1248 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2621
timestamp 1666464484
transform -1 0 1248 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2622
timestamp 1666464484
transform -1 0 1248 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2623
timestamp 1666464484
transform -1 0 1248 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2624
timestamp 1666464484
transform -1 0 2496 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2625
timestamp 1666464484
transform -1 0 2496 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2626
timestamp 1666464484
transform 1 0 1248 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2627
timestamp 1666464484
transform 1 0 1248 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2628
timestamp 1666464484
transform 1 0 1248 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2629
timestamp 1666464484
transform 1 0 1248 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2630
timestamp 1666464484
transform 1 0 1248 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2631
timestamp 1666464484
transform 1 0 1248 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2632
timestamp 1666464484
transform 1 0 1248 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2633
timestamp 1666464484
transform 1 0 1248 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2634
timestamp 1666464484
transform 1 0 1248 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2635
timestamp 1666464484
transform 1 0 1248 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2636
timestamp 1666464484
transform 1 0 1248 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2637
timestamp 1666464484
transform -1 0 2496 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2638
timestamp 1666464484
transform -1 0 2496 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2639
timestamp 1666464484
transform -1 0 2496 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2640
timestamp 1666464484
transform 1 0 3744 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2641
timestamp 1666464484
transform 1 0 3744 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2642
timestamp 1666464484
transform 1 0 3744 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2643
timestamp 1666464484
transform 1 0 3744 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2644
timestamp 1666464484
transform 1 0 3744 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2645
timestamp 1666464484
transform 1 0 3744 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2646
timestamp 1666464484
transform 1 0 3744 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2647
timestamp 1666464484
transform 1 0 3744 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2648
timestamp 1666464484
transform 1 0 3744 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2649
timestamp 1666464484
transform 1 0 3744 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2650
timestamp 1666464484
transform 1 0 3744 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2651
timestamp 1666464484
transform 1 0 3744 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2652
timestamp 1666464484
transform 1 0 2496 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2653
timestamp 1666464484
transform 1 0 2496 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2654
timestamp 1666464484
transform 1 0 2496 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2655
timestamp 1666464484
transform 1 0 2496 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2656
timestamp 1666464484
transform 1 0 2496 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2657
timestamp 1666464484
transform 1 0 2496 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2658
timestamp 1666464484
transform 1 0 2496 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2659
timestamp 1666464484
transform 1 0 2496 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2660
timestamp 1666464484
transform 1 0 2496 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2661
timestamp 1666464484
transform -1 0 2496 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2662
timestamp 1666464484
transform -1 0 2496 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2663
timestamp 1666464484
transform 1 0 3744 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2664
timestamp 1666464484
transform 1 0 3744 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2665
timestamp 1666464484
transform -1 0 2496 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2666
timestamp 1666464484
transform 1 0 0 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2667
timestamp 1666464484
transform 1 0 1248 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2668
timestamp 1666464484
transform 1 0 1248 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2669
timestamp 1666464484
transform 1 0 1248 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2670
timestamp 1666464484
transform 1 0 0 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2671
timestamp 1666464484
transform -1 0 2496 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2672
timestamp 1666464484
transform -1 0 2496 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2673
timestamp 1666464484
transform -1 0 3744 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2674
timestamp 1666464484
transform -1 0 3744 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2675
timestamp 1666464484
transform -1 0 3744 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2676
timestamp 1666464484
transform -1 0 3744 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2677
timestamp 1666464484
transform -1 0 3744 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2678
timestamp 1666464484
transform -1 0 3744 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2679
timestamp 1666464484
transform -1 0 3744 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2680
timestamp 1666464484
transform -1 0 6240 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2681
timestamp 1666464484
transform -1 0 8736 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2682
timestamp 1666464484
transform 1 0 6240 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2683
timestamp 1666464484
transform -1 0 6240 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2684
timestamp 1666464484
transform -1 0 6240 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2685
timestamp 1666464484
transform 1 0 6240 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2686
timestamp 1666464484
transform 1 0 6240 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2687
timestamp 1666464484
transform -1 0 7488 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2688
timestamp 1666464484
transform -1 0 7488 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2689
timestamp 1666464484
transform -1 0 7488 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2690
timestamp 1666464484
transform -1 0 7488 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2691
timestamp 1666464484
transform -1 0 7488 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2692
timestamp 1666464484
transform -1 0 7488 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2693
timestamp 1666464484
transform -1 0 7488 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2694
timestamp 1666464484
transform -1 0 7488 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2695
timestamp 1666464484
transform -1 0 7488 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2696
timestamp 1666464484
transform 1 0 7488 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2697
timestamp 1666464484
transform 1 0 7488 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2698
timestamp 1666464484
transform 1 0 7488 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2699
timestamp 1666464484
transform 1 0 7488 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2700
timestamp 1666464484
transform 1 0 6240 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2701
timestamp 1666464484
transform 1 0 6240 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2702
timestamp 1666464484
transform 1 0 6240 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2703
timestamp 1666464484
transform 1 0 6240 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2704
timestamp 1666464484
transform -1 0 6240 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2705
timestamp 1666464484
transform -1 0 6240 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2706
timestamp 1666464484
transform -1 0 6240 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2707
timestamp 1666464484
transform -1 0 6240 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2708
timestamp 1666464484
transform 1 0 8736 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2709
timestamp 1666464484
transform 1 0 8736 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2710
timestamp 1666464484
transform 1 0 8736 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2711
timestamp 1666464484
transform 1 0 7488 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2712
timestamp 1666464484
transform 1 0 7488 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2713
timestamp 1666464484
transform -1 0 8736 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2714
timestamp 1666464484
transform -1 0 8736 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2715
timestamp 1666464484
transform -1 0 8736 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2716
timestamp 1666464484
transform -1 0 8736 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2717
timestamp 1666464484
transform -1 0 6240 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2718
timestamp 1666464484
transform -1 0 6240 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2719
timestamp 1666464484
transform -1 0 6240 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2720
timestamp 1666464484
transform -1 0 6240 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2721
timestamp 1666464484
transform -1 0 6240 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2722
timestamp 1666464484
transform -1 0 6240 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2723
timestamp 1666464484
transform -1 0 6240 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2724
timestamp 1666464484
transform 1 0 8736 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2725
timestamp 1666464484
transform 1 0 8736 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2726
timestamp 1666464484
transform 1 0 8736 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2727
timestamp 1666464484
transform 1 0 8736 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2728
timestamp 1666464484
transform 1 0 8736 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2729
timestamp 1666464484
transform 1 0 8736 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2730
timestamp 1666464484
transform 1 0 8736 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2731
timestamp 1666464484
transform 1 0 8736 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2732
timestamp 1666464484
transform 1 0 8736 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2733
timestamp 1666464484
transform 1 0 8736 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2734
timestamp 1666464484
transform 1 0 8736 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2735
timestamp 1666464484
transform -1 0 8736 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2736
timestamp 1666464484
transform -1 0 7488 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2737
timestamp 1666464484
transform 1 0 6240 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2738
timestamp 1666464484
transform 1 0 6240 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2739
timestamp 1666464484
transform 1 0 6240 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2740
timestamp 1666464484
transform 1 0 6240 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2741
timestamp 1666464484
transform -1 0 8736 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2742
timestamp 1666464484
transform -1 0 8736 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2743
timestamp 1666464484
transform -1 0 8736 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2744
timestamp 1666464484
transform -1 0 8736 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2745
timestamp 1666464484
transform -1 0 8736 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2746
timestamp 1666464484
transform -1 0 8736 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2747
timestamp 1666464484
transform 1 0 7488 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2748
timestamp 1666464484
transform -1 0 8736 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2749
timestamp 1666464484
transform -1 0 8736 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2750
timestamp 1666464484
transform 1 0 6240 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2751
timestamp 1666464484
transform 1 0 6240 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2752
timestamp 1666464484
transform 1 0 6240 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2753
timestamp 1666464484
transform -1 0 7488 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2754
timestamp 1666464484
transform -1 0 7488 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2755
timestamp 1666464484
transform -1 0 7488 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2756
timestamp 1666464484
transform -1 0 7488 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2757
timestamp 1666464484
transform 1 0 7488 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2758
timestamp 1666464484
transform 1 0 7488 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2759
timestamp 1666464484
transform 1 0 7488 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2760
timestamp 1666464484
transform 1 0 7488 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2761
timestamp 1666464484
transform 1 0 7488 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2762
timestamp 1666464484
transform 1 0 7488 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2763
timestamp 1666464484
transform 1 0 7488 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2764
timestamp 1666464484
transform -1 0 6240 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2765
timestamp 1666464484
transform -1 0 6240 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2766
timestamp 1666464484
transform -1 0 4992 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2767
timestamp 1666464484
transform -1 0 4992 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2768
timestamp 1666464484
transform -1 0 4992 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2769
timestamp 1666464484
transform -1 0 4992 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2770
timestamp 1666464484
transform -1 0 4992 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2771
timestamp 1666464484
transform -1 0 4992 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2772
timestamp 1666464484
transform -1 0 4992 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2773
timestamp 1666464484
transform -1 0 4992 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2774
timestamp 1666464484
transform -1 0 4992 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2775
timestamp 1666464484
transform -1 0 4992 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2776
timestamp 1666464484
transform -1 0 4992 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2777
timestamp 1666464484
transform -1 0 4992 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2778
timestamp 1666464484
transform -1 0 4992 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2779
timestamp 1666464484
transform -1 0 4992 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2780
timestamp 1666464484
transform -1 0 4992 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2781
timestamp 1666464484
transform -1 0 4992 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2782
timestamp 1666464484
transform -1 0 4992 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2783
timestamp 1666464484
transform 1 0 2496 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2784
timestamp 1666464484
transform 1 0 2496 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2785
timestamp 1666464484
transform 1 0 3744 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2786
timestamp 1666464484
transform 1 0 3744 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2787
timestamp 1666464484
transform 1 0 1248 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2788
timestamp 1666464484
transform 1 0 1248 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2789
timestamp 1666464484
transform 1 0 8736 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2790
timestamp 1666464484
transform 1 0 4992 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2791
timestamp 1666464484
transform 1 0 4992 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2792
timestamp 1666464484
transform 1 0 4992 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2793
timestamp 1666464484
transform 1 0 4992 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2794
timestamp 1666464484
transform 1 0 4992 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2795
timestamp 1666464484
transform 1 0 4992 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2796
timestamp 1666464484
transform 1 0 4992 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2797
timestamp 1666464484
transform 1 0 4992 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2798
timestamp 1666464484
transform 1 0 4992 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2799
timestamp 1666464484
transform 1 0 4992 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2800
timestamp 1666464484
transform 1 0 4992 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2801
timestamp 1666464484
transform 1 0 4992 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2802
timestamp 1666464484
transform 1 0 4992 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2803
timestamp 1666464484
transform 1 0 4992 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2804
timestamp 1666464484
transform 1 0 4992 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2805
timestamp 1666464484
transform 1 0 8736 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2806
timestamp 1666464484
transform -1 0 4992 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2807
timestamp 1666464484
transform -1 0 4992 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2808
timestamp 1666464484
transform -1 0 4992 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2809
timestamp 1666464484
transform -1 0 4992 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2810
timestamp 1666464484
transform -1 0 4992 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2811
timestamp 1666464484
transform -1 0 4992 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2812
timestamp 1666464484
transform -1 0 4992 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2813
timestamp 1666464484
transform -1 0 4992 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2814
timestamp 1666464484
transform -1 0 4992 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2815
timestamp 1666464484
transform -1 0 4992 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2816
timestamp 1666464484
transform -1 0 4992 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2817
timestamp 1666464484
transform -1 0 4992 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2818
timestamp 1666464484
transform -1 0 4992 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2819
timestamp 1666464484
transform -1 0 4992 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2820
timestamp 1666464484
transform 1 0 4992 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2821
timestamp 1666464484
transform 1 0 4992 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2822
timestamp 1666464484
transform 1 0 4992 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2823
timestamp 1666464484
transform 1 0 4992 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2824
timestamp 1666464484
transform 1 0 4992 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2825
timestamp 1666464484
transform 1 0 4992 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2826
timestamp 1666464484
transform 1 0 4992 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2827
timestamp 1666464484
transform 1 0 4992 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2828
timestamp 1666464484
transform 1 0 4992 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2829
timestamp 1666464484
transform 1 0 4992 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2830
timestamp 1666464484
transform 1 0 4992 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2831
timestamp 1666464484
transform 1 0 4992 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2832
timestamp 1666464484
transform 1 0 4992 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2833
timestamp 1666464484
transform 1 0 4992 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2834
timestamp 1666464484
transform 1 0 4992 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2835
timestamp 1666464484
transform 1 0 4992 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2836
timestamp 1666464484
transform -1 0 3744 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2837
timestamp 1666464484
transform -1 0 3744 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2838
timestamp 1666464484
transform 1 0 6240 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2839
timestamp 1666464484
transform 1 0 6240 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2840
timestamp 1666464484
transform 1 0 7488 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2841
timestamp 1666464484
transform 1 0 7488 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2842
timestamp 1666464484
transform -1 0 7488 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2843
timestamp 1666464484
transform -1 0 7488 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2844
timestamp 1666464484
transform -1 0 1248 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2845
timestamp 1666464484
transform -1 0 1248 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2846
timestamp 1666464484
transform 1 0 0 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2847
timestamp 1666464484
transform 1 0 0 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2848
timestamp 1666464484
transform -1 0 8736 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2849
timestamp 1666464484
transform -1 0 8736 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2850
timestamp 1666464484
transform -1 0 2496 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2851
timestamp 1666464484
transform -1 0 2496 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2852
timestamp 1666464484
transform 1 0 8736 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2853
timestamp 1666464484
transform 1 0 8736 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2854
timestamp 1666464484
transform 1 0 8736 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2855
timestamp 1666464484
transform 1 0 8736 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2856
timestamp 1666464484
transform 1 0 7488 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2857
timestamp 1666464484
transform 1 0 7488 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2858
timestamp 1666464484
transform 1 0 7488 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2859
timestamp 1666464484
transform -1 0 6240 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2860
timestamp 1666464484
transform -1 0 6240 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2861
timestamp 1666464484
transform -1 0 6240 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2862
timestamp 1666464484
transform 1 0 7488 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2863
timestamp 1666464484
transform 1 0 7488 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2864
timestamp 1666464484
transform 1 0 7488 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2865
timestamp 1666464484
transform 1 0 7488 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2866
timestamp 1666464484
transform 1 0 7488 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2867
timestamp 1666464484
transform 1 0 7488 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2868
timestamp 1666464484
transform 1 0 7488 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2869
timestamp 1666464484
transform 1 0 7488 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2870
timestamp 1666464484
transform 1 0 7488 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2871
timestamp 1666464484
transform 1 0 7488 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2872
timestamp 1666464484
transform -1 0 8736 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2873
timestamp 1666464484
transform -1 0 8736 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2874
timestamp 1666464484
transform -1 0 8736 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2875
timestamp 1666464484
transform -1 0 8736 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2876
timestamp 1666464484
transform -1 0 8736 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2877
timestamp 1666464484
transform -1 0 8736 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2878
timestamp 1666464484
transform -1 0 8736 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2879
timestamp 1666464484
transform -1 0 8736 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2880
timestamp 1666464484
transform -1 0 8736 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2881
timestamp 1666464484
transform -1 0 8736 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2882
timestamp 1666464484
transform -1 0 8736 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2883
timestamp 1666464484
transform -1 0 8736 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2884
timestamp 1666464484
transform -1 0 8736 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2885
timestamp 1666464484
transform -1 0 8736 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2886
timestamp 1666464484
transform 1 0 7488 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2887
timestamp 1666464484
transform 1 0 8736 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2888
timestamp 1666464484
transform -1 0 7488 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2889
timestamp 1666464484
transform -1 0 7488 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2890
timestamp 1666464484
transform -1 0 7488 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2891
timestamp 1666464484
transform -1 0 7488 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2892
timestamp 1666464484
transform -1 0 7488 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2893
timestamp 1666464484
transform -1 0 7488 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2894
timestamp 1666464484
transform -1 0 7488 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2895
timestamp 1666464484
transform -1 0 7488 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2896
timestamp 1666464484
transform -1 0 7488 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2897
timestamp 1666464484
transform -1 0 7488 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2898
timestamp 1666464484
transform -1 0 7488 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2899
timestamp 1666464484
transform -1 0 7488 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2900
timestamp 1666464484
transform -1 0 7488 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2901
timestamp 1666464484
transform -1 0 7488 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2902
timestamp 1666464484
transform 1 0 6240 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2903
timestamp 1666464484
transform 1 0 6240 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2904
timestamp 1666464484
transform 1 0 6240 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2905
timestamp 1666464484
transform 1 0 6240 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2906
timestamp 1666464484
transform 1 0 6240 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2907
timestamp 1666464484
transform 1 0 6240 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2908
timestamp 1666464484
transform 1 0 6240 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2909
timestamp 1666464484
transform 1 0 6240 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2910
timestamp 1666464484
transform 1 0 8736 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2911
timestamp 1666464484
transform 1 0 8736 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2912
timestamp 1666464484
transform -1 0 6240 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2913
timestamp 1666464484
transform -1 0 6240 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2914
timestamp 1666464484
transform -1 0 6240 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2915
timestamp 1666464484
transform -1 0 6240 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2916
timestamp 1666464484
transform -1 0 6240 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2917
timestamp 1666464484
transform -1 0 6240 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2918
timestamp 1666464484
transform -1 0 6240 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2919
timestamp 1666464484
transform -1 0 6240 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2920
timestamp 1666464484
transform -1 0 6240 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2921
timestamp 1666464484
transform -1 0 6240 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2922
timestamp 1666464484
transform -1 0 6240 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2923
timestamp 1666464484
transform 1 0 8736 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2924
timestamp 1666464484
transform 1 0 8736 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2925
timestamp 1666464484
transform 1 0 8736 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2926
timestamp 1666464484
transform 1 0 8736 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2927
timestamp 1666464484
transform 1 0 8736 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2928
timestamp 1666464484
transform 1 0 6240 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2929
timestamp 1666464484
transform 1 0 6240 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2930
timestamp 1666464484
transform 1 0 6240 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2931
timestamp 1666464484
transform 1 0 6240 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2932
timestamp 1666464484
transform 1 0 6240 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2933
timestamp 1666464484
transform 1 0 6240 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2934
timestamp 1666464484
transform 1 0 8736 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2935
timestamp 1666464484
transform 1 0 8736 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2936
timestamp 1666464484
transform 1 0 1248 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2937
timestamp 1666464484
transform 1 0 1248 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2938
timestamp 1666464484
transform -1 0 3744 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2939
timestamp 1666464484
transform -1 0 3744 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2940
timestamp 1666464484
transform -1 0 1248 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2941
timestamp 1666464484
transform -1 0 1248 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2942
timestamp 1666464484
transform -1 0 1248 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2943
timestamp 1666464484
transform -1 0 1248 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2944
timestamp 1666464484
transform 1 0 1248 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2945
timestamp 1666464484
transform 1 0 1248 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2946
timestamp 1666464484
transform 1 0 1248 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2947
timestamp 1666464484
transform 1 0 1248 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2948
timestamp 1666464484
transform -1 0 1248 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2949
timestamp 1666464484
transform -1 0 3744 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2950
timestamp 1666464484
transform -1 0 3744 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2951
timestamp 1666464484
transform -1 0 3744 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2952
timestamp 1666464484
transform 1 0 2496 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2953
timestamp 1666464484
transform 1 0 2496 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2954
timestamp 1666464484
transform 1 0 2496 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2955
timestamp 1666464484
transform 1 0 2496 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2956
timestamp 1666464484
transform 1 0 2496 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2957
timestamp 1666464484
transform 1 0 2496 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2958
timestamp 1666464484
transform 1 0 2496 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2959
timestamp 1666464484
transform 1 0 2496 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2960
timestamp 1666464484
transform 1 0 2496 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2961
timestamp 1666464484
transform 1 0 2496 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2962
timestamp 1666464484
transform 1 0 2496 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2963
timestamp 1666464484
transform 1 0 2496 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2964
timestamp 1666464484
transform 1 0 2496 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2965
timestamp 1666464484
transform 1 0 2496 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2966
timestamp 1666464484
transform -1 0 3744 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2967
timestamp 1666464484
transform -1 0 3744 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2968
timestamp 1666464484
transform -1 0 3744 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2969
timestamp 1666464484
transform -1 0 3744 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2970
timestamp 1666464484
transform -1 0 3744 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2971
timestamp 1666464484
transform -1 0 3744 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2972
timestamp 1666464484
transform -1 0 3744 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2973
timestamp 1666464484
transform -1 0 1248 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2974
timestamp 1666464484
transform -1 0 1248 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2975
timestamp 1666464484
transform -1 0 1248 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2976
timestamp 1666464484
transform -1 0 1248 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2977
timestamp 1666464484
transform -1 0 1248 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2978
timestamp 1666464484
transform -1 0 2496 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2979
timestamp 1666464484
transform -1 0 2496 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2980
timestamp 1666464484
transform -1 0 2496 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2981
timestamp 1666464484
transform -1 0 2496 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2982
timestamp 1666464484
transform -1 0 2496 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2983
timestamp 1666464484
transform -1 0 2496 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2984
timestamp 1666464484
transform -1 0 2496 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2985
timestamp 1666464484
transform -1 0 2496 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2986
timestamp 1666464484
transform -1 0 2496 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2987
timestamp 1666464484
transform -1 0 2496 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2988
timestamp 1666464484
transform -1 0 2496 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2989
timestamp 1666464484
transform -1 0 2496 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2990
timestamp 1666464484
transform -1 0 2496 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2991
timestamp 1666464484
transform -1 0 2496 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2992
timestamp 1666464484
transform -1 0 1248 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2993
timestamp 1666464484
transform -1 0 1248 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2994
timestamp 1666464484
transform -1 0 1248 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2995
timestamp 1666464484
transform -1 0 1248 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2996
timestamp 1666464484
transform 1 0 1248 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2997
timestamp 1666464484
transform 1 0 3744 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2998
timestamp 1666464484
transform 1 0 3744 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_2999
timestamp 1666464484
transform 1 0 3744 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3000
timestamp 1666464484
transform 1 0 3744 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3001
timestamp 1666464484
transform 1 0 3744 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3002
timestamp 1666464484
transform 1 0 0 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3003
timestamp 1666464484
transform 1 0 0 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3004
timestamp 1666464484
transform 1 0 0 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3005
timestamp 1666464484
transform 1 0 0 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3006
timestamp 1666464484
transform 1 0 0 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3007
timestamp 1666464484
transform 1 0 0 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3008
timestamp 1666464484
transform 1 0 0 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3009
timestamp 1666464484
transform 1 0 0 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3010
timestamp 1666464484
transform 1 0 0 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3011
timestamp 1666464484
transform 1 0 0 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3012
timestamp 1666464484
transform 1 0 0 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3013
timestamp 1666464484
transform 1 0 0 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3014
timestamp 1666464484
transform 1 0 0 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3015
timestamp 1666464484
transform 1 0 0 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3016
timestamp 1666464484
transform -1 0 3744 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3017
timestamp 1666464484
transform -1 0 3744 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3018
timestamp 1666464484
transform 1 0 1248 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3019
timestamp 1666464484
transform 1 0 1248 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3020
timestamp 1666464484
transform 1 0 1248 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3021
timestamp 1666464484
transform 1 0 1248 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3022
timestamp 1666464484
transform 1 0 1248 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3023
timestamp 1666464484
transform 1 0 1248 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3024
timestamp 1666464484
transform 1 0 1248 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3025
timestamp 1666464484
transform 1 0 3744 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3026
timestamp 1666464484
transform 1 0 3744 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3027
timestamp 1666464484
transform 1 0 3744 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3028
timestamp 1666464484
transform 1 0 3744 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3029
timestamp 1666464484
transform 1 0 3744 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3030
timestamp 1666464484
transform 1 0 3744 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3031
timestamp 1666464484
transform 1 0 3744 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3032
timestamp 1666464484
transform 1 0 3744 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3033
timestamp 1666464484
transform 1 0 3744 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3034
timestamp 1666464484
transform 1 0 2496 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3035
timestamp 1666464484
transform 1 0 2496 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3036
timestamp 1666464484
transform 1 0 2496 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3037
timestamp 1666464484
transform 1 0 2496 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3038
timestamp 1666464484
transform 1 0 2496 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3039
timestamp 1666464484
transform 1 0 2496 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3040
timestamp 1666464484
transform 1 0 2496 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3041
timestamp 1666464484
transform 1 0 2496 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3042
timestamp 1666464484
transform 1 0 2496 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3043
timestamp 1666464484
transform 1 0 2496 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3044
timestamp 1666464484
transform 1 0 2496 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3045
timestamp 1666464484
transform 1 0 2496 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3046
timestamp 1666464484
transform 1 0 2496 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3047
timestamp 1666464484
transform 1 0 2496 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3048
timestamp 1666464484
transform 1 0 0 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3049
timestamp 1666464484
transform 1 0 0 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3050
timestamp 1666464484
transform 1 0 0 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3051
timestamp 1666464484
transform 1 0 0 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3052
timestamp 1666464484
transform -1 0 2496 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3053
timestamp 1666464484
transform -1 0 1248 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3054
timestamp 1666464484
transform 1 0 3744 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3055
timestamp 1666464484
transform 1 0 3744 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3056
timestamp 1666464484
transform 1 0 3744 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3057
timestamp 1666464484
transform 1 0 3744 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3058
timestamp 1666464484
transform 1 0 3744 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3059
timestamp 1666464484
transform 1 0 3744 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3060
timestamp 1666464484
transform 1 0 3744 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3061
timestamp 1666464484
transform -1 0 1248 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3062
timestamp 1666464484
transform -1 0 1248 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3063
timestamp 1666464484
transform -1 0 1248 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3064
timestamp 1666464484
transform -1 0 1248 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3065
timestamp 1666464484
transform -1 0 1248 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3066
timestamp 1666464484
transform -1 0 2496 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3067
timestamp 1666464484
transform -1 0 2496 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3068
timestamp 1666464484
transform -1 0 2496 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3069
timestamp 1666464484
transform -1 0 2496 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3070
timestamp 1666464484
transform -1 0 2496 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3071
timestamp 1666464484
transform 1 0 1248 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3072
timestamp 1666464484
transform 1 0 1248 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3073
timestamp 1666464484
transform 1 0 1248 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3074
timestamp 1666464484
transform 1 0 1248 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3075
timestamp 1666464484
transform 1 0 1248 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3076
timestamp 1666464484
transform -1 0 3744 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3077
timestamp 1666464484
transform -1 0 3744 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3078
timestamp 1666464484
transform -1 0 3744 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3079
timestamp 1666464484
transform -1 0 3744 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3080
timestamp 1666464484
transform -1 0 3744 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3081
timestamp 1666464484
transform -1 0 3744 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3082
timestamp 1666464484
transform -1 0 3744 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3083
timestamp 1666464484
transform -1 0 3744 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3084
timestamp 1666464484
transform -1 0 3744 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3085
timestamp 1666464484
transform -1 0 3744 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3086
timestamp 1666464484
transform -1 0 3744 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3087
timestamp 1666464484
transform -1 0 3744 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3088
timestamp 1666464484
transform -1 0 3744 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3089
timestamp 1666464484
transform -1 0 3744 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3090
timestamp 1666464484
transform 1 0 1248 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3091
timestamp 1666464484
transform 1 0 1248 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3092
timestamp 1666464484
transform 1 0 1248 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3093
timestamp 1666464484
transform 1 0 1248 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3094
timestamp 1666464484
transform 1 0 1248 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3095
timestamp 1666464484
transform 1 0 1248 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3096
timestamp 1666464484
transform 1 0 1248 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3097
timestamp 1666464484
transform 1 0 1248 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3098
timestamp 1666464484
transform 1 0 1248 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3099
timestamp 1666464484
transform -1 0 1248 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3100
timestamp 1666464484
transform -1 0 1248 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3101
timestamp 1666464484
transform -1 0 1248 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3102
timestamp 1666464484
transform -1 0 1248 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3103
timestamp 1666464484
transform -1 0 1248 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3104
timestamp 1666464484
transform -1 0 1248 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3105
timestamp 1666464484
transform -1 0 1248 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3106
timestamp 1666464484
transform -1 0 1248 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3107
timestamp 1666464484
transform -1 0 2496 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3108
timestamp 1666464484
transform -1 0 2496 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3109
timestamp 1666464484
transform -1 0 2496 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3110
timestamp 1666464484
transform -1 0 2496 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3111
timestamp 1666464484
transform -1 0 2496 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3112
timestamp 1666464484
transform -1 0 2496 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3113
timestamp 1666464484
transform -1 0 2496 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3114
timestamp 1666464484
transform -1 0 2496 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3115
timestamp 1666464484
transform 1 0 3744 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3116
timestamp 1666464484
transform 1 0 3744 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3117
timestamp 1666464484
transform 1 0 3744 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3118
timestamp 1666464484
transform 1 0 3744 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3119
timestamp 1666464484
transform 1 0 3744 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3120
timestamp 1666464484
transform 1 0 3744 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3121
timestamp 1666464484
transform 1 0 3744 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3122
timestamp 1666464484
transform 1 0 0 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3123
timestamp 1666464484
transform 1 0 0 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3124
timestamp 1666464484
transform 1 0 0 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3125
timestamp 1666464484
transform 1 0 0 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3126
timestamp 1666464484
transform 1 0 0 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3127
timestamp 1666464484
transform 1 0 0 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3128
timestamp 1666464484
transform 1 0 0 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3129
timestamp 1666464484
transform 1 0 0 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3130
timestamp 1666464484
transform 1 0 0 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3131
timestamp 1666464484
transform 1 0 0 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3132
timestamp 1666464484
transform 1 0 6240 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3133
timestamp 1666464484
transform 1 0 6240 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3134
timestamp 1666464484
transform -1 0 7488 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3135
timestamp 1666464484
transform -1 0 7488 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3136
timestamp 1666464484
transform -1 0 7488 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3137
timestamp 1666464484
transform -1 0 7488 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3138
timestamp 1666464484
transform -1 0 7488 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3139
timestamp 1666464484
transform -1 0 7488 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3140
timestamp 1666464484
transform -1 0 7488 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3141
timestamp 1666464484
transform -1 0 7488 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3142
timestamp 1666464484
transform -1 0 7488 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3143
timestamp 1666464484
transform -1 0 7488 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3144
timestamp 1666464484
transform -1 0 7488 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3145
timestamp 1666464484
transform 1 0 7488 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3146
timestamp 1666464484
transform -1 0 7488 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3147
timestamp 1666464484
transform -1 0 7488 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3148
timestamp 1666464484
transform -1 0 8736 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3149
timestamp 1666464484
transform -1 0 8736 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3150
timestamp 1666464484
transform -1 0 8736 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3151
timestamp 1666464484
transform -1 0 8736 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3152
timestamp 1666464484
transform -1 0 8736 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3153
timestamp 1666464484
transform -1 0 8736 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3154
timestamp 1666464484
transform 1 0 7488 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3155
timestamp 1666464484
transform 1 0 7488 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3156
timestamp 1666464484
transform 1 0 7488 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3157
timestamp 1666464484
transform 1 0 7488 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3158
timestamp 1666464484
transform 1 0 7488 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3159
timestamp 1666464484
transform 1 0 7488 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3160
timestamp 1666464484
transform 1 0 7488 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3161
timestamp 1666464484
transform 1 0 7488 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3162
timestamp 1666464484
transform 1 0 7488 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3163
timestamp 1666464484
transform 1 0 7488 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3164
timestamp 1666464484
transform 1 0 7488 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3165
timestamp 1666464484
transform 1 0 7488 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3166
timestamp 1666464484
transform 1 0 7488 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3167
timestamp 1666464484
transform 1 0 6240 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3168
timestamp 1666464484
transform 1 0 6240 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3169
timestamp 1666464484
transform 1 0 6240 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3170
timestamp 1666464484
transform 1 0 8736 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3171
timestamp 1666464484
transform 1 0 8736 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3172
timestamp 1666464484
transform 1 0 8736 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3173
timestamp 1666464484
transform 1 0 8736 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3174
timestamp 1666464484
transform 1 0 8736 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3175
timestamp 1666464484
transform 1 0 8736 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3176
timestamp 1666464484
transform 1 0 8736 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3177
timestamp 1666464484
transform 1 0 8736 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3178
timestamp 1666464484
transform 1 0 8736 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3179
timestamp 1666464484
transform 1 0 8736 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3180
timestamp 1666464484
transform 1 0 8736 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3181
timestamp 1666464484
transform 1 0 8736 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3182
timestamp 1666464484
transform 1 0 8736 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3183
timestamp 1666464484
transform 1 0 8736 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3184
timestamp 1666464484
transform -1 0 8736 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3185
timestamp 1666464484
transform -1 0 8736 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3186
timestamp 1666464484
transform -1 0 8736 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3187
timestamp 1666464484
transform -1 0 8736 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3188
timestamp 1666464484
transform -1 0 8736 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3189
timestamp 1666464484
transform -1 0 8736 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3190
timestamp 1666464484
transform -1 0 8736 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3191
timestamp 1666464484
transform -1 0 8736 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3192
timestamp 1666464484
transform 1 0 6240 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3193
timestamp 1666464484
transform 1 0 6240 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3194
timestamp 1666464484
transform 1 0 6240 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3195
timestamp 1666464484
transform 1 0 6240 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3196
timestamp 1666464484
transform -1 0 6240 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3197
timestamp 1666464484
transform -1 0 6240 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3198
timestamp 1666464484
transform -1 0 6240 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3199
timestamp 1666464484
transform -1 0 7488 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3200
timestamp 1666464484
transform 1 0 6240 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3201
timestamp 1666464484
transform 1 0 6240 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3202
timestamp 1666464484
transform 1 0 6240 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3203
timestamp 1666464484
transform -1 0 6240 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3204
timestamp 1666464484
transform -1 0 6240 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3205
timestamp 1666464484
transform -1 0 6240 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3206
timestamp 1666464484
transform -1 0 6240 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3207
timestamp 1666464484
transform -1 0 6240 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3208
timestamp 1666464484
transform -1 0 6240 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3209
timestamp 1666464484
transform -1 0 6240 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3210
timestamp 1666464484
transform -1 0 6240 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3211
timestamp 1666464484
transform -1 0 6240 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3212
timestamp 1666464484
transform -1 0 6240 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3213
timestamp 1666464484
transform -1 0 6240 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3214
timestamp 1666464484
transform 1 0 6240 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3215
timestamp 1666464484
transform 1 0 6240 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3216
timestamp 1666464484
transform 1 0 2496 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3217
timestamp 1666464484
transform 1 0 2496 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3218
timestamp 1666464484
transform -1 0 2496 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3219
timestamp 1666464484
transform 1 0 4992 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3220
timestamp 1666464484
transform 1 0 4992 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3221
timestamp 1666464484
transform 1 0 4992 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3222
timestamp 1666464484
transform 1 0 4992 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3223
timestamp 1666464484
transform 1 0 4992 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3224
timestamp 1666464484
transform 1 0 4992 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3225
timestamp 1666464484
transform 1 0 4992 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3226
timestamp 1666464484
transform 1 0 4992 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3227
timestamp 1666464484
transform 1 0 4992 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3228
timestamp 1666464484
transform 1 0 4992 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3229
timestamp 1666464484
transform 1 0 4992 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3230
timestamp 1666464484
transform 1 0 4992 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3231
timestamp 1666464484
transform 1 0 4992 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3232
timestamp 1666464484
transform 1 0 4992 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3233
timestamp 1666464484
transform 1 0 4992 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3234
timestamp 1666464484
transform 1 0 4992 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3235
timestamp 1666464484
transform 1 0 4992 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3236
timestamp 1666464484
transform 1 0 4992 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3237
timestamp 1666464484
transform 1 0 4992 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3238
timestamp 1666464484
transform 1 0 4992 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3239
timestamp 1666464484
transform 1 0 4992 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3240
timestamp 1666464484
transform 1 0 4992 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3241
timestamp 1666464484
transform 1 0 4992 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3242
timestamp 1666464484
transform 1 0 4992 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3243
timestamp 1666464484
transform 1 0 4992 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3244
timestamp 1666464484
transform 1 0 4992 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3245
timestamp 1666464484
transform 1 0 4992 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3246
timestamp 1666464484
transform 1 0 4992 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3247
timestamp 1666464484
transform 1 0 4992 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3248
timestamp 1666464484
transform 1 0 4992 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3249
timestamp 1666464484
transform -1 0 8736 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3250
timestamp 1666464484
transform -1 0 8736 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3251
timestamp 1666464484
transform -1 0 7488 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3252
timestamp 1666464484
transform -1 0 7488 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3253
timestamp 1666464484
transform 1 0 0 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3254
timestamp 1666464484
transform 1 0 0 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3255
timestamp 1666464484
transform 1 0 3744 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3256
timestamp 1666464484
transform 1 0 3744 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3257
timestamp 1666464484
transform -1 0 6240 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3258
timestamp 1666464484
transform -1 0 6240 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3259
timestamp 1666464484
transform -1 0 3744 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3260
timestamp 1666464484
transform -1 0 3744 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3261
timestamp 1666464484
transform 1 0 7488 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3262
timestamp 1666464484
transform 1 0 7488 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3263
timestamp 1666464484
transform -1 0 4992 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3264
timestamp 1666464484
transform -1 0 4992 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3265
timestamp 1666464484
transform -1 0 4992 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3266
timestamp 1666464484
transform -1 0 4992 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3267
timestamp 1666464484
transform -1 0 4992 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3268
timestamp 1666464484
transform -1 0 4992 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3269
timestamp 1666464484
transform -1 0 4992 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3270
timestamp 1666464484
transform -1 0 4992 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3271
timestamp 1666464484
transform -1 0 4992 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3272
timestamp 1666464484
transform -1 0 4992 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3273
timestamp 1666464484
transform -1 0 4992 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3274
timestamp 1666464484
transform -1 0 4992 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3275
timestamp 1666464484
transform -1 0 4992 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3276
timestamp 1666464484
transform -1 0 4992 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3277
timestamp 1666464484
transform -1 0 4992 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3278
timestamp 1666464484
transform -1 0 4992 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3279
timestamp 1666464484
transform -1 0 4992 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3280
timestamp 1666464484
transform -1 0 4992 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3281
timestamp 1666464484
transform -1 0 4992 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3282
timestamp 1666464484
transform -1 0 4992 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3283
timestamp 1666464484
transform -1 0 4992 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3284
timestamp 1666464484
transform -1 0 4992 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3285
timestamp 1666464484
transform -1 0 4992 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3286
timestamp 1666464484
transform -1 0 4992 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3287
timestamp 1666464484
transform -1 0 4992 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3288
timestamp 1666464484
transform -1 0 4992 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3289
timestamp 1666464484
transform -1 0 4992 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3290
timestamp 1666464484
transform -1 0 4992 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3291
timestamp 1666464484
transform -1 0 4992 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3292
timestamp 1666464484
transform -1 0 4992 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3293
timestamp 1666464484
transform 1 0 8736 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3294
timestamp 1666464484
transform 1 0 8736 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3295
timestamp 1666464484
transform -1 0 1248 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3296
timestamp 1666464484
transform -1 0 1248 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3297
timestamp 1666464484
transform 1 0 1248 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3298
timestamp 1666464484
transform 1 0 1248 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3299
timestamp 1666464484
transform -1 0 2496 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3300
timestamp 1666464484
transform 1 0 6240 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3301
timestamp 1666464484
transform 1 0 6240 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3302
timestamp 1666464484
transform 1 0 16224 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3303
timestamp 1666464484
transform 1 0 16224 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3304
timestamp 1666464484
transform 1 0 16224 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3305
timestamp 1666464484
transform 1 0 16224 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3306
timestamp 1666464484
transform 1 0 16224 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3307
timestamp 1666464484
transform 1 0 16224 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3308
timestamp 1666464484
transform 1 0 16224 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3309
timestamp 1666464484
transform 1 0 16224 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3310
timestamp 1666464484
transform -1 0 16224 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3311
timestamp 1666464484
transform -1 0 16224 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3312
timestamp 1666464484
transform 1 0 17472 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3313
timestamp 1666464484
transform 1 0 17472 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3314
timestamp 1666464484
transform 1 0 17472 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3315
timestamp 1666464484
transform 1 0 17472 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3316
timestamp 1666464484
transform 1 0 17472 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3317
timestamp 1666464484
transform 1 0 17472 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3318
timestamp 1666464484
transform 1 0 17472 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3319
timestamp 1666464484
transform 1 0 17472 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3320
timestamp 1666464484
transform 1 0 17472 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3321
timestamp 1666464484
transform 1 0 17472 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3322
timestamp 1666464484
transform 1 0 17472 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3323
timestamp 1666464484
transform 1 0 17472 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3324
timestamp 1666464484
transform 1 0 17472 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3325
timestamp 1666464484
transform 1 0 17472 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3326
timestamp 1666464484
transform -1 0 16224 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3327
timestamp 1666464484
transform -1 0 16224 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3328
timestamp 1666464484
transform -1 0 16224 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3329
timestamp 1666464484
transform -1 0 16224 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3330
timestamp 1666464484
transform -1 0 16224 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3331
timestamp 1666464484
transform -1 0 16224 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3332
timestamp 1666464484
transform -1 0 16224 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3333
timestamp 1666464484
transform -1 0 16224 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3334
timestamp 1666464484
transform -1 0 16224 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3335
timestamp 1666464484
transform -1 0 16224 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3336
timestamp 1666464484
transform -1 0 16224 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3337
timestamp 1666464484
transform -1 0 16224 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3338
timestamp 1666464484
transform 1 0 16224 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3339
timestamp 1666464484
transform 1 0 16224 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3340
timestamp 1666464484
transform 1 0 16224 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3341
timestamp 1666464484
transform 1 0 16224 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3342
timestamp 1666464484
transform 1 0 16224 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3343
timestamp 1666464484
transform 1 0 16224 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3344
timestamp 1666464484
transform -1 0 17472 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3345
timestamp 1666464484
transform -1 0 17472 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3346
timestamp 1666464484
transform -1 0 18720 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3347
timestamp 1666464484
transform -1 0 18720 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3348
timestamp 1666464484
transform -1 0 18720 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3349
timestamp 1666464484
transform -1 0 18720 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3350
timestamp 1666464484
transform -1 0 18720 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3351
timestamp 1666464484
transform -1 0 18720 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3352
timestamp 1666464484
transform -1 0 18720 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3353
timestamp 1666464484
transform -1 0 18720 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3354
timestamp 1666464484
transform -1 0 18720 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3355
timestamp 1666464484
transform -1 0 18720 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3356
timestamp 1666464484
transform -1 0 18720 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3357
timestamp 1666464484
transform -1 0 18720 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3358
timestamp 1666464484
transform -1 0 18720 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3359
timestamp 1666464484
transform -1 0 18720 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3360
timestamp 1666464484
transform -1 0 17472 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3361
timestamp 1666464484
transform -1 0 17472 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3362
timestamp 1666464484
transform -1 0 17472 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3363
timestamp 1666464484
transform -1 0 17472 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3364
timestamp 1666464484
transform -1 0 17472 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3365
timestamp 1666464484
transform -1 0 17472 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3366
timestamp 1666464484
transform -1 0 17472 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3367
timestamp 1666464484
transform -1 0 17472 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3368
timestamp 1666464484
transform 1 0 18720 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3369
timestamp 1666464484
transform 1 0 18720 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3370
timestamp 1666464484
transform 1 0 18720 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3371
timestamp 1666464484
transform 1 0 18720 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3372
timestamp 1666464484
transform 1 0 18720 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3373
timestamp 1666464484
transform 1 0 18720 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3374
timestamp 1666464484
transform 1 0 18720 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3375
timestamp 1666464484
transform 1 0 18720 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3376
timestamp 1666464484
transform 1 0 18720 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3377
timestamp 1666464484
transform 1 0 18720 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3378
timestamp 1666464484
transform 1 0 18720 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3379
timestamp 1666464484
transform 1 0 18720 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3380
timestamp 1666464484
transform 1 0 18720 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3381
timestamp 1666464484
transform 1 0 18720 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3382
timestamp 1666464484
transform -1 0 17472 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3383
timestamp 1666464484
transform -1 0 17472 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3384
timestamp 1666464484
transform -1 0 17472 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3385
timestamp 1666464484
transform -1 0 17472 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3386
timestamp 1666464484
transform 1 0 11232 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3387
timestamp 1666464484
transform 1 0 11232 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3388
timestamp 1666464484
transform 1 0 11232 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3389
timestamp 1666464484
transform -1 0 12480 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3390
timestamp 1666464484
transform -1 0 12480 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3391
timestamp 1666464484
transform -1 0 12480 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3392
timestamp 1666464484
transform -1 0 12480 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3393
timestamp 1666464484
transform -1 0 12480 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3394
timestamp 1666464484
transform -1 0 12480 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3395
timestamp 1666464484
transform -1 0 12480 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3396
timestamp 1666464484
transform -1 0 12480 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3397
timestamp 1666464484
transform -1 0 13728 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3398
timestamp 1666464484
transform -1 0 13728 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3399
timestamp 1666464484
transform -1 0 13728 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3400
timestamp 1666464484
transform -1 0 13728 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3401
timestamp 1666464484
transform -1 0 13728 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3402
timestamp 1666464484
transform -1 0 13728 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3403
timestamp 1666464484
transform -1 0 13728 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3404
timestamp 1666464484
transform -1 0 11232 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3405
timestamp 1666464484
transform -1 0 11232 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3406
timestamp 1666464484
transform -1 0 11232 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3407
timestamp 1666464484
transform -1 0 11232 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3408
timestamp 1666464484
transform -1 0 11232 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3409
timestamp 1666464484
transform -1 0 11232 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3410
timestamp 1666464484
transform -1 0 11232 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3411
timestamp 1666464484
transform -1 0 11232 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3412
timestamp 1666464484
transform -1 0 11232 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3413
timestamp 1666464484
transform -1 0 11232 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3414
timestamp 1666464484
transform -1 0 11232 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3415
timestamp 1666464484
transform -1 0 11232 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3416
timestamp 1666464484
transform -1 0 11232 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3417
timestamp 1666464484
transform -1 0 11232 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3418
timestamp 1666464484
transform -1 0 13728 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3419
timestamp 1666464484
transform -1 0 13728 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3420
timestamp 1666464484
transform -1 0 13728 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3421
timestamp 1666464484
transform -1 0 13728 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3422
timestamp 1666464484
transform -1 0 13728 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3423
timestamp 1666464484
transform -1 0 13728 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3424
timestamp 1666464484
transform -1 0 13728 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3425
timestamp 1666464484
transform 1 0 11232 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3426
timestamp 1666464484
transform 1 0 11232 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3427
timestamp 1666464484
transform 1 0 11232 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3428
timestamp 1666464484
transform 1 0 11232 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3429
timestamp 1666464484
transform 1 0 11232 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3430
timestamp 1666464484
transform 1 0 12480 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3431
timestamp 1666464484
transform 1 0 12480 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3432
timestamp 1666464484
transform 1 0 12480 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3433
timestamp 1666464484
transform 1 0 12480 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3434
timestamp 1666464484
transform 1 0 12480 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3435
timestamp 1666464484
transform 1 0 12480 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3436
timestamp 1666464484
transform 1 0 12480 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3437
timestamp 1666464484
transform 1 0 12480 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3438
timestamp 1666464484
transform 1 0 12480 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3439
timestamp 1666464484
transform 1 0 12480 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3440
timestamp 1666464484
transform 1 0 11232 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3441
timestamp 1666464484
transform 1 0 11232 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3442
timestamp 1666464484
transform -1 0 12480 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3443
timestamp 1666464484
transform -1 0 12480 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3444
timestamp 1666464484
transform -1 0 12480 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3445
timestamp 1666464484
transform -1 0 12480 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3446
timestamp 1666464484
transform 1 0 12480 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3447
timestamp 1666464484
transform 1 0 12480 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3448
timestamp 1666464484
transform 1 0 13728 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3449
timestamp 1666464484
transform 1 0 13728 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3450
timestamp 1666464484
transform 1 0 13728 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3451
timestamp 1666464484
transform 1 0 13728 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3452
timestamp 1666464484
transform 1 0 13728 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3453
timestamp 1666464484
transform 1 0 13728 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3454
timestamp 1666464484
transform 1 0 13728 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3455
timestamp 1666464484
transform 1 0 13728 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3456
timestamp 1666464484
transform 1 0 13728 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3457
timestamp 1666464484
transform 1 0 13728 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3458
timestamp 1666464484
transform 1 0 13728 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3459
timestamp 1666464484
transform 1 0 13728 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3460
timestamp 1666464484
transform 1 0 13728 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3461
timestamp 1666464484
transform 1 0 13728 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3462
timestamp 1666464484
transform 1 0 12480 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3463
timestamp 1666464484
transform 1 0 12480 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3464
timestamp 1666464484
transform 1 0 11232 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3465
timestamp 1666464484
transform -1 0 12480 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3466
timestamp 1666464484
transform -1 0 12480 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3467
timestamp 1666464484
transform 1 0 11232 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3468
timestamp 1666464484
transform 1 0 11232 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3469
timestamp 1666464484
transform 1 0 11232 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3470
timestamp 1666464484
transform -1 0 12480 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3471
timestamp 1666464484
transform -1 0 12480 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3472
timestamp 1666464484
transform -1 0 11232 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3473
timestamp 1666464484
transform -1 0 11232 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3474
timestamp 1666464484
transform -1 0 11232 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3475
timestamp 1666464484
transform -1 0 11232 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3476
timestamp 1666464484
transform -1 0 11232 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3477
timestamp 1666464484
transform -1 0 11232 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3478
timestamp 1666464484
transform -1 0 11232 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3479
timestamp 1666464484
transform -1 0 11232 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3480
timestamp 1666464484
transform -1 0 11232 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3481
timestamp 1666464484
transform -1 0 11232 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3482
timestamp 1666464484
transform -1 0 11232 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3483
timestamp 1666464484
transform -1 0 11232 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3484
timestamp 1666464484
transform -1 0 11232 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3485
timestamp 1666464484
transform -1 0 11232 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3486
timestamp 1666464484
transform -1 0 12480 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3487
timestamp 1666464484
transform -1 0 12480 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3488
timestamp 1666464484
transform -1 0 12480 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3489
timestamp 1666464484
transform -1 0 12480 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3490
timestamp 1666464484
transform 1 0 11232 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3491
timestamp 1666464484
transform 1 0 11232 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3492
timestamp 1666464484
transform 1 0 11232 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3493
timestamp 1666464484
transform 1 0 11232 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3494
timestamp 1666464484
transform 1 0 11232 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3495
timestamp 1666464484
transform 1 0 11232 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3496
timestamp 1666464484
transform 1 0 11232 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3497
timestamp 1666464484
transform 1 0 11232 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3498
timestamp 1666464484
transform 1 0 11232 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3499
timestamp 1666464484
transform 1 0 11232 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3500
timestamp 1666464484
transform 1 0 11232 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3501
timestamp 1666464484
transform 1 0 11232 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3502
timestamp 1666464484
transform 1 0 13728 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3503
timestamp 1666464484
transform 1 0 13728 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3504
timestamp 1666464484
transform 1 0 13728 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3505
timestamp 1666464484
transform 1 0 13728 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3506
timestamp 1666464484
transform 1 0 13728 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3507
timestamp 1666464484
transform 1 0 13728 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3508
timestamp 1666464484
transform 1 0 13728 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3509
timestamp 1666464484
transform 1 0 13728 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3510
timestamp 1666464484
transform 1 0 13728 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3511
timestamp 1666464484
transform 1 0 13728 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3512
timestamp 1666464484
transform 1 0 13728 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3513
timestamp 1666464484
transform 1 0 13728 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3514
timestamp 1666464484
transform 1 0 13728 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3515
timestamp 1666464484
transform 1 0 13728 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3516
timestamp 1666464484
transform 1 0 11232 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3517
timestamp 1666464484
transform 1 0 11232 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3518
timestamp 1666464484
transform -1 0 12480 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3519
timestamp 1666464484
transform -1 0 12480 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3520
timestamp 1666464484
transform -1 0 13728 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3521
timestamp 1666464484
transform -1 0 13728 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3522
timestamp 1666464484
transform -1 0 13728 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3523
timestamp 1666464484
transform -1 0 13728 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3524
timestamp 1666464484
transform -1 0 13728 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3525
timestamp 1666464484
transform -1 0 13728 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3526
timestamp 1666464484
transform -1 0 13728 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3527
timestamp 1666464484
transform -1 0 13728 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3528
timestamp 1666464484
transform -1 0 13728 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3529
timestamp 1666464484
transform -1 0 13728 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3530
timestamp 1666464484
transform -1 0 13728 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3531
timestamp 1666464484
transform -1 0 13728 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3532
timestamp 1666464484
transform -1 0 13728 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3533
timestamp 1666464484
transform -1 0 13728 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3534
timestamp 1666464484
transform -1 0 12480 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3535
timestamp 1666464484
transform -1 0 12480 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3536
timestamp 1666464484
transform 1 0 12480 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3537
timestamp 1666464484
transform 1 0 12480 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3538
timestamp 1666464484
transform 1 0 12480 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3539
timestamp 1666464484
transform 1 0 12480 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3540
timestamp 1666464484
transform 1 0 12480 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3541
timestamp 1666464484
transform 1 0 12480 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3542
timestamp 1666464484
transform 1 0 12480 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3543
timestamp 1666464484
transform 1 0 12480 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3544
timestamp 1666464484
transform 1 0 12480 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3545
timestamp 1666464484
transform 1 0 12480 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3546
timestamp 1666464484
transform 1 0 12480 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3547
timestamp 1666464484
transform 1 0 12480 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3548
timestamp 1666464484
transform 1 0 12480 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3549
timestamp 1666464484
transform 1 0 12480 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3550
timestamp 1666464484
transform -1 0 12480 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3551
timestamp 1666464484
transform -1 0 12480 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3552
timestamp 1666464484
transform -1 0 12480 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3553
timestamp 1666464484
transform -1 0 12480 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3554
timestamp 1666464484
transform -1 0 16224 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3555
timestamp 1666464484
transform -1 0 16224 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3556
timestamp 1666464484
transform 1 0 16224 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3557
timestamp 1666464484
transform 1 0 16224 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3558
timestamp 1666464484
transform 1 0 16224 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3559
timestamp 1666464484
transform 1 0 16224 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3560
timestamp 1666464484
transform 1 0 16224 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3561
timestamp 1666464484
transform 1 0 16224 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3562
timestamp 1666464484
transform 1 0 16224 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3563
timestamp 1666464484
transform 1 0 16224 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3564
timestamp 1666464484
transform 1 0 16224 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3565
timestamp 1666464484
transform 1 0 16224 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3566
timestamp 1666464484
transform 1 0 16224 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3567
timestamp 1666464484
transform 1 0 16224 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3568
timestamp 1666464484
transform 1 0 16224 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3569
timestamp 1666464484
transform 1 0 16224 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3570
timestamp 1666464484
transform -1 0 16224 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3571
timestamp 1666464484
transform -1 0 16224 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3572
timestamp 1666464484
transform -1 0 16224 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3573
timestamp 1666464484
transform -1 0 16224 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3574
timestamp 1666464484
transform 1 0 18720 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3575
timestamp 1666464484
transform 1 0 18720 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3576
timestamp 1666464484
transform 1 0 18720 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3577
timestamp 1666464484
transform 1 0 18720 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3578
timestamp 1666464484
transform 1 0 18720 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3579
timestamp 1666464484
transform 1 0 18720 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3580
timestamp 1666464484
transform 1 0 18720 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3581
timestamp 1666464484
transform 1 0 18720 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3582
timestamp 1666464484
transform 1 0 18720 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3583
timestamp 1666464484
transform 1 0 18720 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3584
timestamp 1666464484
transform 1 0 18720 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3585
timestamp 1666464484
transform 1 0 18720 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3586
timestamp 1666464484
transform 1 0 18720 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3587
timestamp 1666464484
transform 1 0 18720 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3588
timestamp 1666464484
transform -1 0 16224 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3589
timestamp 1666464484
transform -1 0 16224 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3590
timestamp 1666464484
transform -1 0 16224 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3591
timestamp 1666464484
transform -1 0 16224 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3592
timestamp 1666464484
transform -1 0 18720 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3593
timestamp 1666464484
transform -1 0 18720 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3594
timestamp 1666464484
transform -1 0 18720 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3595
timestamp 1666464484
transform -1 0 18720 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3596
timestamp 1666464484
transform -1 0 18720 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3597
timestamp 1666464484
transform -1 0 18720 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3598
timestamp 1666464484
transform -1 0 18720 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3599
timestamp 1666464484
transform -1 0 18720 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3600
timestamp 1666464484
transform -1 0 18720 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3601
timestamp 1666464484
transform -1 0 18720 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3602
timestamp 1666464484
transform -1 0 18720 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3603
timestamp 1666464484
transform -1 0 18720 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3604
timestamp 1666464484
transform -1 0 18720 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3605
timestamp 1666464484
transform -1 0 18720 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3606
timestamp 1666464484
transform -1 0 16224 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3607
timestamp 1666464484
transform -1 0 16224 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3608
timestamp 1666464484
transform 1 0 17472 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3609
timestamp 1666464484
transform 1 0 17472 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3610
timestamp 1666464484
transform 1 0 17472 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3611
timestamp 1666464484
transform 1 0 17472 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3612
timestamp 1666464484
transform 1 0 17472 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3613
timestamp 1666464484
transform 1 0 17472 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3614
timestamp 1666464484
transform 1 0 17472 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3615
timestamp 1666464484
transform 1 0 17472 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3616
timestamp 1666464484
transform 1 0 17472 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3617
timestamp 1666464484
transform 1 0 17472 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3618
timestamp 1666464484
transform 1 0 17472 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3619
timestamp 1666464484
transform 1 0 17472 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3620
timestamp 1666464484
transform 1 0 17472 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3621
timestamp 1666464484
transform 1 0 17472 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3622
timestamp 1666464484
transform -1 0 16224 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3623
timestamp 1666464484
transform -1 0 16224 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3624
timestamp 1666464484
transform -1 0 17472 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3625
timestamp 1666464484
transform -1 0 17472 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3626
timestamp 1666464484
transform -1 0 17472 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3627
timestamp 1666464484
transform -1 0 17472 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3628
timestamp 1666464484
transform -1 0 17472 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3629
timestamp 1666464484
transform -1 0 17472 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3630
timestamp 1666464484
transform -1 0 17472 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3631
timestamp 1666464484
transform -1 0 17472 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3632
timestamp 1666464484
transform -1 0 17472 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3633
timestamp 1666464484
transform -1 0 17472 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3634
timestamp 1666464484
transform -1 0 17472 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3635
timestamp 1666464484
transform -1 0 17472 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3636
timestamp 1666464484
transform -1 0 17472 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3637
timestamp 1666464484
transform -1 0 17472 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3638
timestamp 1666464484
transform -1 0 14976 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3639
timestamp 1666464484
transform -1 0 14976 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3640
timestamp 1666464484
transform -1 0 11232 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3641
timestamp 1666464484
transform -1 0 11232 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3642
timestamp 1666464484
transform -1 0 14976 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3643
timestamp 1666464484
transform -1 0 14976 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3644
timestamp 1666464484
transform -1 0 14976 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3645
timestamp 1666464484
transform -1 0 14976 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3646
timestamp 1666464484
transform -1 0 14976 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3647
timestamp 1666464484
transform -1 0 14976 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3648
timestamp 1666464484
transform -1 0 14976 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3649
timestamp 1666464484
transform -1 0 14976 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3650
timestamp 1666464484
transform 1 0 13728 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3651
timestamp 1666464484
transform 1 0 13728 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3652
timestamp 1666464484
transform 1 0 11232 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3653
timestamp 1666464484
transform 1 0 11232 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3654
timestamp 1666464484
transform -1 0 13728 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3655
timestamp 1666464484
transform -1 0 13728 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3656
timestamp 1666464484
transform 1 0 12480 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3657
timestamp 1666464484
transform 1 0 12480 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3658
timestamp 1666464484
transform 1 0 18720 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3659
timestamp 1666464484
transform 1 0 18720 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3660
timestamp 1666464484
transform -1 0 12480 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3661
timestamp 1666464484
transform -1 0 12480 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3662
timestamp 1666464484
transform -1 0 18720 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3663
timestamp 1666464484
transform -1 0 18720 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3664
timestamp 1666464484
transform 1 0 17472 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3665
timestamp 1666464484
transform 1 0 17472 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3666
timestamp 1666464484
transform -1 0 17472 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3667
timestamp 1666464484
transform -1 0 17472 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3668
timestamp 1666464484
transform 1 0 16224 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3669
timestamp 1666464484
transform 1 0 16224 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3670
timestamp 1666464484
transform -1 0 16224 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3671
timestamp 1666464484
transform -1 0 16224 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3672
timestamp 1666464484
transform 1 0 14976 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3673
timestamp 1666464484
transform 1 0 14976 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3674
timestamp 1666464484
transform 1 0 14976 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3675
timestamp 1666464484
transform 1 0 14976 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3676
timestamp 1666464484
transform 1 0 14976 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3677
timestamp 1666464484
transform 1 0 14976 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3678
timestamp 1666464484
transform 1 0 14976 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3679
timestamp 1666464484
transform 1 0 14976 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3680
timestamp 1666464484
transform 1 0 14976 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3681
timestamp 1666464484
transform 1 0 14976 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3682
timestamp 1666464484
transform 1 0 14976 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3683
timestamp 1666464484
transform 1 0 14976 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3684
timestamp 1666464484
transform 1 0 14976 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3685
timestamp 1666464484
transform 1 0 14976 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3686
timestamp 1666464484
transform 1 0 14976 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3687
timestamp 1666464484
transform 1 0 14976 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3688
timestamp 1666464484
transform 1 0 14976 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3689
timestamp 1666464484
transform 1 0 14976 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3690
timestamp 1666464484
transform 1 0 14976 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3691
timestamp 1666464484
transform 1 0 14976 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3692
timestamp 1666464484
transform 1 0 14976 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3693
timestamp 1666464484
transform 1 0 14976 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3694
timestamp 1666464484
transform 1 0 14976 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3695
timestamp 1666464484
transform 1 0 14976 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3696
timestamp 1666464484
transform 1 0 14976 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3697
timestamp 1666464484
transform 1 0 14976 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3698
timestamp 1666464484
transform 1 0 14976 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3699
timestamp 1666464484
transform 1 0 14976 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3700
timestamp 1666464484
transform 1 0 14976 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3701
timestamp 1666464484
transform 1 0 14976 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3702
timestamp 1666464484
transform -1 0 14976 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3703
timestamp 1666464484
transform -1 0 14976 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3704
timestamp 1666464484
transform -1 0 14976 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3705
timestamp 1666464484
transform -1 0 14976 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3706
timestamp 1666464484
transform -1 0 14976 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3707
timestamp 1666464484
transform -1 0 14976 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3708
timestamp 1666464484
transform -1 0 14976 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3709
timestamp 1666464484
transform -1 0 14976 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3710
timestamp 1666464484
transform -1 0 14976 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3711
timestamp 1666464484
transform -1 0 14976 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3712
timestamp 1666464484
transform -1 0 14976 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3713
timestamp 1666464484
transform -1 0 14976 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3714
timestamp 1666464484
transform -1 0 14976 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3715
timestamp 1666464484
transform -1 0 14976 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3716
timestamp 1666464484
transform -1 0 14976 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3717
timestamp 1666464484
transform -1 0 14976 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3718
timestamp 1666464484
transform -1 0 14976 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3719
timestamp 1666464484
transform -1 0 14976 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3720
timestamp 1666464484
transform -1 0 14976 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3721
timestamp 1666464484
transform -1 0 14976 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3722
timestamp 1666464484
transform 1 0 2496 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3723
timestamp 1666464484
transform 1 0 2496 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3724
timestamp 1666464484
transform -1 0 11232 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3725
timestamp 1666464484
transform -1 0 11232 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3726
timestamp 1666464484
transform 1 0 4992 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3727
timestamp 1666464484
transform 1 0 4992 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3728
timestamp 1666464484
transform 1 0 9984 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3729
timestamp 1666464484
transform 1 0 9984 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3730
timestamp 1666464484
transform 1 0 9984 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3731
timestamp 1666464484
transform 1 0 9984 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3732
timestamp 1666464484
transform 1 0 9984 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3733
timestamp 1666464484
transform 1 0 9984 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3734
timestamp 1666464484
transform 1 0 9984 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3735
timestamp 1666464484
transform 1 0 9984 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3736
timestamp 1666464484
transform 1 0 9984 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3737
timestamp 1666464484
transform 1 0 9984 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3738
timestamp 1666464484
transform 1 0 9984 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3739
timestamp 1666464484
transform 1 0 9984 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3740
timestamp 1666464484
transform 1 0 9984 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3741
timestamp 1666464484
transform 1 0 9984 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3742
timestamp 1666464484
transform 1 0 9984 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3743
timestamp 1666464484
transform 1 0 9984 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3744
timestamp 1666464484
transform 1 0 9984 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3745
timestamp 1666464484
transform 1 0 9984 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3746
timestamp 1666464484
transform 1 0 9984 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3747
timestamp 1666464484
transform 1 0 9984 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3748
timestamp 1666464484
transform 1 0 9984 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3749
timestamp 1666464484
transform 1 0 9984 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3750
timestamp 1666464484
transform 1 0 9984 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3751
timestamp 1666464484
transform 1 0 9984 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3752
timestamp 1666464484
transform 1 0 9984 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3753
timestamp 1666464484
transform 1 0 9984 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3754
timestamp 1666464484
transform 1 0 9984 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3755
timestamp 1666464484
transform 1 0 9984 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3756
timestamp 1666464484
transform 1 0 9984 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3757
timestamp 1666464484
transform 1 0 9984 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3758
timestamp 1666464484
transform 1 0 9984 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3759
timestamp 1666464484
transform 1 0 9984 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3760
timestamp 1666464484
transform 1 0 9984 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3761
timestamp 1666464484
transform 1 0 9984 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3762
timestamp 1666464484
transform 1 0 9984 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3763
timestamp 1666464484
transform 1 0 9984 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3764
timestamp 1666464484
transform 1 0 9984 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3765
timestamp 1666464484
transform 1 0 9984 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3766
timestamp 1666464484
transform 1 0 9984 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3767
timestamp 1666464484
transform 1 0 9984 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3768
timestamp 1666464484
transform 1 0 9984 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3769
timestamp 1666464484
transform 1 0 9984 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3770
timestamp 1666464484
transform 1 0 9984 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3771
timestamp 1666464484
transform 1 0 9984 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3772
timestamp 1666464484
transform 1 0 9984 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3773
timestamp 1666464484
transform 1 0 9984 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3774
timestamp 1666464484
transform 1 0 9984 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3775
timestamp 1666464484
transform 1 0 9984 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3776
timestamp 1666464484
transform 1 0 9984 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3777
timestamp 1666464484
transform 1 0 9984 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3778
timestamp 1666464484
transform 1 0 9984 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3779
timestamp 1666464484
transform 1 0 9984 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3780
timestamp 1666464484
transform 1 0 9984 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3781
timestamp 1666464484
transform 1 0 9984 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3782
timestamp 1666464484
transform 1 0 9984 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3783
timestamp 1666464484
transform 1 0 9984 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3784
timestamp 1666464484
transform 1 0 9984 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3785
timestamp 1666464484
transform 1 0 9984 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3786
timestamp 1666464484
transform 1 0 9984 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3787
timestamp 1666464484
transform 1 0 9984 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3788
timestamp 1666464484
transform 1 0 9984 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3789
timestamp 1666464484
transform 1 0 9984 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3790
timestamp 1666464484
transform 1 0 9984 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3791
timestamp 1666464484
transform 1 0 0 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3792
timestamp 1666464484
transform 1 0 0 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3793
timestamp 1666464484
transform -1 0 9984 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3794
timestamp 1666464484
transform -1 0 9984 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3795
timestamp 1666464484
transform -1 0 9984 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3796
timestamp 1666464484
transform -1 0 9984 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3797
timestamp 1666464484
transform -1 0 9984 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3798
timestamp 1666464484
transform -1 0 9984 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3799
timestamp 1666464484
transform -1 0 9984 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3800
timestamp 1666464484
transform -1 0 9984 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3801
timestamp 1666464484
transform -1 0 9984 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3802
timestamp 1666464484
transform -1 0 9984 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3803
timestamp 1666464484
transform -1 0 9984 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3804
timestamp 1666464484
transform -1 0 9984 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3805
timestamp 1666464484
transform -1 0 9984 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3806
timestamp 1666464484
transform -1 0 9984 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3807
timestamp 1666464484
transform -1 0 9984 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3808
timestamp 1666464484
transform -1 0 9984 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3809
timestamp 1666464484
transform -1 0 9984 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3810
timestamp 1666464484
transform -1 0 9984 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3811
timestamp 1666464484
transform -1 0 9984 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3812
timestamp 1666464484
transform -1 0 9984 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3813
timestamp 1666464484
transform -1 0 9984 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3814
timestamp 1666464484
transform -1 0 9984 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3815
timestamp 1666464484
transform -1 0 9984 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3816
timestamp 1666464484
transform -1 0 9984 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3817
timestamp 1666464484
transform -1 0 9984 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3818
timestamp 1666464484
transform -1 0 9984 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3819
timestamp 1666464484
transform -1 0 9984 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3820
timestamp 1666464484
transform -1 0 9984 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3821
timestamp 1666464484
transform -1 0 9984 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3822
timestamp 1666464484
transform -1 0 9984 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3823
timestamp 1666464484
transform -1 0 9984 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3824
timestamp 1666464484
transform -1 0 9984 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3825
timestamp 1666464484
transform -1 0 9984 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3826
timestamp 1666464484
transform 1 0 18720 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3827
timestamp 1666464484
transform 1 0 18720 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3828
timestamp 1666464484
transform -1 0 9984 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3829
timestamp 1666464484
transform -1 0 9984 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3830
timestamp 1666464484
transform -1 0 9984 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3831
timestamp 1666464484
transform -1 0 9984 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3832
timestamp 1666464484
transform -1 0 9984 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3833
timestamp 1666464484
transform -1 0 9984 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3834
timestamp 1666464484
transform -1 0 9984 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3835
timestamp 1666464484
transform -1 0 9984 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3836
timestamp 1666464484
transform -1 0 9984 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3837
timestamp 1666464484
transform -1 0 9984 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3838
timestamp 1666464484
transform -1 0 9984 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3839
timestamp 1666464484
transform -1 0 9984 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3840
timestamp 1666464484
transform -1 0 9984 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3841
timestamp 1666464484
transform -1 0 9984 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3842
timestamp 1666464484
transform -1 0 9984 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3843
timestamp 1666464484
transform -1 0 9984 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3844
timestamp 1666464484
transform -1 0 9984 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3845
timestamp 1666464484
transform -1 0 9984 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3846
timestamp 1666464484
transform -1 0 9984 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3847
timestamp 1666464484
transform -1 0 9984 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3848
timestamp 1666464484
transform -1 0 9984 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3849
timestamp 1666464484
transform -1 0 9984 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3850
timestamp 1666464484
transform -1 0 9984 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3851
timestamp 1666464484
transform -1 0 9984 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3852
timestamp 1666464484
transform -1 0 9984 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3853
timestamp 1666464484
transform -1 0 9984 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3854
timestamp 1666464484
transform -1 0 9984 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3855
timestamp 1666464484
transform -1 0 9984 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3856
timestamp 1666464484
transform -1 0 9984 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3857
timestamp 1666464484
transform -1 0 9984 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3858
timestamp 1666464484
transform -1 0 18720 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3859
timestamp 1666464484
transform -1 0 18720 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3860
timestamp 1666464484
transform -1 0 4992 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3861
timestamp 1666464484
transform -1 0 4992 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3862
timestamp 1666464484
transform 1 0 8736 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3863
timestamp 1666464484
transform 1 0 8736 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3864
timestamp 1666464484
transform 1 0 17472 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3865
timestamp 1666464484
transform 1 0 17472 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3866
timestamp 1666464484
transform -1 0 17472 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3867
timestamp 1666464484
transform -1 0 17472 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3868
timestamp 1666464484
transform -1 0 2496 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3869
timestamp 1666464484
transform -1 0 2496 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3870
timestamp 1666464484
transform -1 0 8736 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3871
timestamp 1666464484
transform -1 0 8736 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3872
timestamp 1666464484
transform 1 0 16224 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3873
timestamp 1666464484
transform 1 0 16224 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3874
timestamp 1666464484
transform -1 0 16224 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3875
timestamp 1666464484
transform -1 0 16224 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3876
timestamp 1666464484
transform 1 0 3744 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3877
timestamp 1666464484
transform 1 0 3744 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3878
timestamp 1666464484
transform 1 0 7488 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3879
timestamp 1666464484
transform 1 0 7488 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3880
timestamp 1666464484
transform 1 0 14976 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3881
timestamp 1666464484
transform 1 0 14976 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3882
timestamp 1666464484
transform -1 0 14976 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3883
timestamp 1666464484
transform -1 0 14976 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3884
timestamp 1666464484
transform -1 0 1248 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3885
timestamp 1666464484
transform -1 0 1248 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3886
timestamp 1666464484
transform -1 0 7488 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3887
timestamp 1666464484
transform -1 0 7488 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3888
timestamp 1666464484
transform 1 0 13728 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3889
timestamp 1666464484
transform 1 0 13728 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3890
timestamp 1666464484
transform -1 0 3744 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3891
timestamp 1666464484
transform -1 0 13728 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3892
timestamp 1666464484
transform -1 0 13728 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3893
timestamp 1666464484
transform -1 0 3744 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3894
timestamp 1666464484
transform 1 0 6240 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3895
timestamp 1666464484
transform 1 0 6240 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3896
timestamp 1666464484
transform 1 0 12480 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3897
timestamp 1666464484
transform 1 0 12480 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3898
timestamp 1666464484
transform -1 0 12480 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3899
timestamp 1666464484
transform -1 0 12480 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3900
timestamp 1666464484
transform 1 0 1248 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3901
timestamp 1666464484
transform 1 0 1248 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3902
timestamp 1666464484
transform -1 0 6240 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3903
timestamp 1666464484
transform -1 0 6240 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3904
timestamp 1666464484
transform 1 0 11232 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3905
timestamp 1666464484
transform 1 0 11232 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3906
timestamp 1666464484
transform 1 0 17472 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3907
timestamp 1666464484
transform 1 0 17472 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3908
timestamp 1666464484
transform 1 0 17472 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3909
timestamp 1666464484
transform 1 0 17472 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3910
timestamp 1666464484
transform 1 0 17472 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3911
timestamp 1666464484
transform 1 0 17472 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3912
timestamp 1666464484
transform 1 0 17472 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3913
timestamp 1666464484
transform -1 0 17472 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3914
timestamp 1666464484
transform -1 0 17472 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3915
timestamp 1666464484
transform -1 0 17472 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3916
timestamp 1666464484
transform -1 0 17472 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3917
timestamp 1666464484
transform -1 0 17472 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3918
timestamp 1666464484
transform -1 0 18720 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3919
timestamp 1666464484
transform -1 0 18720 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3920
timestamp 1666464484
transform -1 0 18720 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3921
timestamp 1666464484
transform -1 0 18720 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3922
timestamp 1666464484
transform -1 0 18720 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3923
timestamp 1666464484
transform -1 0 18720 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3924
timestamp 1666464484
transform -1 0 18720 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3925
timestamp 1666464484
transform -1 0 18720 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3926
timestamp 1666464484
transform -1 0 18720 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3927
timestamp 1666464484
transform -1 0 18720 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3928
timestamp 1666464484
transform -1 0 18720 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3929
timestamp 1666464484
transform -1 0 18720 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3930
timestamp 1666464484
transform -1 0 18720 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3931
timestamp 1666464484
transform -1 0 18720 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3932
timestamp 1666464484
transform -1 0 17472 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3933
timestamp 1666464484
transform -1 0 17472 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3934
timestamp 1666464484
transform -1 0 17472 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3935
timestamp 1666464484
transform -1 0 17472 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3936
timestamp 1666464484
transform 1 0 18720 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3937
timestamp 1666464484
transform 1 0 18720 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3938
timestamp 1666464484
transform 1 0 18720 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3939
timestamp 1666464484
transform 1 0 18720 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3940
timestamp 1666464484
transform -1 0 16224 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3941
timestamp 1666464484
transform -1 0 16224 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3942
timestamp 1666464484
transform -1 0 16224 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3943
timestamp 1666464484
transform -1 0 16224 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3944
timestamp 1666464484
transform -1 0 16224 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3945
timestamp 1666464484
transform 1 0 16224 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3946
timestamp 1666464484
transform 1 0 16224 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3947
timestamp 1666464484
transform 1 0 16224 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3948
timestamp 1666464484
transform 1 0 16224 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3949
timestamp 1666464484
transform 1 0 16224 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3950
timestamp 1666464484
transform 1 0 16224 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3951
timestamp 1666464484
transform 1 0 16224 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3952
timestamp 1666464484
transform 1 0 16224 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3953
timestamp 1666464484
transform 1 0 16224 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3954
timestamp 1666464484
transform 1 0 16224 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3955
timestamp 1666464484
transform 1 0 16224 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3956
timestamp 1666464484
transform 1 0 16224 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3957
timestamp 1666464484
transform 1 0 16224 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3958
timestamp 1666464484
transform 1 0 16224 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3959
timestamp 1666464484
transform -1 0 16224 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3960
timestamp 1666464484
transform -1 0 16224 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3961
timestamp 1666464484
transform -1 0 16224 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3962
timestamp 1666464484
transform -1 0 16224 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3963
timestamp 1666464484
transform -1 0 16224 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3964
timestamp 1666464484
transform -1 0 16224 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3965
timestamp 1666464484
transform -1 0 16224 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3966
timestamp 1666464484
transform -1 0 16224 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3967
timestamp 1666464484
transform -1 0 16224 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3968
timestamp 1666464484
transform 1 0 18720 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3969
timestamp 1666464484
transform 1 0 18720 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3970
timestamp 1666464484
transform 1 0 18720 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3971
timestamp 1666464484
transform 1 0 18720 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3972
timestamp 1666464484
transform 1 0 18720 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3973
timestamp 1666464484
transform 1 0 18720 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3974
timestamp 1666464484
transform 1 0 18720 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3975
timestamp 1666464484
transform 1 0 18720 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3976
timestamp 1666464484
transform 1 0 18720 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3977
timestamp 1666464484
transform 1 0 18720 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3978
timestamp 1666464484
transform -1 0 17472 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3979
timestamp 1666464484
transform -1 0 17472 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3980
timestamp 1666464484
transform -1 0 17472 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3981
timestamp 1666464484
transform -1 0 17472 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3982
timestamp 1666464484
transform -1 0 17472 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3983
timestamp 1666464484
transform 1 0 17472 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3984
timestamp 1666464484
transform 1 0 17472 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3985
timestamp 1666464484
transform 1 0 17472 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3986
timestamp 1666464484
transform 1 0 17472 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3987
timestamp 1666464484
transform 1 0 17472 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3988
timestamp 1666464484
transform 1 0 17472 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3989
timestamp 1666464484
transform 1 0 17472 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3990
timestamp 1666464484
transform 1 0 11232 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3991
timestamp 1666464484
transform 1 0 11232 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3992
timestamp 1666464484
transform 1 0 11232 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3993
timestamp 1666464484
transform 1 0 11232 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3994
timestamp 1666464484
transform -1 0 13728 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3995
timestamp 1666464484
transform -1 0 13728 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3996
timestamp 1666464484
transform -1 0 13728 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3997
timestamp 1666464484
transform -1 0 13728 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3998
timestamp 1666464484
transform -1 0 13728 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_3999
timestamp 1666464484
transform -1 0 13728 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4000
timestamp 1666464484
transform -1 0 13728 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4001
timestamp 1666464484
transform -1 0 13728 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4002
timestamp 1666464484
transform -1 0 13728 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4003
timestamp 1666464484
transform -1 0 13728 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4004
timestamp 1666464484
transform -1 0 12480 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4005
timestamp 1666464484
transform -1 0 12480 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4006
timestamp 1666464484
transform -1 0 12480 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4007
timestamp 1666464484
transform -1 0 12480 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4008
timestamp 1666464484
transform -1 0 12480 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4009
timestamp 1666464484
transform -1 0 12480 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4010
timestamp 1666464484
transform 1 0 11232 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4011
timestamp 1666464484
transform 1 0 11232 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4012
timestamp 1666464484
transform 1 0 11232 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4013
timestamp 1666464484
transform 1 0 11232 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4014
timestamp 1666464484
transform 1 0 11232 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4015
timestamp 1666464484
transform -1 0 12480 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4016
timestamp 1666464484
transform -1 0 12480 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4017
timestamp 1666464484
transform -1 0 12480 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4018
timestamp 1666464484
transform -1 0 12480 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4019
timestamp 1666464484
transform 1 0 11232 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4020
timestamp 1666464484
transform 1 0 11232 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4021
timestamp 1666464484
transform 1 0 11232 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4022
timestamp 1666464484
transform 1 0 11232 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4023
timestamp 1666464484
transform 1 0 11232 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4024
timestamp 1666464484
transform -1 0 11232 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4025
timestamp 1666464484
transform -1 0 11232 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4026
timestamp 1666464484
transform -1 0 11232 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4027
timestamp 1666464484
transform -1 0 11232 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4028
timestamp 1666464484
transform -1 0 11232 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4029
timestamp 1666464484
transform -1 0 13728 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4030
timestamp 1666464484
transform -1 0 13728 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4031
timestamp 1666464484
transform 1 0 13728 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4032
timestamp 1666464484
transform 1 0 13728 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4033
timestamp 1666464484
transform 1 0 12480 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4034
timestamp 1666464484
transform 1 0 12480 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4035
timestamp 1666464484
transform 1 0 12480 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4036
timestamp 1666464484
transform 1 0 12480 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4037
timestamp 1666464484
transform 1 0 13728 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4038
timestamp 1666464484
transform 1 0 13728 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4039
timestamp 1666464484
transform 1 0 13728 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4040
timestamp 1666464484
transform 1 0 13728 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4041
timestamp 1666464484
transform 1 0 13728 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4042
timestamp 1666464484
transform 1 0 13728 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4043
timestamp 1666464484
transform 1 0 13728 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4044
timestamp 1666464484
transform 1 0 13728 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4045
timestamp 1666464484
transform 1 0 13728 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4046
timestamp 1666464484
transform 1 0 13728 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4047
timestamp 1666464484
transform 1 0 13728 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4048
timestamp 1666464484
transform 1 0 13728 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4049
timestamp 1666464484
transform -1 0 12480 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4050
timestamp 1666464484
transform -1 0 12480 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4051
timestamp 1666464484
transform -1 0 12480 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4052
timestamp 1666464484
transform -1 0 12480 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4053
timestamp 1666464484
transform 1 0 12480 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4054
timestamp 1666464484
transform 1 0 12480 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4055
timestamp 1666464484
transform 1 0 12480 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4056
timestamp 1666464484
transform 1 0 12480 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4057
timestamp 1666464484
transform 1 0 12480 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4058
timestamp 1666464484
transform 1 0 12480 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4059
timestamp 1666464484
transform 1 0 12480 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4060
timestamp 1666464484
transform 1 0 12480 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4061
timestamp 1666464484
transform 1 0 12480 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4062
timestamp 1666464484
transform 1 0 12480 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4063
timestamp 1666464484
transform -1 0 13728 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4064
timestamp 1666464484
transform -1 0 11232 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4065
timestamp 1666464484
transform -1 0 11232 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4066
timestamp 1666464484
transform -1 0 11232 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4067
timestamp 1666464484
transform -1 0 11232 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4068
timestamp 1666464484
transform -1 0 11232 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4069
timestamp 1666464484
transform -1 0 11232 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4070
timestamp 1666464484
transform -1 0 11232 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4071
timestamp 1666464484
transform -1 0 11232 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4072
timestamp 1666464484
transform -1 0 11232 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4073
timestamp 1666464484
transform -1 0 13728 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4074
timestamp 1666464484
transform 1 0 12480 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4075
timestamp 1666464484
transform 1 0 12480 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4076
timestamp 1666464484
transform 1 0 12480 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4077
timestamp 1666464484
transform 1 0 12480 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4078
timestamp 1666464484
transform 1 0 12480 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4079
timestamp 1666464484
transform -1 0 11232 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4080
timestamp 1666464484
transform -1 0 11232 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4081
timestamp 1666464484
transform 1 0 13728 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4082
timestamp 1666464484
transform 1 0 13728 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4083
timestamp 1666464484
transform 1 0 13728 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4084
timestamp 1666464484
transform 1 0 13728 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4085
timestamp 1666464484
transform 1 0 13728 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4086
timestamp 1666464484
transform 1 0 13728 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4087
timestamp 1666464484
transform 1 0 13728 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4088
timestamp 1666464484
transform 1 0 13728 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4089
timestamp 1666464484
transform 1 0 13728 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4090
timestamp 1666464484
transform -1 0 11232 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4091
timestamp 1666464484
transform -1 0 11232 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4092
timestamp 1666464484
transform 1 0 11232 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4093
timestamp 1666464484
transform 1 0 11232 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4094
timestamp 1666464484
transform 1 0 11232 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4095
timestamp 1666464484
transform 1 0 11232 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4096
timestamp 1666464484
transform -1 0 11232 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4097
timestamp 1666464484
transform -1 0 11232 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4098
timestamp 1666464484
transform -1 0 11232 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4099
timestamp 1666464484
transform -1 0 11232 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4100
timestamp 1666464484
transform -1 0 13728 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4101
timestamp 1666464484
transform -1 0 13728 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4102
timestamp 1666464484
transform -1 0 13728 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4103
timestamp 1666464484
transform -1 0 13728 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4104
timestamp 1666464484
transform -1 0 11232 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4105
timestamp 1666464484
transform -1 0 11232 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4106
timestamp 1666464484
transform -1 0 11232 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4107
timestamp 1666464484
transform -1 0 11232 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4108
timestamp 1666464484
transform -1 0 11232 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4109
timestamp 1666464484
transform -1 0 11232 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4110
timestamp 1666464484
transform 1 0 12480 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4111
timestamp 1666464484
transform 1 0 12480 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4112
timestamp 1666464484
transform 1 0 12480 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4113
timestamp 1666464484
transform 1 0 12480 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4114
timestamp 1666464484
transform -1 0 12480 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4115
timestamp 1666464484
transform -1 0 12480 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4116
timestamp 1666464484
transform -1 0 12480 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4117
timestamp 1666464484
transform -1 0 12480 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4118
timestamp 1666464484
transform -1 0 12480 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4119
timestamp 1666464484
transform -1 0 12480 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4120
timestamp 1666464484
transform -1 0 12480 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4121
timestamp 1666464484
transform -1 0 12480 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4122
timestamp 1666464484
transform -1 0 12480 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4123
timestamp 1666464484
transform -1 0 12480 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4124
timestamp 1666464484
transform -1 0 12480 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4125
timestamp 1666464484
transform -1 0 12480 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4126
timestamp 1666464484
transform -1 0 12480 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4127
timestamp 1666464484
transform -1 0 12480 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4128
timestamp 1666464484
transform 1 0 12480 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4129
timestamp 1666464484
transform 1 0 12480 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4130
timestamp 1666464484
transform -1 0 13728 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4131
timestamp 1666464484
transform -1 0 13728 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4132
timestamp 1666464484
transform -1 0 13728 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4133
timestamp 1666464484
transform -1 0 13728 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4134
timestamp 1666464484
transform 1 0 11232 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4135
timestamp 1666464484
transform 1 0 11232 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4136
timestamp 1666464484
transform 1 0 11232 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4137
timestamp 1666464484
transform 1 0 11232 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4138
timestamp 1666464484
transform 1 0 11232 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4139
timestamp 1666464484
transform 1 0 11232 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4140
timestamp 1666464484
transform 1 0 11232 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4141
timestamp 1666464484
transform 1 0 11232 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4142
timestamp 1666464484
transform 1 0 11232 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4143
timestamp 1666464484
transform 1 0 11232 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4144
timestamp 1666464484
transform 1 0 13728 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4145
timestamp 1666464484
transform 1 0 13728 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4146
timestamp 1666464484
transform 1 0 13728 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4147
timestamp 1666464484
transform 1 0 13728 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4148
timestamp 1666464484
transform 1 0 13728 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4149
timestamp 1666464484
transform -1 0 13728 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4150
timestamp 1666464484
transform -1 0 13728 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4151
timestamp 1666464484
transform -1 0 13728 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4152
timestamp 1666464484
transform -1 0 13728 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4153
timestamp 1666464484
transform -1 0 13728 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4154
timestamp 1666464484
transform -1 0 13728 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4155
timestamp 1666464484
transform 1 0 12480 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4156
timestamp 1666464484
transform 1 0 12480 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4157
timestamp 1666464484
transform 1 0 12480 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4158
timestamp 1666464484
transform -1 0 18720 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4159
timestamp 1666464484
transform -1 0 18720 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4160
timestamp 1666464484
transform -1 0 18720 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4161
timestamp 1666464484
transform -1 0 18720 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4162
timestamp 1666464484
transform -1 0 18720 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4163
timestamp 1666464484
transform -1 0 18720 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4164
timestamp 1666464484
transform -1 0 18720 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4165
timestamp 1666464484
transform -1 0 18720 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4166
timestamp 1666464484
transform -1 0 18720 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4167
timestamp 1666464484
transform -1 0 18720 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4168
timestamp 1666464484
transform 1 0 16224 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4169
timestamp 1666464484
transform 1 0 16224 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4170
timestamp 1666464484
transform 1 0 16224 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4171
timestamp 1666464484
transform 1 0 16224 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4172
timestamp 1666464484
transform 1 0 16224 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4173
timestamp 1666464484
transform 1 0 16224 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4174
timestamp 1666464484
transform 1 0 16224 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4175
timestamp 1666464484
transform 1 0 16224 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4176
timestamp 1666464484
transform 1 0 16224 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4177
timestamp 1666464484
transform 1 0 16224 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4178
timestamp 1666464484
transform -1 0 18720 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4179
timestamp 1666464484
transform -1 0 18720 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4180
timestamp 1666464484
transform 1 0 18720 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4181
timestamp 1666464484
transform 1 0 18720 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4182
timestamp 1666464484
transform -1 0 16224 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4183
timestamp 1666464484
transform -1 0 16224 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4184
timestamp 1666464484
transform -1 0 16224 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4185
timestamp 1666464484
transform -1 0 16224 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4186
timestamp 1666464484
transform -1 0 16224 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4187
timestamp 1666464484
transform -1 0 16224 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4188
timestamp 1666464484
transform -1 0 16224 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4189
timestamp 1666464484
transform -1 0 16224 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4190
timestamp 1666464484
transform -1 0 16224 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4191
timestamp 1666464484
transform -1 0 16224 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4192
timestamp 1666464484
transform -1 0 16224 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4193
timestamp 1666464484
transform -1 0 16224 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4194
timestamp 1666464484
transform -1 0 16224 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4195
timestamp 1666464484
transform -1 0 16224 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4196
timestamp 1666464484
transform 1 0 18720 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4197
timestamp 1666464484
transform 1 0 18720 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4198
timestamp 1666464484
transform 1 0 18720 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4199
timestamp 1666464484
transform 1 0 18720 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4200
timestamp 1666464484
transform 1 0 18720 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4201
timestamp 1666464484
transform 1 0 17472 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4202
timestamp 1666464484
transform 1 0 17472 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4203
timestamp 1666464484
transform 1 0 17472 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4204
timestamp 1666464484
transform 1 0 17472 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4205
timestamp 1666464484
transform 1 0 17472 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4206
timestamp 1666464484
transform 1 0 17472 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4207
timestamp 1666464484
transform 1 0 17472 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4208
timestamp 1666464484
transform 1 0 17472 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4209
timestamp 1666464484
transform 1 0 17472 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4210
timestamp 1666464484
transform 1 0 17472 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4211
timestamp 1666464484
transform 1 0 17472 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4212
timestamp 1666464484
transform 1 0 17472 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4213
timestamp 1666464484
transform 1 0 17472 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4214
timestamp 1666464484
transform 1 0 17472 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4215
timestamp 1666464484
transform 1 0 18720 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4216
timestamp 1666464484
transform 1 0 18720 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4217
timestamp 1666464484
transform 1 0 18720 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4218
timestamp 1666464484
transform -1 0 17472 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4219
timestamp 1666464484
transform -1 0 17472 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4220
timestamp 1666464484
transform -1 0 17472 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4221
timestamp 1666464484
transform -1 0 17472 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4222
timestamp 1666464484
transform -1 0 17472 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4223
timestamp 1666464484
transform -1 0 17472 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4224
timestamp 1666464484
transform -1 0 17472 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4225
timestamp 1666464484
transform -1 0 17472 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4226
timestamp 1666464484
transform -1 0 17472 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4227
timestamp 1666464484
transform -1 0 17472 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4228
timestamp 1666464484
transform -1 0 17472 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4229
timestamp 1666464484
transform -1 0 17472 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4230
timestamp 1666464484
transform -1 0 17472 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4231
timestamp 1666464484
transform -1 0 17472 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4232
timestamp 1666464484
transform 1 0 18720 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4233
timestamp 1666464484
transform 1 0 18720 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4234
timestamp 1666464484
transform 1 0 18720 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4235
timestamp 1666464484
transform 1 0 18720 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4236
timestamp 1666464484
transform -1 0 18720 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4237
timestamp 1666464484
transform -1 0 18720 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4238
timestamp 1666464484
transform 1 0 16224 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4239
timestamp 1666464484
transform 1 0 16224 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4240
timestamp 1666464484
transform 1 0 16224 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4241
timestamp 1666464484
transform 1 0 16224 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4242
timestamp 1666464484
transform -1 0 18720 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4243
timestamp 1666464484
transform -1 0 18720 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4244
timestamp 1666464484
transform -1 0 14976 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4245
timestamp 1666464484
transform -1 0 14976 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4246
timestamp 1666464484
transform -1 0 14976 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4247
timestamp 1666464484
transform -1 0 14976 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4248
timestamp 1666464484
transform -1 0 14976 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4249
timestamp 1666464484
transform -1 0 14976 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4250
timestamp 1666464484
transform -1 0 14976 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4251
timestamp 1666464484
transform -1 0 14976 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4252
timestamp 1666464484
transform -1 0 14976 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4253
timestamp 1666464484
transform -1 0 14976 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4254
timestamp 1666464484
transform -1 0 14976 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4255
timestamp 1666464484
transform -1 0 14976 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4256
timestamp 1666464484
transform -1 0 14976 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4257
timestamp 1666464484
transform -1 0 14976 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4258
timestamp 1666464484
transform -1 0 14976 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4259
timestamp 1666464484
transform -1 0 14976 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4260
timestamp 1666464484
transform -1 0 14976 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4261
timestamp 1666464484
transform -1 0 14976 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4262
timestamp 1666464484
transform -1 0 14976 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4263
timestamp 1666464484
transform -1 0 14976 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4264
timestamp 1666464484
transform -1 0 14976 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4265
timestamp 1666464484
transform -1 0 14976 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4266
timestamp 1666464484
transform -1 0 14976 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4267
timestamp 1666464484
transform -1 0 14976 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4268
timestamp 1666464484
transform -1 0 14976 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4269
timestamp 1666464484
transform -1 0 14976 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4270
timestamp 1666464484
transform -1 0 14976 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4271
timestamp 1666464484
transform -1 0 14976 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4272
timestamp 1666464484
transform -1 0 14976 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4273
timestamp 1666464484
transform -1 0 14976 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4274
timestamp 1666464484
transform 1 0 12480 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4275
timestamp 1666464484
transform 1 0 17472 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4276
timestamp 1666464484
transform 1 0 17472 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4277
timestamp 1666464484
transform -1 0 11232 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4278
timestamp 1666464484
transform -1 0 17472 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4279
timestamp 1666464484
transform -1 0 17472 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4280
timestamp 1666464484
transform 1 0 13728 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4281
timestamp 1666464484
transform 1 0 13728 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4282
timestamp 1666464484
transform 1 0 11232 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4283
timestamp 1666464484
transform 1 0 11232 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4284
timestamp 1666464484
transform 1 0 16224 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4285
timestamp 1666464484
transform 1 0 16224 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4286
timestamp 1666464484
transform -1 0 12480 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4287
timestamp 1666464484
transform -1 0 12480 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4288
timestamp 1666464484
transform -1 0 16224 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4289
timestamp 1666464484
transform -1 0 16224 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4290
timestamp 1666464484
transform -1 0 13728 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4291
timestamp 1666464484
transform -1 0 13728 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4292
timestamp 1666464484
transform 1 0 14976 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4293
timestamp 1666464484
transform 1 0 14976 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4294
timestamp 1666464484
transform 1 0 14976 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4295
timestamp 1666464484
transform 1 0 14976 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4296
timestamp 1666464484
transform 1 0 14976 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4297
timestamp 1666464484
transform 1 0 14976 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4298
timestamp 1666464484
transform 1 0 14976 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4299
timestamp 1666464484
transform 1 0 14976 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4300
timestamp 1666464484
transform 1 0 14976 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4301
timestamp 1666464484
transform 1 0 14976 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4302
timestamp 1666464484
transform 1 0 14976 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4303
timestamp 1666464484
transform 1 0 14976 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4304
timestamp 1666464484
transform 1 0 14976 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4305
timestamp 1666464484
transform 1 0 14976 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4306
timestamp 1666464484
transform 1 0 14976 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4307
timestamp 1666464484
transform 1 0 14976 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4308
timestamp 1666464484
transform 1 0 14976 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4309
timestamp 1666464484
transform 1 0 14976 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4310
timestamp 1666464484
transform 1 0 14976 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4311
timestamp 1666464484
transform 1 0 14976 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4312
timestamp 1666464484
transform 1 0 14976 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4313
timestamp 1666464484
transform 1 0 14976 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4314
timestamp 1666464484
transform 1 0 14976 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4315
timestamp 1666464484
transform 1 0 14976 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4316
timestamp 1666464484
transform 1 0 14976 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4317
timestamp 1666464484
transform 1 0 14976 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4318
timestamp 1666464484
transform 1 0 14976 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4319
timestamp 1666464484
transform 1 0 14976 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4320
timestamp 1666464484
transform 1 0 14976 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4321
timestamp 1666464484
transform 1 0 14976 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4322
timestamp 1666464484
transform 1 0 18720 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4323
timestamp 1666464484
transform 1 0 18720 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4324
timestamp 1666464484
transform -1 0 11232 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4325
timestamp 1666464484
transform 1 0 12480 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4326
timestamp 1666464484
transform 1 0 6240 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4327
timestamp 1666464484
transform 1 0 6240 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4328
timestamp 1666464484
transform 1 0 6240 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4329
timestamp 1666464484
transform 1 0 8736 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4330
timestamp 1666464484
transform 1 0 8736 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4331
timestamp 1666464484
transform 1 0 8736 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4332
timestamp 1666464484
transform 1 0 8736 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4333
timestamp 1666464484
transform 1 0 8736 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4334
timestamp 1666464484
transform 1 0 8736 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4335
timestamp 1666464484
transform 1 0 8736 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4336
timestamp 1666464484
transform 1 0 8736 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4337
timestamp 1666464484
transform 1 0 8736 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4338
timestamp 1666464484
transform 1 0 8736 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4339
timestamp 1666464484
transform 1 0 8736 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4340
timestamp 1666464484
transform 1 0 8736 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4341
timestamp 1666464484
transform 1 0 8736 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4342
timestamp 1666464484
transform 1 0 8736 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4343
timestamp 1666464484
transform 1 0 6240 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4344
timestamp 1666464484
transform 1 0 6240 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4345
timestamp 1666464484
transform 1 0 6240 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4346
timestamp 1666464484
transform 1 0 6240 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4347
timestamp 1666464484
transform 1 0 6240 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4348
timestamp 1666464484
transform -1 0 8736 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4349
timestamp 1666464484
transform -1 0 7488 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4350
timestamp 1666464484
transform -1 0 7488 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4351
timestamp 1666464484
transform -1 0 7488 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4352
timestamp 1666464484
transform -1 0 7488 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4353
timestamp 1666464484
transform -1 0 7488 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4354
timestamp 1666464484
transform -1 0 7488 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4355
timestamp 1666464484
transform -1 0 7488 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4356
timestamp 1666464484
transform -1 0 7488 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4357
timestamp 1666464484
transform -1 0 7488 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4358
timestamp 1666464484
transform 1 0 7488 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4359
timestamp 1666464484
transform 1 0 7488 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4360
timestamp 1666464484
transform 1 0 7488 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4361
timestamp 1666464484
transform 1 0 7488 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4362
timestamp 1666464484
transform 1 0 7488 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4363
timestamp 1666464484
transform 1 0 7488 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4364
timestamp 1666464484
transform 1 0 7488 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4365
timestamp 1666464484
transform -1 0 6240 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4366
timestamp 1666464484
transform -1 0 6240 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4367
timestamp 1666464484
transform -1 0 6240 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4368
timestamp 1666464484
transform -1 0 6240 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4369
timestamp 1666464484
transform -1 0 6240 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4370
timestamp 1666464484
transform -1 0 6240 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4371
timestamp 1666464484
transform -1 0 6240 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4372
timestamp 1666464484
transform -1 0 6240 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4373
timestamp 1666464484
transform -1 0 6240 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4374
timestamp 1666464484
transform -1 0 6240 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4375
timestamp 1666464484
transform -1 0 6240 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4376
timestamp 1666464484
transform -1 0 6240 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4377
timestamp 1666464484
transform -1 0 6240 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4378
timestamp 1666464484
transform 1 0 7488 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4379
timestamp 1666464484
transform 1 0 7488 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4380
timestamp 1666464484
transform 1 0 7488 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4381
timestamp 1666464484
transform -1 0 8736 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4382
timestamp 1666464484
transform -1 0 8736 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4383
timestamp 1666464484
transform -1 0 8736 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4384
timestamp 1666464484
transform -1 0 8736 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4385
timestamp 1666464484
transform -1 0 8736 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4386
timestamp 1666464484
transform -1 0 8736 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4387
timestamp 1666464484
transform -1 0 8736 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4388
timestamp 1666464484
transform -1 0 8736 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4389
timestamp 1666464484
transform -1 0 8736 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4390
timestamp 1666464484
transform -1 0 8736 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4391
timestamp 1666464484
transform -1 0 8736 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4392
timestamp 1666464484
transform -1 0 8736 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4393
timestamp 1666464484
transform -1 0 8736 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4394
timestamp 1666464484
transform 1 0 7488 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4395
timestamp 1666464484
transform 1 0 7488 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4396
timestamp 1666464484
transform -1 0 7488 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4397
timestamp 1666464484
transform -1 0 7488 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4398
timestamp 1666464484
transform -1 0 6240 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4399
timestamp 1666464484
transform -1 0 7488 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4400
timestamp 1666464484
transform -1 0 7488 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4401
timestamp 1666464484
transform -1 0 7488 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4402
timestamp 1666464484
transform 1 0 6240 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4403
timestamp 1666464484
transform 1 0 6240 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4404
timestamp 1666464484
transform 1 0 6240 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4405
timestamp 1666464484
transform 1 0 6240 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4406
timestamp 1666464484
transform 1 0 6240 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4407
timestamp 1666464484
transform 1 0 7488 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4408
timestamp 1666464484
transform 1 0 7488 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4409
timestamp 1666464484
transform 1 0 6240 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4410
timestamp 1666464484
transform 1 0 3744 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4411
timestamp 1666464484
transform 1 0 3744 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4412
timestamp 1666464484
transform 1 0 3744 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4413
timestamp 1666464484
transform 1 0 3744 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4414
timestamp 1666464484
transform 1 0 3744 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4415
timestamp 1666464484
transform 1 0 3744 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4416
timestamp 1666464484
transform 1 0 2496 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4417
timestamp 1666464484
transform 1 0 2496 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4418
timestamp 1666464484
transform 1 0 2496 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4419
timestamp 1666464484
transform 1 0 2496 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4420
timestamp 1666464484
transform 1 0 2496 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4421
timestamp 1666464484
transform 1 0 2496 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4422
timestamp 1666464484
transform 1 0 0 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4423
timestamp 1666464484
transform 1 0 0 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4424
timestamp 1666464484
transform 1 0 1248 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4425
timestamp 1666464484
transform 1 0 1248 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4426
timestamp 1666464484
transform 1 0 1248 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4427
timestamp 1666464484
transform 1 0 1248 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4428
timestamp 1666464484
transform 1 0 1248 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4429
timestamp 1666464484
transform 1 0 1248 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4430
timestamp 1666464484
transform 1 0 0 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4431
timestamp 1666464484
transform 1 0 0 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4432
timestamp 1666464484
transform 1 0 0 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4433
timestamp 1666464484
transform 1 0 0 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4434
timestamp 1666464484
transform -1 0 1248 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4435
timestamp 1666464484
transform -1 0 1248 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4436
timestamp 1666464484
transform -1 0 1248 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4437
timestamp 1666464484
transform -1 0 1248 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4438
timestamp 1666464484
transform -1 0 1248 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4439
timestamp 1666464484
transform -1 0 1248 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4440
timestamp 1666464484
transform -1 0 1248 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4441
timestamp 1666464484
transform -1 0 1248 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4442
timestamp 1666464484
transform -1 0 1248 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4443
timestamp 1666464484
transform -1 0 1248 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4444
timestamp 1666464484
transform -1 0 1248 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4445
timestamp 1666464484
transform -1 0 1248 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4446
timestamp 1666464484
transform -1 0 1248 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4447
timestamp 1666464484
transform -1 0 1248 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4448
timestamp 1666464484
transform -1 0 3744 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4449
timestamp 1666464484
transform -1 0 3744 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4450
timestamp 1666464484
transform -1 0 3744 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4451
timestamp 1666464484
transform -1 0 3744 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4452
timestamp 1666464484
transform -1 0 3744 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4453
timestamp 1666464484
transform -1 0 3744 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4454
timestamp 1666464484
transform -1 0 3744 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4455
timestamp 1666464484
transform -1 0 3744 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4456
timestamp 1666464484
transform -1 0 3744 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4457
timestamp 1666464484
transform -1 0 3744 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4458
timestamp 1666464484
transform -1 0 3744 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4459
timestamp 1666464484
transform -1 0 3744 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4460
timestamp 1666464484
transform -1 0 3744 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4461
timestamp 1666464484
transform -1 0 3744 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4462
timestamp 1666464484
transform 1 0 0 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4463
timestamp 1666464484
transform 1 0 0 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4464
timestamp 1666464484
transform 1 0 0 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4465
timestamp 1666464484
transform 1 0 0 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4466
timestamp 1666464484
transform 1 0 3744 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4467
timestamp 1666464484
transform 1 0 3744 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4468
timestamp 1666464484
transform 1 0 3744 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4469
timestamp 1666464484
transform 1 0 3744 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4470
timestamp 1666464484
transform 1 0 0 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4471
timestamp 1666464484
transform 1 0 3744 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4472
timestamp 1666464484
transform 1 0 3744 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4473
timestamp 1666464484
transform 1 0 3744 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4474
timestamp 1666464484
transform 1 0 1248 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4475
timestamp 1666464484
transform 1 0 1248 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4476
timestamp 1666464484
transform 1 0 1248 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4477
timestamp 1666464484
transform 1 0 1248 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4478
timestamp 1666464484
transform -1 0 2496 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4479
timestamp 1666464484
transform -1 0 2496 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4480
timestamp 1666464484
transform -1 0 2496 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4481
timestamp 1666464484
transform -1 0 2496 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4482
timestamp 1666464484
transform -1 0 2496 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4483
timestamp 1666464484
transform -1 0 2496 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4484
timestamp 1666464484
transform -1 0 2496 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4485
timestamp 1666464484
transform -1 0 2496 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4486
timestamp 1666464484
transform -1 0 2496 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4487
timestamp 1666464484
transform -1 0 2496 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4488
timestamp 1666464484
transform -1 0 2496 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4489
timestamp 1666464484
transform -1 0 2496 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4490
timestamp 1666464484
transform -1 0 2496 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4491
timestamp 1666464484
transform -1 0 2496 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4492
timestamp 1666464484
transform 1 0 0 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4493
timestamp 1666464484
transform 1 0 0 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4494
timestamp 1666464484
transform 1 0 1248 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4495
timestamp 1666464484
transform 1 0 1248 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4496
timestamp 1666464484
transform 1 0 1248 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4497
timestamp 1666464484
transform 1 0 1248 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4498
timestamp 1666464484
transform 1 0 3744 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4499
timestamp 1666464484
transform 1 0 0 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4500
timestamp 1666464484
transform 1 0 2496 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4501
timestamp 1666464484
transform 1 0 2496 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4502
timestamp 1666464484
transform 1 0 2496 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4503
timestamp 1666464484
transform 1 0 2496 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4504
timestamp 1666464484
transform 1 0 2496 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4505
timestamp 1666464484
transform 1 0 2496 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4506
timestamp 1666464484
transform 1 0 2496 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4507
timestamp 1666464484
transform 1 0 2496 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4508
timestamp 1666464484
transform 1 0 0 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4509
timestamp 1666464484
transform 1 0 0 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4510
timestamp 1666464484
transform 1 0 0 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4511
timestamp 1666464484
transform 1 0 0 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4512
timestamp 1666464484
transform 1 0 0 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4513
timestamp 1666464484
transform 1 0 3744 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4514
timestamp 1666464484
transform 1 0 0 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4515
timestamp 1666464484
transform 1 0 0 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4516
timestamp 1666464484
transform 1 0 0 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4517
timestamp 1666464484
transform 1 0 0 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4518
timestamp 1666464484
transform 1 0 3744 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4519
timestamp 1666464484
transform 1 0 3744 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4520
timestamp 1666464484
transform 1 0 3744 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4521
timestamp 1666464484
transform 1 0 3744 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4522
timestamp 1666464484
transform -1 0 1248 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4523
timestamp 1666464484
transform -1 0 1248 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4524
timestamp 1666464484
transform -1 0 3744 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4525
timestamp 1666464484
transform -1 0 3744 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4526
timestamp 1666464484
transform -1 0 3744 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4527
timestamp 1666464484
transform -1 0 3744 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4528
timestamp 1666464484
transform -1 0 3744 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4529
timestamp 1666464484
transform -1 0 3744 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4530
timestamp 1666464484
transform -1 0 3744 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4531
timestamp 1666464484
transform -1 0 3744 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4532
timestamp 1666464484
transform -1 0 3744 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4533
timestamp 1666464484
transform -1 0 3744 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4534
timestamp 1666464484
transform -1 0 3744 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4535
timestamp 1666464484
transform -1 0 3744 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4536
timestamp 1666464484
transform -1 0 3744 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4537
timestamp 1666464484
transform -1 0 3744 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4538
timestamp 1666464484
transform -1 0 1248 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4539
timestamp 1666464484
transform -1 0 1248 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4540
timestamp 1666464484
transform 1 0 0 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4541
timestamp 1666464484
transform 1 0 0 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4542
timestamp 1666464484
transform 1 0 1248 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4543
timestamp 1666464484
transform 1 0 1248 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4544
timestamp 1666464484
transform 1 0 1248 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4545
timestamp 1666464484
transform 1 0 1248 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4546
timestamp 1666464484
transform 1 0 1248 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4547
timestamp 1666464484
transform 1 0 1248 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4548
timestamp 1666464484
transform 1 0 1248 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4549
timestamp 1666464484
transform 1 0 1248 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4550
timestamp 1666464484
transform 1 0 1248 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4551
timestamp 1666464484
transform 1 0 1248 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4552
timestamp 1666464484
transform 1 0 1248 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4553
timestamp 1666464484
transform 1 0 1248 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4554
timestamp 1666464484
transform 1 0 1248 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4555
timestamp 1666464484
transform 1 0 1248 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4556
timestamp 1666464484
transform 1 0 2496 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4557
timestamp 1666464484
transform 1 0 2496 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4558
timestamp 1666464484
transform 1 0 2496 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4559
timestamp 1666464484
transform 1 0 2496 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4560
timestamp 1666464484
transform 1 0 2496 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4561
timestamp 1666464484
transform 1 0 2496 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4562
timestamp 1666464484
transform 1 0 2496 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4563
timestamp 1666464484
transform 1 0 2496 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4564
timestamp 1666464484
transform 1 0 2496 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4565
timestamp 1666464484
transform 1 0 2496 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4566
timestamp 1666464484
transform 1 0 2496 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4567
timestamp 1666464484
transform 1 0 2496 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4568
timestamp 1666464484
transform 1 0 2496 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4569
timestamp 1666464484
transform 1 0 2496 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4570
timestamp 1666464484
transform -1 0 1248 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4571
timestamp 1666464484
transform -1 0 1248 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4572
timestamp 1666464484
transform -1 0 1248 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4573
timestamp 1666464484
transform -1 0 1248 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4574
timestamp 1666464484
transform -1 0 1248 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4575
timestamp 1666464484
transform -1 0 1248 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4576
timestamp 1666464484
transform -1 0 1248 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4577
timestamp 1666464484
transform -1 0 1248 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4578
timestamp 1666464484
transform -1 0 1248 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4579
timestamp 1666464484
transform -1 0 1248 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4580
timestamp 1666464484
transform 1 0 3744 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4581
timestamp 1666464484
transform 1 0 3744 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4582
timestamp 1666464484
transform 1 0 0 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4583
timestamp 1666464484
transform 1 0 0 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4584
timestamp 1666464484
transform 1 0 3744 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4585
timestamp 1666464484
transform 1 0 3744 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4586
timestamp 1666464484
transform 1 0 3744 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4587
timestamp 1666464484
transform 1 0 3744 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4588
timestamp 1666464484
transform 1 0 3744 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4589
timestamp 1666464484
transform 1 0 3744 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4590
timestamp 1666464484
transform -1 0 2496 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4591
timestamp 1666464484
transform -1 0 2496 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4592
timestamp 1666464484
transform -1 0 2496 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4593
timestamp 1666464484
transform -1 0 2496 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4594
timestamp 1666464484
transform -1 0 2496 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4595
timestamp 1666464484
transform -1 0 2496 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4596
timestamp 1666464484
transform -1 0 2496 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4597
timestamp 1666464484
transform -1 0 2496 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4598
timestamp 1666464484
transform -1 0 2496 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4599
timestamp 1666464484
transform -1 0 2496 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4600
timestamp 1666464484
transform -1 0 2496 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4601
timestamp 1666464484
transform -1 0 2496 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4602
timestamp 1666464484
transform -1 0 2496 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4603
timestamp 1666464484
transform -1 0 2496 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4604
timestamp 1666464484
transform 1 0 3744 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4605
timestamp 1666464484
transform 1 0 0 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4606
timestamp 1666464484
transform -1 0 8736 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4607
timestamp 1666464484
transform -1 0 8736 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4608
timestamp 1666464484
transform -1 0 8736 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4609
timestamp 1666464484
transform -1 0 8736 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4610
timestamp 1666464484
transform -1 0 8736 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4611
timestamp 1666464484
transform -1 0 8736 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4612
timestamp 1666464484
transform -1 0 8736 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4613
timestamp 1666464484
transform -1 0 8736 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4614
timestamp 1666464484
transform -1 0 8736 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4615
timestamp 1666464484
transform -1 0 8736 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4616
timestamp 1666464484
transform -1 0 8736 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4617
timestamp 1666464484
transform -1 0 8736 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4618
timestamp 1666464484
transform -1 0 8736 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4619
timestamp 1666464484
transform -1 0 8736 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4620
timestamp 1666464484
transform -1 0 7488 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4621
timestamp 1666464484
transform -1 0 7488 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4622
timestamp 1666464484
transform -1 0 7488 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4623
timestamp 1666464484
transform -1 0 7488 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4624
timestamp 1666464484
transform -1 0 6240 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4625
timestamp 1666464484
transform -1 0 6240 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4626
timestamp 1666464484
transform -1 0 6240 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4627
timestamp 1666464484
transform -1 0 6240 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4628
timestamp 1666464484
transform -1 0 6240 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4629
timestamp 1666464484
transform -1 0 6240 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4630
timestamp 1666464484
transform -1 0 6240 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4631
timestamp 1666464484
transform -1 0 6240 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4632
timestamp 1666464484
transform -1 0 6240 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4633
timestamp 1666464484
transform -1 0 6240 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4634
timestamp 1666464484
transform -1 0 6240 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4635
timestamp 1666464484
transform -1 0 6240 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4636
timestamp 1666464484
transform -1 0 6240 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4637
timestamp 1666464484
transform -1 0 6240 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4638
timestamp 1666464484
transform -1 0 7488 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4639
timestamp 1666464484
transform -1 0 7488 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4640
timestamp 1666464484
transform -1 0 7488 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4641
timestamp 1666464484
transform -1 0 7488 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4642
timestamp 1666464484
transform 1 0 7488 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4643
timestamp 1666464484
transform 1 0 7488 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4644
timestamp 1666464484
transform 1 0 7488 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4645
timestamp 1666464484
transform 1 0 7488 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4646
timestamp 1666464484
transform 1 0 7488 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4647
timestamp 1666464484
transform 1 0 7488 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4648
timestamp 1666464484
transform 1 0 7488 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4649
timestamp 1666464484
transform 1 0 7488 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4650
timestamp 1666464484
transform 1 0 7488 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4651
timestamp 1666464484
transform 1 0 7488 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4652
timestamp 1666464484
transform 1 0 7488 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4653
timestamp 1666464484
transform 1 0 7488 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4654
timestamp 1666464484
transform 1 0 7488 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4655
timestamp 1666464484
transform 1 0 7488 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4656
timestamp 1666464484
transform -1 0 7488 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4657
timestamp 1666464484
transform -1 0 7488 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4658
timestamp 1666464484
transform -1 0 7488 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4659
timestamp 1666464484
transform -1 0 7488 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4660
timestamp 1666464484
transform -1 0 7488 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4661
timestamp 1666464484
transform -1 0 7488 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4662
timestamp 1666464484
transform 1 0 8736 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4663
timestamp 1666464484
transform 1 0 8736 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4664
timestamp 1666464484
transform 1 0 8736 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4665
timestamp 1666464484
transform 1 0 8736 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4666
timestamp 1666464484
transform 1 0 8736 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4667
timestamp 1666464484
transform 1 0 8736 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4668
timestamp 1666464484
transform 1 0 8736 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4669
timestamp 1666464484
transform 1 0 8736 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4670
timestamp 1666464484
transform 1 0 6240 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4671
timestamp 1666464484
transform 1 0 6240 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4672
timestamp 1666464484
transform 1 0 6240 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4673
timestamp 1666464484
transform 1 0 6240 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4674
timestamp 1666464484
transform 1 0 6240 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4675
timestamp 1666464484
transform 1 0 6240 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4676
timestamp 1666464484
transform 1 0 6240 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4677
timestamp 1666464484
transform 1 0 6240 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4678
timestamp 1666464484
transform 1 0 6240 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4679
timestamp 1666464484
transform 1 0 6240 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4680
timestamp 1666464484
transform 1 0 6240 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4681
timestamp 1666464484
transform 1 0 6240 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4682
timestamp 1666464484
transform 1 0 6240 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4683
timestamp 1666464484
transform 1 0 6240 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4684
timestamp 1666464484
transform 1 0 8736 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4685
timestamp 1666464484
transform 1 0 8736 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4686
timestamp 1666464484
transform 1 0 8736 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4687
timestamp 1666464484
transform 1 0 8736 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4688
timestamp 1666464484
transform 1 0 8736 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4689
timestamp 1666464484
transform 1 0 8736 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4690
timestamp 1666464484
transform -1 0 8736 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4691
timestamp 1666464484
transform -1 0 8736 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4692
timestamp 1666464484
transform -1 0 3744 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4693
timestamp 1666464484
transform -1 0 3744 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4694
timestamp 1666464484
transform 1 0 2496 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4695
timestamp 1666464484
transform 1 0 2496 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4696
timestamp 1666464484
transform -1 0 6240 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4697
timestamp 1666464484
transform -1 0 6240 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4698
timestamp 1666464484
transform 1 0 7488 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4699
timestamp 1666464484
transform 1 0 7488 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4700
timestamp 1666464484
transform -1 0 2496 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4701
timestamp 1666464484
transform -1 0 2496 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4702
timestamp 1666464484
transform -1 0 4992 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4703
timestamp 1666464484
transform -1 0 4992 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4704
timestamp 1666464484
transform -1 0 4992 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4705
timestamp 1666464484
transform -1 0 4992 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4706
timestamp 1666464484
transform -1 0 4992 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4707
timestamp 1666464484
transform -1 0 4992 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4708
timestamp 1666464484
transform -1 0 4992 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4709
timestamp 1666464484
transform -1 0 4992 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4710
timestamp 1666464484
transform -1 0 4992 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4711
timestamp 1666464484
transform -1 0 4992 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4712
timestamp 1666464484
transform -1 0 4992 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4713
timestamp 1666464484
transform -1 0 4992 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4714
timestamp 1666464484
transform -1 0 4992 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4715
timestamp 1666464484
transform -1 0 4992 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4716
timestamp 1666464484
transform 1 0 1248 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4717
timestamp 1666464484
transform 1 0 1248 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4718
timestamp 1666464484
transform -1 0 4992 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4719
timestamp 1666464484
transform -1 0 4992 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4720
timestamp 1666464484
transform -1 0 4992 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4721
timestamp 1666464484
transform -1 0 4992 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4722
timestamp 1666464484
transform -1 0 4992 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4723
timestamp 1666464484
transform -1 0 4992 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4724
timestamp 1666464484
transform -1 0 4992 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4725
timestamp 1666464484
transform -1 0 4992 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4726
timestamp 1666464484
transform -1 0 4992 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4727
timestamp 1666464484
transform -1 0 4992 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4728
timestamp 1666464484
transform -1 0 4992 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4729
timestamp 1666464484
transform -1 0 4992 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4730
timestamp 1666464484
transform -1 0 4992 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4731
timestamp 1666464484
transform -1 0 4992 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4732
timestamp 1666464484
transform -1 0 7488 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4733
timestamp 1666464484
transform -1 0 7488 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4734
timestamp 1666464484
transform -1 0 1248 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4735
timestamp 1666464484
transform -1 0 1248 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4736
timestamp 1666464484
transform -1 0 4992 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4737
timestamp 1666464484
transform -1 0 4992 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4738
timestamp 1666464484
transform 1 0 4992 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4739
timestamp 1666464484
transform 1 0 4992 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4740
timestamp 1666464484
transform 1 0 4992 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4741
timestamp 1666464484
transform 1 0 4992 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4742
timestamp 1666464484
transform 1 0 4992 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4743
timestamp 1666464484
transform 1 0 4992 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4744
timestamp 1666464484
transform 1 0 4992 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4745
timestamp 1666464484
transform 1 0 4992 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4746
timestamp 1666464484
transform 1 0 4992 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4747
timestamp 1666464484
transform 1 0 4992 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4748
timestamp 1666464484
transform 1 0 4992 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4749
timestamp 1666464484
transform 1 0 4992 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4750
timestamp 1666464484
transform 1 0 4992 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4751
timestamp 1666464484
transform 1 0 4992 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4752
timestamp 1666464484
transform 1 0 4992 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4753
timestamp 1666464484
transform 1 0 4992 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4754
timestamp 1666464484
transform 1 0 4992 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4755
timestamp 1666464484
transform 1 0 4992 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4756
timestamp 1666464484
transform 1 0 4992 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4757
timestamp 1666464484
transform 1 0 4992 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4758
timestamp 1666464484
transform 1 0 4992 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4759
timestamp 1666464484
transform 1 0 4992 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4760
timestamp 1666464484
transform 1 0 4992 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4761
timestamp 1666464484
transform 1 0 4992 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4762
timestamp 1666464484
transform 1 0 4992 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4763
timestamp 1666464484
transform 1 0 4992 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4764
timestamp 1666464484
transform 1 0 4992 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4765
timestamp 1666464484
transform 1 0 4992 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4766
timestamp 1666464484
transform 1 0 4992 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4767
timestamp 1666464484
transform 1 0 4992 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4768
timestamp 1666464484
transform 1 0 6240 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4769
timestamp 1666464484
transform 1 0 6240 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4770
timestamp 1666464484
transform 1 0 8736 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4771
timestamp 1666464484
transform 1 0 8736 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4772
timestamp 1666464484
transform 1 0 0 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4773
timestamp 1666464484
transform 1 0 0 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4774
timestamp 1666464484
transform 1 0 3744 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4775
timestamp 1666464484
transform 1 0 3744 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4776
timestamp 1666464484
transform 1 0 7488 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4777
timestamp 1666464484
transform 1 0 7488 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4778
timestamp 1666464484
transform 1 0 7488 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4779
timestamp 1666464484
transform 1 0 7488 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4780
timestamp 1666464484
transform 1 0 7488 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4781
timestamp 1666464484
transform 1 0 7488 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4782
timestamp 1666464484
transform 1 0 7488 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4783
timestamp 1666464484
transform 1 0 7488 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4784
timestamp 1666464484
transform 1 0 7488 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4785
timestamp 1666464484
transform 1 0 8736 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4786
timestamp 1666464484
transform 1 0 8736 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4787
timestamp 1666464484
transform 1 0 8736 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4788
timestamp 1666464484
transform 1 0 8736 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4789
timestamp 1666464484
transform 1 0 8736 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4790
timestamp 1666464484
transform 1 0 8736 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4791
timestamp 1666464484
transform 1 0 8736 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4792
timestamp 1666464484
transform 1 0 8736 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4793
timestamp 1666464484
transform 1 0 8736 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4794
timestamp 1666464484
transform 1 0 8736 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4795
timestamp 1666464484
transform 1 0 8736 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4796
timestamp 1666464484
transform 1 0 8736 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4797
timestamp 1666464484
transform 1 0 6240 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4798
timestamp 1666464484
transform 1 0 6240 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4799
timestamp 1666464484
transform 1 0 7488 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4800
timestamp 1666464484
transform 1 0 7488 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4801
timestamp 1666464484
transform 1 0 8736 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4802
timestamp 1666464484
transform 1 0 8736 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4803
timestamp 1666464484
transform 1 0 6240 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4804
timestamp 1666464484
transform 1 0 6240 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4805
timestamp 1666464484
transform 1 0 7488 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4806
timestamp 1666464484
transform 1 0 7488 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4807
timestamp 1666464484
transform -1 0 6240 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4808
timestamp 1666464484
transform -1 0 6240 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4809
timestamp 1666464484
transform 1 0 6240 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4810
timestamp 1666464484
transform 1 0 6240 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4811
timestamp 1666464484
transform -1 0 6240 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4812
timestamp 1666464484
transform -1 0 6240 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4813
timestamp 1666464484
transform -1 0 6240 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4814
timestamp 1666464484
transform -1 0 6240 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4815
timestamp 1666464484
transform -1 0 6240 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4816
timestamp 1666464484
transform -1 0 6240 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4817
timestamp 1666464484
transform -1 0 6240 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4818
timestamp 1666464484
transform -1 0 6240 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4819
timestamp 1666464484
transform -1 0 6240 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4820
timestamp 1666464484
transform -1 0 6240 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4821
timestamp 1666464484
transform 1 0 6240 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4822
timestamp 1666464484
transform -1 0 8736 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4823
timestamp 1666464484
transform -1 0 8736 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4824
timestamp 1666464484
transform -1 0 8736 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4825
timestamp 1666464484
transform -1 0 8736 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4826
timestamp 1666464484
transform -1 0 8736 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4827
timestamp 1666464484
transform -1 0 8736 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4828
timestamp 1666464484
transform -1 0 8736 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4829
timestamp 1666464484
transform -1 0 8736 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4830
timestamp 1666464484
transform -1 0 8736 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4831
timestamp 1666464484
transform -1 0 8736 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4832
timestamp 1666464484
transform -1 0 8736 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4833
timestamp 1666464484
transform -1 0 8736 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4834
timestamp 1666464484
transform 1 0 6240 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4835
timestamp 1666464484
transform 1 0 6240 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4836
timestamp 1666464484
transform 1 0 6240 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4837
timestamp 1666464484
transform 1 0 6240 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4838
timestamp 1666464484
transform -1 0 8736 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4839
timestamp 1666464484
transform -1 0 8736 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4840
timestamp 1666464484
transform -1 0 7488 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4841
timestamp 1666464484
transform -1 0 7488 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4842
timestamp 1666464484
transform -1 0 7488 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4843
timestamp 1666464484
transform -1 0 7488 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4844
timestamp 1666464484
transform -1 0 7488 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4845
timestamp 1666464484
transform -1 0 7488 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4846
timestamp 1666464484
transform -1 0 7488 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4847
timestamp 1666464484
transform -1 0 7488 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4848
timestamp 1666464484
transform 1 0 6240 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4849
timestamp 1666464484
transform -1 0 6240 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4850
timestamp 1666464484
transform -1 0 7488 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4851
timestamp 1666464484
transform -1 0 7488 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4852
timestamp 1666464484
transform -1 0 7488 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4853
timestamp 1666464484
transform -1 0 7488 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4854
timestamp 1666464484
transform -1 0 6240 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4855
timestamp 1666464484
transform 1 0 6240 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4856
timestamp 1666464484
transform -1 0 7488 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4857
timestamp 1666464484
transform -1 0 7488 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4858
timestamp 1666464484
transform 1 0 6240 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4859
timestamp 1666464484
transform 1 0 7488 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4860
timestamp 1666464484
transform -1 0 1248 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4861
timestamp 1666464484
transform -1 0 1248 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4862
timestamp 1666464484
transform -1 0 1248 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4863
timestamp 1666464484
transform 1 0 3744 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4864
timestamp 1666464484
transform 1 0 3744 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4865
timestamp 1666464484
transform 1 0 3744 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4866
timestamp 1666464484
transform 1 0 3744 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4867
timestamp 1666464484
transform -1 0 3744 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4868
timestamp 1666464484
transform -1 0 3744 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4869
timestamp 1666464484
transform -1 0 3744 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4870
timestamp 1666464484
transform -1 0 3744 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4871
timestamp 1666464484
transform -1 0 3744 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4872
timestamp 1666464484
transform -1 0 3744 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4873
timestamp 1666464484
transform -1 0 3744 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4874
timestamp 1666464484
transform -1 0 3744 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4875
timestamp 1666464484
transform -1 0 3744 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4876
timestamp 1666464484
transform -1 0 3744 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4877
timestamp 1666464484
transform -1 0 3744 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4878
timestamp 1666464484
transform -1 0 3744 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4879
timestamp 1666464484
transform -1 0 3744 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4880
timestamp 1666464484
transform -1 0 3744 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4881
timestamp 1666464484
transform 1 0 0 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4882
timestamp 1666464484
transform 1 0 1248 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4883
timestamp 1666464484
transform 1 0 1248 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4884
timestamp 1666464484
transform 1 0 1248 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4885
timestamp 1666464484
transform 1 0 1248 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4886
timestamp 1666464484
transform 1 0 1248 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4887
timestamp 1666464484
transform 1 0 1248 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4888
timestamp 1666464484
transform 1 0 1248 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4889
timestamp 1666464484
transform 1 0 1248 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4890
timestamp 1666464484
transform 1 0 1248 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4891
timestamp 1666464484
transform 1 0 1248 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4892
timestamp 1666464484
transform 1 0 1248 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4893
timestamp 1666464484
transform 1 0 1248 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4894
timestamp 1666464484
transform 1 0 1248 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4895
timestamp 1666464484
transform 1 0 1248 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4896
timestamp 1666464484
transform 1 0 0 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4897
timestamp 1666464484
transform 1 0 0 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4898
timestamp 1666464484
transform 1 0 3744 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4899
timestamp 1666464484
transform 1 0 3744 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4900
timestamp 1666464484
transform 1 0 2496 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4901
timestamp 1666464484
transform 1 0 2496 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4902
timestamp 1666464484
transform 1 0 2496 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4903
timestamp 1666464484
transform 1 0 2496 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4904
timestamp 1666464484
transform 1 0 2496 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4905
timestamp 1666464484
transform 1 0 2496 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4906
timestamp 1666464484
transform 1 0 2496 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4907
timestamp 1666464484
transform 1 0 2496 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4908
timestamp 1666464484
transform 1 0 2496 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4909
timestamp 1666464484
transform 1 0 2496 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4910
timestamp 1666464484
transform 1 0 2496 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4911
timestamp 1666464484
transform 1 0 2496 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4912
timestamp 1666464484
transform 1 0 2496 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4913
timestamp 1666464484
transform 1 0 2496 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4914
timestamp 1666464484
transform 1 0 3744 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4915
timestamp 1666464484
transform 1 0 3744 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4916
timestamp 1666464484
transform 1 0 0 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4917
timestamp 1666464484
transform 1 0 0 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4918
timestamp 1666464484
transform 1 0 0 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4919
timestamp 1666464484
transform 1 0 3744 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4920
timestamp 1666464484
transform 1 0 3744 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4921
timestamp 1666464484
transform 1 0 0 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4922
timestamp 1666464484
transform 1 0 0 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4923
timestamp 1666464484
transform 1 0 0 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4924
timestamp 1666464484
transform 1 0 0 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4925
timestamp 1666464484
transform 1 0 0 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4926
timestamp 1666464484
transform 1 0 0 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4927
timestamp 1666464484
transform 1 0 0 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4928
timestamp 1666464484
transform 1 0 3744 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4929
timestamp 1666464484
transform 1 0 3744 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4930
timestamp 1666464484
transform 1 0 0 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4931
timestamp 1666464484
transform -1 0 1248 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4932
timestamp 1666464484
transform -1 0 1248 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4933
timestamp 1666464484
transform -1 0 2496 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4934
timestamp 1666464484
transform -1 0 2496 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4935
timestamp 1666464484
transform -1 0 2496 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4936
timestamp 1666464484
transform -1 0 2496 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4937
timestamp 1666464484
transform -1 0 2496 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4938
timestamp 1666464484
transform -1 0 2496 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4939
timestamp 1666464484
transform -1 0 2496 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4940
timestamp 1666464484
transform -1 0 2496 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4941
timestamp 1666464484
transform -1 0 2496 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4942
timestamp 1666464484
transform -1 0 2496 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4943
timestamp 1666464484
transform -1 0 2496 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4944
timestamp 1666464484
transform -1 0 2496 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4945
timestamp 1666464484
transform -1 0 2496 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4946
timestamp 1666464484
transform -1 0 2496 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4947
timestamp 1666464484
transform 1 0 3744 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4948
timestamp 1666464484
transform 1 0 3744 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4949
timestamp 1666464484
transform -1 0 1248 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4950
timestamp 1666464484
transform -1 0 1248 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4951
timestamp 1666464484
transform -1 0 1248 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4952
timestamp 1666464484
transform -1 0 1248 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4953
timestamp 1666464484
transform -1 0 1248 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4954
timestamp 1666464484
transform -1 0 1248 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4955
timestamp 1666464484
transform -1 0 1248 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4956
timestamp 1666464484
transform -1 0 1248 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4957
timestamp 1666464484
transform -1 0 1248 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4958
timestamp 1666464484
transform -1 0 3744 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4959
timestamp 1666464484
transform -1 0 3744 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4960
timestamp 1666464484
transform -1 0 3744 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4961
timestamp 1666464484
transform -1 0 3744 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4962
timestamp 1666464484
transform -1 0 3744 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4963
timestamp 1666464484
transform 1 0 3744 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4964
timestamp 1666464484
transform 1 0 3744 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4965
timestamp 1666464484
transform 1 0 3744 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4966
timestamp 1666464484
transform 1 0 3744 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4967
timestamp 1666464484
transform 1 0 3744 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4968
timestamp 1666464484
transform -1 0 3744 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4969
timestamp 1666464484
transform 1 0 3744 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4970
timestamp 1666464484
transform 1 0 1248 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4971
timestamp 1666464484
transform 1 0 0 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4972
timestamp 1666464484
transform 1 0 0 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4973
timestamp 1666464484
transform 1 0 0 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4974
timestamp 1666464484
transform -1 0 1248 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4975
timestamp 1666464484
transform -1 0 1248 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4976
timestamp 1666464484
transform -1 0 1248 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4977
timestamp 1666464484
transform -1 0 1248 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4978
timestamp 1666464484
transform -1 0 1248 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4979
timestamp 1666464484
transform -1 0 1248 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4980
timestamp 1666464484
transform 1 0 0 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4981
timestamp 1666464484
transform 1 0 0 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4982
timestamp 1666464484
transform 1 0 0 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4983
timestamp 1666464484
transform 1 0 1248 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4984
timestamp 1666464484
transform 1 0 1248 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4985
timestamp 1666464484
transform 1 0 1248 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4986
timestamp 1666464484
transform 1 0 1248 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4987
timestamp 1666464484
transform 1 0 1248 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4988
timestamp 1666464484
transform 1 0 1248 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4989
timestamp 1666464484
transform 1 0 0 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4990
timestamp 1666464484
transform 1 0 0 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4991
timestamp 1666464484
transform 1 0 0 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4992
timestamp 1666464484
transform 1 0 0 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4993
timestamp 1666464484
transform -1 0 1248 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4994
timestamp 1666464484
transform -1 0 1248 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4995
timestamp 1666464484
transform -1 0 1248 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4996
timestamp 1666464484
transform -1 0 1248 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4997
timestamp 1666464484
transform -1 0 1248 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4998
timestamp 1666464484
transform -1 0 1248 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_4999
timestamp 1666464484
transform -1 0 1248 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5000
timestamp 1666464484
transform 1 0 0 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5001
timestamp 1666464484
transform 1 0 0 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5002
timestamp 1666464484
transform 1 0 0 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5003
timestamp 1666464484
transform 1 0 1248 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5004
timestamp 1666464484
transform 1 0 1248 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5005
timestamp 1666464484
transform 1 0 1248 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5006
timestamp 1666464484
transform 1 0 1248 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5007
timestamp 1666464484
transform 1 0 1248 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5008
timestamp 1666464484
transform 1 0 1248 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5009
timestamp 1666464484
transform -1 0 3744 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5010
timestamp 1666464484
transform -1 0 3744 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5011
timestamp 1666464484
transform 1 0 3744 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5012
timestamp 1666464484
transform 1 0 3744 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5013
timestamp 1666464484
transform -1 0 3744 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5014
timestamp 1666464484
transform -1 0 3744 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5015
timestamp 1666464484
transform -1 0 3744 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5016
timestamp 1666464484
transform 1 0 3744 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5017
timestamp 1666464484
transform 1 0 3744 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5018
timestamp 1666464484
transform 1 0 3744 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5019
timestamp 1666464484
transform -1 0 3744 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5020
timestamp 1666464484
transform -1 0 3744 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5021
timestamp 1666464484
transform 1 0 3744 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5022
timestamp 1666464484
transform 1 0 3744 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5023
timestamp 1666464484
transform 1 0 2496 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5024
timestamp 1666464484
transform 1 0 2496 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5025
timestamp 1666464484
transform 1 0 2496 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5026
timestamp 1666464484
transform 1 0 2496 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5027
timestamp 1666464484
transform 1 0 2496 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5028
timestamp 1666464484
transform 1 0 2496 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5029
timestamp 1666464484
transform 1 0 2496 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5030
timestamp 1666464484
transform 1 0 2496 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5031
timestamp 1666464484
transform 1 0 2496 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5032
timestamp 1666464484
transform 1 0 2496 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5033
timestamp 1666464484
transform 1 0 2496 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5034
timestamp 1666464484
transform 1 0 2496 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5035
timestamp 1666464484
transform 1 0 2496 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5036
timestamp 1666464484
transform 1 0 2496 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5037
timestamp 1666464484
transform 1 0 2496 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5038
timestamp 1666464484
transform -1 0 2496 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5039
timestamp 1666464484
transform -1 0 2496 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5040
timestamp 1666464484
transform -1 0 2496 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5041
timestamp 1666464484
transform -1 0 2496 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5042
timestamp 1666464484
transform -1 0 2496 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5043
timestamp 1666464484
transform -1 0 2496 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5044
timestamp 1666464484
transform -1 0 2496 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5045
timestamp 1666464484
transform -1 0 2496 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5046
timestamp 1666464484
transform -1 0 2496 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5047
timestamp 1666464484
transform -1 0 2496 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5048
timestamp 1666464484
transform -1 0 2496 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5049
timestamp 1666464484
transform -1 0 2496 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5050
timestamp 1666464484
transform -1 0 2496 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5051
timestamp 1666464484
transform -1 0 2496 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5052
timestamp 1666464484
transform -1 0 2496 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5053
timestamp 1666464484
transform 1 0 1248 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5054
timestamp 1666464484
transform 1 0 1248 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5055
timestamp 1666464484
transform 1 0 3744 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5056
timestamp 1666464484
transform -1 0 1248 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5057
timestamp 1666464484
transform -1 0 1248 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5058
timestamp 1666464484
transform 1 0 3744 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5059
timestamp 1666464484
transform -1 0 3744 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5060
timestamp 1666464484
transform -1 0 3744 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5061
timestamp 1666464484
transform 1 0 0 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5062
timestamp 1666464484
transform 1 0 0 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5063
timestamp 1666464484
transform 1 0 6240 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5064
timestamp 1666464484
transform 1 0 6240 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5065
timestamp 1666464484
transform 1 0 6240 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5066
timestamp 1666464484
transform 1 0 6240 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5067
timestamp 1666464484
transform 1 0 6240 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5068
timestamp 1666464484
transform -1 0 6240 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5069
timestamp 1666464484
transform -1 0 6240 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5070
timestamp 1666464484
transform -1 0 6240 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5071
timestamp 1666464484
transform -1 0 6240 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5072
timestamp 1666464484
transform -1 0 6240 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5073
timestamp 1666464484
transform -1 0 6240 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5074
timestamp 1666464484
transform -1 0 6240 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5075
timestamp 1666464484
transform 1 0 8736 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5076
timestamp 1666464484
transform 1 0 8736 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5077
timestamp 1666464484
transform 1 0 8736 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5078
timestamp 1666464484
transform 1 0 8736 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5079
timestamp 1666464484
transform 1 0 8736 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5080
timestamp 1666464484
transform 1 0 8736 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5081
timestamp 1666464484
transform 1 0 8736 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5082
timestamp 1666464484
transform 1 0 8736 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5083
timestamp 1666464484
transform 1 0 8736 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5084
timestamp 1666464484
transform 1 0 8736 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5085
timestamp 1666464484
transform 1 0 8736 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5086
timestamp 1666464484
transform 1 0 8736 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5087
timestamp 1666464484
transform 1 0 8736 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5088
timestamp 1666464484
transform 1 0 8736 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5089
timestamp 1666464484
transform 1 0 8736 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5090
timestamp 1666464484
transform -1 0 6240 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5091
timestamp 1666464484
transform -1 0 6240 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5092
timestamp 1666464484
transform -1 0 8736 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5093
timestamp 1666464484
transform -1 0 8736 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5094
timestamp 1666464484
transform -1 0 8736 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5095
timestamp 1666464484
transform -1 0 8736 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5096
timestamp 1666464484
transform -1 0 8736 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5097
timestamp 1666464484
transform -1 0 8736 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5098
timestamp 1666464484
transform -1 0 8736 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5099
timestamp 1666464484
transform -1 0 8736 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5100
timestamp 1666464484
transform -1 0 8736 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5101
timestamp 1666464484
transform -1 0 8736 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5102
timestamp 1666464484
transform -1 0 8736 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5103
timestamp 1666464484
transform -1 0 8736 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5104
timestamp 1666464484
transform -1 0 8736 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5105
timestamp 1666464484
transform -1 0 8736 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5106
timestamp 1666464484
transform -1 0 8736 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5107
timestamp 1666464484
transform -1 0 6240 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5108
timestamp 1666464484
transform -1 0 6240 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5109
timestamp 1666464484
transform 1 0 7488 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5110
timestamp 1666464484
transform 1 0 7488 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5111
timestamp 1666464484
transform 1 0 7488 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5112
timestamp 1666464484
transform 1 0 7488 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5113
timestamp 1666464484
transform 1 0 7488 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5114
timestamp 1666464484
transform 1 0 7488 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5115
timestamp 1666464484
transform 1 0 7488 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5116
timestamp 1666464484
transform 1 0 7488 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5117
timestamp 1666464484
transform 1 0 7488 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5118
timestamp 1666464484
transform 1 0 7488 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5119
timestamp 1666464484
transform 1 0 7488 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5120
timestamp 1666464484
transform 1 0 7488 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5121
timestamp 1666464484
transform 1 0 7488 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5122
timestamp 1666464484
transform 1 0 7488 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5123
timestamp 1666464484
transform 1 0 7488 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5124
timestamp 1666464484
transform -1 0 6240 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5125
timestamp 1666464484
transform -1 0 6240 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5126
timestamp 1666464484
transform -1 0 7488 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5127
timestamp 1666464484
transform -1 0 7488 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5128
timestamp 1666464484
transform -1 0 7488 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5129
timestamp 1666464484
transform -1 0 7488 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5130
timestamp 1666464484
transform -1 0 7488 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5131
timestamp 1666464484
transform -1 0 7488 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5132
timestamp 1666464484
transform -1 0 7488 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5133
timestamp 1666464484
transform -1 0 7488 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5134
timestamp 1666464484
transform -1 0 7488 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5135
timestamp 1666464484
transform -1 0 7488 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5136
timestamp 1666464484
transform -1 0 7488 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5137
timestamp 1666464484
transform -1 0 7488 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5138
timestamp 1666464484
transform -1 0 7488 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5139
timestamp 1666464484
transform -1 0 7488 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5140
timestamp 1666464484
transform -1 0 7488 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5141
timestamp 1666464484
transform -1 0 6240 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5142
timestamp 1666464484
transform -1 0 6240 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5143
timestamp 1666464484
transform 1 0 6240 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5144
timestamp 1666464484
transform 1 0 6240 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5145
timestamp 1666464484
transform 1 0 6240 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5146
timestamp 1666464484
transform 1 0 6240 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5147
timestamp 1666464484
transform 1 0 6240 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5148
timestamp 1666464484
transform 1 0 6240 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5149
timestamp 1666464484
transform 1 0 6240 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5150
timestamp 1666464484
transform 1 0 6240 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5151
timestamp 1666464484
transform 1 0 6240 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5152
timestamp 1666464484
transform 1 0 6240 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5153
timestamp 1666464484
transform -1 0 3744 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5154
timestamp 1666464484
transform -1 0 3744 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5155
timestamp 1666464484
transform 1 0 3744 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5156
timestamp 1666464484
transform 1 0 3744 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5157
timestamp 1666464484
transform 1 0 2496 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5158
timestamp 1666464484
transform 1 0 2496 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5159
timestamp 1666464484
transform -1 0 2496 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5160
timestamp 1666464484
transform -1 0 2496 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5161
timestamp 1666464484
transform 1 0 1248 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5162
timestamp 1666464484
transform 1 0 1248 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5163
timestamp 1666464484
transform -1 0 1248 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5164
timestamp 1666464484
transform -1 0 1248 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5165
timestamp 1666464484
transform 1 0 8736 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5166
timestamp 1666464484
transform 1 0 8736 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5167
timestamp 1666464484
transform -1 0 8736 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5168
timestamp 1666464484
transform -1 0 8736 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5169
timestamp 1666464484
transform 1 0 7488 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5170
timestamp 1666464484
transform 1 0 7488 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5171
timestamp 1666464484
transform -1 0 7488 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5172
timestamp 1666464484
transform -1 0 7488 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5173
timestamp 1666464484
transform 1 0 6240 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5174
timestamp 1666464484
transform 1 0 6240 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5175
timestamp 1666464484
transform -1 0 6240 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5176
timestamp 1666464484
transform -1 0 6240 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5177
timestamp 1666464484
transform 1 0 4992 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5178
timestamp 1666464484
transform 1 0 4992 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5179
timestamp 1666464484
transform 1 0 4992 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5180
timestamp 1666464484
transform 1 0 4992 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5181
timestamp 1666464484
transform 1 0 4992 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5182
timestamp 1666464484
transform 1 0 4992 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5183
timestamp 1666464484
transform 1 0 4992 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5184
timestamp 1666464484
transform 1 0 4992 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5185
timestamp 1666464484
transform 1 0 4992 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5186
timestamp 1666464484
transform 1 0 4992 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5187
timestamp 1666464484
transform 1 0 4992 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5188
timestamp 1666464484
transform 1 0 4992 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5189
timestamp 1666464484
transform 1 0 4992 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5190
timestamp 1666464484
transform 1 0 4992 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5191
timestamp 1666464484
transform 1 0 4992 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5192
timestamp 1666464484
transform 1 0 4992 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5193
timestamp 1666464484
transform 1 0 4992 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5194
timestamp 1666464484
transform 1 0 4992 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5195
timestamp 1666464484
transform 1 0 4992 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5196
timestamp 1666464484
transform 1 0 4992 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5197
timestamp 1666464484
transform 1 0 4992 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5198
timestamp 1666464484
transform 1 0 0 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5199
timestamp 1666464484
transform 1 0 0 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5200
timestamp 1666464484
transform 1 0 4992 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5201
timestamp 1666464484
transform 1 0 4992 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5202
timestamp 1666464484
transform 1 0 4992 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5203
timestamp 1666464484
transform 1 0 4992 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5204
timestamp 1666464484
transform 1 0 4992 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5205
timestamp 1666464484
transform 1 0 4992 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5206
timestamp 1666464484
transform 1 0 4992 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5207
timestamp 1666464484
transform 1 0 4992 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5208
timestamp 1666464484
transform 1 0 4992 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5209
timestamp 1666464484
transform 1 0 4992 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5210
timestamp 1666464484
transform -1 0 4992 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5211
timestamp 1666464484
transform -1 0 4992 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5212
timestamp 1666464484
transform -1 0 4992 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5213
timestamp 1666464484
transform -1 0 4992 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5214
timestamp 1666464484
transform -1 0 4992 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5215
timestamp 1666464484
transform -1 0 4992 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5216
timestamp 1666464484
transform -1 0 4992 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5217
timestamp 1666464484
transform -1 0 4992 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5218
timestamp 1666464484
transform -1 0 4992 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5219
timestamp 1666464484
transform -1 0 4992 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5220
timestamp 1666464484
transform -1 0 4992 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5221
timestamp 1666464484
transform -1 0 4992 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5222
timestamp 1666464484
transform -1 0 4992 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5223
timestamp 1666464484
transform -1 0 4992 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5224
timestamp 1666464484
transform -1 0 4992 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5225
timestamp 1666464484
transform -1 0 4992 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5226
timestamp 1666464484
transform -1 0 4992 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5227
timestamp 1666464484
transform -1 0 4992 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5228
timestamp 1666464484
transform -1 0 4992 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5229
timestamp 1666464484
transform -1 0 4992 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5230
timestamp 1666464484
transform -1 0 4992 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5231
timestamp 1666464484
transform -1 0 4992 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5232
timestamp 1666464484
transform -1 0 4992 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5233
timestamp 1666464484
transform -1 0 4992 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5234
timestamp 1666464484
transform -1 0 4992 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5235
timestamp 1666464484
transform -1 0 4992 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5236
timestamp 1666464484
transform -1 0 4992 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5237
timestamp 1666464484
transform -1 0 4992 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5238
timestamp 1666464484
transform -1 0 4992 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5239
timestamp 1666464484
transform -1 0 4992 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5240
timestamp 1666464484
transform -1 0 4992 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5241
timestamp 1666464484
transform 1 0 16224 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5242
timestamp 1666464484
transform 1 0 16224 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5243
timestamp 1666464484
transform 1 0 16224 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5244
timestamp 1666464484
transform 1 0 16224 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5245
timestamp 1666464484
transform 1 0 16224 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5246
timestamp 1666464484
transform -1 0 16224 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5247
timestamp 1666464484
transform -1 0 16224 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5248
timestamp 1666464484
transform -1 0 16224 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5249
timestamp 1666464484
transform -1 0 16224 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5250
timestamp 1666464484
transform 1 0 17472 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5251
timestamp 1666464484
transform 1 0 17472 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5252
timestamp 1666464484
transform 1 0 17472 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5253
timestamp 1666464484
transform 1 0 17472 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5254
timestamp 1666464484
transform 1 0 17472 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5255
timestamp 1666464484
transform 1 0 17472 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5256
timestamp 1666464484
transform 1 0 17472 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5257
timestamp 1666464484
transform 1 0 17472 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5258
timestamp 1666464484
transform 1 0 17472 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5259
timestamp 1666464484
transform 1 0 17472 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5260
timestamp 1666464484
transform 1 0 17472 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5261
timestamp 1666464484
transform 1 0 17472 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5262
timestamp 1666464484
transform 1 0 17472 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5263
timestamp 1666464484
transform 1 0 17472 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5264
timestamp 1666464484
transform -1 0 16224 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5265
timestamp 1666464484
transform -1 0 16224 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5266
timestamp 1666464484
transform -1 0 16224 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5267
timestamp 1666464484
transform -1 0 16224 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5268
timestamp 1666464484
transform 1 0 18720 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5269
timestamp 1666464484
transform 1 0 18720 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5270
timestamp 1666464484
transform 1 0 18720 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5271
timestamp 1666464484
transform 1 0 18720 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5272
timestamp 1666464484
transform 1 0 18720 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5273
timestamp 1666464484
transform 1 0 18720 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5274
timestamp 1666464484
transform 1 0 18720 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5275
timestamp 1666464484
transform 1 0 18720 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5276
timestamp 1666464484
transform 1 0 18720 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5277
timestamp 1666464484
transform 1 0 18720 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5278
timestamp 1666464484
transform 1 0 18720 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5279
timestamp 1666464484
transform 1 0 18720 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5280
timestamp 1666464484
transform 1 0 18720 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5281
timestamp 1666464484
transform 1 0 18720 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5282
timestamp 1666464484
transform -1 0 16224 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5283
timestamp 1666464484
transform -1 0 16224 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5284
timestamp 1666464484
transform -1 0 16224 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5285
timestamp 1666464484
transform -1 0 16224 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5286
timestamp 1666464484
transform -1 0 16224 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5287
timestamp 1666464484
transform -1 0 16224 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5288
timestamp 1666464484
transform 1 0 16224 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5289
timestamp 1666464484
transform 1 0 16224 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5290
timestamp 1666464484
transform 1 0 16224 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5291
timestamp 1666464484
transform 1 0 16224 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5292
timestamp 1666464484
transform 1 0 16224 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5293
timestamp 1666464484
transform 1 0 16224 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5294
timestamp 1666464484
transform 1 0 16224 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5295
timestamp 1666464484
transform 1 0 16224 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5296
timestamp 1666464484
transform 1 0 16224 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5297
timestamp 1666464484
transform -1 0 17472 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5298
timestamp 1666464484
transform -1 0 17472 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5299
timestamp 1666464484
transform -1 0 17472 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5300
timestamp 1666464484
transform -1 0 17472 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5301
timestamp 1666464484
transform -1 0 18720 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5302
timestamp 1666464484
transform -1 0 18720 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5303
timestamp 1666464484
transform -1 0 18720 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5304
timestamp 1666464484
transform -1 0 18720 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5305
timestamp 1666464484
transform -1 0 18720 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5306
timestamp 1666464484
transform -1 0 18720 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5307
timestamp 1666464484
transform -1 0 18720 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5308
timestamp 1666464484
transform -1 0 18720 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5309
timestamp 1666464484
transform -1 0 18720 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5310
timestamp 1666464484
transform -1 0 18720 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5311
timestamp 1666464484
transform -1 0 18720 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5312
timestamp 1666464484
transform -1 0 18720 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5313
timestamp 1666464484
transform -1 0 18720 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5314
timestamp 1666464484
transform -1 0 18720 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5315
timestamp 1666464484
transform -1 0 17472 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5316
timestamp 1666464484
transform -1 0 17472 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5317
timestamp 1666464484
transform -1 0 17472 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5318
timestamp 1666464484
transform -1 0 17472 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5319
timestamp 1666464484
transform -1 0 17472 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5320
timestamp 1666464484
transform -1 0 17472 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5321
timestamp 1666464484
transform -1 0 17472 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5322
timestamp 1666464484
transform -1 0 17472 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5323
timestamp 1666464484
transform -1 0 17472 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5324
timestamp 1666464484
transform -1 0 17472 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5325
timestamp 1666464484
transform 1 0 11232 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5326
timestamp 1666464484
transform 1 0 11232 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5327
timestamp 1666464484
transform 1 0 11232 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5328
timestamp 1666464484
transform -1 0 11232 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5329
timestamp 1666464484
transform -1 0 11232 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5330
timestamp 1666464484
transform -1 0 13728 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5331
timestamp 1666464484
transform -1 0 13728 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5332
timestamp 1666464484
transform -1 0 13728 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5333
timestamp 1666464484
transform -1 0 13728 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5334
timestamp 1666464484
transform -1 0 13728 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5335
timestamp 1666464484
transform -1 0 13728 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5336
timestamp 1666464484
transform -1 0 13728 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5337
timestamp 1666464484
transform -1 0 13728 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5338
timestamp 1666464484
transform -1 0 13728 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5339
timestamp 1666464484
transform -1 0 13728 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5340
timestamp 1666464484
transform -1 0 13728 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5341
timestamp 1666464484
transform -1 0 13728 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5342
timestamp 1666464484
transform -1 0 13728 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5343
timestamp 1666464484
transform -1 0 13728 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5344
timestamp 1666464484
transform -1 0 11232 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5345
timestamp 1666464484
transform -1 0 11232 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5346
timestamp 1666464484
transform 1 0 11232 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5347
timestamp 1666464484
transform 1 0 11232 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5348
timestamp 1666464484
transform 1 0 11232 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5349
timestamp 1666464484
transform 1 0 11232 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5350
timestamp 1666464484
transform 1 0 11232 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5351
timestamp 1666464484
transform 1 0 11232 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5352
timestamp 1666464484
transform 1 0 11232 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5353
timestamp 1666464484
transform -1 0 12480 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5354
timestamp 1666464484
transform -1 0 12480 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5355
timestamp 1666464484
transform -1 0 11232 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5356
timestamp 1666464484
transform -1 0 11232 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5357
timestamp 1666464484
transform -1 0 12480 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5358
timestamp 1666464484
transform -1 0 12480 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5359
timestamp 1666464484
transform -1 0 12480 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5360
timestamp 1666464484
transform -1 0 12480 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5361
timestamp 1666464484
transform -1 0 12480 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5362
timestamp 1666464484
transform -1 0 12480 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5363
timestamp 1666464484
transform -1 0 12480 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5364
timestamp 1666464484
transform -1 0 12480 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5365
timestamp 1666464484
transform 1 0 12480 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5366
timestamp 1666464484
transform 1 0 12480 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5367
timestamp 1666464484
transform 1 0 12480 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5368
timestamp 1666464484
transform 1 0 12480 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5369
timestamp 1666464484
transform 1 0 12480 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5370
timestamp 1666464484
transform 1 0 12480 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5371
timestamp 1666464484
transform 1 0 12480 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5372
timestamp 1666464484
transform 1 0 12480 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5373
timestamp 1666464484
transform 1 0 12480 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5374
timestamp 1666464484
transform 1 0 13728 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5375
timestamp 1666464484
transform 1 0 13728 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5376
timestamp 1666464484
transform 1 0 13728 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5377
timestamp 1666464484
transform 1 0 13728 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5378
timestamp 1666464484
transform 1 0 13728 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5379
timestamp 1666464484
transform 1 0 13728 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5380
timestamp 1666464484
transform 1 0 13728 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5381
timestamp 1666464484
transform 1 0 13728 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5382
timestamp 1666464484
transform 1 0 13728 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5383
timestamp 1666464484
transform 1 0 13728 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5384
timestamp 1666464484
transform 1 0 13728 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5385
timestamp 1666464484
transform 1 0 13728 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5386
timestamp 1666464484
transform 1 0 13728 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5387
timestamp 1666464484
transform 1 0 13728 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5388
timestamp 1666464484
transform -1 0 11232 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5389
timestamp 1666464484
transform -1 0 11232 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5390
timestamp 1666464484
transform 1 0 12480 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5391
timestamp 1666464484
transform 1 0 12480 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5392
timestamp 1666464484
transform 1 0 12480 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5393
timestamp 1666464484
transform 1 0 12480 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5394
timestamp 1666464484
transform 1 0 12480 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5395
timestamp 1666464484
transform -1 0 11232 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5396
timestamp 1666464484
transform -1 0 11232 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5397
timestamp 1666464484
transform -1 0 12480 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5398
timestamp 1666464484
transform -1 0 12480 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5399
timestamp 1666464484
transform -1 0 12480 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5400
timestamp 1666464484
transform -1 0 12480 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5401
timestamp 1666464484
transform -1 0 11232 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5402
timestamp 1666464484
transform -1 0 11232 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5403
timestamp 1666464484
transform -1 0 11232 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5404
timestamp 1666464484
transform -1 0 11232 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5405
timestamp 1666464484
transform 1 0 11232 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5406
timestamp 1666464484
transform 1 0 11232 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5407
timestamp 1666464484
transform 1 0 11232 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5408
timestamp 1666464484
transform 1 0 11232 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5409
timestamp 1666464484
transform -1 0 11232 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5410
timestamp 1666464484
transform -1 0 11232 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5411
timestamp 1666464484
transform -1 0 11232 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5412
timestamp 1666464484
transform -1 0 11232 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5413
timestamp 1666464484
transform -1 0 11232 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5414
timestamp 1666464484
transform -1 0 12480 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5415
timestamp 1666464484
transform -1 0 12480 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5416
timestamp 1666464484
transform -1 0 12480 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5417
timestamp 1666464484
transform -1 0 12480 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5418
timestamp 1666464484
transform -1 0 12480 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5419
timestamp 1666464484
transform 1 0 11232 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5420
timestamp 1666464484
transform 1 0 11232 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5421
timestamp 1666464484
transform 1 0 11232 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5422
timestamp 1666464484
transform -1 0 11232 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5423
timestamp 1666464484
transform -1 0 11232 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5424
timestamp 1666464484
transform 1 0 11232 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5425
timestamp 1666464484
transform 1 0 11232 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5426
timestamp 1666464484
transform 1 0 11232 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5427
timestamp 1666464484
transform 1 0 11232 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5428
timestamp 1666464484
transform 1 0 11232 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5429
timestamp 1666464484
transform 1 0 11232 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5430
timestamp 1666464484
transform 1 0 13728 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5431
timestamp 1666464484
transform -1 0 11232 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5432
timestamp 1666464484
transform -1 0 11232 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5433
timestamp 1666464484
transform 1 0 13728 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5434
timestamp 1666464484
transform 1 0 13728 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5435
timestamp 1666464484
transform 1 0 13728 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5436
timestamp 1666464484
transform 1 0 13728 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5437
timestamp 1666464484
transform 1 0 13728 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5438
timestamp 1666464484
transform 1 0 13728 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5439
timestamp 1666464484
transform 1 0 13728 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5440
timestamp 1666464484
transform 1 0 13728 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5441
timestamp 1666464484
transform 1 0 13728 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5442
timestamp 1666464484
transform 1 0 13728 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5443
timestamp 1666464484
transform 1 0 13728 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5444
timestamp 1666464484
transform 1 0 13728 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5445
timestamp 1666464484
transform 1 0 13728 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5446
timestamp 1666464484
transform 1 0 13728 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5447
timestamp 1666464484
transform 1 0 11232 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5448
timestamp 1666464484
transform 1 0 11232 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5449
timestamp 1666464484
transform -1 0 13728 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5450
timestamp 1666464484
transform -1 0 11232 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5451
timestamp 1666464484
transform -1 0 11232 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5452
timestamp 1666464484
transform -1 0 13728 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5453
timestamp 1666464484
transform -1 0 13728 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5454
timestamp 1666464484
transform -1 0 13728 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5455
timestamp 1666464484
transform -1 0 13728 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5456
timestamp 1666464484
transform -1 0 13728 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5457
timestamp 1666464484
transform -1 0 13728 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5458
timestamp 1666464484
transform -1 0 13728 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5459
timestamp 1666464484
transform -1 0 13728 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5460
timestamp 1666464484
transform -1 0 13728 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5461
timestamp 1666464484
transform -1 0 13728 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5462
timestamp 1666464484
transform -1 0 13728 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5463
timestamp 1666464484
transform -1 0 13728 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5464
timestamp 1666464484
transform -1 0 13728 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5465
timestamp 1666464484
transform -1 0 13728 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5466
timestamp 1666464484
transform 1 0 11232 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5467
timestamp 1666464484
transform 1 0 11232 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5468
timestamp 1666464484
transform 1 0 12480 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5469
timestamp 1666464484
transform -1 0 11232 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5470
timestamp 1666464484
transform -1 0 11232 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5471
timestamp 1666464484
transform 1 0 12480 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5472
timestamp 1666464484
transform 1 0 12480 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5473
timestamp 1666464484
transform 1 0 12480 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5474
timestamp 1666464484
transform 1 0 12480 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5475
timestamp 1666464484
transform 1 0 12480 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5476
timestamp 1666464484
transform 1 0 12480 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5477
timestamp 1666464484
transform 1 0 12480 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5478
timestamp 1666464484
transform 1 0 12480 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5479
timestamp 1666464484
transform 1 0 12480 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5480
timestamp 1666464484
transform 1 0 12480 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5481
timestamp 1666464484
transform 1 0 12480 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5482
timestamp 1666464484
transform 1 0 12480 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5483
timestamp 1666464484
transform 1 0 12480 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5484
timestamp 1666464484
transform 1 0 12480 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5485
timestamp 1666464484
transform 1 0 11232 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5486
timestamp 1666464484
transform 1 0 11232 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5487
timestamp 1666464484
transform -1 0 12480 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5488
timestamp 1666464484
transform -1 0 11232 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5489
timestamp 1666464484
transform -1 0 11232 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5490
timestamp 1666464484
transform -1 0 12480 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5491
timestamp 1666464484
transform -1 0 12480 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5492
timestamp 1666464484
transform -1 0 12480 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5493
timestamp 1666464484
transform -1 0 12480 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5494
timestamp 1666464484
transform -1 0 12480 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5495
timestamp 1666464484
transform -1 0 12480 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5496
timestamp 1666464484
transform -1 0 12480 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5497
timestamp 1666464484
transform -1 0 12480 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5498
timestamp 1666464484
transform -1 0 12480 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5499
timestamp 1666464484
transform 1 0 18720 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5500
timestamp 1666464484
transform 1 0 18720 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5501
timestamp 1666464484
transform 1 0 18720 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5502
timestamp 1666464484
transform 1 0 18720 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5503
timestamp 1666464484
transform 1 0 18720 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5504
timestamp 1666464484
transform 1 0 18720 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5505
timestamp 1666464484
transform 1 0 18720 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5506
timestamp 1666464484
transform 1 0 18720 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5507
timestamp 1666464484
transform 1 0 18720 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5508
timestamp 1666464484
transform 1 0 18720 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5509
timestamp 1666464484
transform 1 0 18720 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5510
timestamp 1666464484
transform 1 0 18720 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5511
timestamp 1666464484
transform 1 0 18720 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5512
timestamp 1666464484
transform 1 0 18720 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5513
timestamp 1666464484
transform 1 0 18720 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5514
timestamp 1666464484
transform -1 0 16224 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5515
timestamp 1666464484
transform -1 0 16224 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5516
timestamp 1666464484
transform -1 0 18720 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5517
timestamp 1666464484
transform -1 0 18720 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5518
timestamp 1666464484
transform -1 0 18720 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5519
timestamp 1666464484
transform -1 0 18720 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5520
timestamp 1666464484
transform -1 0 18720 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5521
timestamp 1666464484
transform -1 0 18720 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5522
timestamp 1666464484
transform -1 0 18720 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5523
timestamp 1666464484
transform -1 0 18720 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5524
timestamp 1666464484
transform -1 0 18720 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5525
timestamp 1666464484
transform -1 0 18720 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5526
timestamp 1666464484
transform -1 0 18720 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5527
timestamp 1666464484
transform -1 0 18720 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5528
timestamp 1666464484
transform -1 0 18720 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5529
timestamp 1666464484
transform -1 0 18720 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5530
timestamp 1666464484
transform -1 0 18720 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5531
timestamp 1666464484
transform -1 0 16224 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5532
timestamp 1666464484
transform -1 0 16224 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5533
timestamp 1666464484
transform 1 0 17472 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5534
timestamp 1666464484
transform 1 0 17472 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5535
timestamp 1666464484
transform 1 0 17472 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5536
timestamp 1666464484
transform 1 0 17472 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5537
timestamp 1666464484
transform 1 0 17472 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5538
timestamp 1666464484
transform 1 0 17472 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5539
timestamp 1666464484
transform 1 0 17472 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5540
timestamp 1666464484
transform 1 0 17472 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5541
timestamp 1666464484
transform 1 0 17472 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5542
timestamp 1666464484
transform 1 0 17472 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5543
timestamp 1666464484
transform 1 0 17472 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5544
timestamp 1666464484
transform 1 0 17472 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5545
timestamp 1666464484
transform 1 0 17472 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5546
timestamp 1666464484
transform 1 0 17472 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5547
timestamp 1666464484
transform 1 0 17472 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5548
timestamp 1666464484
transform -1 0 16224 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5549
timestamp 1666464484
transform -1 0 16224 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5550
timestamp 1666464484
transform -1 0 17472 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5551
timestamp 1666464484
transform -1 0 17472 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5552
timestamp 1666464484
transform -1 0 17472 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5553
timestamp 1666464484
transform -1 0 17472 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5554
timestamp 1666464484
transform -1 0 17472 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5555
timestamp 1666464484
transform -1 0 17472 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5556
timestamp 1666464484
transform -1 0 17472 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5557
timestamp 1666464484
transform -1 0 17472 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5558
timestamp 1666464484
transform -1 0 17472 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5559
timestamp 1666464484
transform -1 0 17472 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5560
timestamp 1666464484
transform -1 0 17472 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5561
timestamp 1666464484
transform -1 0 17472 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5562
timestamp 1666464484
transform -1 0 17472 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5563
timestamp 1666464484
transform -1 0 17472 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5564
timestamp 1666464484
transform -1 0 17472 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5565
timestamp 1666464484
transform -1 0 16224 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5566
timestamp 1666464484
transform -1 0 16224 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5567
timestamp 1666464484
transform 1 0 16224 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5568
timestamp 1666464484
transform 1 0 16224 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5569
timestamp 1666464484
transform 1 0 16224 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5570
timestamp 1666464484
transform 1 0 16224 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5571
timestamp 1666464484
transform 1 0 16224 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5572
timestamp 1666464484
transform 1 0 16224 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5573
timestamp 1666464484
transform 1 0 16224 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5574
timestamp 1666464484
transform 1 0 16224 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5575
timestamp 1666464484
transform 1 0 16224 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5576
timestamp 1666464484
transform 1 0 16224 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5577
timestamp 1666464484
transform 1 0 16224 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5578
timestamp 1666464484
transform 1 0 16224 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5579
timestamp 1666464484
transform 1 0 16224 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5580
timestamp 1666464484
transform 1 0 16224 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5581
timestamp 1666464484
transform 1 0 16224 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5582
timestamp 1666464484
transform -1 0 16224 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5583
timestamp 1666464484
transform -1 0 16224 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5584
timestamp 1666464484
transform -1 0 16224 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5585
timestamp 1666464484
transform -1 0 16224 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5586
timestamp 1666464484
transform -1 0 16224 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5587
timestamp 1666464484
transform -1 0 16224 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5588
timestamp 1666464484
transform -1 0 16224 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5589
timestamp 1666464484
transform 1 0 18720 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5590
timestamp 1666464484
transform 1 0 18720 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5591
timestamp 1666464484
transform -1 0 18720 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5592
timestamp 1666464484
transform -1 0 18720 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5593
timestamp 1666464484
transform 1 0 17472 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5594
timestamp 1666464484
transform 1 0 17472 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5595
timestamp 1666464484
transform -1 0 17472 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5596
timestamp 1666464484
transform -1 0 17472 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5597
timestamp 1666464484
transform 1 0 16224 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5598
timestamp 1666464484
transform 1 0 16224 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5599
timestamp 1666464484
transform -1 0 16224 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5600
timestamp 1666464484
transform -1 0 16224 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5601
timestamp 1666464484
transform -1 0 11232 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5602
timestamp 1666464484
transform -1 0 11232 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5603
timestamp 1666464484
transform 1 0 14976 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5604
timestamp 1666464484
transform 1 0 14976 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5605
timestamp 1666464484
transform 1 0 14976 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5606
timestamp 1666464484
transform 1 0 14976 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5607
timestamp 1666464484
transform 1 0 14976 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5608
timestamp 1666464484
transform 1 0 14976 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5609
timestamp 1666464484
transform 1 0 14976 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5610
timestamp 1666464484
transform 1 0 14976 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5611
timestamp 1666464484
transform 1 0 14976 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5612
timestamp 1666464484
transform 1 0 14976 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5613
timestamp 1666464484
transform 1 0 14976 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5614
timestamp 1666464484
transform 1 0 14976 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5615
timestamp 1666464484
transform 1 0 14976 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5616
timestamp 1666464484
transform 1 0 14976 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5617
timestamp 1666464484
transform 1 0 14976 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5618
timestamp 1666464484
transform 1 0 14976 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5619
timestamp 1666464484
transform 1 0 14976 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5620
timestamp 1666464484
transform 1 0 14976 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5621
timestamp 1666464484
transform 1 0 14976 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5622
timestamp 1666464484
transform 1 0 14976 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5623
timestamp 1666464484
transform 1 0 14976 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5624
timestamp 1666464484
transform 1 0 14976 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5625
timestamp 1666464484
transform 1 0 14976 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5626
timestamp 1666464484
transform 1 0 14976 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5627
timestamp 1666464484
transform 1 0 14976 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5628
timestamp 1666464484
transform 1 0 14976 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5629
timestamp 1666464484
transform 1 0 14976 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5630
timestamp 1666464484
transform 1 0 14976 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5631
timestamp 1666464484
transform 1 0 14976 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5632
timestamp 1666464484
transform 1 0 14976 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5633
timestamp 1666464484
transform 1 0 14976 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5634
timestamp 1666464484
transform -1 0 14976 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5635
timestamp 1666464484
transform -1 0 14976 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5636
timestamp 1666464484
transform -1 0 14976 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5637
timestamp 1666464484
transform -1 0 14976 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5638
timestamp 1666464484
transform -1 0 14976 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5639
timestamp 1666464484
transform -1 0 14976 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5640
timestamp 1666464484
transform -1 0 14976 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5641
timestamp 1666464484
transform -1 0 14976 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5642
timestamp 1666464484
transform -1 0 14976 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5643
timestamp 1666464484
transform -1 0 14976 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5644
timestamp 1666464484
transform -1 0 14976 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5645
timestamp 1666464484
transform -1 0 14976 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5646
timestamp 1666464484
transform -1 0 14976 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5647
timestamp 1666464484
transform -1 0 14976 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5648
timestamp 1666464484
transform -1 0 14976 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5649
timestamp 1666464484
transform -1 0 14976 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5650
timestamp 1666464484
transform -1 0 14976 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5651
timestamp 1666464484
transform -1 0 14976 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5652
timestamp 1666464484
transform -1 0 14976 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5653
timestamp 1666464484
transform -1 0 14976 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5654
timestamp 1666464484
transform -1 0 14976 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5655
timestamp 1666464484
transform -1 0 14976 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5656
timestamp 1666464484
transform -1 0 14976 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5657
timestamp 1666464484
transform -1 0 14976 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5658
timestamp 1666464484
transform -1 0 14976 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5659
timestamp 1666464484
transform -1 0 14976 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5660
timestamp 1666464484
transform -1 0 14976 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5661
timestamp 1666464484
transform -1 0 14976 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5662
timestamp 1666464484
transform -1 0 14976 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5663
timestamp 1666464484
transform -1 0 14976 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5664
timestamp 1666464484
transform -1 0 14976 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5665
timestamp 1666464484
transform 1 0 13728 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5666
timestamp 1666464484
transform 1 0 13728 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5667
timestamp 1666464484
transform -1 0 13728 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5668
timestamp 1666464484
transform -1 0 13728 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5669
timestamp 1666464484
transform 1 0 12480 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5670
timestamp 1666464484
transform 1 0 12480 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5671
timestamp 1666464484
transform -1 0 12480 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5672
timestamp 1666464484
transform -1 0 12480 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5673
timestamp 1666464484
transform 1 0 11232 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5674
timestamp 1666464484
transform 1 0 11232 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5675
timestamp 1666464484
transform -1 0 3744 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5676
timestamp 1666464484
transform -1 0 3744 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5677
timestamp 1666464484
transform 1 0 2496 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5678
timestamp 1666464484
transform 1 0 2496 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5679
timestamp 1666464484
transform -1 0 2496 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5680
timestamp 1666464484
transform -1 0 2496 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5681
timestamp 1666464484
transform 1 0 1248 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5682
timestamp 1666464484
transform 1 0 1248 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5683
timestamp 1666464484
transform -1 0 1248 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5684
timestamp 1666464484
transform -1 0 1248 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5685
timestamp 1666464484
transform 1 0 18720 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5686
timestamp 1666464484
transform 1 0 18720 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5687
timestamp 1666464484
transform -1 0 18720 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5688
timestamp 1666464484
transform -1 0 18720 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5689
timestamp 1666464484
transform 1 0 17472 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5690
timestamp 1666464484
transform 1 0 17472 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5691
timestamp 1666464484
transform -1 0 17472 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5692
timestamp 1666464484
transform -1 0 17472 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5693
timestamp 1666464484
transform 1 0 16224 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5694
timestamp 1666464484
transform 1 0 16224 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5695
timestamp 1666464484
transform -1 0 16224 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5696
timestamp 1666464484
transform -1 0 16224 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5697
timestamp 1666464484
transform 1 0 14976 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5698
timestamp 1666464484
transform 1 0 14976 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5699
timestamp 1666464484
transform -1 0 14976 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5700
timestamp 1666464484
transform -1 0 14976 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5701
timestamp 1666464484
transform 1 0 13728 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5702
timestamp 1666464484
transform 1 0 13728 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5703
timestamp 1666464484
transform -1 0 13728 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5704
timestamp 1666464484
transform -1 0 13728 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5705
timestamp 1666464484
transform 1 0 12480 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5706
timestamp 1666464484
transform 1 0 12480 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5707
timestamp 1666464484
transform -1 0 12480 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5708
timestamp 1666464484
transform -1 0 12480 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5709
timestamp 1666464484
transform 1 0 11232 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5710
timestamp 1666464484
transform 1 0 11232 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5711
timestamp 1666464484
transform -1 0 11232 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5712
timestamp 1666464484
transform -1 0 11232 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5713
timestamp 1666464484
transform 1 0 9984 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5714
timestamp 1666464484
transform 1 0 9984 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5715
timestamp 1666464484
transform 1 0 9984 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5716
timestamp 1666464484
transform 1 0 9984 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5717
timestamp 1666464484
transform 1 0 9984 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5718
timestamp 1666464484
transform 1 0 9984 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5719
timestamp 1666464484
transform 1 0 9984 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5720
timestamp 1666464484
transform 1 0 9984 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5721
timestamp 1666464484
transform 1 0 9984 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5722
timestamp 1666464484
transform 1 0 9984 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5723
timestamp 1666464484
transform 1 0 9984 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5724
timestamp 1666464484
transform 1 0 9984 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5725
timestamp 1666464484
transform 1 0 9984 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5726
timestamp 1666464484
transform 1 0 9984 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5727
timestamp 1666464484
transform 1 0 9984 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5728
timestamp 1666464484
transform 1 0 9984 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5729
timestamp 1666464484
transform 1 0 9984 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5730
timestamp 1666464484
transform 1 0 9984 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5731
timestamp 1666464484
transform 1 0 9984 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5732
timestamp 1666464484
transform 1 0 9984 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5733
timestamp 1666464484
transform 1 0 9984 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5734
timestamp 1666464484
transform 1 0 9984 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5735
timestamp 1666464484
transform 1 0 9984 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5736
timestamp 1666464484
transform 1 0 9984 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5737
timestamp 1666464484
transform 1 0 9984 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5738
timestamp 1666464484
transform 1 0 9984 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5739
timestamp 1666464484
transform 1 0 9984 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5740
timestamp 1666464484
transform 1 0 9984 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5741
timestamp 1666464484
transform 1 0 9984 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5742
timestamp 1666464484
transform 1 0 9984 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5743
timestamp 1666464484
transform 1 0 9984 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5744
timestamp 1666464484
transform 1 0 9984 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5745
timestamp 1666464484
transform 1 0 9984 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5746
timestamp 1666464484
transform 1 0 9984 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5747
timestamp 1666464484
transform 1 0 9984 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5748
timestamp 1666464484
transform 1 0 9984 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5749
timestamp 1666464484
transform 1 0 9984 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5750
timestamp 1666464484
transform 1 0 9984 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5751
timestamp 1666464484
transform 1 0 9984 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5752
timestamp 1666464484
transform 1 0 9984 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5753
timestamp 1666464484
transform 1 0 9984 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5754
timestamp 1666464484
transform 1 0 9984 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5755
timestamp 1666464484
transform 1 0 9984 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5756
timestamp 1666464484
transform 1 0 9984 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5757
timestamp 1666464484
transform 1 0 9984 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5758
timestamp 1666464484
transform 1 0 9984 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5759
timestamp 1666464484
transform 1 0 9984 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5760
timestamp 1666464484
transform 1 0 9984 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5761
timestamp 1666464484
transform 1 0 9984 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5762
timestamp 1666464484
transform 1 0 9984 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5763
timestamp 1666464484
transform 1 0 9984 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5764
timestamp 1666464484
transform 1 0 9984 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5765
timestamp 1666464484
transform 1 0 9984 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5766
timestamp 1666464484
transform 1 0 9984 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5767
timestamp 1666464484
transform 1 0 9984 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5768
timestamp 1666464484
transform 1 0 9984 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5769
timestamp 1666464484
transform 1 0 9984 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5770
timestamp 1666464484
transform 1 0 9984 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5771
timestamp 1666464484
transform 1 0 9984 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5772
timestamp 1666464484
transform 1 0 9984 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5773
timestamp 1666464484
transform 1 0 9984 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5774
timestamp 1666464484
transform 1 0 9984 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5775
timestamp 1666464484
transform 1 0 9984 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5776
timestamp 1666464484
transform 1 0 0 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5777
timestamp 1666464484
transform 1 0 0 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5778
timestamp 1666464484
transform -1 0 9984 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5779
timestamp 1666464484
transform -1 0 9984 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5780
timestamp 1666464484
transform -1 0 9984 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5781
timestamp 1666464484
transform -1 0 9984 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5782
timestamp 1666464484
transform -1 0 9984 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5783
timestamp 1666464484
transform -1 0 9984 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5784
timestamp 1666464484
transform -1 0 9984 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5785
timestamp 1666464484
transform -1 0 9984 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5786
timestamp 1666464484
transform -1 0 9984 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5787
timestamp 1666464484
transform -1 0 9984 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5788
timestamp 1666464484
transform -1 0 9984 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5789
timestamp 1666464484
transform -1 0 9984 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5790
timestamp 1666464484
transform -1 0 9984 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5791
timestamp 1666464484
transform -1 0 9984 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5792
timestamp 1666464484
transform -1 0 9984 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5793
timestamp 1666464484
transform -1 0 9984 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5794
timestamp 1666464484
transform -1 0 9984 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5795
timestamp 1666464484
transform -1 0 9984 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5796
timestamp 1666464484
transform -1 0 9984 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5797
timestamp 1666464484
transform -1 0 9984 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5798
timestamp 1666464484
transform -1 0 9984 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5799
timestamp 1666464484
transform -1 0 9984 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5800
timestamp 1666464484
transform -1 0 9984 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5801
timestamp 1666464484
transform -1 0 9984 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5802
timestamp 1666464484
transform -1 0 9984 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5803
timestamp 1666464484
transform -1 0 9984 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5804
timestamp 1666464484
transform -1 0 9984 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5805
timestamp 1666464484
transform -1 0 9984 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5806
timestamp 1666464484
transform -1 0 9984 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5807
timestamp 1666464484
transform -1 0 9984 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5808
timestamp 1666464484
transform -1 0 9984 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5809
timestamp 1666464484
transform -1 0 9984 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5810
timestamp 1666464484
transform -1 0 9984 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5811
timestamp 1666464484
transform -1 0 9984 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5812
timestamp 1666464484
transform -1 0 9984 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5813
timestamp 1666464484
transform -1 0 9984 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5814
timestamp 1666464484
transform -1 0 9984 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5815
timestamp 1666464484
transform -1 0 9984 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5816
timestamp 1666464484
transform -1 0 9984 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5817
timestamp 1666464484
transform -1 0 9984 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5818
timestamp 1666464484
transform -1 0 9984 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5819
timestamp 1666464484
transform -1 0 9984 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5820
timestamp 1666464484
transform -1 0 9984 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5821
timestamp 1666464484
transform -1 0 9984 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5822
timestamp 1666464484
transform -1 0 9984 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5823
timestamp 1666464484
transform -1 0 9984 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5824
timestamp 1666464484
transform -1 0 9984 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5825
timestamp 1666464484
transform -1 0 9984 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5826
timestamp 1666464484
transform -1 0 9984 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5827
timestamp 1666464484
transform -1 0 9984 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5828
timestamp 1666464484
transform -1 0 9984 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5829
timestamp 1666464484
transform -1 0 9984 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5830
timestamp 1666464484
transform -1 0 9984 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5831
timestamp 1666464484
transform -1 0 9984 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5832
timestamp 1666464484
transform -1 0 9984 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5833
timestamp 1666464484
transform -1 0 9984 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5834
timestamp 1666464484
transform -1 0 9984 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5835
timestamp 1666464484
transform -1 0 9984 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5836
timestamp 1666464484
transform -1 0 9984 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5837
timestamp 1666464484
transform -1 0 9984 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5838
timestamp 1666464484
transform -1 0 9984 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5839
timestamp 1666464484
transform -1 0 9984 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5840
timestamp 1666464484
transform -1 0 9984 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5841
timestamp 1666464484
transform 1 0 8736 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5842
timestamp 1666464484
transform 1 0 8736 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5843
timestamp 1666464484
transform -1 0 8736 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5844
timestamp 1666464484
transform -1 0 8736 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5845
timestamp 1666464484
transform 1 0 7488 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5846
timestamp 1666464484
transform 1 0 7488 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5847
timestamp 1666464484
transform -1 0 7488 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5848
timestamp 1666464484
transform -1 0 7488 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5849
timestamp 1666464484
transform 1 0 6240 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5850
timestamp 1666464484
transform 1 0 6240 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5851
timestamp 1666464484
transform -1 0 6240 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5852
timestamp 1666464484
transform -1 0 6240 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5853
timestamp 1666464484
transform 1 0 4992 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5854
timestamp 1666464484
transform 1 0 4992 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5855
timestamp 1666464484
transform -1 0 4992 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5856
timestamp 1666464484
transform -1 0 4992 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5857
timestamp 1666464484
transform 1 0 3744 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5858
timestamp 1666464484
transform 1 0 3744 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5859
timestamp 1666464484
transform -1 0 36192 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5860
timestamp 1666464484
transform -1 0 36192 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5861
timestamp 1666464484
transform -1 0 36192 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5862
timestamp 1666464484
transform -1 0 38688 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5863
timestamp 1666464484
transform -1 0 38688 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5864
timestamp 1666464484
transform -1 0 38688 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5865
timestamp 1666464484
transform -1 0 38688 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5866
timestamp 1666464484
transform -1 0 38688 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5867
timestamp 1666464484
transform -1 0 38688 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5868
timestamp 1666464484
transform -1 0 38688 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5869
timestamp 1666464484
transform -1 0 38688 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5870
timestamp 1666464484
transform -1 0 38688 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5871
timestamp 1666464484
transform -1 0 38688 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5872
timestamp 1666464484
transform -1 0 38688 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5873
timestamp 1666464484
transform -1 0 38688 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5874
timestamp 1666464484
transform -1 0 38688 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5875
timestamp 1666464484
transform -1 0 38688 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5876
timestamp 1666464484
transform 1 0 37440 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5877
timestamp 1666464484
transform 1 0 37440 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5878
timestamp 1666464484
transform 1 0 38688 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5879
timestamp 1666464484
transform 1 0 38688 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5880
timestamp 1666464484
transform 1 0 38688 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5881
timestamp 1666464484
transform 1 0 38688 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5882
timestamp 1666464484
transform 1 0 38688 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5883
timestamp 1666464484
transform 1 0 38688 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5884
timestamp 1666464484
transform 1 0 38688 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5885
timestamp 1666464484
transform 1 0 38688 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5886
timestamp 1666464484
transform 1 0 38688 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5887
timestamp 1666464484
transform 1 0 38688 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5888
timestamp 1666464484
transform 1 0 38688 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5889
timestamp 1666464484
transform 1 0 38688 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5890
timestamp 1666464484
transform 1 0 38688 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5891
timestamp 1666464484
transform 1 0 38688 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5892
timestamp 1666464484
transform 1 0 37440 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5893
timestamp 1666464484
transform 1 0 37440 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5894
timestamp 1666464484
transform 1 0 37440 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5895
timestamp 1666464484
transform 1 0 37440 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5896
timestamp 1666464484
transform 1 0 37440 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5897
timestamp 1666464484
transform 1 0 37440 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5898
timestamp 1666464484
transform 1 0 37440 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5899
timestamp 1666464484
transform 1 0 37440 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5900
timestamp 1666464484
transform 1 0 37440 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5901
timestamp 1666464484
transform 1 0 37440 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5902
timestamp 1666464484
transform 1 0 36192 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5903
timestamp 1666464484
transform 1 0 36192 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5904
timestamp 1666464484
transform -1 0 36192 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5905
timestamp 1666464484
transform -1 0 36192 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5906
timestamp 1666464484
transform -1 0 36192 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5907
timestamp 1666464484
transform -1 0 36192 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5908
timestamp 1666464484
transform -1 0 39936 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5909
timestamp 1666464484
transform -1 0 39936 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5910
timestamp 1666464484
transform -1 0 39936 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5911
timestamp 1666464484
transform -1 0 39936 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5912
timestamp 1666464484
transform -1 0 39936 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5913
timestamp 1666464484
transform -1 0 39936 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5914
timestamp 1666464484
transform -1 0 39936 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5915
timestamp 1666464484
transform -1 0 39936 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5916
timestamp 1666464484
transform -1 0 39936 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5917
timestamp 1666464484
transform -1 0 39936 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5918
timestamp 1666464484
transform -1 0 39936 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5919
timestamp 1666464484
transform -1 0 39936 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5920
timestamp 1666464484
transform -1 0 39936 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5921
timestamp 1666464484
transform -1 0 39936 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5922
timestamp 1666464484
transform -1 0 36192 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5923
timestamp 1666464484
transform -1 0 36192 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5924
timestamp 1666464484
transform -1 0 36192 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5925
timestamp 1666464484
transform -1 0 36192 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5926
timestamp 1666464484
transform -1 0 36192 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5927
timestamp 1666464484
transform -1 0 36192 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5928
timestamp 1666464484
transform -1 0 37440 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5929
timestamp 1666464484
transform -1 0 37440 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5930
timestamp 1666464484
transform -1 0 37440 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5931
timestamp 1666464484
transform -1 0 37440 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5932
timestamp 1666464484
transform -1 0 37440 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5933
timestamp 1666464484
transform -1 0 37440 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5934
timestamp 1666464484
transform -1 0 37440 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5935
timestamp 1666464484
transform -1 0 37440 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5936
timestamp 1666464484
transform -1 0 37440 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5937
timestamp 1666464484
transform -1 0 37440 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5938
timestamp 1666464484
transform -1 0 37440 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5939
timestamp 1666464484
transform -1 0 37440 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5940
timestamp 1666464484
transform -1 0 37440 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5941
timestamp 1666464484
transform -1 0 37440 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5942
timestamp 1666464484
transform -1 0 36192 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5943
timestamp 1666464484
transform 1 0 36192 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5944
timestamp 1666464484
transform 1 0 36192 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5945
timestamp 1666464484
transform 1 0 36192 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5946
timestamp 1666464484
transform 1 0 36192 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5947
timestamp 1666464484
transform 1 0 36192 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5948
timestamp 1666464484
transform 1 0 36192 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5949
timestamp 1666464484
transform 1 0 36192 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5950
timestamp 1666464484
transform 1 0 36192 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5951
timestamp 1666464484
transform 1 0 36192 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5952
timestamp 1666464484
transform 1 0 36192 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5953
timestamp 1666464484
transform 1 0 36192 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5954
timestamp 1666464484
transform 1 0 36192 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5955
timestamp 1666464484
transform 1 0 37440 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5956
timestamp 1666464484
transform 1 0 37440 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5957
timestamp 1666464484
transform 1 0 33696 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5958
timestamp 1666464484
transform 1 0 33696 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5959
timestamp 1666464484
transform 1 0 33696 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5960
timestamp 1666464484
transform 1 0 33696 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5961
timestamp 1666464484
transform 1 0 33696 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5962
timestamp 1666464484
transform 1 0 33696 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5963
timestamp 1666464484
transform -1 0 33696 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5964
timestamp 1666464484
transform -1 0 33696 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5965
timestamp 1666464484
transform -1 0 33696 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5966
timestamp 1666464484
transform -1 0 33696 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5967
timestamp 1666464484
transform -1 0 33696 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5968
timestamp 1666464484
transform -1 0 33696 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5969
timestamp 1666464484
transform -1 0 33696 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5970
timestamp 1666464484
transform -1 0 33696 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5971
timestamp 1666464484
transform -1 0 33696 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5972
timestamp 1666464484
transform -1 0 33696 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5973
timestamp 1666464484
transform -1 0 33696 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5974
timestamp 1666464484
transform -1 0 33696 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5975
timestamp 1666464484
transform -1 0 33696 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5976
timestamp 1666464484
transform -1 0 33696 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5977
timestamp 1666464484
transform -1 0 32448 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5978
timestamp 1666464484
transform -1 0 32448 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5979
timestamp 1666464484
transform -1 0 32448 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5980
timestamp 1666464484
transform -1 0 32448 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5981
timestamp 1666464484
transform -1 0 32448 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5982
timestamp 1666464484
transform -1 0 32448 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5983
timestamp 1666464484
transform -1 0 32448 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5984
timestamp 1666464484
transform -1 0 32448 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5985
timestamp 1666464484
transform -1 0 32448 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5986
timestamp 1666464484
transform -1 0 32448 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5987
timestamp 1666464484
transform 1 0 33696 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5988
timestamp 1666464484
transform 1 0 33696 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5989
timestamp 1666464484
transform 1 0 33696 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5990
timestamp 1666464484
transform 1 0 33696 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5991
timestamp 1666464484
transform 1 0 32448 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5992
timestamp 1666464484
transform 1 0 32448 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5993
timestamp 1666464484
transform 1 0 32448 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5994
timestamp 1666464484
transform -1 0 31200 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5995
timestamp 1666464484
transform -1 0 31200 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5996
timestamp 1666464484
transform -1 0 31200 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5997
timestamp 1666464484
transform -1 0 31200 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5998
timestamp 1666464484
transform -1 0 31200 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_5999
timestamp 1666464484
transform 1 0 32448 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6000
timestamp 1666464484
transform 1 0 32448 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6001
timestamp 1666464484
transform 1 0 32448 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6002
timestamp 1666464484
transform 1 0 32448 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6003
timestamp 1666464484
transform 1 0 31200 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6004
timestamp 1666464484
transform 1 0 31200 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6005
timestamp 1666464484
transform 1 0 31200 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6006
timestamp 1666464484
transform 1 0 31200 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6007
timestamp 1666464484
transform 1 0 31200 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6008
timestamp 1666464484
transform 1 0 32448 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6009
timestamp 1666464484
transform 1 0 32448 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6010
timestamp 1666464484
transform 1 0 32448 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6011
timestamp 1666464484
transform 1 0 33696 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6012
timestamp 1666464484
transform -1 0 31200 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6013
timestamp 1666464484
transform -1 0 31200 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6014
timestamp 1666464484
transform -1 0 31200 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6015
timestamp 1666464484
transform -1 0 31200 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6016
timestamp 1666464484
transform -1 0 31200 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6017
timestamp 1666464484
transform -1 0 31200 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6018
timestamp 1666464484
transform -1 0 31200 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6019
timestamp 1666464484
transform -1 0 31200 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6020
timestamp 1666464484
transform -1 0 31200 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6021
timestamp 1666464484
transform 1 0 33696 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6022
timestamp 1666464484
transform 1 0 33696 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6023
timestamp 1666464484
transform -1 0 32448 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6024
timestamp 1666464484
transform -1 0 32448 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6025
timestamp 1666464484
transform -1 0 32448 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6026
timestamp 1666464484
transform -1 0 32448 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6027
timestamp 1666464484
transform 1 0 31200 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6028
timestamp 1666464484
transform 1 0 31200 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6029
timestamp 1666464484
transform 1 0 31200 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6030
timestamp 1666464484
transform 1 0 31200 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6031
timestamp 1666464484
transform 1 0 32448 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6032
timestamp 1666464484
transform 1 0 32448 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6033
timestamp 1666464484
transform 1 0 32448 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6034
timestamp 1666464484
transform 1 0 32448 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6035
timestamp 1666464484
transform 1 0 31200 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6036
timestamp 1666464484
transform 1 0 31200 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6037
timestamp 1666464484
transform 1 0 31200 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6038
timestamp 1666464484
transform 1 0 31200 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6039
timestamp 1666464484
transform 1 0 31200 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6040
timestamp 1666464484
transform 1 0 33696 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6041
timestamp 1666464484
transform -1 0 33696 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6042
timestamp 1666464484
transform -1 0 33696 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6043
timestamp 1666464484
transform -1 0 33696 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6044
timestamp 1666464484
transform -1 0 33696 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6045
timestamp 1666464484
transform 1 0 32448 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6046
timestamp 1666464484
transform 1 0 32448 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6047
timestamp 1666464484
transform 1 0 32448 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6048
timestamp 1666464484
transform 1 0 32448 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6049
timestamp 1666464484
transform 1 0 32448 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6050
timestamp 1666464484
transform 1 0 32448 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6051
timestamp 1666464484
transform 1 0 32448 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6052
timestamp 1666464484
transform 1 0 32448 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6053
timestamp 1666464484
transform 1 0 32448 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6054
timestamp 1666464484
transform 1 0 32448 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6055
timestamp 1666464484
transform 1 0 32448 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6056
timestamp 1666464484
transform 1 0 32448 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6057
timestamp 1666464484
transform 1 0 32448 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6058
timestamp 1666464484
transform 1 0 33696 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6059
timestamp 1666464484
transform -1 0 32448 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6060
timestamp 1666464484
transform -1 0 32448 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6061
timestamp 1666464484
transform 1 0 31200 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6062
timestamp 1666464484
transform 1 0 31200 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6063
timestamp 1666464484
transform 1 0 31200 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6064
timestamp 1666464484
transform 1 0 31200 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6065
timestamp 1666464484
transform -1 0 32448 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6066
timestamp 1666464484
transform -1 0 32448 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6067
timestamp 1666464484
transform -1 0 32448 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6068
timestamp 1666464484
transform -1 0 32448 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6069
timestamp 1666464484
transform -1 0 32448 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6070
timestamp 1666464484
transform -1 0 32448 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6071
timestamp 1666464484
transform 1 0 31200 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6072
timestamp 1666464484
transform 1 0 31200 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6073
timestamp 1666464484
transform 1 0 31200 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6074
timestamp 1666464484
transform 1 0 31200 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6075
timestamp 1666464484
transform 1 0 31200 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6076
timestamp 1666464484
transform 1 0 31200 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6077
timestamp 1666464484
transform 1 0 31200 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6078
timestamp 1666464484
transform 1 0 31200 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6079
timestamp 1666464484
transform 1 0 31200 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6080
timestamp 1666464484
transform 1 0 31200 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6081
timestamp 1666464484
transform 1 0 33696 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6082
timestamp 1666464484
transform 1 0 33696 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6083
timestamp 1666464484
transform 1 0 33696 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6084
timestamp 1666464484
transform 1 0 33696 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6085
timestamp 1666464484
transform 1 0 33696 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6086
timestamp 1666464484
transform -1 0 32448 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6087
timestamp 1666464484
transform -1 0 32448 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6088
timestamp 1666464484
transform -1 0 33696 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6089
timestamp 1666464484
transform -1 0 33696 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6090
timestamp 1666464484
transform -1 0 33696 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6091
timestamp 1666464484
transform -1 0 33696 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6092
timestamp 1666464484
transform -1 0 33696 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6093
timestamp 1666464484
transform -1 0 33696 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6094
timestamp 1666464484
transform -1 0 33696 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6095
timestamp 1666464484
transform -1 0 33696 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6096
timestamp 1666464484
transform -1 0 33696 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6097
timestamp 1666464484
transform -1 0 33696 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6098
timestamp 1666464484
transform -1 0 32448 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6099
timestamp 1666464484
transform -1 0 32448 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6100
timestamp 1666464484
transform -1 0 32448 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6101
timestamp 1666464484
transform -1 0 32448 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6102
timestamp 1666464484
transform 1 0 33696 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6103
timestamp 1666464484
transform 1 0 33696 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6104
timestamp 1666464484
transform 1 0 33696 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6105
timestamp 1666464484
transform 1 0 33696 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6106
timestamp 1666464484
transform 1 0 33696 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6107
timestamp 1666464484
transform 1 0 33696 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6108
timestamp 1666464484
transform 1 0 33696 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6109
timestamp 1666464484
transform -1 0 31200 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6110
timestamp 1666464484
transform -1 0 31200 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6111
timestamp 1666464484
transform -1 0 31200 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6112
timestamp 1666464484
transform -1 0 31200 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6113
timestamp 1666464484
transform -1 0 31200 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6114
timestamp 1666464484
transform -1 0 31200 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6115
timestamp 1666464484
transform -1 0 31200 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6116
timestamp 1666464484
transform -1 0 31200 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6117
timestamp 1666464484
transform -1 0 31200 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6118
timestamp 1666464484
transform -1 0 31200 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6119
timestamp 1666464484
transform -1 0 31200 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6120
timestamp 1666464484
transform -1 0 31200 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6121
timestamp 1666464484
transform -1 0 31200 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6122
timestamp 1666464484
transform -1 0 31200 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6123
timestamp 1666464484
transform 1 0 33696 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6124
timestamp 1666464484
transform 1 0 32448 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6125
timestamp 1666464484
transform 1 0 36192 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6126
timestamp 1666464484
transform 1 0 36192 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6127
timestamp 1666464484
transform -1 0 39936 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6128
timestamp 1666464484
transform -1 0 39936 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6129
timestamp 1666464484
transform -1 0 39936 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6130
timestamp 1666464484
transform -1 0 39936 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6131
timestamp 1666464484
transform -1 0 39936 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6132
timestamp 1666464484
transform -1 0 39936 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6133
timestamp 1666464484
transform -1 0 39936 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6134
timestamp 1666464484
transform -1 0 39936 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6135
timestamp 1666464484
transform -1 0 39936 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6136
timestamp 1666464484
transform -1 0 39936 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6137
timestamp 1666464484
transform -1 0 39936 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6138
timestamp 1666464484
transform -1 0 39936 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6139
timestamp 1666464484
transform -1 0 39936 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6140
timestamp 1666464484
transform -1 0 39936 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6141
timestamp 1666464484
transform 1 0 36192 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6142
timestamp 1666464484
transform 1 0 36192 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6143
timestamp 1666464484
transform 1 0 36192 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6144
timestamp 1666464484
transform 1 0 36192 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6145
timestamp 1666464484
transform 1 0 36192 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6146
timestamp 1666464484
transform 1 0 36192 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6147
timestamp 1666464484
transform 1 0 36192 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6148
timestamp 1666464484
transform 1 0 36192 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6149
timestamp 1666464484
transform -1 0 36192 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6150
timestamp 1666464484
transform -1 0 36192 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6151
timestamp 1666464484
transform -1 0 36192 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6152
timestamp 1666464484
transform -1 0 36192 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6153
timestamp 1666464484
transform -1 0 36192 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6154
timestamp 1666464484
transform 1 0 37440 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6155
timestamp 1666464484
transform 1 0 37440 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6156
timestamp 1666464484
transform 1 0 37440 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6157
timestamp 1666464484
transform 1 0 37440 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6158
timestamp 1666464484
transform 1 0 37440 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6159
timestamp 1666464484
transform 1 0 37440 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6160
timestamp 1666464484
transform 1 0 37440 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6161
timestamp 1666464484
transform 1 0 37440 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6162
timestamp 1666464484
transform 1 0 37440 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6163
timestamp 1666464484
transform 1 0 37440 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6164
timestamp 1666464484
transform 1 0 37440 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6165
timestamp 1666464484
transform 1 0 37440 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6166
timestamp 1666464484
transform 1 0 37440 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6167
timestamp 1666464484
transform 1 0 37440 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6168
timestamp 1666464484
transform -1 0 36192 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6169
timestamp 1666464484
transform -1 0 36192 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6170
timestamp 1666464484
transform -1 0 36192 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6171
timestamp 1666464484
transform -1 0 37440 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6172
timestamp 1666464484
transform -1 0 37440 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6173
timestamp 1666464484
transform 1 0 38688 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6174
timestamp 1666464484
transform 1 0 38688 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6175
timestamp 1666464484
transform 1 0 38688 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6176
timestamp 1666464484
transform 1 0 38688 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6177
timestamp 1666464484
transform 1 0 38688 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6178
timestamp 1666464484
transform 1 0 38688 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6179
timestamp 1666464484
transform 1 0 38688 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6180
timestamp 1666464484
transform 1 0 38688 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6181
timestamp 1666464484
transform 1 0 38688 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6182
timestamp 1666464484
transform 1 0 38688 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6183
timestamp 1666464484
transform 1 0 38688 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6184
timestamp 1666464484
transform 1 0 38688 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6185
timestamp 1666464484
transform 1 0 38688 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6186
timestamp 1666464484
transform 1 0 38688 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6187
timestamp 1666464484
transform -1 0 37440 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6188
timestamp 1666464484
transform -1 0 37440 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6189
timestamp 1666464484
transform -1 0 37440 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6190
timestamp 1666464484
transform -1 0 37440 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6191
timestamp 1666464484
transform -1 0 38688 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6192
timestamp 1666464484
transform -1 0 38688 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6193
timestamp 1666464484
transform -1 0 38688 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6194
timestamp 1666464484
transform -1 0 38688 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6195
timestamp 1666464484
transform -1 0 38688 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6196
timestamp 1666464484
transform -1 0 38688 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6197
timestamp 1666464484
transform -1 0 38688 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6198
timestamp 1666464484
transform -1 0 38688 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6199
timestamp 1666464484
transform -1 0 38688 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6200
timestamp 1666464484
transform -1 0 38688 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6201
timestamp 1666464484
transform -1 0 38688 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6202
timestamp 1666464484
transform -1 0 38688 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6203
timestamp 1666464484
transform -1 0 38688 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6204
timestamp 1666464484
transform -1 0 38688 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6205
timestamp 1666464484
transform -1 0 37440 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6206
timestamp 1666464484
transform -1 0 37440 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6207
timestamp 1666464484
transform -1 0 37440 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6208
timestamp 1666464484
transform -1 0 37440 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6209
timestamp 1666464484
transform -1 0 37440 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6210
timestamp 1666464484
transform -1 0 37440 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6211
timestamp 1666464484
transform -1 0 37440 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6212
timestamp 1666464484
transform -1 0 37440 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6213
timestamp 1666464484
transform -1 0 36192 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6214
timestamp 1666464484
transform -1 0 36192 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6215
timestamp 1666464484
transform -1 0 36192 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6216
timestamp 1666464484
transform -1 0 36192 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6217
timestamp 1666464484
transform -1 0 36192 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6218
timestamp 1666464484
transform -1 0 36192 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6219
timestamp 1666464484
transform 1 0 36192 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6220
timestamp 1666464484
transform 1 0 36192 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6221
timestamp 1666464484
transform 1 0 36192 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6222
timestamp 1666464484
transform 1 0 36192 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6223
timestamp 1666464484
transform -1 0 33696 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6224
timestamp 1666464484
transform -1 0 33696 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6225
timestamp 1666464484
transform -1 0 39936 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6226
timestamp 1666464484
transform -1 0 39936 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6227
timestamp 1666464484
transform 1 0 34944 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6228
timestamp 1666464484
transform 1 0 34944 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6229
timestamp 1666464484
transform 1 0 34944 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6230
timestamp 1666464484
transform 1 0 34944 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6231
timestamp 1666464484
transform 1 0 34944 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6232
timestamp 1666464484
transform 1 0 34944 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6233
timestamp 1666464484
transform 1 0 34944 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6234
timestamp 1666464484
transform 1 0 34944 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6235
timestamp 1666464484
transform 1 0 34944 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6236
timestamp 1666464484
transform 1 0 34944 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6237
timestamp 1666464484
transform 1 0 34944 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6238
timestamp 1666464484
transform 1 0 34944 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6239
timestamp 1666464484
transform 1 0 34944 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6240
timestamp 1666464484
transform 1 0 34944 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6241
timestamp 1666464484
transform 1 0 34944 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6242
timestamp 1666464484
transform 1 0 34944 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6243
timestamp 1666464484
transform 1 0 34944 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6244
timestamp 1666464484
transform 1 0 34944 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6245
timestamp 1666464484
transform 1 0 34944 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6246
timestamp 1666464484
transform 1 0 34944 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6247
timestamp 1666464484
transform 1 0 34944 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6248
timestamp 1666464484
transform 1 0 34944 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6249
timestamp 1666464484
transform 1 0 34944 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6250
timestamp 1666464484
transform 1 0 34944 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6251
timestamp 1666464484
transform 1 0 34944 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6252
timestamp 1666464484
transform 1 0 34944 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6253
timestamp 1666464484
transform 1 0 34944 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6254
timestamp 1666464484
transform 1 0 34944 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6255
timestamp 1666464484
transform 1 0 34944 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6256
timestamp 1666464484
transform 1 0 34944 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6257
timestamp 1666464484
transform 1 0 38688 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6258
timestamp 1666464484
transform 1 0 38688 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6259
timestamp 1666464484
transform -1 0 31200 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6260
timestamp 1666464484
transform 1 0 32448 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6261
timestamp 1666464484
transform -1 0 38688 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6262
timestamp 1666464484
transform -1 0 38688 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6263
timestamp 1666464484
transform -1 0 34944 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6264
timestamp 1666464484
transform -1 0 34944 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6265
timestamp 1666464484
transform -1 0 34944 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6266
timestamp 1666464484
transform -1 0 34944 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6267
timestamp 1666464484
transform -1 0 34944 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6268
timestamp 1666464484
transform -1 0 34944 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6269
timestamp 1666464484
transform -1 0 34944 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6270
timestamp 1666464484
transform -1 0 34944 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6271
timestamp 1666464484
transform -1 0 34944 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6272
timestamp 1666464484
transform -1 0 34944 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6273
timestamp 1666464484
transform -1 0 34944 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6274
timestamp 1666464484
transform -1 0 34944 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6275
timestamp 1666464484
transform -1 0 34944 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6276
timestamp 1666464484
transform -1 0 34944 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6277
timestamp 1666464484
transform -1 0 34944 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6278
timestamp 1666464484
transform -1 0 34944 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6279
timestamp 1666464484
transform -1 0 34944 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6280
timestamp 1666464484
transform -1 0 34944 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6281
timestamp 1666464484
transform -1 0 34944 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6282
timestamp 1666464484
transform -1 0 34944 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6283
timestamp 1666464484
transform -1 0 34944 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6284
timestamp 1666464484
transform -1 0 34944 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6285
timestamp 1666464484
transform -1 0 34944 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6286
timestamp 1666464484
transform -1 0 34944 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6287
timestamp 1666464484
transform -1 0 34944 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6288
timestamp 1666464484
transform -1 0 34944 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6289
timestamp 1666464484
transform -1 0 34944 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6290
timestamp 1666464484
transform -1 0 34944 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6291
timestamp 1666464484
transform -1 0 34944 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6292
timestamp 1666464484
transform -1 0 34944 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6293
timestamp 1666464484
transform 1 0 32448 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6294
timestamp 1666464484
transform 1 0 37440 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6295
timestamp 1666464484
transform 1 0 37440 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6296
timestamp 1666464484
transform -1 0 31200 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6297
timestamp 1666464484
transform -1 0 37440 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6298
timestamp 1666464484
transform -1 0 37440 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6299
timestamp 1666464484
transform 1 0 33696 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6300
timestamp 1666464484
transform 1 0 33696 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6301
timestamp 1666464484
transform 1 0 31200 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6302
timestamp 1666464484
transform 1 0 31200 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6303
timestamp 1666464484
transform 1 0 36192 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6304
timestamp 1666464484
transform 1 0 36192 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6305
timestamp 1666464484
transform -1 0 32448 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6306
timestamp 1666464484
transform -1 0 32448 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6307
timestamp 1666464484
transform -1 0 36192 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6308
timestamp 1666464484
transform -1 0 36192 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6309
timestamp 1666464484
transform 1 0 27456 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6310
timestamp 1666464484
transform 1 0 27456 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6311
timestamp 1666464484
transform 1 0 27456 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6312
timestamp 1666464484
transform 1 0 27456 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6313
timestamp 1666464484
transform 1 0 27456 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6314
timestamp 1666464484
transform 1 0 27456 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6315
timestamp 1666464484
transform 1 0 27456 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6316
timestamp 1666464484
transform 1 0 27456 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6317
timestamp 1666464484
transform -1 0 26208 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6318
timestamp 1666464484
transform -1 0 26208 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6319
timestamp 1666464484
transform -1 0 26208 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6320
timestamp 1666464484
transform -1 0 26208 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6321
timestamp 1666464484
transform -1 0 26208 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6322
timestamp 1666464484
transform -1 0 26208 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6323
timestamp 1666464484
transform -1 0 26208 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6324
timestamp 1666464484
transform -1 0 26208 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6325
timestamp 1666464484
transform -1 0 26208 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6326
timestamp 1666464484
transform -1 0 26208 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6327
timestamp 1666464484
transform -1 0 26208 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6328
timestamp 1666464484
transform 1 0 27456 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6329
timestamp 1666464484
transform 1 0 27456 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6330
timestamp 1666464484
transform -1 0 28704 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6331
timestamp 1666464484
transform -1 0 28704 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6332
timestamp 1666464484
transform -1 0 28704 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6333
timestamp 1666464484
transform -1 0 28704 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6334
timestamp 1666464484
transform -1 0 28704 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6335
timestamp 1666464484
transform -1 0 28704 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6336
timestamp 1666464484
transform -1 0 28704 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6337
timestamp 1666464484
transform -1 0 28704 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6338
timestamp 1666464484
transform -1 0 28704 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6339
timestamp 1666464484
transform 1 0 28704 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6340
timestamp 1666464484
transform 1 0 28704 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6341
timestamp 1666464484
transform 1 0 28704 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6342
timestamp 1666464484
transform 1 0 28704 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6343
timestamp 1666464484
transform 1 0 28704 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6344
timestamp 1666464484
transform 1 0 28704 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6345
timestamp 1666464484
transform 1 0 28704 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6346
timestamp 1666464484
transform 1 0 28704 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6347
timestamp 1666464484
transform 1 0 28704 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6348
timestamp 1666464484
transform 1 0 28704 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6349
timestamp 1666464484
transform 1 0 28704 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6350
timestamp 1666464484
transform 1 0 28704 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6351
timestamp 1666464484
transform 1 0 28704 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6352
timestamp 1666464484
transform 1 0 28704 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6353
timestamp 1666464484
transform -1 0 28704 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6354
timestamp 1666464484
transform -1 0 28704 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6355
timestamp 1666464484
transform -1 0 28704 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6356
timestamp 1666464484
transform -1 0 28704 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6357
timestamp 1666464484
transform 1 0 26208 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6358
timestamp 1666464484
transform 1 0 26208 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6359
timestamp 1666464484
transform 1 0 26208 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6360
timestamp 1666464484
transform 1 0 26208 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6361
timestamp 1666464484
transform 1 0 26208 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6362
timestamp 1666464484
transform 1 0 26208 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6363
timestamp 1666464484
transform 1 0 26208 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6364
timestamp 1666464484
transform 1 0 26208 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6365
timestamp 1666464484
transform 1 0 26208 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6366
timestamp 1666464484
transform 1 0 26208 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6367
timestamp 1666464484
transform 1 0 26208 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6368
timestamp 1666464484
transform -1 0 27456 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6369
timestamp 1666464484
transform -1 0 27456 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6370
timestamp 1666464484
transform -1 0 27456 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6371
timestamp 1666464484
transform -1 0 27456 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6372
timestamp 1666464484
transform -1 0 27456 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6373
timestamp 1666464484
transform -1 0 27456 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6374
timestamp 1666464484
transform -1 0 27456 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6375
timestamp 1666464484
transform -1 0 27456 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6376
timestamp 1666464484
transform -1 0 27456 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6377
timestamp 1666464484
transform -1 0 27456 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6378
timestamp 1666464484
transform -1 0 27456 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6379
timestamp 1666464484
transform -1 0 27456 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6380
timestamp 1666464484
transform -1 0 27456 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6381
timestamp 1666464484
transform -1 0 27456 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6382
timestamp 1666464484
transform 1 0 26208 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6383
timestamp 1666464484
transform 1 0 26208 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6384
timestamp 1666464484
transform 1 0 26208 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6385
timestamp 1666464484
transform -1 0 28704 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6386
timestamp 1666464484
transform 1 0 27456 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6387
timestamp 1666464484
transform 1 0 27456 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6388
timestamp 1666464484
transform 1 0 27456 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6389
timestamp 1666464484
transform 1 0 27456 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6390
timestamp 1666464484
transform -1 0 26208 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6391
timestamp 1666464484
transform -1 0 26208 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6392
timestamp 1666464484
transform -1 0 26208 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6393
timestamp 1666464484
transform 1 0 23712 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6394
timestamp 1666464484
transform 1 0 23712 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6395
timestamp 1666464484
transform 1 0 21216 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6396
timestamp 1666464484
transform -1 0 21216 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6397
timestamp 1666464484
transform -1 0 23712 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6398
timestamp 1666464484
transform -1 0 21216 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6399
timestamp 1666464484
transform -1 0 21216 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6400
timestamp 1666464484
transform -1 0 22464 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6401
timestamp 1666464484
transform -1 0 22464 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6402
timestamp 1666464484
transform -1 0 21216 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6403
timestamp 1666464484
transform -1 0 23712 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6404
timestamp 1666464484
transform -1 0 23712 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6405
timestamp 1666464484
transform -1 0 23712 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6406
timestamp 1666464484
transform -1 0 23712 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6407
timestamp 1666464484
transform -1 0 23712 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6408
timestamp 1666464484
transform -1 0 22464 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6409
timestamp 1666464484
transform -1 0 22464 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6410
timestamp 1666464484
transform -1 0 23712 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6411
timestamp 1666464484
transform -1 0 23712 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6412
timestamp 1666464484
transform -1 0 23712 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6413
timestamp 1666464484
transform -1 0 23712 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6414
timestamp 1666464484
transform -1 0 23712 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6415
timestamp 1666464484
transform -1 0 23712 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6416
timestamp 1666464484
transform -1 0 23712 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6417
timestamp 1666464484
transform -1 0 22464 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6418
timestamp 1666464484
transform 1 0 23712 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6419
timestamp 1666464484
transform 1 0 22464 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6420
timestamp 1666464484
transform 1 0 22464 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6421
timestamp 1666464484
transform 1 0 22464 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6422
timestamp 1666464484
transform 1 0 22464 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6423
timestamp 1666464484
transform 1 0 22464 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6424
timestamp 1666464484
transform 1 0 22464 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6425
timestamp 1666464484
transform 1 0 22464 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6426
timestamp 1666464484
transform 1 0 22464 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6427
timestamp 1666464484
transform 1 0 22464 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6428
timestamp 1666464484
transform 1 0 23712 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6429
timestamp 1666464484
transform -1 0 21216 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6430
timestamp 1666464484
transform -1 0 21216 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6431
timestamp 1666464484
transform -1 0 21216 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6432
timestamp 1666464484
transform -1 0 21216 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6433
timestamp 1666464484
transform -1 0 21216 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6434
timestamp 1666464484
transform -1 0 21216 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6435
timestamp 1666464484
transform 1 0 21216 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6436
timestamp 1666464484
transform 1 0 21216 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6437
timestamp 1666464484
transform 1 0 21216 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6438
timestamp 1666464484
transform 1 0 21216 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6439
timestamp 1666464484
transform -1 0 22464 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6440
timestamp 1666464484
transform -1 0 22464 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6441
timestamp 1666464484
transform -1 0 22464 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6442
timestamp 1666464484
transform -1 0 22464 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6443
timestamp 1666464484
transform -1 0 22464 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6444
timestamp 1666464484
transform -1 0 22464 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6445
timestamp 1666464484
transform -1 0 22464 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6446
timestamp 1666464484
transform 1 0 22464 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6447
timestamp 1666464484
transform 1 0 22464 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6448
timestamp 1666464484
transform 1 0 22464 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6449
timestamp 1666464484
transform 1 0 22464 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6450
timestamp 1666464484
transform 1 0 22464 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6451
timestamp 1666464484
transform -1 0 22464 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6452
timestamp 1666464484
transform -1 0 22464 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6453
timestamp 1666464484
transform -1 0 21216 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6454
timestamp 1666464484
transform -1 0 21216 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6455
timestamp 1666464484
transform -1 0 23712 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6456
timestamp 1666464484
transform 1 0 21216 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6457
timestamp 1666464484
transform 1 0 21216 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6458
timestamp 1666464484
transform 1 0 21216 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6459
timestamp 1666464484
transform 1 0 21216 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6460
timestamp 1666464484
transform -1 0 21216 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6461
timestamp 1666464484
transform -1 0 21216 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6462
timestamp 1666464484
transform 1 0 21216 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6463
timestamp 1666464484
transform 1 0 21216 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6464
timestamp 1666464484
transform 1 0 21216 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6465
timestamp 1666464484
transform 1 0 21216 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6466
timestamp 1666464484
transform 1 0 21216 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6467
timestamp 1666464484
transform 1 0 23712 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6468
timestamp 1666464484
transform 1 0 23712 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6469
timestamp 1666464484
transform 1 0 23712 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6470
timestamp 1666464484
transform 1 0 23712 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6471
timestamp 1666464484
transform 1 0 23712 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6472
timestamp 1666464484
transform 1 0 23712 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6473
timestamp 1666464484
transform 1 0 23712 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6474
timestamp 1666464484
transform 1 0 23712 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6475
timestamp 1666464484
transform 1 0 23712 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6476
timestamp 1666464484
transform 1 0 23712 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6477
timestamp 1666464484
transform -1 0 21216 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6478
timestamp 1666464484
transform -1 0 21216 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6479
timestamp 1666464484
transform 1 0 21216 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6480
timestamp 1666464484
transform 1 0 21216 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6481
timestamp 1666464484
transform 1 0 21216 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6482
timestamp 1666464484
transform 1 0 22464 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6483
timestamp 1666464484
transform 1 0 22464 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6484
timestamp 1666464484
transform 1 0 22464 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6485
timestamp 1666464484
transform 1 0 22464 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6486
timestamp 1666464484
transform 1 0 22464 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6487
timestamp 1666464484
transform 1 0 22464 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6488
timestamp 1666464484
transform 1 0 22464 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6489
timestamp 1666464484
transform 1 0 22464 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6490
timestamp 1666464484
transform 1 0 22464 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6491
timestamp 1666464484
transform 1 0 22464 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6492
timestamp 1666464484
transform 1 0 22464 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6493
timestamp 1666464484
transform 1 0 22464 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6494
timestamp 1666464484
transform 1 0 22464 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6495
timestamp 1666464484
transform 1 0 22464 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6496
timestamp 1666464484
transform -1 0 22464 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6497
timestamp 1666464484
transform -1 0 22464 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6498
timestamp 1666464484
transform -1 0 21216 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6499
timestamp 1666464484
transform -1 0 21216 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6500
timestamp 1666464484
transform -1 0 21216 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6501
timestamp 1666464484
transform -1 0 21216 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6502
timestamp 1666464484
transform -1 0 22464 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6503
timestamp 1666464484
transform -1 0 22464 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6504
timestamp 1666464484
transform -1 0 22464 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6505
timestamp 1666464484
transform -1 0 22464 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6506
timestamp 1666464484
transform -1 0 22464 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6507
timestamp 1666464484
transform -1 0 22464 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6508
timestamp 1666464484
transform -1 0 21216 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6509
timestamp 1666464484
transform -1 0 21216 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6510
timestamp 1666464484
transform -1 0 22464 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6511
timestamp 1666464484
transform -1 0 22464 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6512
timestamp 1666464484
transform -1 0 21216 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6513
timestamp 1666464484
transform -1 0 21216 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6514
timestamp 1666464484
transform -1 0 21216 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6515
timestamp 1666464484
transform -1 0 21216 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6516
timestamp 1666464484
transform 1 0 23712 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6517
timestamp 1666464484
transform 1 0 23712 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6518
timestamp 1666464484
transform 1 0 23712 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6519
timestamp 1666464484
transform 1 0 23712 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6520
timestamp 1666464484
transform 1 0 23712 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6521
timestamp 1666464484
transform 1 0 23712 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6522
timestamp 1666464484
transform 1 0 23712 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6523
timestamp 1666464484
transform 1 0 23712 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6524
timestamp 1666464484
transform 1 0 23712 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6525
timestamp 1666464484
transform 1 0 23712 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6526
timestamp 1666464484
transform 1 0 23712 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6527
timestamp 1666464484
transform 1 0 23712 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6528
timestamp 1666464484
transform 1 0 23712 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6529
timestamp 1666464484
transform 1 0 23712 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6530
timestamp 1666464484
transform -1 0 22464 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6531
timestamp 1666464484
transform -1 0 22464 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6532
timestamp 1666464484
transform -1 0 22464 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6533
timestamp 1666464484
transform -1 0 22464 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6534
timestamp 1666464484
transform -1 0 23712 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6535
timestamp 1666464484
transform -1 0 23712 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6536
timestamp 1666464484
transform -1 0 23712 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6537
timestamp 1666464484
transform -1 0 23712 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6538
timestamp 1666464484
transform -1 0 23712 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6539
timestamp 1666464484
transform -1 0 23712 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6540
timestamp 1666464484
transform -1 0 23712 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6541
timestamp 1666464484
transform -1 0 23712 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6542
timestamp 1666464484
transform -1 0 23712 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6543
timestamp 1666464484
transform -1 0 23712 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6544
timestamp 1666464484
transform -1 0 23712 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6545
timestamp 1666464484
transform -1 0 23712 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6546
timestamp 1666464484
transform -1 0 23712 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6547
timestamp 1666464484
transform -1 0 23712 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6548
timestamp 1666464484
transform -1 0 21216 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6549
timestamp 1666464484
transform -1 0 21216 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6550
timestamp 1666464484
transform 1 0 21216 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6551
timestamp 1666464484
transform 1 0 21216 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6552
timestamp 1666464484
transform 1 0 21216 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6553
timestamp 1666464484
transform 1 0 21216 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6554
timestamp 1666464484
transform 1 0 21216 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6555
timestamp 1666464484
transform 1 0 21216 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6556
timestamp 1666464484
transform 1 0 21216 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6557
timestamp 1666464484
transform 1 0 21216 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6558
timestamp 1666464484
transform 1 0 21216 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6559
timestamp 1666464484
transform 1 0 21216 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6560
timestamp 1666464484
transform 1 0 21216 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6561
timestamp 1666464484
transform 1 0 27456 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6562
timestamp 1666464484
transform 1 0 27456 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6563
timestamp 1666464484
transform 1 0 27456 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6564
timestamp 1666464484
transform 1 0 28704 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6565
timestamp 1666464484
transform 1 0 28704 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6566
timestamp 1666464484
transform -1 0 27456 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6567
timestamp 1666464484
transform -1 0 27456 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6568
timestamp 1666464484
transform -1 0 27456 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6569
timestamp 1666464484
transform -1 0 27456 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6570
timestamp 1666464484
transform -1 0 27456 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6571
timestamp 1666464484
transform -1 0 27456 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6572
timestamp 1666464484
transform -1 0 27456 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6573
timestamp 1666464484
transform -1 0 27456 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6574
timestamp 1666464484
transform -1 0 27456 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6575
timestamp 1666464484
transform -1 0 27456 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6576
timestamp 1666464484
transform -1 0 27456 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6577
timestamp 1666464484
transform -1 0 27456 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6578
timestamp 1666464484
transform -1 0 27456 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6579
timestamp 1666464484
transform -1 0 27456 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6580
timestamp 1666464484
transform 1 0 28704 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6581
timestamp 1666464484
transform 1 0 28704 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6582
timestamp 1666464484
transform 1 0 28704 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6583
timestamp 1666464484
transform 1 0 28704 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6584
timestamp 1666464484
transform 1 0 26208 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6585
timestamp 1666464484
transform 1 0 26208 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6586
timestamp 1666464484
transform 1 0 26208 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6587
timestamp 1666464484
transform 1 0 26208 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6588
timestamp 1666464484
transform 1 0 26208 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6589
timestamp 1666464484
transform 1 0 26208 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6590
timestamp 1666464484
transform 1 0 26208 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6591
timestamp 1666464484
transform 1 0 26208 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6592
timestamp 1666464484
transform 1 0 26208 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6593
timestamp 1666464484
transform 1 0 26208 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6594
timestamp 1666464484
transform 1 0 26208 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6595
timestamp 1666464484
transform 1 0 26208 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6596
timestamp 1666464484
transform 1 0 26208 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6597
timestamp 1666464484
transform 1 0 26208 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6598
timestamp 1666464484
transform 1 0 28704 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6599
timestamp 1666464484
transform 1 0 28704 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6600
timestamp 1666464484
transform 1 0 28704 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6601
timestamp 1666464484
transform 1 0 28704 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6602
timestamp 1666464484
transform -1 0 26208 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6603
timestamp 1666464484
transform -1 0 26208 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6604
timestamp 1666464484
transform -1 0 26208 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6605
timestamp 1666464484
transform -1 0 26208 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6606
timestamp 1666464484
transform -1 0 26208 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6607
timestamp 1666464484
transform -1 0 26208 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6608
timestamp 1666464484
transform -1 0 26208 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6609
timestamp 1666464484
transform -1 0 26208 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6610
timestamp 1666464484
transform -1 0 26208 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6611
timestamp 1666464484
transform -1 0 26208 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6612
timestamp 1666464484
transform -1 0 26208 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6613
timestamp 1666464484
transform -1 0 26208 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6614
timestamp 1666464484
transform -1 0 26208 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6615
timestamp 1666464484
transform -1 0 26208 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6616
timestamp 1666464484
transform 1 0 28704 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6617
timestamp 1666464484
transform 1 0 28704 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6618
timestamp 1666464484
transform 1 0 28704 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6619
timestamp 1666464484
transform 1 0 28704 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6620
timestamp 1666464484
transform 1 0 27456 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6621
timestamp 1666464484
transform 1 0 27456 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6622
timestamp 1666464484
transform 1 0 27456 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6623
timestamp 1666464484
transform 1 0 27456 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6624
timestamp 1666464484
transform 1 0 27456 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6625
timestamp 1666464484
transform 1 0 27456 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6626
timestamp 1666464484
transform 1 0 27456 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6627
timestamp 1666464484
transform 1 0 27456 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6628
timestamp 1666464484
transform -1 0 28704 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6629
timestamp 1666464484
transform -1 0 28704 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6630
timestamp 1666464484
transform -1 0 28704 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6631
timestamp 1666464484
transform -1 0 28704 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6632
timestamp 1666464484
transform -1 0 28704 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6633
timestamp 1666464484
transform -1 0 28704 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6634
timestamp 1666464484
transform -1 0 28704 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6635
timestamp 1666464484
transform -1 0 28704 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6636
timestamp 1666464484
transform -1 0 28704 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6637
timestamp 1666464484
transform -1 0 28704 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6638
timestamp 1666464484
transform -1 0 28704 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6639
timestamp 1666464484
transform -1 0 28704 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6640
timestamp 1666464484
transform -1 0 28704 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6641
timestamp 1666464484
transform -1 0 28704 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6642
timestamp 1666464484
transform 1 0 27456 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6643
timestamp 1666464484
transform 1 0 27456 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6644
timestamp 1666464484
transform 1 0 27456 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6645
timestamp 1666464484
transform -1 0 24960 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6646
timestamp 1666464484
transform -1 0 24960 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6647
timestamp 1666464484
transform -1 0 24960 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6648
timestamp 1666464484
transform 1 0 22464 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6649
timestamp 1666464484
transform 1 0 22464 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6650
timestamp 1666464484
transform -1 0 27456 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6651
timestamp 1666464484
transform -1 0 27456 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6652
timestamp 1666464484
transform 1 0 23712 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6653
timestamp 1666464484
transform 1 0 23712 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6654
timestamp 1666464484
transform 1 0 26208 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6655
timestamp 1666464484
transform 1 0 26208 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6656
timestamp 1666464484
transform 1 0 21216 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6657
timestamp 1666464484
transform 1 0 21216 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6658
timestamp 1666464484
transform -1 0 26208 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6659
timestamp 1666464484
transform -1 0 26208 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6660
timestamp 1666464484
transform -1 0 21216 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6661
timestamp 1666464484
transform -1 0 21216 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6662
timestamp 1666464484
transform -1 0 23712 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6663
timestamp 1666464484
transform -1 0 23712 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6664
timestamp 1666464484
transform 1 0 24960 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6665
timestamp 1666464484
transform 1 0 24960 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6666
timestamp 1666464484
transform 1 0 24960 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6667
timestamp 1666464484
transform 1 0 24960 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6668
timestamp 1666464484
transform 1 0 24960 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6669
timestamp 1666464484
transform 1 0 24960 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6670
timestamp 1666464484
transform 1 0 24960 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6671
timestamp 1666464484
transform 1 0 24960 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6672
timestamp 1666464484
transform 1 0 24960 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6673
timestamp 1666464484
transform 1 0 24960 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6674
timestamp 1666464484
transform 1 0 24960 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6675
timestamp 1666464484
transform 1 0 24960 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6676
timestamp 1666464484
transform 1 0 24960 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6677
timestamp 1666464484
transform 1 0 24960 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6678
timestamp 1666464484
transform 1 0 24960 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6679
timestamp 1666464484
transform 1 0 24960 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6680
timestamp 1666464484
transform 1 0 24960 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6681
timestamp 1666464484
transform 1 0 24960 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6682
timestamp 1666464484
transform 1 0 24960 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6683
timestamp 1666464484
transform 1 0 24960 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6684
timestamp 1666464484
transform 1 0 24960 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6685
timestamp 1666464484
transform 1 0 24960 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6686
timestamp 1666464484
transform 1 0 24960 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6687
timestamp 1666464484
transform 1 0 24960 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6688
timestamp 1666464484
transform 1 0 24960 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6689
timestamp 1666464484
transform 1 0 24960 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6690
timestamp 1666464484
transform 1 0 28704 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6691
timestamp 1666464484
transform 1 0 28704 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6692
timestamp 1666464484
transform 1 0 24960 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6693
timestamp 1666464484
transform 1 0 24960 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6694
timestamp 1666464484
transform 1 0 24960 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6695
timestamp 1666464484
transform 1 0 24960 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6696
timestamp 1666464484
transform -1 0 22464 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6697
timestamp 1666464484
transform -1 0 22464 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6698
timestamp 1666464484
transform -1 0 28704 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6699
timestamp 1666464484
transform -1 0 28704 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6700
timestamp 1666464484
transform -1 0 24960 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6701
timestamp 1666464484
transform -1 0 24960 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6702
timestamp 1666464484
transform -1 0 24960 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6703
timestamp 1666464484
transform -1 0 24960 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6704
timestamp 1666464484
transform -1 0 24960 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6705
timestamp 1666464484
transform -1 0 24960 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6706
timestamp 1666464484
transform -1 0 24960 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6707
timestamp 1666464484
transform -1 0 24960 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6708
timestamp 1666464484
transform -1 0 24960 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6709
timestamp 1666464484
transform -1 0 24960 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6710
timestamp 1666464484
transform -1 0 24960 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6711
timestamp 1666464484
transform -1 0 24960 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6712
timestamp 1666464484
transform -1 0 24960 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6713
timestamp 1666464484
transform -1 0 24960 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6714
timestamp 1666464484
transform -1 0 24960 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6715
timestamp 1666464484
transform -1 0 24960 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6716
timestamp 1666464484
transform -1 0 24960 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6717
timestamp 1666464484
transform -1 0 24960 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6718
timestamp 1666464484
transform -1 0 24960 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6719
timestamp 1666464484
transform -1 0 24960 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6720
timestamp 1666464484
transform -1 0 24960 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6721
timestamp 1666464484
transform -1 0 24960 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6722
timestamp 1666464484
transform -1 0 24960 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6723
timestamp 1666464484
transform -1 0 24960 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6724
timestamp 1666464484
transform -1 0 24960 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6725
timestamp 1666464484
transform -1 0 24960 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6726
timestamp 1666464484
transform -1 0 24960 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6727
timestamp 1666464484
transform 1 0 27456 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6728
timestamp 1666464484
transform 1 0 27456 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6729
timestamp 1666464484
transform -1 0 26208 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6730
timestamp 1666464484
transform -1 0 26208 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6731
timestamp 1666464484
transform -1 0 26208 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6732
timestamp 1666464484
transform 1 0 27456 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6733
timestamp 1666464484
transform 1 0 27456 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6734
timestamp 1666464484
transform 1 0 28704 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6735
timestamp 1666464484
transform 1 0 28704 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6736
timestamp 1666464484
transform 1 0 28704 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6737
timestamp 1666464484
transform 1 0 28704 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6738
timestamp 1666464484
transform 1 0 28704 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6739
timestamp 1666464484
transform 1 0 28704 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6740
timestamp 1666464484
transform 1 0 28704 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6741
timestamp 1666464484
transform 1 0 28704 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6742
timestamp 1666464484
transform 1 0 28704 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6743
timestamp 1666464484
transform 1 0 28704 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6744
timestamp 1666464484
transform 1 0 28704 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6745
timestamp 1666464484
transform 1 0 28704 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6746
timestamp 1666464484
transform 1 0 28704 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6747
timestamp 1666464484
transform 1 0 28704 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6748
timestamp 1666464484
transform 1 0 27456 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6749
timestamp 1666464484
transform 1 0 27456 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6750
timestamp 1666464484
transform 1 0 27456 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6751
timestamp 1666464484
transform 1 0 26208 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6752
timestamp 1666464484
transform 1 0 26208 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6753
timestamp 1666464484
transform 1 0 26208 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6754
timestamp 1666464484
transform 1 0 26208 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6755
timestamp 1666464484
transform 1 0 26208 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6756
timestamp 1666464484
transform 1 0 26208 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6757
timestamp 1666464484
transform -1 0 26208 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6758
timestamp 1666464484
transform -1 0 26208 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6759
timestamp 1666464484
transform -1 0 26208 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6760
timestamp 1666464484
transform -1 0 26208 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6761
timestamp 1666464484
transform -1 0 26208 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6762
timestamp 1666464484
transform -1 0 26208 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6763
timestamp 1666464484
transform -1 0 26208 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6764
timestamp 1666464484
transform -1 0 26208 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6765
timestamp 1666464484
transform -1 0 26208 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6766
timestamp 1666464484
transform -1 0 26208 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6767
timestamp 1666464484
transform -1 0 26208 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6768
timestamp 1666464484
transform 1 0 26208 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6769
timestamp 1666464484
transform -1 0 28704 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6770
timestamp 1666464484
transform -1 0 28704 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6771
timestamp 1666464484
transform -1 0 28704 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6772
timestamp 1666464484
transform -1 0 28704 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6773
timestamp 1666464484
transform -1 0 28704 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6774
timestamp 1666464484
transform -1 0 28704 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6775
timestamp 1666464484
transform -1 0 28704 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6776
timestamp 1666464484
transform -1 0 28704 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6777
timestamp 1666464484
transform -1 0 28704 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6778
timestamp 1666464484
transform -1 0 28704 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6779
timestamp 1666464484
transform -1 0 28704 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6780
timestamp 1666464484
transform -1 0 28704 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6781
timestamp 1666464484
transform -1 0 28704 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6782
timestamp 1666464484
transform -1 0 28704 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6783
timestamp 1666464484
transform 1 0 26208 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6784
timestamp 1666464484
transform 1 0 26208 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6785
timestamp 1666464484
transform 1 0 26208 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6786
timestamp 1666464484
transform -1 0 27456 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6787
timestamp 1666464484
transform -1 0 27456 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6788
timestamp 1666464484
transform -1 0 27456 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6789
timestamp 1666464484
transform -1 0 27456 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6790
timestamp 1666464484
transform -1 0 27456 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6791
timestamp 1666464484
transform -1 0 27456 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6792
timestamp 1666464484
transform -1 0 27456 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6793
timestamp 1666464484
transform -1 0 27456 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6794
timestamp 1666464484
transform -1 0 27456 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6795
timestamp 1666464484
transform -1 0 27456 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6796
timestamp 1666464484
transform -1 0 27456 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6797
timestamp 1666464484
transform -1 0 27456 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6798
timestamp 1666464484
transform -1 0 27456 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6799
timestamp 1666464484
transform -1 0 27456 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6800
timestamp 1666464484
transform 1 0 26208 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6801
timestamp 1666464484
transform 1 0 26208 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6802
timestamp 1666464484
transform 1 0 26208 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6803
timestamp 1666464484
transform 1 0 26208 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6804
timestamp 1666464484
transform 1 0 27456 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6805
timestamp 1666464484
transform 1 0 27456 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6806
timestamp 1666464484
transform 1 0 27456 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6807
timestamp 1666464484
transform 1 0 27456 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6808
timestamp 1666464484
transform 1 0 27456 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6809
timestamp 1666464484
transform 1 0 27456 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6810
timestamp 1666464484
transform 1 0 27456 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6811
timestamp 1666464484
transform 1 0 27456 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6812
timestamp 1666464484
transform 1 0 27456 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6813
timestamp 1666464484
transform 1 0 21216 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6814
timestamp 1666464484
transform 1 0 21216 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6815
timestamp 1666464484
transform -1 0 22464 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6816
timestamp 1666464484
transform -1 0 22464 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6817
timestamp 1666464484
transform -1 0 22464 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6818
timestamp 1666464484
transform -1 0 22464 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6819
timestamp 1666464484
transform -1 0 22464 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6820
timestamp 1666464484
transform 1 0 22464 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6821
timestamp 1666464484
transform 1 0 22464 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6822
timestamp 1666464484
transform 1 0 22464 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6823
timestamp 1666464484
transform 1 0 22464 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6824
timestamp 1666464484
transform 1 0 23712 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6825
timestamp 1666464484
transform 1 0 23712 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6826
timestamp 1666464484
transform 1 0 23712 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6827
timestamp 1666464484
transform 1 0 23712 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6828
timestamp 1666464484
transform 1 0 23712 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6829
timestamp 1666464484
transform -1 0 21216 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6830
timestamp 1666464484
transform -1 0 21216 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6831
timestamp 1666464484
transform 1 0 23712 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6832
timestamp 1666464484
transform 1 0 23712 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6833
timestamp 1666464484
transform 1 0 22464 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6834
timestamp 1666464484
transform 1 0 22464 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6835
timestamp 1666464484
transform 1 0 23712 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6836
timestamp 1666464484
transform 1 0 23712 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6837
timestamp 1666464484
transform 1 0 23712 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6838
timestamp 1666464484
transform 1 0 23712 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6839
timestamp 1666464484
transform 1 0 23712 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6840
timestamp 1666464484
transform 1 0 23712 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6841
timestamp 1666464484
transform 1 0 23712 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6842
timestamp 1666464484
transform 1 0 21216 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6843
timestamp 1666464484
transform 1 0 21216 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6844
timestamp 1666464484
transform 1 0 22464 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6845
timestamp 1666464484
transform -1 0 21216 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6846
timestamp 1666464484
transform -1 0 21216 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6847
timestamp 1666464484
transform 1 0 22464 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6848
timestamp 1666464484
transform 1 0 22464 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6849
timestamp 1666464484
transform 1 0 22464 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6850
timestamp 1666464484
transform 1 0 21216 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6851
timestamp 1666464484
transform 1 0 21216 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6852
timestamp 1666464484
transform 1 0 22464 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6853
timestamp 1666464484
transform 1 0 22464 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6854
timestamp 1666464484
transform 1 0 22464 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6855
timestamp 1666464484
transform 1 0 22464 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6856
timestamp 1666464484
transform 1 0 21216 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6857
timestamp 1666464484
transform -1 0 22464 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6858
timestamp 1666464484
transform -1 0 22464 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6859
timestamp 1666464484
transform -1 0 22464 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6860
timestamp 1666464484
transform -1 0 22464 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6861
timestamp 1666464484
transform -1 0 22464 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6862
timestamp 1666464484
transform -1 0 22464 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6863
timestamp 1666464484
transform -1 0 23712 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6864
timestamp 1666464484
transform -1 0 23712 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6865
timestamp 1666464484
transform -1 0 23712 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6866
timestamp 1666464484
transform -1 0 21216 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6867
timestamp 1666464484
transform -1 0 21216 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6868
timestamp 1666464484
transform -1 0 23712 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6869
timestamp 1666464484
transform -1 0 23712 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6870
timestamp 1666464484
transform -1 0 23712 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6871
timestamp 1666464484
transform -1 0 23712 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6872
timestamp 1666464484
transform -1 0 22464 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6873
timestamp 1666464484
transform -1 0 21216 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6874
timestamp 1666464484
transform -1 0 23712 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6875
timestamp 1666464484
transform -1 0 23712 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6876
timestamp 1666464484
transform -1 0 23712 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6877
timestamp 1666464484
transform -1 0 23712 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6878
timestamp 1666464484
transform -1 0 23712 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6879
timestamp 1666464484
transform -1 0 23712 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6880
timestamp 1666464484
transform -1 0 23712 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6881
timestamp 1666464484
transform 1 0 21216 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6882
timestamp 1666464484
transform 1 0 21216 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6883
timestamp 1666464484
transform 1 0 21216 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6884
timestamp 1666464484
transform -1 0 21216 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6885
timestamp 1666464484
transform 1 0 21216 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6886
timestamp 1666464484
transform -1 0 21216 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6887
timestamp 1666464484
transform 1 0 21216 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6888
timestamp 1666464484
transform 1 0 21216 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6889
timestamp 1666464484
transform -1 0 21216 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6890
timestamp 1666464484
transform -1 0 21216 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6891
timestamp 1666464484
transform 1 0 21216 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6892
timestamp 1666464484
transform -1 0 21216 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6893
timestamp 1666464484
transform -1 0 21216 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6894
timestamp 1666464484
transform -1 0 21216 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6895
timestamp 1666464484
transform -1 0 22464 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6896
timestamp 1666464484
transform -1 0 22464 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6897
timestamp 1666464484
transform -1 0 23712 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6898
timestamp 1666464484
transform -1 0 23712 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6899
timestamp 1666464484
transform -1 0 23712 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6900
timestamp 1666464484
transform -1 0 23712 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6901
timestamp 1666464484
transform -1 0 23712 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6902
timestamp 1666464484
transform -1 0 23712 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6903
timestamp 1666464484
transform -1 0 23712 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6904
timestamp 1666464484
transform -1 0 23712 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6905
timestamp 1666464484
transform -1 0 23712 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6906
timestamp 1666464484
transform -1 0 23712 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6907
timestamp 1666464484
transform 1 0 21216 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6908
timestamp 1666464484
transform 1 0 21216 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6909
timestamp 1666464484
transform -1 0 21216 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6910
timestamp 1666464484
transform -1 0 21216 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6911
timestamp 1666464484
transform 1 0 22464 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6912
timestamp 1666464484
transform 1 0 22464 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6913
timestamp 1666464484
transform 1 0 22464 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6914
timestamp 1666464484
transform 1 0 22464 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6915
timestamp 1666464484
transform 1 0 22464 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6916
timestamp 1666464484
transform 1 0 22464 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6917
timestamp 1666464484
transform 1 0 22464 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6918
timestamp 1666464484
transform 1 0 22464 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6919
timestamp 1666464484
transform 1 0 22464 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6920
timestamp 1666464484
transform 1 0 22464 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6921
timestamp 1666464484
transform 1 0 22464 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6922
timestamp 1666464484
transform 1 0 22464 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6923
timestamp 1666464484
transform -1 0 21216 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6924
timestamp 1666464484
transform -1 0 21216 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6925
timestamp 1666464484
transform 1 0 22464 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6926
timestamp 1666464484
transform 1 0 22464 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6927
timestamp 1666464484
transform 1 0 22464 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6928
timestamp 1666464484
transform 1 0 21216 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6929
timestamp 1666464484
transform 1 0 21216 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6930
timestamp 1666464484
transform -1 0 21216 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6931
timestamp 1666464484
transform -1 0 21216 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6932
timestamp 1666464484
transform -1 0 21216 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6933
timestamp 1666464484
transform -1 0 22464 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6934
timestamp 1666464484
transform -1 0 22464 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6935
timestamp 1666464484
transform -1 0 22464 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6936
timestamp 1666464484
transform -1 0 22464 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6937
timestamp 1666464484
transform -1 0 22464 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6938
timestamp 1666464484
transform -1 0 22464 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6939
timestamp 1666464484
transform -1 0 22464 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6940
timestamp 1666464484
transform -1 0 22464 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6941
timestamp 1666464484
transform -1 0 22464 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6942
timestamp 1666464484
transform -1 0 22464 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6943
timestamp 1666464484
transform -1 0 22464 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6944
timestamp 1666464484
transform -1 0 22464 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6945
timestamp 1666464484
transform -1 0 22464 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6946
timestamp 1666464484
transform -1 0 22464 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6947
timestamp 1666464484
transform -1 0 22464 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6948
timestamp 1666464484
transform 1 0 21216 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6949
timestamp 1666464484
transform 1 0 21216 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6950
timestamp 1666464484
transform -1 0 21216 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6951
timestamp 1666464484
transform -1 0 21216 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6952
timestamp 1666464484
transform -1 0 21216 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6953
timestamp 1666464484
transform -1 0 21216 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6954
timestamp 1666464484
transform -1 0 21216 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6955
timestamp 1666464484
transform -1 0 21216 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6956
timestamp 1666464484
transform 1 0 21216 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6957
timestamp 1666464484
transform 1 0 21216 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6958
timestamp 1666464484
transform 1 0 21216 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6959
timestamp 1666464484
transform 1 0 21216 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6960
timestamp 1666464484
transform 1 0 21216 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6961
timestamp 1666464484
transform 1 0 21216 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6962
timestamp 1666464484
transform 1 0 21216 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6963
timestamp 1666464484
transform 1 0 23712 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6964
timestamp 1666464484
transform 1 0 23712 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6965
timestamp 1666464484
transform 1 0 23712 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6966
timestamp 1666464484
transform 1 0 23712 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6967
timestamp 1666464484
transform 1 0 23712 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6968
timestamp 1666464484
transform 1 0 23712 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6969
timestamp 1666464484
transform 1 0 23712 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6970
timestamp 1666464484
transform 1 0 23712 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6971
timestamp 1666464484
transform 1 0 23712 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6972
timestamp 1666464484
transform 1 0 23712 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6973
timestamp 1666464484
transform 1 0 23712 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6974
timestamp 1666464484
transform 1 0 23712 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6975
timestamp 1666464484
transform 1 0 23712 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6976
timestamp 1666464484
transform 1 0 23712 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6977
timestamp 1666464484
transform 1 0 23712 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6978
timestamp 1666464484
transform 1 0 21216 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6979
timestamp 1666464484
transform 1 0 21216 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6980
timestamp 1666464484
transform -1 0 21216 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6981
timestamp 1666464484
transform -1 0 21216 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6982
timestamp 1666464484
transform -1 0 23712 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6983
timestamp 1666464484
transform -1 0 23712 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6984
timestamp 1666464484
transform -1 0 23712 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6985
timestamp 1666464484
transform -1 0 23712 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6986
timestamp 1666464484
transform -1 0 23712 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6987
timestamp 1666464484
transform -1 0 28704 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6988
timestamp 1666464484
transform -1 0 28704 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6989
timestamp 1666464484
transform -1 0 28704 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6990
timestamp 1666464484
transform -1 0 28704 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6991
timestamp 1666464484
transform -1 0 28704 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6992
timestamp 1666464484
transform -1 0 28704 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6993
timestamp 1666464484
transform -1 0 28704 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6994
timestamp 1666464484
transform -1 0 28704 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6995
timestamp 1666464484
transform -1 0 28704 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6996
timestamp 1666464484
transform -1 0 28704 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6997
timestamp 1666464484
transform -1 0 28704 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6998
timestamp 1666464484
transform -1 0 28704 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_6999
timestamp 1666464484
transform -1 0 28704 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7000
timestamp 1666464484
transform -1 0 28704 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7001
timestamp 1666464484
transform -1 0 26208 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7002
timestamp 1666464484
transform -1 0 26208 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7003
timestamp 1666464484
transform 1 0 27456 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7004
timestamp 1666464484
transform 1 0 27456 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7005
timestamp 1666464484
transform 1 0 27456 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7006
timestamp 1666464484
transform 1 0 27456 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7007
timestamp 1666464484
transform 1 0 27456 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7008
timestamp 1666464484
transform 1 0 27456 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7009
timestamp 1666464484
transform 1 0 27456 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7010
timestamp 1666464484
transform 1 0 27456 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7011
timestamp 1666464484
transform 1 0 27456 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7012
timestamp 1666464484
transform 1 0 27456 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7013
timestamp 1666464484
transform 1 0 27456 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7014
timestamp 1666464484
transform 1 0 27456 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7015
timestamp 1666464484
transform 1 0 27456 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7016
timestamp 1666464484
transform 1 0 27456 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7017
timestamp 1666464484
transform 1 0 27456 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7018
timestamp 1666464484
transform -1 0 26208 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7019
timestamp 1666464484
transform -1 0 26208 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7020
timestamp 1666464484
transform -1 0 26208 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7021
timestamp 1666464484
transform -1 0 27456 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7022
timestamp 1666464484
transform -1 0 27456 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7023
timestamp 1666464484
transform -1 0 27456 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7024
timestamp 1666464484
transform -1 0 27456 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7025
timestamp 1666464484
transform -1 0 27456 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7026
timestamp 1666464484
transform -1 0 27456 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7027
timestamp 1666464484
transform -1 0 27456 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7028
timestamp 1666464484
transform -1 0 27456 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7029
timestamp 1666464484
transform -1 0 27456 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7030
timestamp 1666464484
transform -1 0 27456 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7031
timestamp 1666464484
transform -1 0 27456 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7032
timestamp 1666464484
transform -1 0 27456 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7033
timestamp 1666464484
transform -1 0 27456 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7034
timestamp 1666464484
transform -1 0 27456 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7035
timestamp 1666464484
transform -1 0 27456 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7036
timestamp 1666464484
transform -1 0 26208 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7037
timestamp 1666464484
transform -1 0 26208 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7038
timestamp 1666464484
transform -1 0 26208 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7039
timestamp 1666464484
transform 1 0 26208 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7040
timestamp 1666464484
transform 1 0 26208 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7041
timestamp 1666464484
transform 1 0 26208 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7042
timestamp 1666464484
transform 1 0 26208 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7043
timestamp 1666464484
transform 1 0 26208 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7044
timestamp 1666464484
transform 1 0 26208 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7045
timestamp 1666464484
transform 1 0 26208 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7046
timestamp 1666464484
transform 1 0 26208 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7047
timestamp 1666464484
transform 1 0 26208 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7048
timestamp 1666464484
transform 1 0 26208 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7049
timestamp 1666464484
transform 1 0 26208 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7050
timestamp 1666464484
transform 1 0 26208 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7051
timestamp 1666464484
transform 1 0 26208 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7052
timestamp 1666464484
transform 1 0 26208 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7053
timestamp 1666464484
transform 1 0 26208 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7054
timestamp 1666464484
transform -1 0 26208 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7055
timestamp 1666464484
transform -1 0 26208 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7056
timestamp 1666464484
transform -1 0 26208 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7057
timestamp 1666464484
transform 1 0 28704 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7058
timestamp 1666464484
transform 1 0 28704 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7059
timestamp 1666464484
transform 1 0 28704 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7060
timestamp 1666464484
transform 1 0 28704 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7061
timestamp 1666464484
transform 1 0 28704 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7062
timestamp 1666464484
transform 1 0 28704 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7063
timestamp 1666464484
transform 1 0 28704 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7064
timestamp 1666464484
transform 1 0 28704 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7065
timestamp 1666464484
transform 1 0 28704 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7066
timestamp 1666464484
transform 1 0 28704 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7067
timestamp 1666464484
transform 1 0 28704 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7068
timestamp 1666464484
transform 1 0 28704 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7069
timestamp 1666464484
transform 1 0 28704 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7070
timestamp 1666464484
transform 1 0 28704 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7071
timestamp 1666464484
transform -1 0 26208 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7072
timestamp 1666464484
transform -1 0 26208 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7073
timestamp 1666464484
transform 1 0 28704 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7074
timestamp 1666464484
transform -1 0 26208 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7075
timestamp 1666464484
transform -1 0 26208 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7076
timestamp 1666464484
transform -1 0 28704 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7077
timestamp 1666464484
transform 1 0 24960 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7078
timestamp 1666464484
transform 1 0 24960 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7079
timestamp 1666464484
transform 1 0 24960 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7080
timestamp 1666464484
transform 1 0 24960 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7081
timestamp 1666464484
transform 1 0 24960 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7082
timestamp 1666464484
transform 1 0 24960 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7083
timestamp 1666464484
transform 1 0 24960 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7084
timestamp 1666464484
transform 1 0 24960 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7085
timestamp 1666464484
transform 1 0 24960 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7086
timestamp 1666464484
transform 1 0 24960 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7087
timestamp 1666464484
transform 1 0 24960 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7088
timestamp 1666464484
transform 1 0 24960 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7089
timestamp 1666464484
transform 1 0 24960 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7090
timestamp 1666464484
transform 1 0 24960 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7091
timestamp 1666464484
transform 1 0 24960 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7092
timestamp 1666464484
transform 1 0 24960 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7093
timestamp 1666464484
transform 1 0 24960 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7094
timestamp 1666464484
transform 1 0 24960 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7095
timestamp 1666464484
transform 1 0 24960 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7096
timestamp 1666464484
transform 1 0 24960 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7097
timestamp 1666464484
transform 1 0 24960 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7098
timestamp 1666464484
transform 1 0 24960 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7099
timestamp 1666464484
transform 1 0 24960 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7100
timestamp 1666464484
transform 1 0 24960 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7101
timestamp 1666464484
transform 1 0 24960 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7102
timestamp 1666464484
transform 1 0 24960 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7103
timestamp 1666464484
transform 1 0 24960 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7104
timestamp 1666464484
transform 1 0 24960 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7105
timestamp 1666464484
transform 1 0 24960 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7106
timestamp 1666464484
transform 1 0 24960 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7107
timestamp 1666464484
transform 1 0 24960 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7108
timestamp 1666464484
transform -1 0 24960 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7109
timestamp 1666464484
transform -1 0 24960 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7110
timestamp 1666464484
transform -1 0 24960 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7111
timestamp 1666464484
transform -1 0 24960 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7112
timestamp 1666464484
transform -1 0 24960 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7113
timestamp 1666464484
transform -1 0 24960 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7114
timestamp 1666464484
transform -1 0 24960 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7115
timestamp 1666464484
transform -1 0 24960 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7116
timestamp 1666464484
transform -1 0 24960 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7117
timestamp 1666464484
transform -1 0 24960 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7118
timestamp 1666464484
transform -1 0 24960 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7119
timestamp 1666464484
transform -1 0 24960 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7120
timestamp 1666464484
transform -1 0 24960 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7121
timestamp 1666464484
transform -1 0 24960 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7122
timestamp 1666464484
transform -1 0 24960 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7123
timestamp 1666464484
transform -1 0 24960 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7124
timestamp 1666464484
transform -1 0 24960 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7125
timestamp 1666464484
transform -1 0 24960 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7126
timestamp 1666464484
transform -1 0 24960 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7127
timestamp 1666464484
transform -1 0 24960 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7128
timestamp 1666464484
transform -1 0 24960 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7129
timestamp 1666464484
transform -1 0 24960 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7130
timestamp 1666464484
transform -1 0 24960 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7131
timestamp 1666464484
transform -1 0 24960 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7132
timestamp 1666464484
transform -1 0 24960 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7133
timestamp 1666464484
transform -1 0 24960 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7134
timestamp 1666464484
transform -1 0 24960 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7135
timestamp 1666464484
transform -1 0 24960 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7136
timestamp 1666464484
transform -1 0 24960 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7137
timestamp 1666464484
transform -1 0 24960 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7138
timestamp 1666464484
transform -1 0 24960 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7139
timestamp 1666464484
transform 1 0 23712 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7140
timestamp 1666464484
transform 1 0 23712 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7141
timestamp 1666464484
transform -1 0 23712 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7142
timestamp 1666464484
transform -1 0 23712 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7143
timestamp 1666464484
transform 1 0 22464 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7144
timestamp 1666464484
transform 1 0 22464 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7145
timestamp 1666464484
transform -1 0 22464 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7146
timestamp 1666464484
transform -1 0 22464 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7147
timestamp 1666464484
transform -1 0 21216 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7148
timestamp 1666464484
transform -1 0 21216 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7149
timestamp 1666464484
transform 1 0 28704 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7150
timestamp 1666464484
transform 1 0 28704 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7151
timestamp 1666464484
transform -1 0 28704 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7152
timestamp 1666464484
transform -1 0 28704 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7153
timestamp 1666464484
transform 1 0 27456 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7154
timestamp 1666464484
transform 1 0 27456 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7155
timestamp 1666464484
transform 1 0 21216 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7156
timestamp 1666464484
transform -1 0 27456 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7157
timestamp 1666464484
transform -1 0 27456 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7158
timestamp 1666464484
transform 1 0 21216 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7159
timestamp 1666464484
transform 1 0 26208 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7160
timestamp 1666464484
transform 1 0 26208 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7161
timestamp 1666464484
transform -1 0 26208 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7162
timestamp 1666464484
transform -1 0 26208 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7163
timestamp 1666464484
transform -1 0 37440 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7164
timestamp 1666464484
transform -1 0 37440 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7165
timestamp 1666464484
transform -1 0 37440 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7166
timestamp 1666464484
transform -1 0 37440 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7167
timestamp 1666464484
transform -1 0 37440 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7168
timestamp 1666464484
transform -1 0 37440 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7169
timestamp 1666464484
transform -1 0 37440 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7170
timestamp 1666464484
transform -1 0 37440 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7171
timestamp 1666464484
transform -1 0 37440 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7172
timestamp 1666464484
transform 1 0 36192 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7173
timestamp 1666464484
transform 1 0 36192 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7174
timestamp 1666464484
transform 1 0 36192 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7175
timestamp 1666464484
transform 1 0 36192 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7176
timestamp 1666464484
transform 1 0 36192 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7177
timestamp 1666464484
transform -1 0 36192 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7178
timestamp 1666464484
transform -1 0 36192 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7179
timestamp 1666464484
transform -1 0 36192 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7180
timestamp 1666464484
transform -1 0 39936 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7181
timestamp 1666464484
transform -1 0 39936 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7182
timestamp 1666464484
transform -1 0 39936 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7183
timestamp 1666464484
transform -1 0 39936 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7184
timestamp 1666464484
transform -1 0 39936 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7185
timestamp 1666464484
transform -1 0 39936 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7186
timestamp 1666464484
transform -1 0 39936 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7187
timestamp 1666464484
transform -1 0 39936 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7188
timestamp 1666464484
transform -1 0 39936 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7189
timestamp 1666464484
transform -1 0 39936 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7190
timestamp 1666464484
transform -1 0 39936 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7191
timestamp 1666464484
transform -1 0 39936 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7192
timestamp 1666464484
transform -1 0 39936 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7193
timestamp 1666464484
transform -1 0 39936 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7194
timestamp 1666464484
transform -1 0 36192 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7195
timestamp 1666464484
transform 1 0 37440 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7196
timestamp 1666464484
transform 1 0 37440 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7197
timestamp 1666464484
transform 1 0 37440 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7198
timestamp 1666464484
transform 1 0 37440 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7199
timestamp 1666464484
transform 1 0 37440 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7200
timestamp 1666464484
transform 1 0 37440 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7201
timestamp 1666464484
transform 1 0 37440 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7202
timestamp 1666464484
transform 1 0 37440 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7203
timestamp 1666464484
transform 1 0 37440 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7204
timestamp 1666464484
transform 1 0 37440 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7205
timestamp 1666464484
transform 1 0 37440 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7206
timestamp 1666464484
transform 1 0 37440 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7207
timestamp 1666464484
transform 1 0 37440 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7208
timestamp 1666464484
transform 1 0 37440 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7209
timestamp 1666464484
transform -1 0 36192 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7210
timestamp 1666464484
transform -1 0 36192 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7211
timestamp 1666464484
transform -1 0 36192 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7212
timestamp 1666464484
transform -1 0 36192 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7213
timestamp 1666464484
transform 1 0 38688 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7214
timestamp 1666464484
transform 1 0 38688 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7215
timestamp 1666464484
transform 1 0 38688 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7216
timestamp 1666464484
transform 1 0 38688 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7217
timestamp 1666464484
transform 1 0 38688 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7218
timestamp 1666464484
transform 1 0 38688 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7219
timestamp 1666464484
transform 1 0 38688 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7220
timestamp 1666464484
transform 1 0 38688 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7221
timestamp 1666464484
transform 1 0 38688 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7222
timestamp 1666464484
transform 1 0 38688 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7223
timestamp 1666464484
transform 1 0 38688 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7224
timestamp 1666464484
transform 1 0 38688 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7225
timestamp 1666464484
transform 1 0 38688 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7226
timestamp 1666464484
transform 1 0 38688 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7227
timestamp 1666464484
transform -1 0 36192 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7228
timestamp 1666464484
transform -1 0 36192 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7229
timestamp 1666464484
transform -1 0 36192 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7230
timestamp 1666464484
transform -1 0 36192 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7231
timestamp 1666464484
transform -1 0 36192 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7232
timestamp 1666464484
transform -1 0 36192 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7233
timestamp 1666464484
transform 1 0 36192 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7234
timestamp 1666464484
transform 1 0 36192 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7235
timestamp 1666464484
transform 1 0 36192 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7236
timestamp 1666464484
transform 1 0 36192 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7237
timestamp 1666464484
transform 1 0 36192 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7238
timestamp 1666464484
transform 1 0 36192 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7239
timestamp 1666464484
transform 1 0 36192 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7240
timestamp 1666464484
transform 1 0 36192 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7241
timestamp 1666464484
transform 1 0 36192 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7242
timestamp 1666464484
transform -1 0 37440 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7243
timestamp 1666464484
transform -1 0 37440 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7244
timestamp 1666464484
transform -1 0 37440 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7245
timestamp 1666464484
transform -1 0 37440 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7246
timestamp 1666464484
transform -1 0 38688 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7247
timestamp 1666464484
transform -1 0 38688 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7248
timestamp 1666464484
transform -1 0 38688 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7249
timestamp 1666464484
transform -1 0 38688 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7250
timestamp 1666464484
transform -1 0 38688 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7251
timestamp 1666464484
transform -1 0 38688 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7252
timestamp 1666464484
transform -1 0 38688 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7253
timestamp 1666464484
transform -1 0 38688 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7254
timestamp 1666464484
transform -1 0 38688 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7255
timestamp 1666464484
transform -1 0 38688 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7256
timestamp 1666464484
transform -1 0 38688 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7257
timestamp 1666464484
transform -1 0 38688 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7258
timestamp 1666464484
transform -1 0 38688 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7259
timestamp 1666464484
transform -1 0 38688 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7260
timestamp 1666464484
transform -1 0 37440 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7261
timestamp 1666464484
transform -1 0 33696 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7262
timestamp 1666464484
transform -1 0 33696 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7263
timestamp 1666464484
transform -1 0 33696 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7264
timestamp 1666464484
transform -1 0 33696 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7265
timestamp 1666464484
transform -1 0 33696 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7266
timestamp 1666464484
transform -1 0 33696 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7267
timestamp 1666464484
transform -1 0 33696 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7268
timestamp 1666464484
transform -1 0 33696 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7269
timestamp 1666464484
transform -1 0 33696 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7270
timestamp 1666464484
transform -1 0 33696 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7271
timestamp 1666464484
transform -1 0 33696 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7272
timestamp 1666464484
transform -1 0 33696 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7273
timestamp 1666464484
transform -1 0 33696 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7274
timestamp 1666464484
transform -1 0 31200 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7275
timestamp 1666464484
transform -1 0 31200 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7276
timestamp 1666464484
transform 1 0 31200 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7277
timestamp 1666464484
transform -1 0 31200 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7278
timestamp 1666464484
transform -1 0 32448 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7279
timestamp 1666464484
transform -1 0 32448 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7280
timestamp 1666464484
transform -1 0 32448 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7281
timestamp 1666464484
transform -1 0 32448 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7282
timestamp 1666464484
transform -1 0 32448 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7283
timestamp 1666464484
transform -1 0 32448 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7284
timestamp 1666464484
transform -1 0 32448 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7285
timestamp 1666464484
transform -1 0 32448 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7286
timestamp 1666464484
transform -1 0 32448 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7287
timestamp 1666464484
transform -1 0 32448 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7288
timestamp 1666464484
transform -1 0 32448 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7289
timestamp 1666464484
transform -1 0 32448 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7290
timestamp 1666464484
transform -1 0 31200 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7291
timestamp 1666464484
transform -1 0 31200 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7292
timestamp 1666464484
transform -1 0 32448 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7293
timestamp 1666464484
transform -1 0 32448 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7294
timestamp 1666464484
transform -1 0 31200 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7295
timestamp 1666464484
transform 1 0 32448 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7296
timestamp 1666464484
transform 1 0 32448 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7297
timestamp 1666464484
transform 1 0 32448 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7298
timestamp 1666464484
transform 1 0 32448 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7299
timestamp 1666464484
transform 1 0 32448 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7300
timestamp 1666464484
transform 1 0 32448 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7301
timestamp 1666464484
transform 1 0 32448 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7302
timestamp 1666464484
transform 1 0 32448 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7303
timestamp 1666464484
transform 1 0 32448 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7304
timestamp 1666464484
transform 1 0 32448 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7305
timestamp 1666464484
transform 1 0 32448 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7306
timestamp 1666464484
transform 1 0 32448 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7307
timestamp 1666464484
transform 1 0 32448 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7308
timestamp 1666464484
transform 1 0 32448 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7309
timestamp 1666464484
transform 1 0 33696 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7310
timestamp 1666464484
transform 1 0 33696 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7311
timestamp 1666464484
transform 1 0 33696 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7312
timestamp 1666464484
transform 1 0 33696 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7313
timestamp 1666464484
transform 1 0 33696 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7314
timestamp 1666464484
transform 1 0 33696 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7315
timestamp 1666464484
transform 1 0 33696 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7316
timestamp 1666464484
transform 1 0 33696 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7317
timestamp 1666464484
transform 1 0 33696 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7318
timestamp 1666464484
transform 1 0 33696 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7319
timestamp 1666464484
transform 1 0 33696 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7320
timestamp 1666464484
transform 1 0 33696 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7321
timestamp 1666464484
transform 1 0 33696 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7322
timestamp 1666464484
transform 1 0 33696 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7323
timestamp 1666464484
transform -1 0 31200 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7324
timestamp 1666464484
transform -1 0 31200 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7325
timestamp 1666464484
transform -1 0 31200 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7326
timestamp 1666464484
transform -1 0 31200 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7327
timestamp 1666464484
transform -1 0 31200 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7328
timestamp 1666464484
transform -1 0 31200 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7329
timestamp 1666464484
transform 1 0 31200 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7330
timestamp 1666464484
transform 1 0 31200 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7331
timestamp 1666464484
transform 1 0 31200 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7332
timestamp 1666464484
transform 1 0 31200 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7333
timestamp 1666464484
transform 1 0 31200 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7334
timestamp 1666464484
transform 1 0 31200 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7335
timestamp 1666464484
transform 1 0 31200 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7336
timestamp 1666464484
transform 1 0 31200 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7337
timestamp 1666464484
transform 1 0 31200 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7338
timestamp 1666464484
transform 1 0 31200 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7339
timestamp 1666464484
transform 1 0 31200 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7340
timestamp 1666464484
transform 1 0 31200 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7341
timestamp 1666464484
transform -1 0 31200 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7342
timestamp 1666464484
transform -1 0 31200 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7343
timestamp 1666464484
transform 1 0 31200 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7344
timestamp 1666464484
transform -1 0 33696 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7345
timestamp 1666464484
transform -1 0 32448 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7346
timestamp 1666464484
transform -1 0 32448 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7347
timestamp 1666464484
transform -1 0 32448 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7348
timestamp 1666464484
transform -1 0 31200 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7349
timestamp 1666464484
transform -1 0 31200 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7350
timestamp 1666464484
transform -1 0 32448 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7351
timestamp 1666464484
transform -1 0 32448 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7352
timestamp 1666464484
transform -1 0 32448 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7353
timestamp 1666464484
transform -1 0 32448 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7354
timestamp 1666464484
transform -1 0 32448 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7355
timestamp 1666464484
transform -1 0 32448 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7356
timestamp 1666464484
transform -1 0 32448 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7357
timestamp 1666464484
transform -1 0 32448 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7358
timestamp 1666464484
transform -1 0 31200 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7359
timestamp 1666464484
transform -1 0 31200 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7360
timestamp 1666464484
transform 1 0 31200 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7361
timestamp 1666464484
transform 1 0 31200 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7362
timestamp 1666464484
transform -1 0 31200 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7363
timestamp 1666464484
transform -1 0 31200 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7364
timestamp 1666464484
transform 1 0 31200 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7365
timestamp 1666464484
transform 1 0 31200 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7366
timestamp 1666464484
transform 1 0 31200 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7367
timestamp 1666464484
transform 1 0 31200 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7368
timestamp 1666464484
transform 1 0 31200 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7369
timestamp 1666464484
transform -1 0 31200 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7370
timestamp 1666464484
transform -1 0 31200 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7371
timestamp 1666464484
transform 1 0 31200 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7372
timestamp 1666464484
transform 1 0 31200 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7373
timestamp 1666464484
transform 1 0 31200 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7374
timestamp 1666464484
transform 1 0 33696 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7375
timestamp 1666464484
transform 1 0 33696 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7376
timestamp 1666464484
transform 1 0 33696 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7377
timestamp 1666464484
transform 1 0 33696 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7378
timestamp 1666464484
transform 1 0 33696 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7379
timestamp 1666464484
transform 1 0 33696 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7380
timestamp 1666464484
transform 1 0 33696 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7381
timestamp 1666464484
transform -1 0 31200 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7382
timestamp 1666464484
transform -1 0 31200 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7383
timestamp 1666464484
transform 1 0 33696 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7384
timestamp 1666464484
transform 1 0 33696 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7385
timestamp 1666464484
transform 1 0 33696 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7386
timestamp 1666464484
transform 1 0 33696 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7387
timestamp 1666464484
transform 1 0 33696 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7388
timestamp 1666464484
transform 1 0 33696 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7389
timestamp 1666464484
transform 1 0 33696 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7390
timestamp 1666464484
transform 1 0 33696 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7391
timestamp 1666464484
transform 1 0 31200 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7392
timestamp 1666464484
transform 1 0 31200 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7393
timestamp 1666464484
transform -1 0 33696 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7394
timestamp 1666464484
transform -1 0 33696 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7395
timestamp 1666464484
transform -1 0 33696 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7396
timestamp 1666464484
transform -1 0 33696 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7397
timestamp 1666464484
transform -1 0 33696 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7398
timestamp 1666464484
transform -1 0 33696 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7399
timestamp 1666464484
transform -1 0 33696 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7400
timestamp 1666464484
transform -1 0 31200 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7401
timestamp 1666464484
transform -1 0 31200 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7402
timestamp 1666464484
transform -1 0 33696 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7403
timestamp 1666464484
transform -1 0 33696 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7404
timestamp 1666464484
transform -1 0 33696 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7405
timestamp 1666464484
transform -1 0 33696 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7406
timestamp 1666464484
transform -1 0 33696 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7407
timestamp 1666464484
transform -1 0 33696 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7408
timestamp 1666464484
transform -1 0 33696 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7409
timestamp 1666464484
transform -1 0 33696 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7410
timestamp 1666464484
transform 1 0 31200 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7411
timestamp 1666464484
transform 1 0 31200 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7412
timestamp 1666464484
transform 1 0 32448 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7413
timestamp 1666464484
transform 1 0 32448 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7414
timestamp 1666464484
transform 1 0 32448 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7415
timestamp 1666464484
transform 1 0 32448 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7416
timestamp 1666464484
transform 1 0 32448 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7417
timestamp 1666464484
transform 1 0 32448 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7418
timestamp 1666464484
transform 1 0 32448 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7419
timestamp 1666464484
transform -1 0 31200 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7420
timestamp 1666464484
transform -1 0 31200 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7421
timestamp 1666464484
transform 1 0 32448 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7422
timestamp 1666464484
transform 1 0 32448 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7423
timestamp 1666464484
transform 1 0 32448 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7424
timestamp 1666464484
transform 1 0 32448 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7425
timestamp 1666464484
transform 1 0 32448 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7426
timestamp 1666464484
transform 1 0 32448 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7427
timestamp 1666464484
transform 1 0 32448 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7428
timestamp 1666464484
transform 1 0 32448 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7429
timestamp 1666464484
transform 1 0 31200 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7430
timestamp 1666464484
transform -1 0 31200 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7431
timestamp 1666464484
transform -1 0 32448 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7432
timestamp 1666464484
transform -1 0 32448 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7433
timestamp 1666464484
transform -1 0 32448 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7434
timestamp 1666464484
transform -1 0 32448 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7435
timestamp 1666464484
transform 1 0 38688 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7436
timestamp 1666464484
transform 1 0 38688 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7437
timestamp 1666464484
transform -1 0 38688 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7438
timestamp 1666464484
transform -1 0 38688 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7439
timestamp 1666464484
transform -1 0 38688 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7440
timestamp 1666464484
transform -1 0 38688 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7441
timestamp 1666464484
transform -1 0 38688 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7442
timestamp 1666464484
transform -1 0 38688 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7443
timestamp 1666464484
transform 1 0 38688 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7444
timestamp 1666464484
transform -1 0 39936 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7445
timestamp 1666464484
transform -1 0 39936 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7446
timestamp 1666464484
transform -1 0 39936 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7447
timestamp 1666464484
transform -1 0 39936 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7448
timestamp 1666464484
transform -1 0 39936 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7449
timestamp 1666464484
transform -1 0 39936 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7450
timestamp 1666464484
transform 1 0 38688 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7451
timestamp 1666464484
transform 1 0 38688 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7452
timestamp 1666464484
transform 1 0 38688 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7453
timestamp 1666464484
transform -1 0 36192 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7454
timestamp 1666464484
transform -1 0 36192 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7455
timestamp 1666464484
transform 1 0 36192 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7456
timestamp 1666464484
transform 1 0 36192 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7457
timestamp 1666464484
transform 1 0 36192 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7458
timestamp 1666464484
transform 1 0 36192 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7459
timestamp 1666464484
transform -1 0 36192 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7460
timestamp 1666464484
transform -1 0 36192 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7461
timestamp 1666464484
transform -1 0 36192 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7462
timestamp 1666464484
transform -1 0 36192 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7463
timestamp 1666464484
transform 1 0 36192 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7464
timestamp 1666464484
transform 1 0 36192 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7465
timestamp 1666464484
transform 1 0 36192 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7466
timestamp 1666464484
transform 1 0 36192 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7467
timestamp 1666464484
transform 1 0 36192 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7468
timestamp 1666464484
transform 1 0 36192 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7469
timestamp 1666464484
transform -1 0 36192 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7470
timestamp 1666464484
transform -1 0 36192 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7471
timestamp 1666464484
transform -1 0 36192 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7472
timestamp 1666464484
transform -1 0 36192 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7473
timestamp 1666464484
transform -1 0 36192 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7474
timestamp 1666464484
transform -1 0 36192 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7475
timestamp 1666464484
transform -1 0 36192 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7476
timestamp 1666464484
transform 1 0 36192 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7477
timestamp 1666464484
transform 1 0 36192 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7478
timestamp 1666464484
transform 1 0 36192 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7479
timestamp 1666464484
transform -1 0 39936 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7480
timestamp 1666464484
transform -1 0 39936 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7481
timestamp 1666464484
transform -1 0 39936 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7482
timestamp 1666464484
transform -1 0 39936 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7483
timestamp 1666464484
transform -1 0 39936 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7484
timestamp 1666464484
transform -1 0 39936 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7485
timestamp 1666464484
transform -1 0 39936 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7486
timestamp 1666464484
transform -1 0 38688 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7487
timestamp 1666464484
transform -1 0 38688 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7488
timestamp 1666464484
transform 1 0 38688 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7489
timestamp 1666464484
transform 1 0 38688 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7490
timestamp 1666464484
transform 1 0 38688 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7491
timestamp 1666464484
transform 1 0 38688 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7492
timestamp 1666464484
transform 1 0 38688 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7493
timestamp 1666464484
transform 1 0 38688 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7494
timestamp 1666464484
transform 1 0 38688 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7495
timestamp 1666464484
transform -1 0 38688 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7496
timestamp 1666464484
transform -1 0 38688 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7497
timestamp 1666464484
transform -1 0 38688 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7498
timestamp 1666464484
transform -1 0 38688 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7499
timestamp 1666464484
transform -1 0 38688 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7500
timestamp 1666464484
transform -1 0 39936 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7501
timestamp 1666464484
transform -1 0 39936 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7502
timestamp 1666464484
transform 1 0 38688 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7503
timestamp 1666464484
transform 1 0 38688 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7504
timestamp 1666464484
transform -1 0 38688 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7505
timestamp 1666464484
transform -1 0 38688 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7506
timestamp 1666464484
transform -1 0 36192 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7507
timestamp 1666464484
transform -1 0 36192 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7508
timestamp 1666464484
transform 1 0 37440 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7509
timestamp 1666464484
transform 1 0 37440 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7510
timestamp 1666464484
transform 1 0 37440 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7511
timestamp 1666464484
transform 1 0 37440 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7512
timestamp 1666464484
transform 1 0 37440 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7513
timestamp 1666464484
transform 1 0 37440 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7514
timestamp 1666464484
transform 1 0 37440 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7515
timestamp 1666464484
transform 1 0 37440 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7516
timestamp 1666464484
transform 1 0 37440 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7517
timestamp 1666464484
transform 1 0 37440 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7518
timestamp 1666464484
transform 1 0 37440 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7519
timestamp 1666464484
transform 1 0 37440 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7520
timestamp 1666464484
transform 1 0 37440 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7521
timestamp 1666464484
transform 1 0 37440 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7522
timestamp 1666464484
transform 1 0 37440 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7523
timestamp 1666464484
transform -1 0 37440 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7524
timestamp 1666464484
transform -1 0 37440 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7525
timestamp 1666464484
transform -1 0 37440 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7526
timestamp 1666464484
transform -1 0 37440 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7527
timestamp 1666464484
transform -1 0 37440 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7528
timestamp 1666464484
transform -1 0 37440 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7529
timestamp 1666464484
transform -1 0 37440 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7530
timestamp 1666464484
transform -1 0 37440 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7531
timestamp 1666464484
transform -1 0 37440 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7532
timestamp 1666464484
transform -1 0 37440 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7533
timestamp 1666464484
transform -1 0 37440 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7534
timestamp 1666464484
transform -1 0 37440 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7535
timestamp 1666464484
transform -1 0 37440 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7536
timestamp 1666464484
transform -1 0 37440 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7537
timestamp 1666464484
transform -1 0 37440 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7538
timestamp 1666464484
transform 1 0 36192 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7539
timestamp 1666464484
transform 1 0 36192 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7540
timestamp 1666464484
transform -1 0 39936 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7541
timestamp 1666464484
transform -1 0 39936 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7542
timestamp 1666464484
transform 1 0 38688 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7543
timestamp 1666464484
transform 1 0 38688 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7544
timestamp 1666464484
transform -1 0 38688 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7545
timestamp 1666464484
transform -1 0 38688 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7546
timestamp 1666464484
transform 1 0 37440 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7547
timestamp 1666464484
transform 1 0 37440 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7548
timestamp 1666464484
transform -1 0 37440 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7549
timestamp 1666464484
transform -1 0 37440 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7550
timestamp 1666464484
transform 1 0 36192 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7551
timestamp 1666464484
transform 1 0 36192 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7552
timestamp 1666464484
transform -1 0 36192 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7553
timestamp 1666464484
transform -1 0 36192 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7554
timestamp 1666464484
transform -1 0 31200 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7555
timestamp 1666464484
transform -1 0 31200 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7556
timestamp 1666464484
transform 1 0 34944 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7557
timestamp 1666464484
transform 1 0 34944 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7558
timestamp 1666464484
transform 1 0 34944 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7559
timestamp 1666464484
transform 1 0 34944 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7560
timestamp 1666464484
transform 1 0 34944 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7561
timestamp 1666464484
transform 1 0 34944 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7562
timestamp 1666464484
transform 1 0 34944 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7563
timestamp 1666464484
transform 1 0 34944 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7564
timestamp 1666464484
transform 1 0 34944 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7565
timestamp 1666464484
transform 1 0 34944 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7566
timestamp 1666464484
transform 1 0 34944 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7567
timestamp 1666464484
transform 1 0 34944 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7568
timestamp 1666464484
transform 1 0 34944 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7569
timestamp 1666464484
transform 1 0 34944 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7570
timestamp 1666464484
transform 1 0 34944 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7571
timestamp 1666464484
transform 1 0 34944 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7572
timestamp 1666464484
transform 1 0 34944 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7573
timestamp 1666464484
transform 1 0 34944 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7574
timestamp 1666464484
transform 1 0 34944 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7575
timestamp 1666464484
transform 1 0 34944 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7576
timestamp 1666464484
transform 1 0 34944 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7577
timestamp 1666464484
transform 1 0 34944 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7578
timestamp 1666464484
transform 1 0 34944 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7579
timestamp 1666464484
transform 1 0 34944 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7580
timestamp 1666464484
transform 1 0 34944 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7581
timestamp 1666464484
transform 1 0 34944 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7582
timestamp 1666464484
transform 1 0 34944 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7583
timestamp 1666464484
transform 1 0 34944 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7584
timestamp 1666464484
transform 1 0 34944 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7585
timestamp 1666464484
transform 1 0 34944 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7586
timestamp 1666464484
transform 1 0 34944 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7587
timestamp 1666464484
transform -1 0 34944 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7588
timestamp 1666464484
transform -1 0 34944 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7589
timestamp 1666464484
transform -1 0 34944 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7590
timestamp 1666464484
transform -1 0 34944 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7591
timestamp 1666464484
transform -1 0 34944 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7592
timestamp 1666464484
transform -1 0 34944 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7593
timestamp 1666464484
transform -1 0 34944 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7594
timestamp 1666464484
transform -1 0 34944 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7595
timestamp 1666464484
transform -1 0 34944 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7596
timestamp 1666464484
transform -1 0 34944 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7597
timestamp 1666464484
transform -1 0 34944 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7598
timestamp 1666464484
transform -1 0 34944 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7599
timestamp 1666464484
transform -1 0 34944 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7600
timestamp 1666464484
transform -1 0 34944 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7601
timestamp 1666464484
transform -1 0 34944 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7602
timestamp 1666464484
transform -1 0 34944 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7603
timestamp 1666464484
transform -1 0 34944 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7604
timestamp 1666464484
transform -1 0 34944 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7605
timestamp 1666464484
transform -1 0 34944 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7606
timestamp 1666464484
transform -1 0 34944 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7607
timestamp 1666464484
transform -1 0 34944 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7608
timestamp 1666464484
transform -1 0 34944 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7609
timestamp 1666464484
transform -1 0 34944 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7610
timestamp 1666464484
transform -1 0 34944 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7611
timestamp 1666464484
transform -1 0 34944 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7612
timestamp 1666464484
transform -1 0 34944 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7613
timestamp 1666464484
transform -1 0 34944 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7614
timestamp 1666464484
transform -1 0 34944 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7615
timestamp 1666464484
transform -1 0 34944 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7616
timestamp 1666464484
transform -1 0 34944 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7617
timestamp 1666464484
transform -1 0 34944 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7618
timestamp 1666464484
transform 1 0 33696 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7619
timestamp 1666464484
transform 1 0 33696 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7620
timestamp 1666464484
transform -1 0 33696 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7621
timestamp 1666464484
transform -1 0 33696 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7622
timestamp 1666464484
transform 1 0 32448 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7623
timestamp 1666464484
transform 1 0 32448 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7624
timestamp 1666464484
transform -1 0 32448 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7625
timestamp 1666464484
transform -1 0 32448 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7626
timestamp 1666464484
transform 1 0 31200 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7627
timestamp 1666464484
transform 1 0 31200 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7628
timestamp 1666464484
transform -1 0 39936 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7629
timestamp 1666464484
transform -1 0 39936 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7630
timestamp 1666464484
transform 1 0 38688 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7631
timestamp 1666464484
transform 1 0 38688 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7632
timestamp 1666464484
transform -1 0 38688 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7633
timestamp 1666464484
transform -1 0 38688 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7634
timestamp 1666464484
transform 1 0 37440 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7635
timestamp 1666464484
transform 1 0 37440 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7636
timestamp 1666464484
transform -1 0 37440 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7637
timestamp 1666464484
transform -1 0 37440 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7638
timestamp 1666464484
transform 1 0 36192 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7639
timestamp 1666464484
transform 1 0 36192 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7640
timestamp 1666464484
transform -1 0 36192 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7641
timestamp 1666464484
transform -1 0 36192 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7642
timestamp 1666464484
transform 1 0 34944 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7643
timestamp 1666464484
transform 1 0 34944 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7644
timestamp 1666464484
transform -1 0 34944 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7645
timestamp 1666464484
transform -1 0 34944 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7646
timestamp 1666464484
transform 1 0 33696 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7647
timestamp 1666464484
transform 1 0 33696 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7648
timestamp 1666464484
transform -1 0 33696 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7649
timestamp 1666464484
transform -1 0 33696 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7650
timestamp 1666464484
transform 1 0 32448 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7651
timestamp 1666464484
transform 1 0 32448 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7652
timestamp 1666464484
transform -1 0 32448 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7653
timestamp 1666464484
transform -1 0 32448 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7654
timestamp 1666464484
transform 1 0 31200 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7655
timestamp 1666464484
transform 1 0 31200 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7656
timestamp 1666464484
transform -1 0 31200 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7657
timestamp 1666464484
transform -1 0 31200 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7658
timestamp 1666464484
transform -1 0 21216 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7659
timestamp 1666464484
transform -1 0 21216 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7660
timestamp 1666464484
transform 1 0 29952 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7661
timestamp 1666464484
transform 1 0 29952 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7662
timestamp 1666464484
transform 1 0 29952 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7663
timestamp 1666464484
transform 1 0 29952 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7664
timestamp 1666464484
transform 1 0 29952 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7665
timestamp 1666464484
transform 1 0 29952 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7666
timestamp 1666464484
transform 1 0 29952 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7667
timestamp 1666464484
transform 1 0 29952 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7668
timestamp 1666464484
transform 1 0 29952 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7669
timestamp 1666464484
transform 1 0 29952 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7670
timestamp 1666464484
transform 1 0 29952 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7671
timestamp 1666464484
transform 1 0 29952 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7672
timestamp 1666464484
transform 1 0 29952 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7673
timestamp 1666464484
transform 1 0 29952 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7674
timestamp 1666464484
transform 1 0 29952 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7675
timestamp 1666464484
transform 1 0 29952 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7676
timestamp 1666464484
transform 1 0 29952 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7677
timestamp 1666464484
transform 1 0 29952 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7678
timestamp 1666464484
transform 1 0 29952 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7679
timestamp 1666464484
transform 1 0 29952 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7680
timestamp 1666464484
transform 1 0 29952 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7681
timestamp 1666464484
transform 1 0 29952 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7682
timestamp 1666464484
transform 1 0 29952 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7683
timestamp 1666464484
transform 1 0 29952 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7684
timestamp 1666464484
transform 1 0 29952 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7685
timestamp 1666464484
transform 1 0 29952 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7686
timestamp 1666464484
transform 1 0 29952 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7687
timestamp 1666464484
transform 1 0 29952 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7688
timestamp 1666464484
transform 1 0 29952 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7689
timestamp 1666464484
transform 1 0 29952 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7690
timestamp 1666464484
transform 1 0 29952 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7691
timestamp 1666464484
transform 1 0 29952 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7692
timestamp 1666464484
transform 1 0 29952 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7693
timestamp 1666464484
transform 1 0 29952 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7694
timestamp 1666464484
transform 1 0 29952 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7695
timestamp 1666464484
transform 1 0 29952 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7696
timestamp 1666464484
transform 1 0 29952 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7697
timestamp 1666464484
transform 1 0 29952 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7698
timestamp 1666464484
transform 1 0 29952 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7699
timestamp 1666464484
transform 1 0 29952 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7700
timestamp 1666464484
transform 1 0 29952 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7701
timestamp 1666464484
transform 1 0 29952 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7702
timestamp 1666464484
transform 1 0 29952 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7703
timestamp 1666464484
transform 1 0 29952 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7704
timestamp 1666464484
transform 1 0 29952 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7705
timestamp 1666464484
transform 1 0 29952 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7706
timestamp 1666464484
transform 1 0 29952 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7707
timestamp 1666464484
transform 1 0 29952 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7708
timestamp 1666464484
transform 1 0 29952 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7709
timestamp 1666464484
transform 1 0 29952 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7710
timestamp 1666464484
transform 1 0 29952 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7711
timestamp 1666464484
transform 1 0 29952 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7712
timestamp 1666464484
transform 1 0 29952 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7713
timestamp 1666464484
transform 1 0 29952 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7714
timestamp 1666464484
transform 1 0 29952 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7715
timestamp 1666464484
transform 1 0 29952 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7716
timestamp 1666464484
transform 1 0 29952 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7717
timestamp 1666464484
transform 1 0 29952 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7718
timestamp 1666464484
transform 1 0 29952 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7719
timestamp 1666464484
transform 1 0 29952 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7720
timestamp 1666464484
transform 1 0 29952 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7721
timestamp 1666464484
transform 1 0 29952 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7722
timestamp 1666464484
transform 1 0 29952 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7723
timestamp 1666464484
transform -1 0 29952 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7724
timestamp 1666464484
transform -1 0 29952 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7725
timestamp 1666464484
transform -1 0 29952 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7726
timestamp 1666464484
transform -1 0 29952 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7727
timestamp 1666464484
transform -1 0 29952 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7728
timestamp 1666464484
transform -1 0 29952 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7729
timestamp 1666464484
transform -1 0 29952 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7730
timestamp 1666464484
transform -1 0 29952 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7731
timestamp 1666464484
transform -1 0 29952 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7732
timestamp 1666464484
transform -1 0 29952 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7733
timestamp 1666464484
transform -1 0 29952 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7734
timestamp 1666464484
transform -1 0 29952 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7735
timestamp 1666464484
transform -1 0 29952 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7736
timestamp 1666464484
transform -1 0 29952 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7737
timestamp 1666464484
transform -1 0 29952 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7738
timestamp 1666464484
transform -1 0 29952 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7739
timestamp 1666464484
transform -1 0 29952 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7740
timestamp 1666464484
transform -1 0 29952 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7741
timestamp 1666464484
transform -1 0 29952 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7742
timestamp 1666464484
transform -1 0 29952 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7743
timestamp 1666464484
transform -1 0 29952 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7744
timestamp 1666464484
transform -1 0 29952 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7745
timestamp 1666464484
transform -1 0 29952 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7746
timestamp 1666464484
transform -1 0 29952 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7747
timestamp 1666464484
transform -1 0 29952 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7748
timestamp 1666464484
transform -1 0 29952 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7749
timestamp 1666464484
transform -1 0 29952 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7750
timestamp 1666464484
transform -1 0 29952 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7751
timestamp 1666464484
transform -1 0 29952 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7752
timestamp 1666464484
transform -1 0 29952 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7753
timestamp 1666464484
transform -1 0 29952 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7754
timestamp 1666464484
transform -1 0 29952 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7755
timestamp 1666464484
transform -1 0 29952 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7756
timestamp 1666464484
transform -1 0 29952 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7757
timestamp 1666464484
transform -1 0 29952 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7758
timestamp 1666464484
transform -1 0 29952 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7759
timestamp 1666464484
transform -1 0 29952 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7760
timestamp 1666464484
transform -1 0 29952 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7761
timestamp 1666464484
transform -1 0 29952 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7762
timestamp 1666464484
transform -1 0 29952 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7763
timestamp 1666464484
transform -1 0 29952 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7764
timestamp 1666464484
transform -1 0 29952 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7765
timestamp 1666464484
transform -1 0 29952 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7766
timestamp 1666464484
transform -1 0 29952 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7767
timestamp 1666464484
transform -1 0 29952 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7768
timestamp 1666464484
transform -1 0 29952 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7769
timestamp 1666464484
transform -1 0 29952 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7770
timestamp 1666464484
transform -1 0 29952 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7771
timestamp 1666464484
transform -1 0 29952 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7772
timestamp 1666464484
transform -1 0 29952 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7773
timestamp 1666464484
transform -1 0 29952 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7774
timestamp 1666464484
transform -1 0 29952 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7775
timestamp 1666464484
transform -1 0 29952 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7776
timestamp 1666464484
transform -1 0 29952 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7777
timestamp 1666464484
transform -1 0 29952 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7778
timestamp 1666464484
transform -1 0 29952 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7779
timestamp 1666464484
transform -1 0 29952 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7780
timestamp 1666464484
transform -1 0 29952 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7781
timestamp 1666464484
transform -1 0 29952 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7782
timestamp 1666464484
transform -1 0 29952 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7783
timestamp 1666464484
transform -1 0 29952 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7784
timestamp 1666464484
transform -1 0 29952 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7785
timestamp 1666464484
transform -1 0 29952 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7786
timestamp 1666464484
transform 1 0 28704 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7787
timestamp 1666464484
transform 1 0 28704 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7788
timestamp 1666464484
transform -1 0 28704 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7789
timestamp 1666464484
transform -1 0 28704 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7790
timestamp 1666464484
transform 1 0 27456 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7791
timestamp 1666464484
transform 1 0 27456 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7792
timestamp 1666464484
transform -1 0 27456 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7793
timestamp 1666464484
transform -1 0 27456 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7794
timestamp 1666464484
transform 1 0 26208 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7795
timestamp 1666464484
transform 1 0 26208 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7796
timestamp 1666464484
transform -1 0 26208 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7797
timestamp 1666464484
transform -1 0 26208 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7798
timestamp 1666464484
transform 1 0 24960 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7799
timestamp 1666464484
transform 1 0 24960 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7800
timestamp 1666464484
transform -1 0 24960 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7801
timestamp 1666464484
transform -1 0 24960 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7802
timestamp 1666464484
transform 1 0 23712 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7803
timestamp 1666464484
transform 1 0 23712 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7804
timestamp 1666464484
transform -1 0 23712 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7805
timestamp 1666464484
transform -1 0 23712 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7806
timestamp 1666464484
transform 1 0 22464 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7807
timestamp 1666464484
transform 1 0 22464 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7808
timestamp 1666464484
transform -1 0 22464 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7809
timestamp 1666464484
transform -1 0 22464 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7810
timestamp 1666464484
transform 1 0 21216 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7811
timestamp 1666464484
transform 1 0 21216 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7812
timestamp 1666464484
transform -1 0 39936 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7813
timestamp 1666464484
transform -1 0 39936 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7814
timestamp 1666464484
transform 1 0 38688 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7815
timestamp 1666464484
transform 1 0 38688 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7816
timestamp 1666464484
transform -1 0 38688 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7817
timestamp 1666464484
transform -1 0 38688 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7818
timestamp 1666464484
transform 1 0 37440 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7819
timestamp 1666464484
transform 1 0 37440 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7820
timestamp 1666464484
transform -1 0 37440 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7821
timestamp 1666464484
transform -1 0 37440 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7822
timestamp 1666464484
transform 1 0 36192 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7823
timestamp 1666464484
transform 1 0 36192 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7824
timestamp 1666464484
transform -1 0 36192 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7825
timestamp 1666464484
transform -1 0 36192 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7826
timestamp 1666464484
transform 1 0 34944 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7827
timestamp 1666464484
transform 1 0 34944 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7828
timestamp 1666464484
transform -1 0 34944 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7829
timestamp 1666464484
transform -1 0 34944 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7830
timestamp 1666464484
transform 1 0 33696 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7831
timestamp 1666464484
transform 1 0 33696 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7832
timestamp 1666464484
transform -1 0 33696 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7833
timestamp 1666464484
transform -1 0 33696 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7834
timestamp 1666464484
transform 1 0 32448 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7835
timestamp 1666464484
transform 1 0 32448 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7836
timestamp 1666464484
transform -1 0 32448 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7837
timestamp 1666464484
transform -1 0 32448 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7838
timestamp 1666464484
transform 1 0 31200 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7839
timestamp 1666464484
transform 1 0 31200 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7840
timestamp 1666464484
transform -1 0 31200 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7841
timestamp 1666464484
transform -1 0 31200 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7842
timestamp 1666464484
transform 1 0 29952 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7843
timestamp 1666464484
transform 1 0 29952 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7844
timestamp 1666464484
transform -1 0 29952 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7845
timestamp 1666464484
transform -1 0 29952 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7846
timestamp 1666464484
transform 1 0 28704 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7847
timestamp 1666464484
transform 1 0 28704 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7848
timestamp 1666464484
transform -1 0 28704 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7849
timestamp 1666464484
transform -1 0 28704 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7850
timestamp 1666464484
transform 1 0 27456 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7851
timestamp 1666464484
transform 1 0 27456 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7852
timestamp 1666464484
transform -1 0 27456 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7853
timestamp 1666464484
transform -1 0 27456 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7854
timestamp 1666464484
transform 1 0 26208 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7855
timestamp 1666464484
transform 1 0 26208 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7856
timestamp 1666464484
transform -1 0 26208 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7857
timestamp 1666464484
transform -1 0 26208 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7858
timestamp 1666464484
transform 1 0 24960 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7859
timestamp 1666464484
transform 1 0 24960 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7860
timestamp 1666464484
transform -1 0 24960 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7861
timestamp 1666464484
transform -1 0 24960 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7862
timestamp 1666464484
transform 1 0 23712 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7863
timestamp 1666464484
transform 1 0 23712 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7864
timestamp 1666464484
transform -1 0 23712 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7865
timestamp 1666464484
transform -1 0 23712 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7866
timestamp 1666464484
transform 1 0 22464 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7867
timestamp 1666464484
transform 1 0 22464 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7868
timestamp 1666464484
transform -1 0 22464 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7869
timestamp 1666464484
transform -1 0 22464 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7870
timestamp 1666464484
transform 1 0 21216 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7871
timestamp 1666464484
transform 1 0 21216 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7872
timestamp 1666464484
transform -1 0 21216 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7873
timestamp 1666464484
transform -1 0 21216 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7874
timestamp 1666464484
transform 1 0 19968 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7875
timestamp 1666464484
transform 1 0 19968 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7876
timestamp 1666464484
transform 1 0 19968 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7877
timestamp 1666464484
transform 1 0 19968 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7878
timestamp 1666464484
transform 1 0 19968 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7879
timestamp 1666464484
transform 1 0 19968 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7880
timestamp 1666464484
transform 1 0 19968 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7881
timestamp 1666464484
transform 1 0 19968 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7882
timestamp 1666464484
transform 1 0 19968 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7883
timestamp 1666464484
transform 1 0 19968 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7884
timestamp 1666464484
transform 1 0 19968 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7885
timestamp 1666464484
transform 1 0 19968 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7886
timestamp 1666464484
transform 1 0 19968 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7887
timestamp 1666464484
transform 1 0 19968 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7888
timestamp 1666464484
transform 1 0 19968 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7889
timestamp 1666464484
transform 1 0 19968 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7890
timestamp 1666464484
transform 1 0 19968 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7891
timestamp 1666464484
transform 1 0 19968 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7892
timestamp 1666464484
transform 1 0 19968 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7893
timestamp 1666464484
transform 1 0 19968 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7894
timestamp 1666464484
transform 1 0 19968 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7895
timestamp 1666464484
transform 1 0 19968 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7896
timestamp 1666464484
transform 1 0 19968 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7897
timestamp 1666464484
transform 1 0 19968 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7898
timestamp 1666464484
transform 1 0 19968 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7899
timestamp 1666464484
transform 1 0 19968 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7900
timestamp 1666464484
transform 1 0 19968 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7901
timestamp 1666464484
transform 1 0 19968 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7902
timestamp 1666464484
transform 1 0 19968 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7903
timestamp 1666464484
transform 1 0 19968 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7904
timestamp 1666464484
transform 1 0 19968 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7905
timestamp 1666464484
transform 1 0 19968 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7906
timestamp 1666464484
transform 1 0 19968 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7907
timestamp 1666464484
transform 1 0 19968 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7908
timestamp 1666464484
transform 1 0 19968 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7909
timestamp 1666464484
transform 1 0 19968 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7910
timestamp 1666464484
transform 1 0 19968 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7911
timestamp 1666464484
transform 1 0 19968 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7912
timestamp 1666464484
transform 1 0 19968 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7913
timestamp 1666464484
transform 1 0 19968 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7914
timestamp 1666464484
transform 1 0 19968 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7915
timestamp 1666464484
transform 1 0 19968 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7916
timestamp 1666464484
transform 1 0 19968 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7917
timestamp 1666464484
transform 1 0 19968 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7918
timestamp 1666464484
transform 1 0 19968 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7919
timestamp 1666464484
transform 1 0 19968 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7920
timestamp 1666464484
transform 1 0 19968 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7921
timestamp 1666464484
transform 1 0 19968 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7922
timestamp 1666464484
transform 1 0 19968 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7923
timestamp 1666464484
transform 1 0 19968 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7924
timestamp 1666464484
transform 1 0 19968 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7925
timestamp 1666464484
transform 1 0 19968 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7926
timestamp 1666464484
transform 1 0 19968 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7927
timestamp 1666464484
transform 1 0 19968 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7928
timestamp 1666464484
transform 1 0 19968 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7929
timestamp 1666464484
transform 1 0 19968 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7930
timestamp 1666464484
transform 1 0 19968 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7931
timestamp 1666464484
transform 1 0 19968 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7932
timestamp 1666464484
transform 1 0 19968 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7933
timestamp 1666464484
transform 1 0 19968 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7934
timestamp 1666464484
transform 1 0 19968 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7935
timestamp 1666464484
transform 1 0 19968 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7936
timestamp 1666464484
transform 1 0 19968 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7937
timestamp 1666464484
transform 1 0 19968 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7938
timestamp 1666464484
transform 1 0 19968 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7939
timestamp 1666464484
transform 1 0 19968 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7940
timestamp 1666464484
transform 1 0 19968 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7941
timestamp 1666464484
transform 1 0 19968 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7942
timestamp 1666464484
transform 1 0 19968 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7943
timestamp 1666464484
transform 1 0 19968 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7944
timestamp 1666464484
transform 1 0 19968 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7945
timestamp 1666464484
transform 1 0 19968 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7946
timestamp 1666464484
transform 1 0 19968 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7947
timestamp 1666464484
transform 1 0 19968 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7948
timestamp 1666464484
transform 1 0 19968 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7949
timestamp 1666464484
transform 1 0 19968 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7950
timestamp 1666464484
transform 1 0 19968 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7951
timestamp 1666464484
transform 1 0 19968 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7952
timestamp 1666464484
transform 1 0 19968 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7953
timestamp 1666464484
transform 1 0 19968 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7954
timestamp 1666464484
transform 1 0 19968 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7955
timestamp 1666464484
transform 1 0 19968 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7956
timestamp 1666464484
transform 1 0 19968 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7957
timestamp 1666464484
transform 1 0 19968 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7958
timestamp 1666464484
transform 1 0 19968 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7959
timestamp 1666464484
transform 1 0 19968 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7960
timestamp 1666464484
transform 1 0 19968 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7961
timestamp 1666464484
transform 1 0 19968 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7962
timestamp 1666464484
transform 1 0 19968 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7963
timestamp 1666464484
transform 1 0 19968 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7964
timestamp 1666464484
transform 1 0 19968 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7965
timestamp 1666464484
transform 1 0 19968 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7966
timestamp 1666464484
transform 1 0 19968 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7967
timestamp 1666464484
transform 1 0 19968 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7968
timestamp 1666464484
transform 1 0 19968 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7969
timestamp 1666464484
transform 1 0 19968 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7970
timestamp 1666464484
transform 1 0 19968 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7971
timestamp 1666464484
transform 1 0 19968 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7972
timestamp 1666464484
transform 1 0 19968 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7973
timestamp 1666464484
transform 1 0 19968 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7974
timestamp 1666464484
transform 1 0 19968 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7975
timestamp 1666464484
transform 1 0 19968 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7976
timestamp 1666464484
transform 1 0 19968 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7977
timestamp 1666464484
transform 1 0 19968 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7978
timestamp 1666464484
transform 1 0 19968 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7979
timestamp 1666464484
transform 1 0 19968 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7980
timestamp 1666464484
transform 1 0 19968 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7981
timestamp 1666464484
transform 1 0 19968 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7982
timestamp 1666464484
transform 1 0 19968 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7983
timestamp 1666464484
transform 1 0 19968 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7984
timestamp 1666464484
transform 1 0 19968 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7985
timestamp 1666464484
transform 1 0 19968 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7986
timestamp 1666464484
transform 1 0 19968 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7987
timestamp 1666464484
transform 1 0 19968 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7988
timestamp 1666464484
transform 1 0 19968 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7989
timestamp 1666464484
transform 1 0 19968 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7990
timestamp 1666464484
transform 1 0 19968 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7991
timestamp 1666464484
transform 1 0 19968 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7992
timestamp 1666464484
transform 1 0 19968 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7993
timestamp 1666464484
transform 1 0 19968 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7994
timestamp 1666464484
transform 1 0 19968 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7995
timestamp 1666464484
transform 1 0 19968 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7996
timestamp 1666464484
transform 1 0 19968 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7997
timestamp 1666464484
transform 1 0 19968 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7998
timestamp 1666464484
transform 1 0 19968 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_7999
timestamp 1666464484
transform 1 0 19968 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8000
timestamp 1666464484
transform 1 0 19968 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8001
timestamp 1666464484
transform 1 0 19968 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8002
timestamp 1666464484
transform -1 0 19968 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8003
timestamp 1666464484
transform -1 0 19968 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8004
timestamp 1666464484
transform -1 0 19968 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8005
timestamp 1666464484
transform -1 0 19968 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8006
timestamp 1666464484
transform -1 0 19968 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8007
timestamp 1666464484
transform -1 0 19968 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8008
timestamp 1666464484
transform -1 0 19968 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8009
timestamp 1666464484
transform -1 0 19968 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8010
timestamp 1666464484
transform -1 0 19968 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8011
timestamp 1666464484
transform -1 0 19968 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8012
timestamp 1666464484
transform -1 0 19968 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8013
timestamp 1666464484
transform -1 0 19968 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8014
timestamp 1666464484
transform -1 0 19968 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8015
timestamp 1666464484
transform -1 0 19968 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8016
timestamp 1666464484
transform -1 0 19968 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8017
timestamp 1666464484
transform -1 0 19968 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8018
timestamp 1666464484
transform -1 0 19968 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8019
timestamp 1666464484
transform -1 0 19968 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8020
timestamp 1666464484
transform -1 0 19968 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8021
timestamp 1666464484
transform -1 0 19968 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8022
timestamp 1666464484
transform -1 0 19968 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8023
timestamp 1666464484
transform -1 0 19968 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8024
timestamp 1666464484
transform -1 0 19968 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8025
timestamp 1666464484
transform -1 0 19968 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8026
timestamp 1666464484
transform -1 0 19968 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8027
timestamp 1666464484
transform -1 0 19968 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8028
timestamp 1666464484
transform -1 0 19968 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8029
timestamp 1666464484
transform -1 0 19968 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8030
timestamp 1666464484
transform -1 0 19968 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8031
timestamp 1666464484
transform -1 0 19968 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8032
timestamp 1666464484
transform -1 0 19968 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8033
timestamp 1666464484
transform -1 0 19968 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8034
timestamp 1666464484
transform -1 0 19968 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8035
timestamp 1666464484
transform -1 0 19968 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8036
timestamp 1666464484
transform -1 0 19968 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8037
timestamp 1666464484
transform -1 0 19968 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8038
timestamp 1666464484
transform -1 0 19968 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8039
timestamp 1666464484
transform -1 0 19968 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8040
timestamp 1666464484
transform -1 0 19968 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8041
timestamp 1666464484
transform -1 0 19968 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8042
timestamp 1666464484
transform -1 0 19968 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8043
timestamp 1666464484
transform -1 0 19968 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8044
timestamp 1666464484
transform -1 0 19968 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8045
timestamp 1666464484
transform -1 0 19968 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8046
timestamp 1666464484
transform -1 0 19968 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8047
timestamp 1666464484
transform -1 0 19968 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8048
timestamp 1666464484
transform -1 0 19968 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8049
timestamp 1666464484
transform -1 0 19968 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8050
timestamp 1666464484
transform -1 0 19968 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8051
timestamp 1666464484
transform -1 0 19968 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8052
timestamp 1666464484
transform -1 0 19968 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8053
timestamp 1666464484
transform -1 0 19968 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8054
timestamp 1666464484
transform -1 0 19968 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8055
timestamp 1666464484
transform -1 0 19968 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8056
timestamp 1666464484
transform -1 0 19968 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8057
timestamp 1666464484
transform -1 0 19968 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8058
timestamp 1666464484
transform -1 0 19968 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8059
timestamp 1666464484
transform -1 0 19968 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8060
timestamp 1666464484
transform -1 0 19968 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8061
timestamp 1666464484
transform -1 0 19968 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8062
timestamp 1666464484
transform -1 0 19968 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8063
timestamp 1666464484
transform -1 0 19968 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8064
timestamp 1666464484
transform -1 0 19968 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8065
timestamp 1666464484
transform -1 0 19968 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8066
timestamp 1666464484
transform -1 0 19968 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8067
timestamp 1666464484
transform -1 0 19968 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8068
timestamp 1666464484
transform -1 0 19968 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8069
timestamp 1666464484
transform -1 0 19968 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8070
timestamp 1666464484
transform -1 0 19968 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8071
timestamp 1666464484
transform -1 0 19968 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8072
timestamp 1666464484
transform -1 0 19968 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8073
timestamp 1666464484
transform -1 0 19968 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8074
timestamp 1666464484
transform -1 0 19968 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8075
timestamp 1666464484
transform -1 0 19968 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8076
timestamp 1666464484
transform -1 0 19968 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8077
timestamp 1666464484
transform -1 0 19968 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8078
timestamp 1666464484
transform -1 0 19968 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8079
timestamp 1666464484
transform -1 0 19968 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8080
timestamp 1666464484
transform -1 0 19968 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8081
timestamp 1666464484
transform -1 0 19968 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8082
timestamp 1666464484
transform -1 0 19968 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8083
timestamp 1666464484
transform -1 0 19968 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8084
timestamp 1666464484
transform -1 0 19968 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8085
timestamp 1666464484
transform -1 0 19968 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8086
timestamp 1666464484
transform -1 0 19968 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8087
timestamp 1666464484
transform -1 0 19968 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8088
timestamp 1666464484
transform -1 0 19968 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8089
timestamp 1666464484
transform -1 0 19968 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8090
timestamp 1666464484
transform -1 0 19968 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8091
timestamp 1666464484
transform -1 0 19968 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8092
timestamp 1666464484
transform -1 0 19968 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8093
timestamp 1666464484
transform -1 0 19968 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8094
timestamp 1666464484
transform -1 0 19968 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8095
timestamp 1666464484
transform -1 0 19968 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8096
timestamp 1666464484
transform -1 0 19968 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8097
timestamp 1666464484
transform -1 0 19968 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8098
timestamp 1666464484
transform -1 0 19968 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8099
timestamp 1666464484
transform -1 0 19968 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8100
timestamp 1666464484
transform -1 0 19968 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8101
timestamp 1666464484
transform -1 0 19968 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8102
timestamp 1666464484
transform -1 0 19968 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8103
timestamp 1666464484
transform -1 0 19968 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8104
timestamp 1666464484
transform -1 0 19968 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8105
timestamp 1666464484
transform -1 0 19968 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8106
timestamp 1666464484
transform -1 0 19968 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8107
timestamp 1666464484
transform -1 0 19968 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8108
timestamp 1666464484
transform -1 0 19968 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8109
timestamp 1666464484
transform -1 0 19968 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8110
timestamp 1666464484
transform -1 0 19968 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8111
timestamp 1666464484
transform -1 0 19968 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8112
timestamp 1666464484
transform -1 0 19968 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8113
timestamp 1666464484
transform -1 0 19968 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8114
timestamp 1666464484
transform -1 0 19968 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8115
timestamp 1666464484
transform -1 0 19968 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8116
timestamp 1666464484
transform -1 0 19968 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8117
timestamp 1666464484
transform -1 0 19968 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8118
timestamp 1666464484
transform -1 0 19968 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8119
timestamp 1666464484
transform -1 0 19968 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8120
timestamp 1666464484
transform -1 0 19968 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8121
timestamp 1666464484
transform -1 0 19968 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8122
timestamp 1666464484
transform -1 0 19968 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8123
timestamp 1666464484
transform -1 0 19968 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8124
timestamp 1666464484
transform -1 0 19968 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8125
timestamp 1666464484
transform -1 0 19968 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8126
timestamp 1666464484
transform -1 0 19968 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8127
timestamp 1666464484
transform -1 0 19968 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8128
timestamp 1666464484
transform -1 0 19968 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8129
timestamp 1666464484
transform -1 0 19968 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8130
timestamp 1666464484
transform 1 0 18720 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8131
timestamp 1666464484
transform 1 0 18720 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8132
timestamp 1666464484
transform -1 0 18720 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8133
timestamp 1666464484
transform -1 0 18720 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8134
timestamp 1666464484
transform 1 0 17472 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8135
timestamp 1666464484
transform 1 0 17472 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8136
timestamp 1666464484
transform -1 0 17472 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8137
timestamp 1666464484
transform -1 0 17472 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8138
timestamp 1666464484
transform 1 0 16224 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8139
timestamp 1666464484
transform 1 0 16224 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8140
timestamp 1666464484
transform -1 0 16224 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8141
timestamp 1666464484
transform -1 0 16224 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8142
timestamp 1666464484
transform 1 0 14976 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8143
timestamp 1666464484
transform 1 0 14976 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8144
timestamp 1666464484
transform -1 0 14976 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8145
timestamp 1666464484
transform -1 0 14976 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8146
timestamp 1666464484
transform 1 0 13728 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8147
timestamp 1666464484
transform 1 0 13728 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8148
timestamp 1666464484
transform -1 0 13728 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8149
timestamp 1666464484
transform -1 0 13728 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8150
timestamp 1666464484
transform 1 0 12480 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8151
timestamp 1666464484
transform 1 0 12480 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8152
timestamp 1666464484
transform -1 0 12480 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8153
timestamp 1666464484
transform -1 0 12480 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8154
timestamp 1666464484
transform 1 0 11232 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8155
timestamp 1666464484
transform 1 0 11232 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8156
timestamp 1666464484
transform -1 0 11232 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8157
timestamp 1666464484
transform -1 0 11232 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8158
timestamp 1666464484
transform 1 0 9984 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8159
timestamp 1666464484
transform 1 0 9984 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8160
timestamp 1666464484
transform -1 0 9984 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8161
timestamp 1666464484
transform -1 0 9984 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8162
timestamp 1666464484
transform 1 0 8736 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8163
timestamp 1666464484
transform 1 0 8736 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8164
timestamp 1666464484
transform -1 0 8736 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8165
timestamp 1666464484
transform -1 0 8736 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8166
timestamp 1666464484
transform 1 0 7488 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8167
timestamp 1666464484
transform 1 0 7488 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8168
timestamp 1666464484
transform -1 0 7488 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8169
timestamp 1666464484
transform -1 0 7488 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8170
timestamp 1666464484
transform 1 0 6240 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8171
timestamp 1666464484
transform 1 0 6240 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8172
timestamp 1666464484
transform -1 0 6240 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8173
timestamp 1666464484
transform -1 0 6240 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8174
timestamp 1666464484
transform 1 0 4992 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8175
timestamp 1666464484
transform 1 0 4992 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8176
timestamp 1666464484
transform -1 0 4992 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8177
timestamp 1666464484
transform -1 0 4992 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8178
timestamp 1666464484
transform 1 0 3744 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8179
timestamp 1666464484
transform 1 0 3744 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8180
timestamp 1666464484
transform -1 0 3744 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8181
timestamp 1666464484
transform -1 0 3744 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8182
timestamp 1666464484
transform 1 0 2496 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8183
timestamp 1666464484
transform 1 0 2496 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8184
timestamp 1666464484
transform -1 0 2496 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8185
timestamp 1666464484
transform -1 0 2496 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8186
timestamp 1666464484
transform 1 0 1248 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8187
timestamp 1666464484
transform 1 0 1248 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8188
timestamp 1666464484
transform -1 0 1248 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8189
timestamp 1666464484
transform -1 0 1248 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8190
timestamp 1666464484
transform 1 0 0 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_1  sky130_fd_bd_sram__openram_dp_cell_8191
timestamp 1666464484
transform 1 0 0 0 -1 25280
box -42 -105 650 421
<< labels >>
rlabel metal1 s 37680 48439 37680 48439 4 vdd
port 513 nsew
rlabel metal1 s 37680 49229 37680 49229 4 vdd
port 513 nsew
rlabel metal1 s 37680 50310 37680 50310 4 vdd
port 513 nsew
rlabel metal1 s 39696 47940 39696 47940 4 vdd
port 513 nsew
rlabel metal1 s 38928 47940 38928 47940 4 vdd
port 513 nsew
rlabel metal1 s 38448 47940 38448 47940 4 vdd
port 513 nsew
rlabel metal1 s 38928 49229 38928 49229 4 vdd
port 513 nsew
rlabel metal1 s 39696 48439 39696 48439 4 vdd
port 513 nsew
rlabel metal1 s 38928 47649 38928 47649 4 vdd
port 513 nsew
rlabel metal1 s 39696 49520 39696 49520 4 vdd
port 513 nsew
rlabel metal1 s 38928 48730 38928 48730 4 vdd
port 513 nsew
rlabel metal1 s 37680 50019 37680 50019 4 vdd
port 513 nsew
rlabel metal1 s 38448 48439 38448 48439 4 vdd
port 513 nsew
rlabel metal1 s 37680 47649 37680 47649 4 vdd
port 513 nsew
rlabel metal1 s 38448 48730 38448 48730 4 vdd
port 513 nsew
rlabel metal1 s 39696 48730 39696 48730 4 vdd
port 513 nsew
rlabel metal1 s 39696 50019 39696 50019 4 vdd
port 513 nsew
rlabel metal1 s 38448 50019 38448 50019 4 vdd
port 513 nsew
rlabel metal1 s 38928 50019 38928 50019 4 vdd
port 513 nsew
rlabel metal1 s 39696 50310 39696 50310 4 vdd
port 513 nsew
rlabel metal1 s 37680 49520 37680 49520 4 vdd
port 513 nsew
rlabel metal1 s 38928 49520 38928 49520 4 vdd
port 513 nsew
rlabel metal1 s 38928 50310 38928 50310 4 vdd
port 513 nsew
rlabel metal1 s 39696 47649 39696 47649 4 vdd
port 513 nsew
rlabel metal1 s 37680 47940 37680 47940 4 vdd
port 513 nsew
rlabel metal1 s 38928 48439 38928 48439 4 vdd
port 513 nsew
rlabel metal1 s 38448 50310 38448 50310 4 vdd
port 513 nsew
rlabel metal1 s 39696 49229 39696 49229 4 vdd
port 513 nsew
rlabel metal1 s 38448 49520 38448 49520 4 vdd
port 513 nsew
rlabel metal1 s 38448 49229 38448 49229 4 vdd
port 513 nsew
rlabel metal1 s 38448 47649 38448 47649 4 vdd
port 513 nsew
rlabel metal1 s 37680 48730 37680 48730 4 vdd
port 513 nsew
rlabel metal1 s 37200 47649 37200 47649 4 vdd
port 513 nsew
rlabel metal1 s 36432 50019 36432 50019 4 vdd
port 513 nsew
rlabel metal1 s 35184 47940 35184 47940 4 vdd
port 513 nsew
rlabel metal1 s 36432 48730 36432 48730 4 vdd
port 513 nsew
rlabel metal1 s 36432 49229 36432 49229 4 vdd
port 513 nsew
rlabel metal1 s 35184 50310 35184 50310 4 vdd
port 513 nsew
rlabel metal1 s 36432 47940 36432 47940 4 vdd
port 513 nsew
rlabel metal1 s 35952 47940 35952 47940 4 vdd
port 513 nsew
rlabel metal1 s 36432 47649 36432 47649 4 vdd
port 513 nsew
rlabel metal1 s 35952 47649 35952 47649 4 vdd
port 513 nsew
rlabel metal1 s 35184 50019 35184 50019 4 vdd
port 513 nsew
rlabel metal1 s 37200 48730 37200 48730 4 vdd
port 513 nsew
rlabel metal1 s 35952 50310 35952 50310 4 vdd
port 513 nsew
rlabel metal1 s 35952 48730 35952 48730 4 vdd
port 513 nsew
rlabel metal1 s 35184 49520 35184 49520 4 vdd
port 513 nsew
rlabel metal1 s 35184 48730 35184 48730 4 vdd
port 513 nsew
rlabel metal1 s 37200 49229 37200 49229 4 vdd
port 513 nsew
rlabel metal1 s 37200 50310 37200 50310 4 vdd
port 513 nsew
rlabel metal1 s 35952 50019 35952 50019 4 vdd
port 513 nsew
rlabel metal1 s 35952 49520 35952 49520 4 vdd
port 513 nsew
rlabel metal1 s 37200 48439 37200 48439 4 vdd
port 513 nsew
rlabel metal1 s 36432 49520 36432 49520 4 vdd
port 513 nsew
rlabel metal1 s 35184 47649 35184 47649 4 vdd
port 513 nsew
rlabel metal1 s 35184 48439 35184 48439 4 vdd
port 513 nsew
rlabel metal1 s 35952 48439 35952 48439 4 vdd
port 513 nsew
rlabel metal1 s 36432 50310 36432 50310 4 vdd
port 513 nsew
rlabel metal1 s 37200 50019 37200 50019 4 vdd
port 513 nsew
rlabel metal1 s 37200 49520 37200 49520 4 vdd
port 513 nsew
rlabel metal1 s 35952 49229 35952 49229 4 vdd
port 513 nsew
rlabel metal1 s 35184 49229 35184 49229 4 vdd
port 513 nsew
rlabel metal1 s 36432 48439 36432 48439 4 vdd
port 513 nsew
rlabel metal1 s 37200 47940 37200 47940 4 vdd
port 513 nsew
rlabel metal1 s 35184 45279 35184 45279 4 vdd
port 513 nsew
rlabel metal1 s 37200 45279 37200 45279 4 vdd
port 513 nsew
rlabel metal1 s 36432 46069 36432 46069 4 vdd
port 513 nsew
rlabel metal1 s 35184 46859 35184 46859 4 vdd
port 513 nsew
rlabel metal1 s 37200 46859 37200 46859 4 vdd
port 513 nsew
rlabel metal1 s 36432 45279 36432 45279 4 vdd
port 513 nsew
rlabel metal1 s 35184 44780 35184 44780 4 vdd
port 513 nsew
rlabel metal1 s 35184 47150 35184 47150 4 vdd
port 513 nsew
rlabel metal1 s 35184 45570 35184 45570 4 vdd
port 513 nsew
rlabel metal1 s 35952 44489 35952 44489 4 vdd
port 513 nsew
rlabel metal1 s 35184 46360 35184 46360 4 vdd
port 513 nsew
rlabel metal1 s 37200 44489 37200 44489 4 vdd
port 513 nsew
rlabel metal1 s 37200 46069 37200 46069 4 vdd
port 513 nsew
rlabel metal1 s 37200 47150 37200 47150 4 vdd
port 513 nsew
rlabel metal1 s 36432 44489 36432 44489 4 vdd
port 513 nsew
rlabel metal1 s 36432 47150 36432 47150 4 vdd
port 513 nsew
rlabel metal1 s 37200 44780 37200 44780 4 vdd
port 513 nsew
rlabel metal1 s 35952 45279 35952 45279 4 vdd
port 513 nsew
rlabel metal1 s 35952 46069 35952 46069 4 vdd
port 513 nsew
rlabel metal1 s 36432 46360 36432 46360 4 vdd
port 513 nsew
rlabel metal1 s 37200 46360 37200 46360 4 vdd
port 513 nsew
rlabel metal1 s 35952 45570 35952 45570 4 vdd
port 513 nsew
rlabel metal1 s 36432 45570 36432 45570 4 vdd
port 513 nsew
rlabel metal1 s 35952 47150 35952 47150 4 vdd
port 513 nsew
rlabel metal1 s 36432 44780 36432 44780 4 vdd
port 513 nsew
rlabel metal1 s 35184 46069 35184 46069 4 vdd
port 513 nsew
rlabel metal1 s 35952 44780 35952 44780 4 vdd
port 513 nsew
rlabel metal1 s 35952 46360 35952 46360 4 vdd
port 513 nsew
rlabel metal1 s 35184 44489 35184 44489 4 vdd
port 513 nsew
rlabel metal1 s 36432 46859 36432 46859 4 vdd
port 513 nsew
rlabel metal1 s 35952 46859 35952 46859 4 vdd
port 513 nsew
rlabel metal1 s 37200 45570 37200 45570 4 vdd
port 513 nsew
rlabel metal1 s 38928 46360 38928 46360 4 vdd
port 513 nsew
rlabel metal1 s 39696 46859 39696 46859 4 vdd
port 513 nsew
rlabel metal1 s 38928 45570 38928 45570 4 vdd
port 513 nsew
rlabel metal1 s 39696 46360 39696 46360 4 vdd
port 513 nsew
rlabel metal1 s 38928 45279 38928 45279 4 vdd
port 513 nsew
rlabel metal1 s 38928 46069 38928 46069 4 vdd
port 513 nsew
rlabel metal1 s 37680 45570 37680 45570 4 vdd
port 513 nsew
rlabel metal1 s 37680 47150 37680 47150 4 vdd
port 513 nsew
rlabel metal1 s 38448 45279 38448 45279 4 vdd
port 513 nsew
rlabel metal1 s 38928 47150 38928 47150 4 vdd
port 513 nsew
rlabel metal1 s 37680 44489 37680 44489 4 vdd
port 513 nsew
rlabel metal1 s 39696 45570 39696 45570 4 vdd
port 513 nsew
rlabel metal1 s 38928 44780 38928 44780 4 vdd
port 513 nsew
rlabel metal1 s 37680 45279 37680 45279 4 vdd
port 513 nsew
rlabel metal1 s 37680 46360 37680 46360 4 vdd
port 513 nsew
rlabel metal1 s 38928 46859 38928 46859 4 vdd
port 513 nsew
rlabel metal1 s 38448 44780 38448 44780 4 vdd
port 513 nsew
rlabel metal1 s 38448 44489 38448 44489 4 vdd
port 513 nsew
rlabel metal1 s 37680 46069 37680 46069 4 vdd
port 513 nsew
rlabel metal1 s 38448 46360 38448 46360 4 vdd
port 513 nsew
rlabel metal1 s 38928 44489 38928 44489 4 vdd
port 513 nsew
rlabel metal1 s 38448 46069 38448 46069 4 vdd
port 513 nsew
rlabel metal1 s 38448 46859 38448 46859 4 vdd
port 513 nsew
rlabel metal1 s 39696 47150 39696 47150 4 vdd
port 513 nsew
rlabel metal1 s 37680 46859 37680 46859 4 vdd
port 513 nsew
rlabel metal1 s 38448 47150 38448 47150 4 vdd
port 513 nsew
rlabel metal1 s 38448 45570 38448 45570 4 vdd
port 513 nsew
rlabel metal1 s 39696 46069 39696 46069 4 vdd
port 513 nsew
rlabel metal1 s 39696 44780 39696 44780 4 vdd
port 513 nsew
rlabel metal1 s 37680 44780 37680 44780 4 vdd
port 513 nsew
rlabel metal1 s 39696 44489 39696 44489 4 vdd
port 513 nsew
rlabel metal1 s 39696 45279 39696 45279 4 vdd
port 513 nsew
rlabel metal1 s 33456 48439 33456 48439 4 vdd
port 513 nsew
rlabel metal1 s 34704 50019 34704 50019 4 vdd
port 513 nsew
rlabel metal1 s 34704 47649 34704 47649 4 vdd
port 513 nsew
rlabel metal1 s 33936 47649 33936 47649 4 vdd
port 513 nsew
rlabel metal1 s 33456 47940 33456 47940 4 vdd
port 513 nsew
rlabel metal1 s 34704 50310 34704 50310 4 vdd
port 513 nsew
rlabel metal1 s 33456 48730 33456 48730 4 vdd
port 513 nsew
rlabel metal1 s 33456 49520 33456 49520 4 vdd
port 513 nsew
rlabel metal1 s 32688 48439 32688 48439 4 vdd
port 513 nsew
rlabel metal1 s 34704 48439 34704 48439 4 vdd
port 513 nsew
rlabel metal1 s 33936 48730 33936 48730 4 vdd
port 513 nsew
rlabel metal1 s 33456 49229 33456 49229 4 vdd
port 513 nsew
rlabel metal1 s 33936 49520 33936 49520 4 vdd
port 513 nsew
rlabel metal1 s 33456 50310 33456 50310 4 vdd
port 513 nsew
rlabel metal1 s 33456 47649 33456 47649 4 vdd
port 513 nsew
rlabel metal1 s 32688 48730 32688 48730 4 vdd
port 513 nsew
rlabel metal1 s 34704 47940 34704 47940 4 vdd
port 513 nsew
rlabel metal1 s 32688 50310 32688 50310 4 vdd
port 513 nsew
rlabel metal1 s 34704 48730 34704 48730 4 vdd
port 513 nsew
rlabel metal1 s 34704 49520 34704 49520 4 vdd
port 513 nsew
rlabel metal1 s 32688 49229 32688 49229 4 vdd
port 513 nsew
rlabel metal1 s 34704 49229 34704 49229 4 vdd
port 513 nsew
rlabel metal1 s 32688 49520 32688 49520 4 vdd
port 513 nsew
rlabel metal1 s 32688 50019 32688 50019 4 vdd
port 513 nsew
rlabel metal1 s 33936 50310 33936 50310 4 vdd
port 513 nsew
rlabel metal1 s 33936 49229 33936 49229 4 vdd
port 513 nsew
rlabel metal1 s 33456 50019 33456 50019 4 vdd
port 513 nsew
rlabel metal1 s 32688 47940 32688 47940 4 vdd
port 513 nsew
rlabel metal1 s 33936 47940 33936 47940 4 vdd
port 513 nsew
rlabel metal1 s 33936 50019 33936 50019 4 vdd
port 513 nsew
rlabel metal1 s 32688 47649 32688 47649 4 vdd
port 513 nsew
rlabel metal1 s 33936 48439 33936 48439 4 vdd
port 513 nsew
rlabel metal1 s 30192 49520 30192 49520 4 vdd
port 513 nsew
rlabel metal1 s 30192 47940 30192 47940 4 vdd
port 513 nsew
rlabel metal1 s 30960 50310 30960 50310 4 vdd
port 513 nsew
rlabel metal1 s 32208 47940 32208 47940 4 vdd
port 513 nsew
rlabel metal1 s 32208 49520 32208 49520 4 vdd
port 513 nsew
rlabel metal1 s 30960 48439 30960 48439 4 vdd
port 513 nsew
rlabel metal1 s 32208 50019 32208 50019 4 vdd
port 513 nsew
rlabel metal1 s 31440 49520 31440 49520 4 vdd
port 513 nsew
rlabel metal1 s 30960 50019 30960 50019 4 vdd
port 513 nsew
rlabel metal1 s 32208 49229 32208 49229 4 vdd
port 513 nsew
rlabel metal1 s 30960 48730 30960 48730 4 vdd
port 513 nsew
rlabel metal1 s 31440 50310 31440 50310 4 vdd
port 513 nsew
rlabel metal1 s 31440 50019 31440 50019 4 vdd
port 513 nsew
rlabel metal1 s 32208 48439 32208 48439 4 vdd
port 513 nsew
rlabel metal1 s 32208 47649 32208 47649 4 vdd
port 513 nsew
rlabel metal1 s 30960 49229 30960 49229 4 vdd
port 513 nsew
rlabel metal1 s 31440 49229 31440 49229 4 vdd
port 513 nsew
rlabel metal1 s 30192 47649 30192 47649 4 vdd
port 513 nsew
rlabel metal1 s 31440 48439 31440 48439 4 vdd
port 513 nsew
rlabel metal1 s 30960 49520 30960 49520 4 vdd
port 513 nsew
rlabel metal1 s 30192 50310 30192 50310 4 vdd
port 513 nsew
rlabel metal1 s 32208 48730 32208 48730 4 vdd
port 513 nsew
rlabel metal1 s 30192 50019 30192 50019 4 vdd
port 513 nsew
rlabel metal1 s 32208 50310 32208 50310 4 vdd
port 513 nsew
rlabel metal1 s 30960 47649 30960 47649 4 vdd
port 513 nsew
rlabel metal1 s 31440 47649 31440 47649 4 vdd
port 513 nsew
rlabel metal1 s 30192 48439 30192 48439 4 vdd
port 513 nsew
rlabel metal1 s 31440 47940 31440 47940 4 vdd
port 513 nsew
rlabel metal1 s 30960 47940 30960 47940 4 vdd
port 513 nsew
rlabel metal1 s 31440 48730 31440 48730 4 vdd
port 513 nsew
rlabel metal1 s 30192 49229 30192 49229 4 vdd
port 513 nsew
rlabel metal1 s 30192 48730 30192 48730 4 vdd
port 513 nsew
rlabel metal1 s 30192 44780 30192 44780 4 vdd
port 513 nsew
rlabel metal1 s 32208 44780 32208 44780 4 vdd
port 513 nsew
rlabel metal1 s 31440 46360 31440 46360 4 vdd
port 513 nsew
rlabel metal1 s 30960 44489 30960 44489 4 vdd
port 513 nsew
rlabel metal1 s 31440 47150 31440 47150 4 vdd
port 513 nsew
rlabel metal1 s 30960 46859 30960 46859 4 vdd
port 513 nsew
rlabel metal1 s 30192 46360 30192 46360 4 vdd
port 513 nsew
rlabel metal1 s 30960 46360 30960 46360 4 vdd
port 513 nsew
rlabel metal1 s 31440 46859 31440 46859 4 vdd
port 513 nsew
rlabel metal1 s 32208 44489 32208 44489 4 vdd
port 513 nsew
rlabel metal1 s 30192 44489 30192 44489 4 vdd
port 513 nsew
rlabel metal1 s 32208 46360 32208 46360 4 vdd
port 513 nsew
rlabel metal1 s 32208 45570 32208 45570 4 vdd
port 513 nsew
rlabel metal1 s 31440 45570 31440 45570 4 vdd
port 513 nsew
rlabel metal1 s 30192 47150 30192 47150 4 vdd
port 513 nsew
rlabel metal1 s 30192 45570 30192 45570 4 vdd
port 513 nsew
rlabel metal1 s 30960 44780 30960 44780 4 vdd
port 513 nsew
rlabel metal1 s 30960 45570 30960 45570 4 vdd
port 513 nsew
rlabel metal1 s 30192 46859 30192 46859 4 vdd
port 513 nsew
rlabel metal1 s 30960 47150 30960 47150 4 vdd
port 513 nsew
rlabel metal1 s 32208 46859 32208 46859 4 vdd
port 513 nsew
rlabel metal1 s 32208 46069 32208 46069 4 vdd
port 513 nsew
rlabel metal1 s 31440 46069 31440 46069 4 vdd
port 513 nsew
rlabel metal1 s 30960 46069 30960 46069 4 vdd
port 513 nsew
rlabel metal1 s 31440 44780 31440 44780 4 vdd
port 513 nsew
rlabel metal1 s 30192 46069 30192 46069 4 vdd
port 513 nsew
rlabel metal1 s 31440 45279 31440 45279 4 vdd
port 513 nsew
rlabel metal1 s 32208 47150 32208 47150 4 vdd
port 513 nsew
rlabel metal1 s 30960 45279 30960 45279 4 vdd
port 513 nsew
rlabel metal1 s 32208 45279 32208 45279 4 vdd
port 513 nsew
rlabel metal1 s 30192 45279 30192 45279 4 vdd
port 513 nsew
rlabel metal1 s 31440 44489 31440 44489 4 vdd
port 513 nsew
rlabel metal1 s 34704 45279 34704 45279 4 vdd
port 513 nsew
rlabel metal1 s 33456 45279 33456 45279 4 vdd
port 513 nsew
rlabel metal1 s 33936 44780 33936 44780 4 vdd
port 513 nsew
rlabel metal1 s 34704 44489 34704 44489 4 vdd
port 513 nsew
rlabel metal1 s 32688 46859 32688 46859 4 vdd
port 513 nsew
rlabel metal1 s 33456 47150 33456 47150 4 vdd
port 513 nsew
rlabel metal1 s 32688 45570 32688 45570 4 vdd
port 513 nsew
rlabel metal1 s 32688 45279 32688 45279 4 vdd
port 513 nsew
rlabel metal1 s 33936 47150 33936 47150 4 vdd
port 513 nsew
rlabel metal1 s 33936 44489 33936 44489 4 vdd
port 513 nsew
rlabel metal1 s 33456 46069 33456 46069 4 vdd
port 513 nsew
rlabel metal1 s 32688 46360 32688 46360 4 vdd
port 513 nsew
rlabel metal1 s 32688 47150 32688 47150 4 vdd
port 513 nsew
rlabel metal1 s 33456 46859 33456 46859 4 vdd
port 513 nsew
rlabel metal1 s 32688 44780 32688 44780 4 vdd
port 513 nsew
rlabel metal1 s 33936 45279 33936 45279 4 vdd
port 513 nsew
rlabel metal1 s 34704 45570 34704 45570 4 vdd
port 513 nsew
rlabel metal1 s 33456 44780 33456 44780 4 vdd
port 513 nsew
rlabel metal1 s 33936 46069 33936 46069 4 vdd
port 513 nsew
rlabel metal1 s 34704 44780 34704 44780 4 vdd
port 513 nsew
rlabel metal1 s 32688 44489 32688 44489 4 vdd
port 513 nsew
rlabel metal1 s 34704 46859 34704 46859 4 vdd
port 513 nsew
rlabel metal1 s 33456 44489 33456 44489 4 vdd
port 513 nsew
rlabel metal1 s 33936 45570 33936 45570 4 vdd
port 513 nsew
rlabel metal1 s 33456 46360 33456 46360 4 vdd
port 513 nsew
rlabel metal1 s 34704 46069 34704 46069 4 vdd
port 513 nsew
rlabel metal1 s 34704 47150 34704 47150 4 vdd
port 513 nsew
rlabel metal1 s 33456 45570 33456 45570 4 vdd
port 513 nsew
rlabel metal1 s 32688 46069 32688 46069 4 vdd
port 513 nsew
rlabel metal1 s 33936 46859 33936 46859 4 vdd
port 513 nsew
rlabel metal1 s 34704 46360 34704 46360 4 vdd
port 513 nsew
rlabel metal1 s 33936 46360 33936 46360 4 vdd
port 513 nsew
rlabel metal1 s 33936 43200 33936 43200 4 vdd
port 513 nsew
rlabel metal1 s 33456 41620 33456 41620 4 vdd
port 513 nsew
rlabel metal1 s 33936 41620 33936 41620 4 vdd
port 513 nsew
rlabel metal1 s 33936 43990 33936 43990 4 vdd
port 513 nsew
rlabel metal1 s 34704 43699 34704 43699 4 vdd
port 513 nsew
rlabel metal1 s 33456 43699 33456 43699 4 vdd
port 513 nsew
rlabel metal1 s 34704 43990 34704 43990 4 vdd
port 513 nsew
rlabel metal1 s 33936 42909 33936 42909 4 vdd
port 513 nsew
rlabel metal1 s 32688 43699 32688 43699 4 vdd
port 513 nsew
rlabel metal1 s 33456 43990 33456 43990 4 vdd
port 513 nsew
rlabel metal1 s 32688 41329 32688 41329 4 vdd
port 513 nsew
rlabel metal1 s 32688 42909 32688 42909 4 vdd
port 513 nsew
rlabel metal1 s 32688 43200 32688 43200 4 vdd
port 513 nsew
rlabel metal1 s 32688 41620 32688 41620 4 vdd
port 513 nsew
rlabel metal1 s 33936 42410 33936 42410 4 vdd
port 513 nsew
rlabel metal1 s 33936 43699 33936 43699 4 vdd
port 513 nsew
rlabel metal1 s 33456 41329 33456 41329 4 vdd
port 513 nsew
rlabel metal1 s 34704 42119 34704 42119 4 vdd
port 513 nsew
rlabel metal1 s 34704 43200 34704 43200 4 vdd
port 513 nsew
rlabel metal1 s 34704 41329 34704 41329 4 vdd
port 513 nsew
rlabel metal1 s 34704 42410 34704 42410 4 vdd
port 513 nsew
rlabel metal1 s 34704 42909 34704 42909 4 vdd
port 513 nsew
rlabel metal1 s 32688 42119 32688 42119 4 vdd
port 513 nsew
rlabel metal1 s 33456 43200 33456 43200 4 vdd
port 513 nsew
rlabel metal1 s 33456 42410 33456 42410 4 vdd
port 513 nsew
rlabel metal1 s 33456 42909 33456 42909 4 vdd
port 513 nsew
rlabel metal1 s 33456 42119 33456 42119 4 vdd
port 513 nsew
rlabel metal1 s 33936 41329 33936 41329 4 vdd
port 513 nsew
rlabel metal1 s 32688 43990 32688 43990 4 vdd
port 513 nsew
rlabel metal1 s 34704 41620 34704 41620 4 vdd
port 513 nsew
rlabel metal1 s 33936 42119 33936 42119 4 vdd
port 513 nsew
rlabel metal1 s 32688 42410 32688 42410 4 vdd
port 513 nsew
rlabel metal1 s 32208 41620 32208 41620 4 vdd
port 513 nsew
rlabel metal1 s 30192 43990 30192 43990 4 vdd
port 513 nsew
rlabel metal1 s 30192 42909 30192 42909 4 vdd
port 513 nsew
rlabel metal1 s 31440 43699 31440 43699 4 vdd
port 513 nsew
rlabel metal1 s 30192 42410 30192 42410 4 vdd
port 513 nsew
rlabel metal1 s 32208 42410 32208 42410 4 vdd
port 513 nsew
rlabel metal1 s 30192 41620 30192 41620 4 vdd
port 513 nsew
rlabel metal1 s 31440 42119 31440 42119 4 vdd
port 513 nsew
rlabel metal1 s 30960 43990 30960 43990 4 vdd
port 513 nsew
rlabel metal1 s 32208 42909 32208 42909 4 vdd
port 513 nsew
rlabel metal1 s 30960 43699 30960 43699 4 vdd
port 513 nsew
rlabel metal1 s 31440 43200 31440 43200 4 vdd
port 513 nsew
rlabel metal1 s 30960 43200 30960 43200 4 vdd
port 513 nsew
rlabel metal1 s 30192 43200 30192 43200 4 vdd
port 513 nsew
rlabel metal1 s 32208 43200 32208 43200 4 vdd
port 513 nsew
rlabel metal1 s 30960 42119 30960 42119 4 vdd
port 513 nsew
rlabel metal1 s 30960 41329 30960 41329 4 vdd
port 513 nsew
rlabel metal1 s 31440 41329 31440 41329 4 vdd
port 513 nsew
rlabel metal1 s 32208 43699 32208 43699 4 vdd
port 513 nsew
rlabel metal1 s 32208 43990 32208 43990 4 vdd
port 513 nsew
rlabel metal1 s 30960 42410 30960 42410 4 vdd
port 513 nsew
rlabel metal1 s 31440 43990 31440 43990 4 vdd
port 513 nsew
rlabel metal1 s 30192 42119 30192 42119 4 vdd
port 513 nsew
rlabel metal1 s 30192 41329 30192 41329 4 vdd
port 513 nsew
rlabel metal1 s 31440 41620 31440 41620 4 vdd
port 513 nsew
rlabel metal1 s 31440 42410 31440 42410 4 vdd
port 513 nsew
rlabel metal1 s 30192 43699 30192 43699 4 vdd
port 513 nsew
rlabel metal1 s 30960 41620 30960 41620 4 vdd
port 513 nsew
rlabel metal1 s 30960 42909 30960 42909 4 vdd
port 513 nsew
rlabel metal1 s 31440 42909 31440 42909 4 vdd
port 513 nsew
rlabel metal1 s 32208 41329 32208 41329 4 vdd
port 513 nsew
rlabel metal1 s 32208 42119 32208 42119 4 vdd
port 513 nsew
rlabel metal1 s 30192 39250 30192 39250 4 vdd
port 513 nsew
rlabel metal1 s 32208 39749 32208 39749 4 vdd
port 513 nsew
rlabel metal1 s 32208 39250 32208 39250 4 vdd
port 513 nsew
rlabel metal1 s 30192 38959 30192 38959 4 vdd
port 513 nsew
rlabel metal1 s 31440 40539 31440 40539 4 vdd
port 513 nsew
rlabel metal1 s 31440 38460 31440 38460 4 vdd
port 513 nsew
rlabel metal1 s 32208 38959 32208 38959 4 vdd
port 513 nsew
rlabel metal1 s 32208 38169 32208 38169 4 vdd
port 513 nsew
rlabel metal1 s 30960 40539 30960 40539 4 vdd
port 513 nsew
rlabel metal1 s 31440 38959 31440 38959 4 vdd
port 513 nsew
rlabel metal1 s 30960 40040 30960 40040 4 vdd
port 513 nsew
rlabel metal1 s 30960 39250 30960 39250 4 vdd
port 513 nsew
rlabel metal1 s 30192 40539 30192 40539 4 vdd
port 513 nsew
rlabel metal1 s 30960 38460 30960 38460 4 vdd
port 513 nsew
rlabel metal1 s 32208 38460 32208 38460 4 vdd
port 513 nsew
rlabel metal1 s 30960 39749 30960 39749 4 vdd
port 513 nsew
rlabel metal1 s 30192 38460 30192 38460 4 vdd
port 513 nsew
rlabel metal1 s 32208 40830 32208 40830 4 vdd
port 513 nsew
rlabel metal1 s 32208 40040 32208 40040 4 vdd
port 513 nsew
rlabel metal1 s 31440 38169 31440 38169 4 vdd
port 513 nsew
rlabel metal1 s 30192 40040 30192 40040 4 vdd
port 513 nsew
rlabel metal1 s 30192 40830 30192 40830 4 vdd
port 513 nsew
rlabel metal1 s 30960 38169 30960 38169 4 vdd
port 513 nsew
rlabel metal1 s 31440 40830 31440 40830 4 vdd
port 513 nsew
rlabel metal1 s 30192 39749 30192 39749 4 vdd
port 513 nsew
rlabel metal1 s 32208 40539 32208 40539 4 vdd
port 513 nsew
rlabel metal1 s 30192 38169 30192 38169 4 vdd
port 513 nsew
rlabel metal1 s 31440 39749 31440 39749 4 vdd
port 513 nsew
rlabel metal1 s 31440 39250 31440 39250 4 vdd
port 513 nsew
rlabel metal1 s 30960 40830 30960 40830 4 vdd
port 513 nsew
rlabel metal1 s 31440 40040 31440 40040 4 vdd
port 513 nsew
rlabel metal1 s 30960 38959 30960 38959 4 vdd
port 513 nsew
rlabel metal1 s 32688 38169 32688 38169 4 vdd
port 513 nsew
rlabel metal1 s 34704 39250 34704 39250 4 vdd
port 513 nsew
rlabel metal1 s 33936 38460 33936 38460 4 vdd
port 513 nsew
rlabel metal1 s 33936 40040 33936 40040 4 vdd
port 513 nsew
rlabel metal1 s 33936 38169 33936 38169 4 vdd
port 513 nsew
rlabel metal1 s 33456 40040 33456 40040 4 vdd
port 513 nsew
rlabel metal1 s 34704 40040 34704 40040 4 vdd
port 513 nsew
rlabel metal1 s 32688 40539 32688 40539 4 vdd
port 513 nsew
rlabel metal1 s 34704 39749 34704 39749 4 vdd
port 513 nsew
rlabel metal1 s 32688 39749 32688 39749 4 vdd
port 513 nsew
rlabel metal1 s 34704 40539 34704 40539 4 vdd
port 513 nsew
rlabel metal1 s 34704 40830 34704 40830 4 vdd
port 513 nsew
rlabel metal1 s 33456 39250 33456 39250 4 vdd
port 513 nsew
rlabel metal1 s 33936 40539 33936 40539 4 vdd
port 513 nsew
rlabel metal1 s 33456 38959 33456 38959 4 vdd
port 513 nsew
rlabel metal1 s 32688 40040 32688 40040 4 vdd
port 513 nsew
rlabel metal1 s 33936 40830 33936 40830 4 vdd
port 513 nsew
rlabel metal1 s 33936 39250 33936 39250 4 vdd
port 513 nsew
rlabel metal1 s 32688 38959 32688 38959 4 vdd
port 513 nsew
rlabel metal1 s 33456 38460 33456 38460 4 vdd
port 513 nsew
rlabel metal1 s 32688 39250 32688 39250 4 vdd
port 513 nsew
rlabel metal1 s 33936 39749 33936 39749 4 vdd
port 513 nsew
rlabel metal1 s 33936 38959 33936 38959 4 vdd
port 513 nsew
rlabel metal1 s 33456 40830 33456 40830 4 vdd
port 513 nsew
rlabel metal1 s 32688 40830 32688 40830 4 vdd
port 513 nsew
rlabel metal1 s 34704 38959 34704 38959 4 vdd
port 513 nsew
rlabel metal1 s 33456 38169 33456 38169 4 vdd
port 513 nsew
rlabel metal1 s 33456 39749 33456 39749 4 vdd
port 513 nsew
rlabel metal1 s 34704 38169 34704 38169 4 vdd
port 513 nsew
rlabel metal1 s 33456 40539 33456 40539 4 vdd
port 513 nsew
rlabel metal1 s 32688 38460 32688 38460 4 vdd
port 513 nsew
rlabel metal1 s 34704 38460 34704 38460 4 vdd
port 513 nsew
rlabel metal1 s 38448 41329 38448 41329 4 vdd
port 513 nsew
rlabel metal1 s 38448 42410 38448 42410 4 vdd
port 513 nsew
rlabel metal1 s 38928 42410 38928 42410 4 vdd
port 513 nsew
rlabel metal1 s 39696 43699 39696 43699 4 vdd
port 513 nsew
rlabel metal1 s 38928 41620 38928 41620 4 vdd
port 513 nsew
rlabel metal1 s 37680 43699 37680 43699 4 vdd
port 513 nsew
rlabel metal1 s 37680 42119 37680 42119 4 vdd
port 513 nsew
rlabel metal1 s 38448 43699 38448 43699 4 vdd
port 513 nsew
rlabel metal1 s 38448 43200 38448 43200 4 vdd
port 513 nsew
rlabel metal1 s 37680 41329 37680 41329 4 vdd
port 513 nsew
rlabel metal1 s 39696 43200 39696 43200 4 vdd
port 513 nsew
rlabel metal1 s 39696 42119 39696 42119 4 vdd
port 513 nsew
rlabel metal1 s 39696 41620 39696 41620 4 vdd
port 513 nsew
rlabel metal1 s 38928 43200 38928 43200 4 vdd
port 513 nsew
rlabel metal1 s 38928 42119 38928 42119 4 vdd
port 513 nsew
rlabel metal1 s 37680 42909 37680 42909 4 vdd
port 513 nsew
rlabel metal1 s 38928 43990 38928 43990 4 vdd
port 513 nsew
rlabel metal1 s 39696 41329 39696 41329 4 vdd
port 513 nsew
rlabel metal1 s 39696 42410 39696 42410 4 vdd
port 513 nsew
rlabel metal1 s 38448 43990 38448 43990 4 vdd
port 513 nsew
rlabel metal1 s 38928 43699 38928 43699 4 vdd
port 513 nsew
rlabel metal1 s 39696 43990 39696 43990 4 vdd
port 513 nsew
rlabel metal1 s 37680 41620 37680 41620 4 vdd
port 513 nsew
rlabel metal1 s 38928 42909 38928 42909 4 vdd
port 513 nsew
rlabel metal1 s 39696 42909 39696 42909 4 vdd
port 513 nsew
rlabel metal1 s 38448 42909 38448 42909 4 vdd
port 513 nsew
rlabel metal1 s 38448 42119 38448 42119 4 vdd
port 513 nsew
rlabel metal1 s 37680 43200 37680 43200 4 vdd
port 513 nsew
rlabel metal1 s 38448 41620 38448 41620 4 vdd
port 513 nsew
rlabel metal1 s 37680 43990 37680 43990 4 vdd
port 513 nsew
rlabel metal1 s 38928 41329 38928 41329 4 vdd
port 513 nsew
rlabel metal1 s 37680 42410 37680 42410 4 vdd
port 513 nsew
rlabel metal1 s 35952 41329 35952 41329 4 vdd
port 513 nsew
rlabel metal1 s 36432 43990 36432 43990 4 vdd
port 513 nsew
rlabel metal1 s 37200 42119 37200 42119 4 vdd
port 513 nsew
rlabel metal1 s 36432 41329 36432 41329 4 vdd
port 513 nsew
rlabel metal1 s 37200 41620 37200 41620 4 vdd
port 513 nsew
rlabel metal1 s 36432 43699 36432 43699 4 vdd
port 513 nsew
rlabel metal1 s 35952 42119 35952 42119 4 vdd
port 513 nsew
rlabel metal1 s 36432 41620 36432 41620 4 vdd
port 513 nsew
rlabel metal1 s 36432 42119 36432 42119 4 vdd
port 513 nsew
rlabel metal1 s 35952 43699 35952 43699 4 vdd
port 513 nsew
rlabel metal1 s 36432 43200 36432 43200 4 vdd
port 513 nsew
rlabel metal1 s 37200 41329 37200 41329 4 vdd
port 513 nsew
rlabel metal1 s 35184 42909 35184 42909 4 vdd
port 513 nsew
rlabel metal1 s 35184 42410 35184 42410 4 vdd
port 513 nsew
rlabel metal1 s 35952 43200 35952 43200 4 vdd
port 513 nsew
rlabel metal1 s 36432 42909 36432 42909 4 vdd
port 513 nsew
rlabel metal1 s 37200 43990 37200 43990 4 vdd
port 513 nsew
rlabel metal1 s 35184 43990 35184 43990 4 vdd
port 513 nsew
rlabel metal1 s 35952 41620 35952 41620 4 vdd
port 513 nsew
rlabel metal1 s 37200 42909 37200 42909 4 vdd
port 513 nsew
rlabel metal1 s 36432 42410 36432 42410 4 vdd
port 513 nsew
rlabel metal1 s 37200 43200 37200 43200 4 vdd
port 513 nsew
rlabel metal1 s 37200 42410 37200 42410 4 vdd
port 513 nsew
rlabel metal1 s 35184 41620 35184 41620 4 vdd
port 513 nsew
rlabel metal1 s 35952 42909 35952 42909 4 vdd
port 513 nsew
rlabel metal1 s 35184 43200 35184 43200 4 vdd
port 513 nsew
rlabel metal1 s 35184 43699 35184 43699 4 vdd
port 513 nsew
rlabel metal1 s 35184 41329 35184 41329 4 vdd
port 513 nsew
rlabel metal1 s 35184 42119 35184 42119 4 vdd
port 513 nsew
rlabel metal1 s 37200 43699 37200 43699 4 vdd
port 513 nsew
rlabel metal1 s 35952 42410 35952 42410 4 vdd
port 513 nsew
rlabel metal1 s 35952 43990 35952 43990 4 vdd
port 513 nsew
rlabel metal1 s 35184 38169 35184 38169 4 vdd
port 513 nsew
rlabel metal1 s 37200 38169 37200 38169 4 vdd
port 513 nsew
rlabel metal1 s 35184 39749 35184 39749 4 vdd
port 513 nsew
rlabel metal1 s 36432 40040 36432 40040 4 vdd
port 513 nsew
rlabel metal1 s 37200 40830 37200 40830 4 vdd
port 513 nsew
rlabel metal1 s 35184 40539 35184 40539 4 vdd
port 513 nsew
rlabel metal1 s 35184 38460 35184 38460 4 vdd
port 513 nsew
rlabel metal1 s 36432 40539 36432 40539 4 vdd
port 513 nsew
rlabel metal1 s 35184 38959 35184 38959 4 vdd
port 513 nsew
rlabel metal1 s 35952 38169 35952 38169 4 vdd
port 513 nsew
rlabel metal1 s 37200 40539 37200 40539 4 vdd
port 513 nsew
rlabel metal1 s 35952 40830 35952 40830 4 vdd
port 513 nsew
rlabel metal1 s 35184 39250 35184 39250 4 vdd
port 513 nsew
rlabel metal1 s 37200 38959 37200 38959 4 vdd
port 513 nsew
rlabel metal1 s 35952 38460 35952 38460 4 vdd
port 513 nsew
rlabel metal1 s 35952 38959 35952 38959 4 vdd
port 513 nsew
rlabel metal1 s 36432 38460 36432 38460 4 vdd
port 513 nsew
rlabel metal1 s 37200 39250 37200 39250 4 vdd
port 513 nsew
rlabel metal1 s 37200 40040 37200 40040 4 vdd
port 513 nsew
rlabel metal1 s 35952 39749 35952 39749 4 vdd
port 513 nsew
rlabel metal1 s 36432 40830 36432 40830 4 vdd
port 513 nsew
rlabel metal1 s 36432 38959 36432 38959 4 vdd
port 513 nsew
rlabel metal1 s 36432 39749 36432 39749 4 vdd
port 513 nsew
rlabel metal1 s 35184 40830 35184 40830 4 vdd
port 513 nsew
rlabel metal1 s 35952 40040 35952 40040 4 vdd
port 513 nsew
rlabel metal1 s 37200 39749 37200 39749 4 vdd
port 513 nsew
rlabel metal1 s 35952 40539 35952 40539 4 vdd
port 513 nsew
rlabel metal1 s 36432 38169 36432 38169 4 vdd
port 513 nsew
rlabel metal1 s 35952 39250 35952 39250 4 vdd
port 513 nsew
rlabel metal1 s 36432 39250 36432 39250 4 vdd
port 513 nsew
rlabel metal1 s 37200 38460 37200 38460 4 vdd
port 513 nsew
rlabel metal1 s 35184 40040 35184 40040 4 vdd
port 513 nsew
rlabel metal1 s 38928 40830 38928 40830 4 vdd
port 513 nsew
rlabel metal1 s 38928 39749 38928 39749 4 vdd
port 513 nsew
rlabel metal1 s 37680 40539 37680 40539 4 vdd
port 513 nsew
rlabel metal1 s 38928 39250 38928 39250 4 vdd
port 513 nsew
rlabel metal1 s 39696 38460 39696 38460 4 vdd
port 513 nsew
rlabel metal1 s 39696 38959 39696 38959 4 vdd
port 513 nsew
rlabel metal1 s 39696 40040 39696 40040 4 vdd
port 513 nsew
rlabel metal1 s 38448 39749 38448 39749 4 vdd
port 513 nsew
rlabel metal1 s 38928 40040 38928 40040 4 vdd
port 513 nsew
rlabel metal1 s 38448 38959 38448 38959 4 vdd
port 513 nsew
rlabel metal1 s 39696 38169 39696 38169 4 vdd
port 513 nsew
rlabel metal1 s 38448 39250 38448 39250 4 vdd
port 513 nsew
rlabel metal1 s 37680 38169 37680 38169 4 vdd
port 513 nsew
rlabel metal1 s 38448 38460 38448 38460 4 vdd
port 513 nsew
rlabel metal1 s 37680 40830 37680 40830 4 vdd
port 513 nsew
rlabel metal1 s 37680 40040 37680 40040 4 vdd
port 513 nsew
rlabel metal1 s 38928 38959 38928 38959 4 vdd
port 513 nsew
rlabel metal1 s 37680 39250 37680 39250 4 vdd
port 513 nsew
rlabel metal1 s 38448 40040 38448 40040 4 vdd
port 513 nsew
rlabel metal1 s 39696 39749 39696 39749 4 vdd
port 513 nsew
rlabel metal1 s 38928 38169 38928 38169 4 vdd
port 513 nsew
rlabel metal1 s 38448 40830 38448 40830 4 vdd
port 513 nsew
rlabel metal1 s 37680 38959 37680 38959 4 vdd
port 513 nsew
rlabel metal1 s 38448 40539 38448 40539 4 vdd
port 513 nsew
rlabel metal1 s 39696 40830 39696 40830 4 vdd
port 513 nsew
rlabel metal1 s 39696 40539 39696 40539 4 vdd
port 513 nsew
rlabel metal1 s 38928 38460 38928 38460 4 vdd
port 513 nsew
rlabel metal1 s 39696 39250 39696 39250 4 vdd
port 513 nsew
rlabel metal1 s 38928 40539 38928 40539 4 vdd
port 513 nsew
rlabel metal1 s 37680 39749 37680 39749 4 vdd
port 513 nsew
rlabel metal1 s 38448 38169 38448 38169 4 vdd
port 513 nsew
rlabel metal1 s 37680 38460 37680 38460 4 vdd
port 513 nsew
rlabel metal1 s 29712 48439 29712 48439 4 vdd
port 513 nsew
rlabel metal1 s 28464 47940 28464 47940 4 vdd
port 513 nsew
rlabel metal1 s 28944 47940 28944 47940 4 vdd
port 513 nsew
rlabel metal1 s 28944 49229 28944 49229 4 vdd
port 513 nsew
rlabel metal1 s 28944 50019 28944 50019 4 vdd
port 513 nsew
rlabel metal1 s 28464 50310 28464 50310 4 vdd
port 513 nsew
rlabel metal1 s 27696 47649 27696 47649 4 vdd
port 513 nsew
rlabel metal1 s 29712 47940 29712 47940 4 vdd
port 513 nsew
rlabel metal1 s 28944 48730 28944 48730 4 vdd
port 513 nsew
rlabel metal1 s 29712 47649 29712 47649 4 vdd
port 513 nsew
rlabel metal1 s 29712 48730 29712 48730 4 vdd
port 513 nsew
rlabel metal1 s 28464 49520 28464 49520 4 vdd
port 513 nsew
rlabel metal1 s 29712 50310 29712 50310 4 vdd
port 513 nsew
rlabel metal1 s 28464 48439 28464 48439 4 vdd
port 513 nsew
rlabel metal1 s 29712 49229 29712 49229 4 vdd
port 513 nsew
rlabel metal1 s 28464 48730 28464 48730 4 vdd
port 513 nsew
rlabel metal1 s 28464 47649 28464 47649 4 vdd
port 513 nsew
rlabel metal1 s 29712 49520 29712 49520 4 vdd
port 513 nsew
rlabel metal1 s 27696 50019 27696 50019 4 vdd
port 513 nsew
rlabel metal1 s 27696 49229 27696 49229 4 vdd
port 513 nsew
rlabel metal1 s 27696 48730 27696 48730 4 vdd
port 513 nsew
rlabel metal1 s 28944 47649 28944 47649 4 vdd
port 513 nsew
rlabel metal1 s 28944 48439 28944 48439 4 vdd
port 513 nsew
rlabel metal1 s 27696 47940 27696 47940 4 vdd
port 513 nsew
rlabel metal1 s 28944 49520 28944 49520 4 vdd
port 513 nsew
rlabel metal1 s 28944 50310 28944 50310 4 vdd
port 513 nsew
rlabel metal1 s 29712 50019 29712 50019 4 vdd
port 513 nsew
rlabel metal1 s 27696 49520 27696 49520 4 vdd
port 513 nsew
rlabel metal1 s 27696 48439 27696 48439 4 vdd
port 513 nsew
rlabel metal1 s 27696 50310 27696 50310 4 vdd
port 513 nsew
rlabel metal1 s 28464 50019 28464 50019 4 vdd
port 513 nsew
rlabel metal1 s 28464 49229 28464 49229 4 vdd
port 513 nsew
rlabel metal1 s 26448 49229 26448 49229 4 vdd
port 513 nsew
rlabel metal1 s 27216 48730 27216 48730 4 vdd
port 513 nsew
rlabel metal1 s 26448 48730 26448 48730 4 vdd
port 513 nsew
rlabel metal1 s 26448 50019 26448 50019 4 vdd
port 513 nsew
rlabel metal1 s 26448 48439 26448 48439 4 vdd
port 513 nsew
rlabel metal1 s 25968 47940 25968 47940 4 vdd
port 513 nsew
rlabel metal1 s 25200 49229 25200 49229 4 vdd
port 513 nsew
rlabel metal1 s 25200 49520 25200 49520 4 vdd
port 513 nsew
rlabel metal1 s 27216 48439 27216 48439 4 vdd
port 513 nsew
rlabel metal1 s 25200 47649 25200 47649 4 vdd
port 513 nsew
rlabel metal1 s 25968 49229 25968 49229 4 vdd
port 513 nsew
rlabel metal1 s 25200 48439 25200 48439 4 vdd
port 513 nsew
rlabel metal1 s 25200 47940 25200 47940 4 vdd
port 513 nsew
rlabel metal1 s 25968 48439 25968 48439 4 vdd
port 513 nsew
rlabel metal1 s 27216 47649 27216 47649 4 vdd
port 513 nsew
rlabel metal1 s 25968 50019 25968 50019 4 vdd
port 513 nsew
rlabel metal1 s 26448 47940 26448 47940 4 vdd
port 513 nsew
rlabel metal1 s 26448 47649 26448 47649 4 vdd
port 513 nsew
rlabel metal1 s 25200 50310 25200 50310 4 vdd
port 513 nsew
rlabel metal1 s 25968 50310 25968 50310 4 vdd
port 513 nsew
rlabel metal1 s 25200 50019 25200 50019 4 vdd
port 513 nsew
rlabel metal1 s 27216 50019 27216 50019 4 vdd
port 513 nsew
rlabel metal1 s 25968 47649 25968 47649 4 vdd
port 513 nsew
rlabel metal1 s 25968 48730 25968 48730 4 vdd
port 513 nsew
rlabel metal1 s 27216 49229 27216 49229 4 vdd
port 513 nsew
rlabel metal1 s 25968 49520 25968 49520 4 vdd
port 513 nsew
rlabel metal1 s 27216 47940 27216 47940 4 vdd
port 513 nsew
rlabel metal1 s 25200 48730 25200 48730 4 vdd
port 513 nsew
rlabel metal1 s 26448 50310 26448 50310 4 vdd
port 513 nsew
rlabel metal1 s 27216 50310 27216 50310 4 vdd
port 513 nsew
rlabel metal1 s 26448 49520 26448 49520 4 vdd
port 513 nsew
rlabel metal1 s 27216 49520 27216 49520 4 vdd
port 513 nsew
rlabel metal1 s 25200 46360 25200 46360 4 vdd
port 513 nsew
rlabel metal1 s 27216 46360 27216 46360 4 vdd
port 513 nsew
rlabel metal1 s 25968 44489 25968 44489 4 vdd
port 513 nsew
rlabel metal1 s 27216 44489 27216 44489 4 vdd
port 513 nsew
rlabel metal1 s 25200 47150 25200 47150 4 vdd
port 513 nsew
rlabel metal1 s 26448 45570 26448 45570 4 vdd
port 513 nsew
rlabel metal1 s 25200 44489 25200 44489 4 vdd
port 513 nsew
rlabel metal1 s 27216 47150 27216 47150 4 vdd
port 513 nsew
rlabel metal1 s 26448 46859 26448 46859 4 vdd
port 513 nsew
rlabel metal1 s 27216 45279 27216 45279 4 vdd
port 513 nsew
rlabel metal1 s 25968 44780 25968 44780 4 vdd
port 513 nsew
rlabel metal1 s 27216 44780 27216 44780 4 vdd
port 513 nsew
rlabel metal1 s 27216 46859 27216 46859 4 vdd
port 513 nsew
rlabel metal1 s 25968 47150 25968 47150 4 vdd
port 513 nsew
rlabel metal1 s 25200 45279 25200 45279 4 vdd
port 513 nsew
rlabel metal1 s 25200 45570 25200 45570 4 vdd
port 513 nsew
rlabel metal1 s 26448 47150 26448 47150 4 vdd
port 513 nsew
rlabel metal1 s 25968 46069 25968 46069 4 vdd
port 513 nsew
rlabel metal1 s 25200 46859 25200 46859 4 vdd
port 513 nsew
rlabel metal1 s 27216 46069 27216 46069 4 vdd
port 513 nsew
rlabel metal1 s 26448 46069 26448 46069 4 vdd
port 513 nsew
rlabel metal1 s 25968 45279 25968 45279 4 vdd
port 513 nsew
rlabel metal1 s 26448 44489 26448 44489 4 vdd
port 513 nsew
rlabel metal1 s 25968 45570 25968 45570 4 vdd
port 513 nsew
rlabel metal1 s 25968 46859 25968 46859 4 vdd
port 513 nsew
rlabel metal1 s 26448 44780 26448 44780 4 vdd
port 513 nsew
rlabel metal1 s 26448 46360 26448 46360 4 vdd
port 513 nsew
rlabel metal1 s 25200 46069 25200 46069 4 vdd
port 513 nsew
rlabel metal1 s 27216 45570 27216 45570 4 vdd
port 513 nsew
rlabel metal1 s 26448 45279 26448 45279 4 vdd
port 513 nsew
rlabel metal1 s 25968 46360 25968 46360 4 vdd
port 513 nsew
rlabel metal1 s 25200 44780 25200 44780 4 vdd
port 513 nsew
rlabel metal1 s 28944 46069 28944 46069 4 vdd
port 513 nsew
rlabel metal1 s 28464 46859 28464 46859 4 vdd
port 513 nsew
rlabel metal1 s 28464 44489 28464 44489 4 vdd
port 513 nsew
rlabel metal1 s 28944 44489 28944 44489 4 vdd
port 513 nsew
rlabel metal1 s 27696 46069 27696 46069 4 vdd
port 513 nsew
rlabel metal1 s 29712 44780 29712 44780 4 vdd
port 513 nsew
rlabel metal1 s 28464 46360 28464 46360 4 vdd
port 513 nsew
rlabel metal1 s 29712 45570 29712 45570 4 vdd
port 513 nsew
rlabel metal1 s 28464 46069 28464 46069 4 vdd
port 513 nsew
rlabel metal1 s 28944 45570 28944 45570 4 vdd
port 513 nsew
rlabel metal1 s 27696 44489 27696 44489 4 vdd
port 513 nsew
rlabel metal1 s 28944 46360 28944 46360 4 vdd
port 513 nsew
rlabel metal1 s 29712 46069 29712 46069 4 vdd
port 513 nsew
rlabel metal1 s 29712 46360 29712 46360 4 vdd
port 513 nsew
rlabel metal1 s 28944 44780 28944 44780 4 vdd
port 513 nsew
rlabel metal1 s 28944 46859 28944 46859 4 vdd
port 513 nsew
rlabel metal1 s 28944 47150 28944 47150 4 vdd
port 513 nsew
rlabel metal1 s 28464 47150 28464 47150 4 vdd
port 513 nsew
rlabel metal1 s 27696 45570 27696 45570 4 vdd
port 513 nsew
rlabel metal1 s 27696 44780 27696 44780 4 vdd
port 513 nsew
rlabel metal1 s 28464 44780 28464 44780 4 vdd
port 513 nsew
rlabel metal1 s 29712 45279 29712 45279 4 vdd
port 513 nsew
rlabel metal1 s 27696 47150 27696 47150 4 vdd
port 513 nsew
rlabel metal1 s 29712 44489 29712 44489 4 vdd
port 513 nsew
rlabel metal1 s 28464 45570 28464 45570 4 vdd
port 513 nsew
rlabel metal1 s 27696 46360 27696 46360 4 vdd
port 513 nsew
rlabel metal1 s 28464 45279 28464 45279 4 vdd
port 513 nsew
rlabel metal1 s 29712 46859 29712 46859 4 vdd
port 513 nsew
rlabel metal1 s 27696 45279 27696 45279 4 vdd
port 513 nsew
rlabel metal1 s 28944 45279 28944 45279 4 vdd
port 513 nsew
rlabel metal1 s 27696 46859 27696 46859 4 vdd
port 513 nsew
rlabel metal1 s 29712 47150 29712 47150 4 vdd
port 513 nsew
rlabel metal1 s 23952 50310 23952 50310 4 vdd
port 513 nsew
rlabel metal1 s 23472 47940 23472 47940 4 vdd
port 513 nsew
rlabel metal1 s 24720 48439 24720 48439 4 vdd
port 513 nsew
rlabel metal1 s 23952 47649 23952 47649 4 vdd
port 513 nsew
rlabel metal1 s 23472 50019 23472 50019 4 vdd
port 513 nsew
rlabel metal1 s 23952 50019 23952 50019 4 vdd
port 513 nsew
rlabel metal1 s 22704 50310 22704 50310 4 vdd
port 513 nsew
rlabel metal1 s 22704 48439 22704 48439 4 vdd
port 513 nsew
rlabel metal1 s 23952 49229 23952 49229 4 vdd
port 513 nsew
rlabel metal1 s 24720 50019 24720 50019 4 vdd
port 513 nsew
rlabel metal1 s 24720 49520 24720 49520 4 vdd
port 513 nsew
rlabel metal1 s 22704 49520 22704 49520 4 vdd
port 513 nsew
rlabel metal1 s 24720 47649 24720 47649 4 vdd
port 513 nsew
rlabel metal1 s 22704 47649 22704 47649 4 vdd
port 513 nsew
rlabel metal1 s 24720 47940 24720 47940 4 vdd
port 513 nsew
rlabel metal1 s 23952 49520 23952 49520 4 vdd
port 513 nsew
rlabel metal1 s 22704 49229 22704 49229 4 vdd
port 513 nsew
rlabel metal1 s 24720 49229 24720 49229 4 vdd
port 513 nsew
rlabel metal1 s 23472 47649 23472 47649 4 vdd
port 513 nsew
rlabel metal1 s 23952 48439 23952 48439 4 vdd
port 513 nsew
rlabel metal1 s 22704 47940 22704 47940 4 vdd
port 513 nsew
rlabel metal1 s 23952 48730 23952 48730 4 vdd
port 513 nsew
rlabel metal1 s 24720 50310 24720 50310 4 vdd
port 513 nsew
rlabel metal1 s 23952 47940 23952 47940 4 vdd
port 513 nsew
rlabel metal1 s 23472 50310 23472 50310 4 vdd
port 513 nsew
rlabel metal1 s 24720 48730 24720 48730 4 vdd
port 513 nsew
rlabel metal1 s 23472 48730 23472 48730 4 vdd
port 513 nsew
rlabel metal1 s 22704 50019 22704 50019 4 vdd
port 513 nsew
rlabel metal1 s 22704 48730 22704 48730 4 vdd
port 513 nsew
rlabel metal1 s 23472 49229 23472 49229 4 vdd
port 513 nsew
rlabel metal1 s 23472 49520 23472 49520 4 vdd
port 513 nsew
rlabel metal1 s 23472 48439 23472 48439 4 vdd
port 513 nsew
rlabel metal1 s 22224 48730 22224 48730 4 vdd
port 513 nsew
rlabel metal1 s 21456 47940 21456 47940 4 vdd
port 513 nsew
rlabel metal1 s 22224 49520 22224 49520 4 vdd
port 513 nsew
rlabel metal1 s 20976 48439 20976 48439 4 vdd
port 513 nsew
rlabel metal1 s 20208 49520 20208 49520 4 vdd
port 513 nsew
rlabel metal1 s 20208 48439 20208 48439 4 vdd
port 513 nsew
rlabel metal1 s 20208 50310 20208 50310 4 vdd
port 513 nsew
rlabel metal1 s 21456 49229 21456 49229 4 vdd
port 513 nsew
rlabel metal1 s 22224 47649 22224 47649 4 vdd
port 513 nsew
rlabel metal1 s 22224 50019 22224 50019 4 vdd
port 513 nsew
rlabel metal1 s 20208 48730 20208 48730 4 vdd
port 513 nsew
rlabel metal1 s 22224 50310 22224 50310 4 vdd
port 513 nsew
rlabel metal1 s 20976 47940 20976 47940 4 vdd
port 513 nsew
rlabel metal1 s 20976 48730 20976 48730 4 vdd
port 513 nsew
rlabel metal1 s 20208 47649 20208 47649 4 vdd
port 513 nsew
rlabel metal1 s 20976 49520 20976 49520 4 vdd
port 513 nsew
rlabel metal1 s 21456 50019 21456 50019 4 vdd
port 513 nsew
rlabel metal1 s 20208 50019 20208 50019 4 vdd
port 513 nsew
rlabel metal1 s 21456 49520 21456 49520 4 vdd
port 513 nsew
rlabel metal1 s 21456 48439 21456 48439 4 vdd
port 513 nsew
rlabel metal1 s 22224 49229 22224 49229 4 vdd
port 513 nsew
rlabel metal1 s 20976 47649 20976 47649 4 vdd
port 513 nsew
rlabel metal1 s 21456 50310 21456 50310 4 vdd
port 513 nsew
rlabel metal1 s 21456 48730 21456 48730 4 vdd
port 513 nsew
rlabel metal1 s 20976 50019 20976 50019 4 vdd
port 513 nsew
rlabel metal1 s 22224 48439 22224 48439 4 vdd
port 513 nsew
rlabel metal1 s 22224 47940 22224 47940 4 vdd
port 513 nsew
rlabel metal1 s 20976 50310 20976 50310 4 vdd
port 513 nsew
rlabel metal1 s 21456 47649 21456 47649 4 vdd
port 513 nsew
rlabel metal1 s 20208 47940 20208 47940 4 vdd
port 513 nsew
rlabel metal1 s 20976 49229 20976 49229 4 vdd
port 513 nsew
rlabel metal1 s 20208 49229 20208 49229 4 vdd
port 513 nsew
rlabel metal1 s 20208 45570 20208 45570 4 vdd
port 513 nsew
rlabel metal1 s 22224 46360 22224 46360 4 vdd
port 513 nsew
rlabel metal1 s 20976 47150 20976 47150 4 vdd
port 513 nsew
rlabel metal1 s 22224 46859 22224 46859 4 vdd
port 513 nsew
rlabel metal1 s 21456 44780 21456 44780 4 vdd
port 513 nsew
rlabel metal1 s 21456 47150 21456 47150 4 vdd
port 513 nsew
rlabel metal1 s 20208 46069 20208 46069 4 vdd
port 513 nsew
rlabel metal1 s 20976 46859 20976 46859 4 vdd
port 513 nsew
rlabel metal1 s 20208 46859 20208 46859 4 vdd
port 513 nsew
rlabel metal1 s 20208 44780 20208 44780 4 vdd
port 513 nsew
rlabel metal1 s 20208 44489 20208 44489 4 vdd
port 513 nsew
rlabel metal1 s 20976 46069 20976 46069 4 vdd
port 513 nsew
rlabel metal1 s 21456 46360 21456 46360 4 vdd
port 513 nsew
rlabel metal1 s 20976 45570 20976 45570 4 vdd
port 513 nsew
rlabel metal1 s 21456 45279 21456 45279 4 vdd
port 513 nsew
rlabel metal1 s 20208 45279 20208 45279 4 vdd
port 513 nsew
rlabel metal1 s 21456 46069 21456 46069 4 vdd
port 513 nsew
rlabel metal1 s 22224 46069 22224 46069 4 vdd
port 513 nsew
rlabel metal1 s 20976 44780 20976 44780 4 vdd
port 513 nsew
rlabel metal1 s 21456 45570 21456 45570 4 vdd
port 513 nsew
rlabel metal1 s 22224 45279 22224 45279 4 vdd
port 513 nsew
rlabel metal1 s 22224 45570 22224 45570 4 vdd
port 513 nsew
rlabel metal1 s 22224 44489 22224 44489 4 vdd
port 513 nsew
rlabel metal1 s 22224 44780 22224 44780 4 vdd
port 513 nsew
rlabel metal1 s 20208 46360 20208 46360 4 vdd
port 513 nsew
rlabel metal1 s 20208 47150 20208 47150 4 vdd
port 513 nsew
rlabel metal1 s 20976 46360 20976 46360 4 vdd
port 513 nsew
rlabel metal1 s 20976 45279 20976 45279 4 vdd
port 513 nsew
rlabel metal1 s 21456 46859 21456 46859 4 vdd
port 513 nsew
rlabel metal1 s 22224 47150 22224 47150 4 vdd
port 513 nsew
rlabel metal1 s 21456 44489 21456 44489 4 vdd
port 513 nsew
rlabel metal1 s 20976 44489 20976 44489 4 vdd
port 513 nsew
rlabel metal1 s 24720 44489 24720 44489 4 vdd
port 513 nsew
rlabel metal1 s 23472 44489 23472 44489 4 vdd
port 513 nsew
rlabel metal1 s 22704 44489 22704 44489 4 vdd
port 513 nsew
rlabel metal1 s 23952 46859 23952 46859 4 vdd
port 513 nsew
rlabel metal1 s 23952 46069 23952 46069 4 vdd
port 513 nsew
rlabel metal1 s 23952 45279 23952 45279 4 vdd
port 513 nsew
rlabel metal1 s 23952 46360 23952 46360 4 vdd
port 513 nsew
rlabel metal1 s 22704 45279 22704 45279 4 vdd
port 513 nsew
rlabel metal1 s 23472 46859 23472 46859 4 vdd
port 513 nsew
rlabel metal1 s 23952 44780 23952 44780 4 vdd
port 513 nsew
rlabel metal1 s 23472 45279 23472 45279 4 vdd
port 513 nsew
rlabel metal1 s 24720 47150 24720 47150 4 vdd
port 513 nsew
rlabel metal1 s 22704 45570 22704 45570 4 vdd
port 513 nsew
rlabel metal1 s 22704 46360 22704 46360 4 vdd
port 513 nsew
rlabel metal1 s 23472 46360 23472 46360 4 vdd
port 513 nsew
rlabel metal1 s 22704 47150 22704 47150 4 vdd
port 513 nsew
rlabel metal1 s 23472 45570 23472 45570 4 vdd
port 513 nsew
rlabel metal1 s 23472 47150 23472 47150 4 vdd
port 513 nsew
rlabel metal1 s 24720 46069 24720 46069 4 vdd
port 513 nsew
rlabel metal1 s 22704 44780 22704 44780 4 vdd
port 513 nsew
rlabel metal1 s 23472 46069 23472 46069 4 vdd
port 513 nsew
rlabel metal1 s 22704 46069 22704 46069 4 vdd
port 513 nsew
rlabel metal1 s 24720 46360 24720 46360 4 vdd
port 513 nsew
rlabel metal1 s 23952 45570 23952 45570 4 vdd
port 513 nsew
rlabel metal1 s 23472 44780 23472 44780 4 vdd
port 513 nsew
rlabel metal1 s 24720 44780 24720 44780 4 vdd
port 513 nsew
rlabel metal1 s 23952 44489 23952 44489 4 vdd
port 513 nsew
rlabel metal1 s 23952 47150 23952 47150 4 vdd
port 513 nsew
rlabel metal1 s 24720 46859 24720 46859 4 vdd
port 513 nsew
rlabel metal1 s 24720 45279 24720 45279 4 vdd
port 513 nsew
rlabel metal1 s 22704 46859 22704 46859 4 vdd
port 513 nsew
rlabel metal1 s 24720 45570 24720 45570 4 vdd
port 513 nsew
rlabel metal1 s 23952 41620 23952 41620 4 vdd
port 513 nsew
rlabel metal1 s 23472 43200 23472 43200 4 vdd
port 513 nsew
rlabel metal1 s 22704 42909 22704 42909 4 vdd
port 513 nsew
rlabel metal1 s 23472 42119 23472 42119 4 vdd
port 513 nsew
rlabel metal1 s 22704 42119 22704 42119 4 vdd
port 513 nsew
rlabel metal1 s 22704 43699 22704 43699 4 vdd
port 513 nsew
rlabel metal1 s 24720 42119 24720 42119 4 vdd
port 513 nsew
rlabel metal1 s 23472 43990 23472 43990 4 vdd
port 513 nsew
rlabel metal1 s 24720 43699 24720 43699 4 vdd
port 513 nsew
rlabel metal1 s 24720 41620 24720 41620 4 vdd
port 513 nsew
rlabel metal1 s 23952 41329 23952 41329 4 vdd
port 513 nsew
rlabel metal1 s 23952 43200 23952 43200 4 vdd
port 513 nsew
rlabel metal1 s 23472 41620 23472 41620 4 vdd
port 513 nsew
rlabel metal1 s 24720 43990 24720 43990 4 vdd
port 513 nsew
rlabel metal1 s 24720 43200 24720 43200 4 vdd
port 513 nsew
rlabel metal1 s 24720 42909 24720 42909 4 vdd
port 513 nsew
rlabel metal1 s 24720 41329 24720 41329 4 vdd
port 513 nsew
rlabel metal1 s 24720 42410 24720 42410 4 vdd
port 513 nsew
rlabel metal1 s 22704 41620 22704 41620 4 vdd
port 513 nsew
rlabel metal1 s 23952 42909 23952 42909 4 vdd
port 513 nsew
rlabel metal1 s 23472 43699 23472 43699 4 vdd
port 513 nsew
rlabel metal1 s 23952 43990 23952 43990 4 vdd
port 513 nsew
rlabel metal1 s 23952 43699 23952 43699 4 vdd
port 513 nsew
rlabel metal1 s 22704 42410 22704 42410 4 vdd
port 513 nsew
rlabel metal1 s 22704 43200 22704 43200 4 vdd
port 513 nsew
rlabel metal1 s 23952 42119 23952 42119 4 vdd
port 513 nsew
rlabel metal1 s 22704 41329 22704 41329 4 vdd
port 513 nsew
rlabel metal1 s 23952 42410 23952 42410 4 vdd
port 513 nsew
rlabel metal1 s 23472 41329 23472 41329 4 vdd
port 513 nsew
rlabel metal1 s 23472 42410 23472 42410 4 vdd
port 513 nsew
rlabel metal1 s 22704 43990 22704 43990 4 vdd
port 513 nsew
rlabel metal1 s 23472 42909 23472 42909 4 vdd
port 513 nsew
rlabel metal1 s 22224 42410 22224 42410 4 vdd
port 513 nsew
rlabel metal1 s 20976 42909 20976 42909 4 vdd
port 513 nsew
rlabel metal1 s 20976 41620 20976 41620 4 vdd
port 513 nsew
rlabel metal1 s 20208 43699 20208 43699 4 vdd
port 513 nsew
rlabel metal1 s 21456 42909 21456 42909 4 vdd
port 513 nsew
rlabel metal1 s 20208 42909 20208 42909 4 vdd
port 513 nsew
rlabel metal1 s 20976 42410 20976 42410 4 vdd
port 513 nsew
rlabel metal1 s 20208 43200 20208 43200 4 vdd
port 513 nsew
rlabel metal1 s 20976 43699 20976 43699 4 vdd
port 513 nsew
rlabel metal1 s 22224 43200 22224 43200 4 vdd
port 513 nsew
rlabel metal1 s 20208 43990 20208 43990 4 vdd
port 513 nsew
rlabel metal1 s 20976 43200 20976 43200 4 vdd
port 513 nsew
rlabel metal1 s 20976 41329 20976 41329 4 vdd
port 513 nsew
rlabel metal1 s 21456 43200 21456 43200 4 vdd
port 513 nsew
rlabel metal1 s 22224 42119 22224 42119 4 vdd
port 513 nsew
rlabel metal1 s 20208 41329 20208 41329 4 vdd
port 513 nsew
rlabel metal1 s 21456 41329 21456 41329 4 vdd
port 513 nsew
rlabel metal1 s 22224 43699 22224 43699 4 vdd
port 513 nsew
rlabel metal1 s 20208 42119 20208 42119 4 vdd
port 513 nsew
rlabel metal1 s 22224 43990 22224 43990 4 vdd
port 513 nsew
rlabel metal1 s 21456 42119 21456 42119 4 vdd
port 513 nsew
rlabel metal1 s 21456 42410 21456 42410 4 vdd
port 513 nsew
rlabel metal1 s 22224 41620 22224 41620 4 vdd
port 513 nsew
rlabel metal1 s 20976 42119 20976 42119 4 vdd
port 513 nsew
rlabel metal1 s 20208 42410 20208 42410 4 vdd
port 513 nsew
rlabel metal1 s 21456 43990 21456 43990 4 vdd
port 513 nsew
rlabel metal1 s 21456 41620 21456 41620 4 vdd
port 513 nsew
rlabel metal1 s 20976 43990 20976 43990 4 vdd
port 513 nsew
rlabel metal1 s 21456 43699 21456 43699 4 vdd
port 513 nsew
rlabel metal1 s 22224 42909 22224 42909 4 vdd
port 513 nsew
rlabel metal1 s 22224 41329 22224 41329 4 vdd
port 513 nsew
rlabel metal1 s 20208 41620 20208 41620 4 vdd
port 513 nsew
rlabel metal1 s 21456 38460 21456 38460 4 vdd
port 513 nsew
rlabel metal1 s 20208 38169 20208 38169 4 vdd
port 513 nsew
rlabel metal1 s 20208 38959 20208 38959 4 vdd
port 513 nsew
rlabel metal1 s 20976 38169 20976 38169 4 vdd
port 513 nsew
rlabel metal1 s 21456 40830 21456 40830 4 vdd
port 513 nsew
rlabel metal1 s 22224 40040 22224 40040 4 vdd
port 513 nsew
rlabel metal1 s 21456 38169 21456 38169 4 vdd
port 513 nsew
rlabel metal1 s 22224 40830 22224 40830 4 vdd
port 513 nsew
rlabel metal1 s 20976 38959 20976 38959 4 vdd
port 513 nsew
rlabel metal1 s 20976 40040 20976 40040 4 vdd
port 513 nsew
rlabel metal1 s 20208 39749 20208 39749 4 vdd
port 513 nsew
rlabel metal1 s 20208 40830 20208 40830 4 vdd
port 513 nsew
rlabel metal1 s 20976 39749 20976 39749 4 vdd
port 513 nsew
rlabel metal1 s 21456 40040 21456 40040 4 vdd
port 513 nsew
rlabel metal1 s 20208 40539 20208 40539 4 vdd
port 513 nsew
rlabel metal1 s 20208 40040 20208 40040 4 vdd
port 513 nsew
rlabel metal1 s 20208 38460 20208 38460 4 vdd
port 513 nsew
rlabel metal1 s 22224 38169 22224 38169 4 vdd
port 513 nsew
rlabel metal1 s 22224 39250 22224 39250 4 vdd
port 513 nsew
rlabel metal1 s 21456 38959 21456 38959 4 vdd
port 513 nsew
rlabel metal1 s 22224 38460 22224 38460 4 vdd
port 513 nsew
rlabel metal1 s 21456 40539 21456 40539 4 vdd
port 513 nsew
rlabel metal1 s 20208 39250 20208 39250 4 vdd
port 513 nsew
rlabel metal1 s 21456 39250 21456 39250 4 vdd
port 513 nsew
rlabel metal1 s 20976 39250 20976 39250 4 vdd
port 513 nsew
rlabel metal1 s 20976 40830 20976 40830 4 vdd
port 513 nsew
rlabel metal1 s 20976 40539 20976 40539 4 vdd
port 513 nsew
rlabel metal1 s 21456 39749 21456 39749 4 vdd
port 513 nsew
rlabel metal1 s 20976 38460 20976 38460 4 vdd
port 513 nsew
rlabel metal1 s 22224 39749 22224 39749 4 vdd
port 513 nsew
rlabel metal1 s 22224 40539 22224 40539 4 vdd
port 513 nsew
rlabel metal1 s 22224 38959 22224 38959 4 vdd
port 513 nsew
rlabel metal1 s 23472 39250 23472 39250 4 vdd
port 513 nsew
rlabel metal1 s 22704 38460 22704 38460 4 vdd
port 513 nsew
rlabel metal1 s 23952 38959 23952 38959 4 vdd
port 513 nsew
rlabel metal1 s 22704 38959 22704 38959 4 vdd
port 513 nsew
rlabel metal1 s 24720 38169 24720 38169 4 vdd
port 513 nsew
rlabel metal1 s 22704 39749 22704 39749 4 vdd
port 513 nsew
rlabel metal1 s 22704 38169 22704 38169 4 vdd
port 513 nsew
rlabel metal1 s 22704 40830 22704 40830 4 vdd
port 513 nsew
rlabel metal1 s 24720 39749 24720 39749 4 vdd
port 513 nsew
rlabel metal1 s 22704 39250 22704 39250 4 vdd
port 513 nsew
rlabel metal1 s 23472 38169 23472 38169 4 vdd
port 513 nsew
rlabel metal1 s 23472 38460 23472 38460 4 vdd
port 513 nsew
rlabel metal1 s 24720 39250 24720 39250 4 vdd
port 513 nsew
rlabel metal1 s 24720 40539 24720 40539 4 vdd
port 513 nsew
rlabel metal1 s 22704 40040 22704 40040 4 vdd
port 513 nsew
rlabel metal1 s 24720 38460 24720 38460 4 vdd
port 513 nsew
rlabel metal1 s 24720 40830 24720 40830 4 vdd
port 513 nsew
rlabel metal1 s 23952 39749 23952 39749 4 vdd
port 513 nsew
rlabel metal1 s 24720 40040 24720 40040 4 vdd
port 513 nsew
rlabel metal1 s 24720 38959 24720 38959 4 vdd
port 513 nsew
rlabel metal1 s 23472 40040 23472 40040 4 vdd
port 513 nsew
rlabel metal1 s 22704 40539 22704 40539 4 vdd
port 513 nsew
rlabel metal1 s 23952 38460 23952 38460 4 vdd
port 513 nsew
rlabel metal1 s 23472 40539 23472 40539 4 vdd
port 513 nsew
rlabel metal1 s 23952 39250 23952 39250 4 vdd
port 513 nsew
rlabel metal1 s 23952 40830 23952 40830 4 vdd
port 513 nsew
rlabel metal1 s 23952 38169 23952 38169 4 vdd
port 513 nsew
rlabel metal1 s 23952 40539 23952 40539 4 vdd
port 513 nsew
rlabel metal1 s 23472 40830 23472 40830 4 vdd
port 513 nsew
rlabel metal1 s 23472 39749 23472 39749 4 vdd
port 513 nsew
rlabel metal1 s 23472 38959 23472 38959 4 vdd
port 513 nsew
rlabel metal1 s 23952 40040 23952 40040 4 vdd
port 513 nsew
rlabel metal1 s 28944 43699 28944 43699 4 vdd
port 513 nsew
rlabel metal1 s 28464 43990 28464 43990 4 vdd
port 513 nsew
rlabel metal1 s 29712 42909 29712 42909 4 vdd
port 513 nsew
rlabel metal1 s 29712 43990 29712 43990 4 vdd
port 513 nsew
rlabel metal1 s 27696 43200 27696 43200 4 vdd
port 513 nsew
rlabel metal1 s 28464 42410 28464 42410 4 vdd
port 513 nsew
rlabel metal1 s 27696 43990 27696 43990 4 vdd
port 513 nsew
rlabel metal1 s 28464 43200 28464 43200 4 vdd
port 513 nsew
rlabel metal1 s 28944 41329 28944 41329 4 vdd
port 513 nsew
rlabel metal1 s 27696 41620 27696 41620 4 vdd
port 513 nsew
rlabel metal1 s 29712 43200 29712 43200 4 vdd
port 513 nsew
rlabel metal1 s 28464 42909 28464 42909 4 vdd
port 513 nsew
rlabel metal1 s 28944 43200 28944 43200 4 vdd
port 513 nsew
rlabel metal1 s 29712 42410 29712 42410 4 vdd
port 513 nsew
rlabel metal1 s 27696 43699 27696 43699 4 vdd
port 513 nsew
rlabel metal1 s 28464 42119 28464 42119 4 vdd
port 513 nsew
rlabel metal1 s 29712 43699 29712 43699 4 vdd
port 513 nsew
rlabel metal1 s 28464 43699 28464 43699 4 vdd
port 513 nsew
rlabel metal1 s 28944 42410 28944 42410 4 vdd
port 513 nsew
rlabel metal1 s 27696 42119 27696 42119 4 vdd
port 513 nsew
rlabel metal1 s 27696 41329 27696 41329 4 vdd
port 513 nsew
rlabel metal1 s 29712 41620 29712 41620 4 vdd
port 513 nsew
rlabel metal1 s 28944 43990 28944 43990 4 vdd
port 513 nsew
rlabel metal1 s 29712 41329 29712 41329 4 vdd
port 513 nsew
rlabel metal1 s 28944 42909 28944 42909 4 vdd
port 513 nsew
rlabel metal1 s 28464 41620 28464 41620 4 vdd
port 513 nsew
rlabel metal1 s 27696 42410 27696 42410 4 vdd
port 513 nsew
rlabel metal1 s 28464 41329 28464 41329 4 vdd
port 513 nsew
rlabel metal1 s 28944 42119 28944 42119 4 vdd
port 513 nsew
rlabel metal1 s 28944 41620 28944 41620 4 vdd
port 513 nsew
rlabel metal1 s 29712 42119 29712 42119 4 vdd
port 513 nsew
rlabel metal1 s 27696 42909 27696 42909 4 vdd
port 513 nsew
rlabel metal1 s 27216 42410 27216 42410 4 vdd
port 513 nsew
rlabel metal1 s 26448 41329 26448 41329 4 vdd
port 513 nsew
rlabel metal1 s 27216 43699 27216 43699 4 vdd
port 513 nsew
rlabel metal1 s 25200 42909 25200 42909 4 vdd
port 513 nsew
rlabel metal1 s 25968 43200 25968 43200 4 vdd
port 513 nsew
rlabel metal1 s 27216 43990 27216 43990 4 vdd
port 513 nsew
rlabel metal1 s 27216 43200 27216 43200 4 vdd
port 513 nsew
rlabel metal1 s 25200 43200 25200 43200 4 vdd
port 513 nsew
rlabel metal1 s 26448 42410 26448 42410 4 vdd
port 513 nsew
rlabel metal1 s 25968 42119 25968 42119 4 vdd
port 513 nsew
rlabel metal1 s 25968 41329 25968 41329 4 vdd
port 513 nsew
rlabel metal1 s 26448 43990 26448 43990 4 vdd
port 513 nsew
rlabel metal1 s 25200 42410 25200 42410 4 vdd
port 513 nsew
rlabel metal1 s 25200 43990 25200 43990 4 vdd
port 513 nsew
rlabel metal1 s 26448 42909 26448 42909 4 vdd
port 513 nsew
rlabel metal1 s 27216 42909 27216 42909 4 vdd
port 513 nsew
rlabel metal1 s 25968 41620 25968 41620 4 vdd
port 513 nsew
rlabel metal1 s 25200 41329 25200 41329 4 vdd
port 513 nsew
rlabel metal1 s 25200 42119 25200 42119 4 vdd
port 513 nsew
rlabel metal1 s 27216 41620 27216 41620 4 vdd
port 513 nsew
rlabel metal1 s 26448 42119 26448 42119 4 vdd
port 513 nsew
rlabel metal1 s 26448 41620 26448 41620 4 vdd
port 513 nsew
rlabel metal1 s 25200 41620 25200 41620 4 vdd
port 513 nsew
rlabel metal1 s 25968 42909 25968 42909 4 vdd
port 513 nsew
rlabel metal1 s 25968 43990 25968 43990 4 vdd
port 513 nsew
rlabel metal1 s 26448 43699 26448 43699 4 vdd
port 513 nsew
rlabel metal1 s 25968 43699 25968 43699 4 vdd
port 513 nsew
rlabel metal1 s 25968 42410 25968 42410 4 vdd
port 513 nsew
rlabel metal1 s 27216 41329 27216 41329 4 vdd
port 513 nsew
rlabel metal1 s 27216 42119 27216 42119 4 vdd
port 513 nsew
rlabel metal1 s 26448 43200 26448 43200 4 vdd
port 513 nsew
rlabel metal1 s 25200 43699 25200 43699 4 vdd
port 513 nsew
rlabel metal1 s 25968 38460 25968 38460 4 vdd
port 513 nsew
rlabel metal1 s 25200 38959 25200 38959 4 vdd
port 513 nsew
rlabel metal1 s 25200 39250 25200 39250 4 vdd
port 513 nsew
rlabel metal1 s 25968 40830 25968 40830 4 vdd
port 513 nsew
rlabel metal1 s 27216 38959 27216 38959 4 vdd
port 513 nsew
rlabel metal1 s 25200 38169 25200 38169 4 vdd
port 513 nsew
rlabel metal1 s 26448 39749 26448 39749 4 vdd
port 513 nsew
rlabel metal1 s 26448 39250 26448 39250 4 vdd
port 513 nsew
rlabel metal1 s 25968 38169 25968 38169 4 vdd
port 513 nsew
rlabel metal1 s 25968 39250 25968 39250 4 vdd
port 513 nsew
rlabel metal1 s 25968 40539 25968 40539 4 vdd
port 513 nsew
rlabel metal1 s 26448 40539 26448 40539 4 vdd
port 513 nsew
rlabel metal1 s 27216 40830 27216 40830 4 vdd
port 513 nsew
rlabel metal1 s 25200 38460 25200 38460 4 vdd
port 513 nsew
rlabel metal1 s 25200 40040 25200 40040 4 vdd
port 513 nsew
rlabel metal1 s 27216 40539 27216 40539 4 vdd
port 513 nsew
rlabel metal1 s 27216 40040 27216 40040 4 vdd
port 513 nsew
rlabel metal1 s 25200 40830 25200 40830 4 vdd
port 513 nsew
rlabel metal1 s 26448 38460 26448 38460 4 vdd
port 513 nsew
rlabel metal1 s 25968 39749 25968 39749 4 vdd
port 513 nsew
rlabel metal1 s 27216 39749 27216 39749 4 vdd
port 513 nsew
rlabel metal1 s 26448 40830 26448 40830 4 vdd
port 513 nsew
rlabel metal1 s 27216 39250 27216 39250 4 vdd
port 513 nsew
rlabel metal1 s 26448 38169 26448 38169 4 vdd
port 513 nsew
rlabel metal1 s 27216 38460 27216 38460 4 vdd
port 513 nsew
rlabel metal1 s 26448 40040 26448 40040 4 vdd
port 513 nsew
rlabel metal1 s 25200 39749 25200 39749 4 vdd
port 513 nsew
rlabel metal1 s 25968 38959 25968 38959 4 vdd
port 513 nsew
rlabel metal1 s 26448 38959 26448 38959 4 vdd
port 513 nsew
rlabel metal1 s 25200 40539 25200 40539 4 vdd
port 513 nsew
rlabel metal1 s 27216 38169 27216 38169 4 vdd
port 513 nsew
rlabel metal1 s 25968 40040 25968 40040 4 vdd
port 513 nsew
rlabel metal1 s 28944 40539 28944 40539 4 vdd
port 513 nsew
rlabel metal1 s 28944 40040 28944 40040 4 vdd
port 513 nsew
rlabel metal1 s 28464 39250 28464 39250 4 vdd
port 513 nsew
rlabel metal1 s 27696 38959 27696 38959 4 vdd
port 513 nsew
rlabel metal1 s 27696 39250 27696 39250 4 vdd
port 513 nsew
rlabel metal1 s 28464 38959 28464 38959 4 vdd
port 513 nsew
rlabel metal1 s 28944 40830 28944 40830 4 vdd
port 513 nsew
rlabel metal1 s 28464 40830 28464 40830 4 vdd
port 513 nsew
rlabel metal1 s 27696 38169 27696 38169 4 vdd
port 513 nsew
rlabel metal1 s 29712 39250 29712 39250 4 vdd
port 513 nsew
rlabel metal1 s 28464 39749 28464 39749 4 vdd
port 513 nsew
rlabel metal1 s 28944 39749 28944 39749 4 vdd
port 513 nsew
rlabel metal1 s 29712 40040 29712 40040 4 vdd
port 513 nsew
rlabel metal1 s 28944 38959 28944 38959 4 vdd
port 513 nsew
rlabel metal1 s 29712 40539 29712 40539 4 vdd
port 513 nsew
rlabel metal1 s 28464 40539 28464 40539 4 vdd
port 513 nsew
rlabel metal1 s 27696 38460 27696 38460 4 vdd
port 513 nsew
rlabel metal1 s 28464 38169 28464 38169 4 vdd
port 513 nsew
rlabel metal1 s 28464 38460 28464 38460 4 vdd
port 513 nsew
rlabel metal1 s 28944 38169 28944 38169 4 vdd
port 513 nsew
rlabel metal1 s 28464 40040 28464 40040 4 vdd
port 513 nsew
rlabel metal1 s 27696 40830 27696 40830 4 vdd
port 513 nsew
rlabel metal1 s 27696 40539 27696 40539 4 vdd
port 513 nsew
rlabel metal1 s 29712 38460 29712 38460 4 vdd
port 513 nsew
rlabel metal1 s 28944 38460 28944 38460 4 vdd
port 513 nsew
rlabel metal1 s 29712 38959 29712 38959 4 vdd
port 513 nsew
rlabel metal1 s 29712 40830 29712 40830 4 vdd
port 513 nsew
rlabel metal1 s 27696 39749 27696 39749 4 vdd
port 513 nsew
rlabel metal1 s 29712 38169 29712 38169 4 vdd
port 513 nsew
rlabel metal1 s 28944 39250 28944 39250 4 vdd
port 513 nsew
rlabel metal1 s 29712 39749 29712 39749 4 vdd
port 513 nsew
rlabel metal1 s 27696 40040 27696 40040 4 vdd
port 513 nsew
rlabel metal1 s 29712 37379 29712 37379 4 vdd
port 513 nsew
rlabel metal1 s 28944 35300 28944 35300 4 vdd
port 513 nsew
rlabel metal1 s 29712 36880 29712 36880 4 vdd
port 513 nsew
rlabel metal1 s 27696 36090 27696 36090 4 vdd
port 513 nsew
rlabel metal1 s 28944 35009 28944 35009 4 vdd
port 513 nsew
rlabel metal1 s 27696 37670 27696 37670 4 vdd
port 513 nsew
rlabel metal1 s 29712 35300 29712 35300 4 vdd
port 513 nsew
rlabel metal1 s 27696 36589 27696 36589 4 vdd
port 513 nsew
rlabel metal1 s 28944 37379 28944 37379 4 vdd
port 513 nsew
rlabel metal1 s 27696 35009 27696 35009 4 vdd
port 513 nsew
rlabel metal1 s 27696 35799 27696 35799 4 vdd
port 513 nsew
rlabel metal1 s 27696 37379 27696 37379 4 vdd
port 513 nsew
rlabel metal1 s 28464 36589 28464 36589 4 vdd
port 513 nsew
rlabel metal1 s 29712 35009 29712 35009 4 vdd
port 513 nsew
rlabel metal1 s 29712 37670 29712 37670 4 vdd
port 513 nsew
rlabel metal1 s 28464 36090 28464 36090 4 vdd
port 513 nsew
rlabel metal1 s 28944 36589 28944 36589 4 vdd
port 513 nsew
rlabel metal1 s 28944 36880 28944 36880 4 vdd
port 513 nsew
rlabel metal1 s 28464 35009 28464 35009 4 vdd
port 513 nsew
rlabel metal1 s 28464 36880 28464 36880 4 vdd
port 513 nsew
rlabel metal1 s 28464 35300 28464 35300 4 vdd
port 513 nsew
rlabel metal1 s 28944 37670 28944 37670 4 vdd
port 513 nsew
rlabel metal1 s 27696 35300 27696 35300 4 vdd
port 513 nsew
rlabel metal1 s 28464 35799 28464 35799 4 vdd
port 513 nsew
rlabel metal1 s 29712 36090 29712 36090 4 vdd
port 513 nsew
rlabel metal1 s 29712 36589 29712 36589 4 vdd
port 513 nsew
rlabel metal1 s 28944 36090 28944 36090 4 vdd
port 513 nsew
rlabel metal1 s 27696 36880 27696 36880 4 vdd
port 513 nsew
rlabel metal1 s 29712 35799 29712 35799 4 vdd
port 513 nsew
rlabel metal1 s 28464 37379 28464 37379 4 vdd
port 513 nsew
rlabel metal1 s 28464 37670 28464 37670 4 vdd
port 513 nsew
rlabel metal1 s 28944 35799 28944 35799 4 vdd
port 513 nsew
rlabel metal1 s 27216 35799 27216 35799 4 vdd
port 513 nsew
rlabel metal1 s 25968 35799 25968 35799 4 vdd
port 513 nsew
rlabel metal1 s 25200 37670 25200 37670 4 vdd
port 513 nsew
rlabel metal1 s 27216 35009 27216 35009 4 vdd
port 513 nsew
rlabel metal1 s 27216 36090 27216 36090 4 vdd
port 513 nsew
rlabel metal1 s 26448 37379 26448 37379 4 vdd
port 513 nsew
rlabel metal1 s 26448 35799 26448 35799 4 vdd
port 513 nsew
rlabel metal1 s 26448 36090 26448 36090 4 vdd
port 513 nsew
rlabel metal1 s 25200 36589 25200 36589 4 vdd
port 513 nsew
rlabel metal1 s 26448 37670 26448 37670 4 vdd
port 513 nsew
rlabel metal1 s 27216 35300 27216 35300 4 vdd
port 513 nsew
rlabel metal1 s 26448 35009 26448 35009 4 vdd
port 513 nsew
rlabel metal1 s 25200 37379 25200 37379 4 vdd
port 513 nsew
rlabel metal1 s 25200 35300 25200 35300 4 vdd
port 513 nsew
rlabel metal1 s 26448 36880 26448 36880 4 vdd
port 513 nsew
rlabel metal1 s 27216 37379 27216 37379 4 vdd
port 513 nsew
rlabel metal1 s 27216 36589 27216 36589 4 vdd
port 513 nsew
rlabel metal1 s 27216 37670 27216 37670 4 vdd
port 513 nsew
rlabel metal1 s 25200 35009 25200 35009 4 vdd
port 513 nsew
rlabel metal1 s 25968 37379 25968 37379 4 vdd
port 513 nsew
rlabel metal1 s 26448 35300 26448 35300 4 vdd
port 513 nsew
rlabel metal1 s 27216 36880 27216 36880 4 vdd
port 513 nsew
rlabel metal1 s 25968 36090 25968 36090 4 vdd
port 513 nsew
rlabel metal1 s 25200 36880 25200 36880 4 vdd
port 513 nsew
rlabel metal1 s 25968 35300 25968 35300 4 vdd
port 513 nsew
rlabel metal1 s 26448 36589 26448 36589 4 vdd
port 513 nsew
rlabel metal1 s 25200 35799 25200 35799 4 vdd
port 513 nsew
rlabel metal1 s 25968 36589 25968 36589 4 vdd
port 513 nsew
rlabel metal1 s 25200 36090 25200 36090 4 vdd
port 513 nsew
rlabel metal1 s 25968 37670 25968 37670 4 vdd
port 513 nsew
rlabel metal1 s 25968 36880 25968 36880 4 vdd
port 513 nsew
rlabel metal1 s 25968 35009 25968 35009 4 vdd
port 513 nsew
rlabel metal1 s 25968 32140 25968 32140 4 vdd
port 513 nsew
rlabel metal1 s 27216 32639 27216 32639 4 vdd
port 513 nsew
rlabel metal1 s 26448 33429 26448 33429 4 vdd
port 513 nsew
rlabel metal1 s 25200 32930 25200 32930 4 vdd
port 513 nsew
rlabel metal1 s 25200 34219 25200 34219 4 vdd
port 513 nsew
rlabel metal1 s 27216 34510 27216 34510 4 vdd
port 513 nsew
rlabel metal1 s 27216 34219 27216 34219 4 vdd
port 513 nsew
rlabel metal1 s 25968 34510 25968 34510 4 vdd
port 513 nsew
rlabel metal1 s 25968 32930 25968 32930 4 vdd
port 513 nsew
rlabel metal1 s 25200 34510 25200 34510 4 vdd
port 513 nsew
rlabel metal1 s 26448 32140 26448 32140 4 vdd
port 513 nsew
rlabel metal1 s 26448 31849 26448 31849 4 vdd
port 513 nsew
rlabel metal1 s 25200 33720 25200 33720 4 vdd
port 513 nsew
rlabel metal1 s 26448 34219 26448 34219 4 vdd
port 513 nsew
rlabel metal1 s 27216 33720 27216 33720 4 vdd
port 513 nsew
rlabel metal1 s 27216 31849 27216 31849 4 vdd
port 513 nsew
rlabel metal1 s 25200 32140 25200 32140 4 vdd
port 513 nsew
rlabel metal1 s 27216 32140 27216 32140 4 vdd
port 513 nsew
rlabel metal1 s 26448 32930 26448 32930 4 vdd
port 513 nsew
rlabel metal1 s 25968 31849 25968 31849 4 vdd
port 513 nsew
rlabel metal1 s 26448 34510 26448 34510 4 vdd
port 513 nsew
rlabel metal1 s 25200 31849 25200 31849 4 vdd
port 513 nsew
rlabel metal1 s 26448 32639 26448 32639 4 vdd
port 513 nsew
rlabel metal1 s 25968 32639 25968 32639 4 vdd
port 513 nsew
rlabel metal1 s 27216 33429 27216 33429 4 vdd
port 513 nsew
rlabel metal1 s 26448 33720 26448 33720 4 vdd
port 513 nsew
rlabel metal1 s 25200 32639 25200 32639 4 vdd
port 513 nsew
rlabel metal1 s 25200 33429 25200 33429 4 vdd
port 513 nsew
rlabel metal1 s 25968 34219 25968 34219 4 vdd
port 513 nsew
rlabel metal1 s 27216 32930 27216 32930 4 vdd
port 513 nsew
rlabel metal1 s 25968 33429 25968 33429 4 vdd
port 513 nsew
rlabel metal1 s 25968 33720 25968 33720 4 vdd
port 513 nsew
rlabel metal1 s 29712 34510 29712 34510 4 vdd
port 513 nsew
rlabel metal1 s 27696 31849 27696 31849 4 vdd
port 513 nsew
rlabel metal1 s 28944 32930 28944 32930 4 vdd
port 513 nsew
rlabel metal1 s 28944 32639 28944 32639 4 vdd
port 513 nsew
rlabel metal1 s 28464 32140 28464 32140 4 vdd
port 513 nsew
rlabel metal1 s 28944 31849 28944 31849 4 vdd
port 513 nsew
rlabel metal1 s 28464 34219 28464 34219 4 vdd
port 513 nsew
rlabel metal1 s 27696 33720 27696 33720 4 vdd
port 513 nsew
rlabel metal1 s 29712 31849 29712 31849 4 vdd
port 513 nsew
rlabel metal1 s 27696 32930 27696 32930 4 vdd
port 513 nsew
rlabel metal1 s 27696 34510 27696 34510 4 vdd
port 513 nsew
rlabel metal1 s 28464 31849 28464 31849 4 vdd
port 513 nsew
rlabel metal1 s 27696 33429 27696 33429 4 vdd
port 513 nsew
rlabel metal1 s 29712 33429 29712 33429 4 vdd
port 513 nsew
rlabel metal1 s 28944 34510 28944 34510 4 vdd
port 513 nsew
rlabel metal1 s 29712 32639 29712 32639 4 vdd
port 513 nsew
rlabel metal1 s 28464 34510 28464 34510 4 vdd
port 513 nsew
rlabel metal1 s 28944 32140 28944 32140 4 vdd
port 513 nsew
rlabel metal1 s 28944 33429 28944 33429 4 vdd
port 513 nsew
rlabel metal1 s 28464 32930 28464 32930 4 vdd
port 513 nsew
rlabel metal1 s 29712 32140 29712 32140 4 vdd
port 513 nsew
rlabel metal1 s 28464 33720 28464 33720 4 vdd
port 513 nsew
rlabel metal1 s 28944 34219 28944 34219 4 vdd
port 513 nsew
rlabel metal1 s 29712 34219 29712 34219 4 vdd
port 513 nsew
rlabel metal1 s 27696 32639 27696 32639 4 vdd
port 513 nsew
rlabel metal1 s 28464 32639 28464 32639 4 vdd
port 513 nsew
rlabel metal1 s 27696 32140 27696 32140 4 vdd
port 513 nsew
rlabel metal1 s 28944 33720 28944 33720 4 vdd
port 513 nsew
rlabel metal1 s 28464 33429 28464 33429 4 vdd
port 513 nsew
rlabel metal1 s 27696 34219 27696 34219 4 vdd
port 513 nsew
rlabel metal1 s 29712 32930 29712 32930 4 vdd
port 513 nsew
rlabel metal1 s 29712 33720 29712 33720 4 vdd
port 513 nsew
rlabel metal1 s 23952 37670 23952 37670 4 vdd
port 513 nsew
rlabel metal1 s 22704 37379 22704 37379 4 vdd
port 513 nsew
rlabel metal1 s 23472 37379 23472 37379 4 vdd
port 513 nsew
rlabel metal1 s 22704 36090 22704 36090 4 vdd
port 513 nsew
rlabel metal1 s 23952 36090 23952 36090 4 vdd
port 513 nsew
rlabel metal1 s 23952 35300 23952 35300 4 vdd
port 513 nsew
rlabel metal1 s 23472 37670 23472 37670 4 vdd
port 513 nsew
rlabel metal1 s 22704 35300 22704 35300 4 vdd
port 513 nsew
rlabel metal1 s 22704 37670 22704 37670 4 vdd
port 513 nsew
rlabel metal1 s 22704 35009 22704 35009 4 vdd
port 513 nsew
rlabel metal1 s 23952 35799 23952 35799 4 vdd
port 513 nsew
rlabel metal1 s 22704 36880 22704 36880 4 vdd
port 513 nsew
rlabel metal1 s 24720 35799 24720 35799 4 vdd
port 513 nsew
rlabel metal1 s 23472 35009 23472 35009 4 vdd
port 513 nsew
rlabel metal1 s 24720 36589 24720 36589 4 vdd
port 513 nsew
rlabel metal1 s 23952 35009 23952 35009 4 vdd
port 513 nsew
rlabel metal1 s 23472 36880 23472 36880 4 vdd
port 513 nsew
rlabel metal1 s 24720 36880 24720 36880 4 vdd
port 513 nsew
rlabel metal1 s 23952 36880 23952 36880 4 vdd
port 513 nsew
rlabel metal1 s 23952 37379 23952 37379 4 vdd
port 513 nsew
rlabel metal1 s 23472 35300 23472 35300 4 vdd
port 513 nsew
rlabel metal1 s 23952 36589 23952 36589 4 vdd
port 513 nsew
rlabel metal1 s 24720 35300 24720 35300 4 vdd
port 513 nsew
rlabel metal1 s 24720 35009 24720 35009 4 vdd
port 513 nsew
rlabel metal1 s 24720 37379 24720 37379 4 vdd
port 513 nsew
rlabel metal1 s 24720 37670 24720 37670 4 vdd
port 513 nsew
rlabel metal1 s 23472 35799 23472 35799 4 vdd
port 513 nsew
rlabel metal1 s 24720 36090 24720 36090 4 vdd
port 513 nsew
rlabel metal1 s 22704 35799 22704 35799 4 vdd
port 513 nsew
rlabel metal1 s 23472 36589 23472 36589 4 vdd
port 513 nsew
rlabel metal1 s 23472 36090 23472 36090 4 vdd
port 513 nsew
rlabel metal1 s 22704 36589 22704 36589 4 vdd
port 513 nsew
rlabel metal1 s 21456 37379 21456 37379 4 vdd
port 513 nsew
rlabel metal1 s 21456 35009 21456 35009 4 vdd
port 513 nsew
rlabel metal1 s 21456 36090 21456 36090 4 vdd
port 513 nsew
rlabel metal1 s 22224 36090 22224 36090 4 vdd
port 513 nsew
rlabel metal1 s 20976 36090 20976 36090 4 vdd
port 513 nsew
rlabel metal1 s 20976 35799 20976 35799 4 vdd
port 513 nsew
rlabel metal1 s 22224 37379 22224 37379 4 vdd
port 513 nsew
rlabel metal1 s 21456 35799 21456 35799 4 vdd
port 513 nsew
rlabel metal1 s 20976 37670 20976 37670 4 vdd
port 513 nsew
rlabel metal1 s 22224 35300 22224 35300 4 vdd
port 513 nsew
rlabel metal1 s 22224 35799 22224 35799 4 vdd
port 513 nsew
rlabel metal1 s 20976 35300 20976 35300 4 vdd
port 513 nsew
rlabel metal1 s 21456 35300 21456 35300 4 vdd
port 513 nsew
rlabel metal1 s 20208 35300 20208 35300 4 vdd
port 513 nsew
rlabel metal1 s 21456 37670 21456 37670 4 vdd
port 513 nsew
rlabel metal1 s 20976 35009 20976 35009 4 vdd
port 513 nsew
rlabel metal1 s 21456 36880 21456 36880 4 vdd
port 513 nsew
rlabel metal1 s 20976 37379 20976 37379 4 vdd
port 513 nsew
rlabel metal1 s 20976 36589 20976 36589 4 vdd
port 513 nsew
rlabel metal1 s 22224 35009 22224 35009 4 vdd
port 513 nsew
rlabel metal1 s 20976 36880 20976 36880 4 vdd
port 513 nsew
rlabel metal1 s 20208 37670 20208 37670 4 vdd
port 513 nsew
rlabel metal1 s 20208 35799 20208 35799 4 vdd
port 513 nsew
rlabel metal1 s 22224 37670 22224 37670 4 vdd
port 513 nsew
rlabel metal1 s 20208 35009 20208 35009 4 vdd
port 513 nsew
rlabel metal1 s 22224 36589 22224 36589 4 vdd
port 513 nsew
rlabel metal1 s 21456 36589 21456 36589 4 vdd
port 513 nsew
rlabel metal1 s 20208 37379 20208 37379 4 vdd
port 513 nsew
rlabel metal1 s 20208 36090 20208 36090 4 vdd
port 513 nsew
rlabel metal1 s 22224 36880 22224 36880 4 vdd
port 513 nsew
rlabel metal1 s 20208 36880 20208 36880 4 vdd
port 513 nsew
rlabel metal1 s 20208 36589 20208 36589 4 vdd
port 513 nsew
rlabel metal1 s 22224 34510 22224 34510 4 vdd
port 513 nsew
rlabel metal1 s 20208 33720 20208 33720 4 vdd
port 513 nsew
rlabel metal1 s 22224 34219 22224 34219 4 vdd
port 513 nsew
rlabel metal1 s 22224 31849 22224 31849 4 vdd
port 513 nsew
rlabel metal1 s 20976 34219 20976 34219 4 vdd
port 513 nsew
rlabel metal1 s 22224 33429 22224 33429 4 vdd
port 513 nsew
rlabel metal1 s 21456 34510 21456 34510 4 vdd
port 513 nsew
rlabel metal1 s 20208 34510 20208 34510 4 vdd
port 513 nsew
rlabel metal1 s 21456 33720 21456 33720 4 vdd
port 513 nsew
rlabel metal1 s 21456 32930 21456 32930 4 vdd
port 513 nsew
rlabel metal1 s 21456 33429 21456 33429 4 vdd
port 513 nsew
rlabel metal1 s 20976 32140 20976 32140 4 vdd
port 513 nsew
rlabel metal1 s 20208 31849 20208 31849 4 vdd
port 513 nsew
rlabel metal1 s 22224 32639 22224 32639 4 vdd
port 513 nsew
rlabel metal1 s 20208 32639 20208 32639 4 vdd
port 513 nsew
rlabel metal1 s 22224 32930 22224 32930 4 vdd
port 513 nsew
rlabel metal1 s 20976 33720 20976 33720 4 vdd
port 513 nsew
rlabel metal1 s 20208 34219 20208 34219 4 vdd
port 513 nsew
rlabel metal1 s 20208 32930 20208 32930 4 vdd
port 513 nsew
rlabel metal1 s 21456 31849 21456 31849 4 vdd
port 513 nsew
rlabel metal1 s 21456 32140 21456 32140 4 vdd
port 513 nsew
rlabel metal1 s 22224 33720 22224 33720 4 vdd
port 513 nsew
rlabel metal1 s 21456 32639 21456 32639 4 vdd
port 513 nsew
rlabel metal1 s 20976 32930 20976 32930 4 vdd
port 513 nsew
rlabel metal1 s 20208 32140 20208 32140 4 vdd
port 513 nsew
rlabel metal1 s 22224 32140 22224 32140 4 vdd
port 513 nsew
rlabel metal1 s 20208 33429 20208 33429 4 vdd
port 513 nsew
rlabel metal1 s 21456 34219 21456 34219 4 vdd
port 513 nsew
rlabel metal1 s 20976 34510 20976 34510 4 vdd
port 513 nsew
rlabel metal1 s 20976 32639 20976 32639 4 vdd
port 513 nsew
rlabel metal1 s 20976 33429 20976 33429 4 vdd
port 513 nsew
rlabel metal1 s 20976 31849 20976 31849 4 vdd
port 513 nsew
rlabel metal1 s 24720 33720 24720 33720 4 vdd
port 513 nsew
rlabel metal1 s 24720 32930 24720 32930 4 vdd
port 513 nsew
rlabel metal1 s 23472 31849 23472 31849 4 vdd
port 513 nsew
rlabel metal1 s 23472 34219 23472 34219 4 vdd
port 513 nsew
rlabel metal1 s 24720 31849 24720 31849 4 vdd
port 513 nsew
rlabel metal1 s 23952 33720 23952 33720 4 vdd
port 513 nsew
rlabel metal1 s 23472 32639 23472 32639 4 vdd
port 513 nsew
rlabel metal1 s 24720 32140 24720 32140 4 vdd
port 513 nsew
rlabel metal1 s 23952 32639 23952 32639 4 vdd
port 513 nsew
rlabel metal1 s 22704 32930 22704 32930 4 vdd
port 513 nsew
rlabel metal1 s 23952 33429 23952 33429 4 vdd
port 513 nsew
rlabel metal1 s 22704 34510 22704 34510 4 vdd
port 513 nsew
rlabel metal1 s 24720 34510 24720 34510 4 vdd
port 513 nsew
rlabel metal1 s 24720 34219 24720 34219 4 vdd
port 513 nsew
rlabel metal1 s 23952 32140 23952 32140 4 vdd
port 513 nsew
rlabel metal1 s 23472 32140 23472 32140 4 vdd
port 513 nsew
rlabel metal1 s 23952 34510 23952 34510 4 vdd
port 513 nsew
rlabel metal1 s 23472 33720 23472 33720 4 vdd
port 513 nsew
rlabel metal1 s 24720 32639 24720 32639 4 vdd
port 513 nsew
rlabel metal1 s 23952 31849 23952 31849 4 vdd
port 513 nsew
rlabel metal1 s 23472 33429 23472 33429 4 vdd
port 513 nsew
rlabel metal1 s 23952 32930 23952 32930 4 vdd
port 513 nsew
rlabel metal1 s 22704 32140 22704 32140 4 vdd
port 513 nsew
rlabel metal1 s 22704 34219 22704 34219 4 vdd
port 513 nsew
rlabel metal1 s 22704 33720 22704 33720 4 vdd
port 513 nsew
rlabel metal1 s 22704 32639 22704 32639 4 vdd
port 513 nsew
rlabel metal1 s 23952 34219 23952 34219 4 vdd
port 513 nsew
rlabel metal1 s 23472 34510 23472 34510 4 vdd
port 513 nsew
rlabel metal1 s 22704 31849 22704 31849 4 vdd
port 513 nsew
rlabel metal1 s 23472 32930 23472 32930 4 vdd
port 513 nsew
rlabel metal1 s 24720 33429 24720 33429 4 vdd
port 513 nsew
rlabel metal1 s 22704 33429 22704 33429 4 vdd
port 513 nsew
rlabel metal1 s 23952 30269 23952 30269 4 vdd
port 513 nsew
rlabel metal1 s 22704 29770 22704 29770 4 vdd
port 513 nsew
rlabel metal1 s 23472 30560 23472 30560 4 vdd
port 513 nsew
rlabel metal1 s 23952 30560 23952 30560 4 vdd
port 513 nsew
rlabel metal1 s 22704 31350 22704 31350 4 vdd
port 513 nsew
rlabel metal1 s 22704 28980 22704 28980 4 vdd
port 513 nsew
rlabel metal1 s 23472 31059 23472 31059 4 vdd
port 513 nsew
rlabel metal1 s 22704 28689 22704 28689 4 vdd
port 513 nsew
rlabel metal1 s 23952 29770 23952 29770 4 vdd
port 513 nsew
rlabel metal1 s 24720 30269 24720 30269 4 vdd
port 513 nsew
rlabel metal1 s 23472 28980 23472 28980 4 vdd
port 513 nsew
rlabel metal1 s 23472 30269 23472 30269 4 vdd
port 513 nsew
rlabel metal1 s 23472 29770 23472 29770 4 vdd
port 513 nsew
rlabel metal1 s 23952 29479 23952 29479 4 vdd
port 513 nsew
rlabel metal1 s 23952 31350 23952 31350 4 vdd
port 513 nsew
rlabel metal1 s 23952 31059 23952 31059 4 vdd
port 513 nsew
rlabel metal1 s 24720 31350 24720 31350 4 vdd
port 513 nsew
rlabel metal1 s 23952 28980 23952 28980 4 vdd
port 513 nsew
rlabel metal1 s 24720 29770 24720 29770 4 vdd
port 513 nsew
rlabel metal1 s 23952 28689 23952 28689 4 vdd
port 513 nsew
rlabel metal1 s 24720 28689 24720 28689 4 vdd
port 513 nsew
rlabel metal1 s 24720 30560 24720 30560 4 vdd
port 513 nsew
rlabel metal1 s 22704 30560 22704 30560 4 vdd
port 513 nsew
rlabel metal1 s 23472 29479 23472 29479 4 vdd
port 513 nsew
rlabel metal1 s 24720 28980 24720 28980 4 vdd
port 513 nsew
rlabel metal1 s 22704 30269 22704 30269 4 vdd
port 513 nsew
rlabel metal1 s 23472 28689 23472 28689 4 vdd
port 513 nsew
rlabel metal1 s 22704 29479 22704 29479 4 vdd
port 513 nsew
rlabel metal1 s 24720 31059 24720 31059 4 vdd
port 513 nsew
rlabel metal1 s 24720 29479 24720 29479 4 vdd
port 513 nsew
rlabel metal1 s 22704 31059 22704 31059 4 vdd
port 513 nsew
rlabel metal1 s 23472 31350 23472 31350 4 vdd
port 513 nsew
rlabel metal1 s 21456 28689 21456 28689 4 vdd
port 513 nsew
rlabel metal1 s 20208 29479 20208 29479 4 vdd
port 513 nsew
rlabel metal1 s 22224 29479 22224 29479 4 vdd
port 513 nsew
rlabel metal1 s 21456 29479 21456 29479 4 vdd
port 513 nsew
rlabel metal1 s 22224 28689 22224 28689 4 vdd
port 513 nsew
rlabel metal1 s 20208 30560 20208 30560 4 vdd
port 513 nsew
rlabel metal1 s 21456 31350 21456 31350 4 vdd
port 513 nsew
rlabel metal1 s 22224 28980 22224 28980 4 vdd
port 513 nsew
rlabel metal1 s 20976 29479 20976 29479 4 vdd
port 513 nsew
rlabel metal1 s 21456 31059 21456 31059 4 vdd
port 513 nsew
rlabel metal1 s 20976 30269 20976 30269 4 vdd
port 513 nsew
rlabel metal1 s 21456 30269 21456 30269 4 vdd
port 513 nsew
rlabel metal1 s 22224 30269 22224 30269 4 vdd
port 513 nsew
rlabel metal1 s 20208 29770 20208 29770 4 vdd
port 513 nsew
rlabel metal1 s 22224 29770 22224 29770 4 vdd
port 513 nsew
rlabel metal1 s 22224 31059 22224 31059 4 vdd
port 513 nsew
rlabel metal1 s 20976 31350 20976 31350 4 vdd
port 513 nsew
rlabel metal1 s 20976 28980 20976 28980 4 vdd
port 513 nsew
rlabel metal1 s 20976 30560 20976 30560 4 vdd
port 513 nsew
rlabel metal1 s 20208 28980 20208 28980 4 vdd
port 513 nsew
rlabel metal1 s 20208 28689 20208 28689 4 vdd
port 513 nsew
rlabel metal1 s 22224 30560 22224 30560 4 vdd
port 513 nsew
rlabel metal1 s 22224 31350 22224 31350 4 vdd
port 513 nsew
rlabel metal1 s 20976 31059 20976 31059 4 vdd
port 513 nsew
rlabel metal1 s 21456 28980 21456 28980 4 vdd
port 513 nsew
rlabel metal1 s 20976 29770 20976 29770 4 vdd
port 513 nsew
rlabel metal1 s 20208 30269 20208 30269 4 vdd
port 513 nsew
rlabel metal1 s 20976 28689 20976 28689 4 vdd
port 513 nsew
rlabel metal1 s 21456 30560 21456 30560 4 vdd
port 513 nsew
rlabel metal1 s 20208 31059 20208 31059 4 vdd
port 513 nsew
rlabel metal1 s 21456 29770 21456 29770 4 vdd
port 513 nsew
rlabel metal1 s 20208 31350 20208 31350 4 vdd
port 513 nsew
rlabel metal1 s 20976 27400 20976 27400 4 vdd
port 513 nsew
rlabel metal1 s 22224 28190 22224 28190 4 vdd
port 513 nsew
rlabel metal1 s 22224 27109 22224 27109 4 vdd
port 513 nsew
rlabel metal1 s 21456 27400 21456 27400 4 vdd
port 513 nsew
rlabel metal1 s 20976 28190 20976 28190 4 vdd
port 513 nsew
rlabel metal1 s 20208 28190 20208 28190 4 vdd
port 513 nsew
rlabel metal1 s 20976 26610 20976 26610 4 vdd
port 513 nsew
rlabel metal1 s 22224 25529 22224 25529 4 vdd
port 513 nsew
rlabel metal1 s 21456 27109 21456 27109 4 vdd
port 513 nsew
rlabel metal1 s 20976 26319 20976 26319 4 vdd
port 513 nsew
rlabel metal1 s 22224 27899 22224 27899 4 vdd
port 513 nsew
rlabel metal1 s 21456 26319 21456 26319 4 vdd
port 513 nsew
rlabel metal1 s 20976 27899 20976 27899 4 vdd
port 513 nsew
rlabel metal1 s 21456 26610 21456 26610 4 vdd
port 513 nsew
rlabel metal1 s 20208 25529 20208 25529 4 vdd
port 513 nsew
rlabel metal1 s 21456 25820 21456 25820 4 vdd
port 513 nsew
rlabel metal1 s 21456 27899 21456 27899 4 vdd
port 513 nsew
rlabel metal1 s 20208 27899 20208 27899 4 vdd
port 513 nsew
rlabel metal1 s 20208 27400 20208 27400 4 vdd
port 513 nsew
rlabel metal1 s 22224 27400 22224 27400 4 vdd
port 513 nsew
rlabel metal1 s 20208 25820 20208 25820 4 vdd
port 513 nsew
rlabel metal1 s 20976 25529 20976 25529 4 vdd
port 513 nsew
rlabel metal1 s 20208 26319 20208 26319 4 vdd
port 513 nsew
rlabel metal1 s 20208 26610 20208 26610 4 vdd
port 513 nsew
rlabel metal1 s 21456 28190 21456 28190 4 vdd
port 513 nsew
rlabel metal1 s 22224 26319 22224 26319 4 vdd
port 513 nsew
rlabel metal1 s 21456 25529 21456 25529 4 vdd
port 513 nsew
rlabel metal1 s 22224 26610 22224 26610 4 vdd
port 513 nsew
rlabel metal1 s 20208 27109 20208 27109 4 vdd
port 513 nsew
rlabel metal1 s 22224 25820 22224 25820 4 vdd
port 513 nsew
rlabel metal1 s 20976 25820 20976 25820 4 vdd
port 513 nsew
rlabel metal1 s 20976 27109 20976 27109 4 vdd
port 513 nsew
rlabel metal1 s 22704 27899 22704 27899 4 vdd
port 513 nsew
rlabel metal1 s 24720 28190 24720 28190 4 vdd
port 513 nsew
rlabel metal1 s 22704 26319 22704 26319 4 vdd
port 513 nsew
rlabel metal1 s 23952 27400 23952 27400 4 vdd
port 513 nsew
rlabel metal1 s 23472 27899 23472 27899 4 vdd
port 513 nsew
rlabel metal1 s 23472 27109 23472 27109 4 vdd
port 513 nsew
rlabel metal1 s 23952 26610 23952 26610 4 vdd
port 513 nsew
rlabel metal1 s 22704 25820 22704 25820 4 vdd
port 513 nsew
rlabel metal1 s 22704 26610 22704 26610 4 vdd
port 513 nsew
rlabel metal1 s 23472 25529 23472 25529 4 vdd
port 513 nsew
rlabel metal1 s 23952 27109 23952 27109 4 vdd
port 513 nsew
rlabel metal1 s 23952 25529 23952 25529 4 vdd
port 513 nsew
rlabel metal1 s 22704 25529 22704 25529 4 vdd
port 513 nsew
rlabel metal1 s 24720 25820 24720 25820 4 vdd
port 513 nsew
rlabel metal1 s 22704 28190 22704 28190 4 vdd
port 513 nsew
rlabel metal1 s 23952 26319 23952 26319 4 vdd
port 513 nsew
rlabel metal1 s 22704 27400 22704 27400 4 vdd
port 513 nsew
rlabel metal1 s 22704 27109 22704 27109 4 vdd
port 513 nsew
rlabel metal1 s 23472 25820 23472 25820 4 vdd
port 513 nsew
rlabel metal1 s 23952 27899 23952 27899 4 vdd
port 513 nsew
rlabel metal1 s 23952 28190 23952 28190 4 vdd
port 513 nsew
rlabel metal1 s 24720 25529 24720 25529 4 vdd
port 513 nsew
rlabel metal1 s 23952 25820 23952 25820 4 vdd
port 513 nsew
rlabel metal1 s 24720 27400 24720 27400 4 vdd
port 513 nsew
rlabel metal1 s 23472 27400 23472 27400 4 vdd
port 513 nsew
rlabel metal1 s 24720 26610 24720 26610 4 vdd
port 513 nsew
rlabel metal1 s 23472 26319 23472 26319 4 vdd
port 513 nsew
rlabel metal1 s 24720 26319 24720 26319 4 vdd
port 513 nsew
rlabel metal1 s 23472 26610 23472 26610 4 vdd
port 513 nsew
rlabel metal1 s 23472 28190 23472 28190 4 vdd
port 513 nsew
rlabel metal1 s 24720 27899 24720 27899 4 vdd
port 513 nsew
rlabel metal1 s 24720 27109 24720 27109 4 vdd
port 513 nsew
rlabel metal1 s 28464 29479 28464 29479 4 vdd
port 513 nsew
rlabel metal1 s 28464 28980 28464 28980 4 vdd
port 513 nsew
rlabel metal1 s 28464 28689 28464 28689 4 vdd
port 513 nsew
rlabel metal1 s 28944 29770 28944 29770 4 vdd
port 513 nsew
rlabel metal1 s 28944 30269 28944 30269 4 vdd
port 513 nsew
rlabel metal1 s 27696 28980 27696 28980 4 vdd
port 513 nsew
rlabel metal1 s 29712 28980 29712 28980 4 vdd
port 513 nsew
rlabel metal1 s 28944 31059 28944 31059 4 vdd
port 513 nsew
rlabel metal1 s 29712 29770 29712 29770 4 vdd
port 513 nsew
rlabel metal1 s 28464 31350 28464 31350 4 vdd
port 513 nsew
rlabel metal1 s 27696 31059 27696 31059 4 vdd
port 513 nsew
rlabel metal1 s 27696 30269 27696 30269 4 vdd
port 513 nsew
rlabel metal1 s 28944 29479 28944 29479 4 vdd
port 513 nsew
rlabel metal1 s 28464 30560 28464 30560 4 vdd
port 513 nsew
rlabel metal1 s 28944 28980 28944 28980 4 vdd
port 513 nsew
rlabel metal1 s 27696 29770 27696 29770 4 vdd
port 513 nsew
rlabel metal1 s 29712 31350 29712 31350 4 vdd
port 513 nsew
rlabel metal1 s 27696 29479 27696 29479 4 vdd
port 513 nsew
rlabel metal1 s 28464 29770 28464 29770 4 vdd
port 513 nsew
rlabel metal1 s 28944 31350 28944 31350 4 vdd
port 513 nsew
rlabel metal1 s 28944 28689 28944 28689 4 vdd
port 513 nsew
rlabel metal1 s 27696 30560 27696 30560 4 vdd
port 513 nsew
rlabel metal1 s 27696 31350 27696 31350 4 vdd
port 513 nsew
rlabel metal1 s 28944 30560 28944 30560 4 vdd
port 513 nsew
rlabel metal1 s 29712 30269 29712 30269 4 vdd
port 513 nsew
rlabel metal1 s 28464 31059 28464 31059 4 vdd
port 513 nsew
rlabel metal1 s 27696 28689 27696 28689 4 vdd
port 513 nsew
rlabel metal1 s 29712 30560 29712 30560 4 vdd
port 513 nsew
rlabel metal1 s 28464 30269 28464 30269 4 vdd
port 513 nsew
rlabel metal1 s 29712 29479 29712 29479 4 vdd
port 513 nsew
rlabel metal1 s 29712 28689 29712 28689 4 vdd
port 513 nsew
rlabel metal1 s 29712 31059 29712 31059 4 vdd
port 513 nsew
rlabel metal1 s 27216 29770 27216 29770 4 vdd
port 513 nsew
rlabel metal1 s 25968 30560 25968 30560 4 vdd
port 513 nsew
rlabel metal1 s 27216 31350 27216 31350 4 vdd
port 513 nsew
rlabel metal1 s 25200 28689 25200 28689 4 vdd
port 513 nsew
rlabel metal1 s 25968 30269 25968 30269 4 vdd
port 513 nsew
rlabel metal1 s 27216 28689 27216 28689 4 vdd
port 513 nsew
rlabel metal1 s 25968 29479 25968 29479 4 vdd
port 513 nsew
rlabel metal1 s 25200 29479 25200 29479 4 vdd
port 513 nsew
rlabel metal1 s 25200 30269 25200 30269 4 vdd
port 513 nsew
rlabel metal1 s 25968 31059 25968 31059 4 vdd
port 513 nsew
rlabel metal1 s 26448 31350 26448 31350 4 vdd
port 513 nsew
rlabel metal1 s 27216 31059 27216 31059 4 vdd
port 513 nsew
rlabel metal1 s 25200 30560 25200 30560 4 vdd
port 513 nsew
rlabel metal1 s 26448 29479 26448 29479 4 vdd
port 513 nsew
rlabel metal1 s 27216 29479 27216 29479 4 vdd
port 513 nsew
rlabel metal1 s 27216 30269 27216 30269 4 vdd
port 513 nsew
rlabel metal1 s 25200 29770 25200 29770 4 vdd
port 513 nsew
rlabel metal1 s 25200 28980 25200 28980 4 vdd
port 513 nsew
rlabel metal1 s 26448 29770 26448 29770 4 vdd
port 513 nsew
rlabel metal1 s 25200 31350 25200 31350 4 vdd
port 513 nsew
rlabel metal1 s 26448 28980 26448 28980 4 vdd
port 513 nsew
rlabel metal1 s 25968 28689 25968 28689 4 vdd
port 513 nsew
rlabel metal1 s 25968 29770 25968 29770 4 vdd
port 513 nsew
rlabel metal1 s 25968 28980 25968 28980 4 vdd
port 513 nsew
rlabel metal1 s 25200 31059 25200 31059 4 vdd
port 513 nsew
rlabel metal1 s 26448 30269 26448 30269 4 vdd
port 513 nsew
rlabel metal1 s 25968 31350 25968 31350 4 vdd
port 513 nsew
rlabel metal1 s 26448 31059 26448 31059 4 vdd
port 513 nsew
rlabel metal1 s 27216 28980 27216 28980 4 vdd
port 513 nsew
rlabel metal1 s 27216 30560 27216 30560 4 vdd
port 513 nsew
rlabel metal1 s 26448 28689 26448 28689 4 vdd
port 513 nsew
rlabel metal1 s 26448 30560 26448 30560 4 vdd
port 513 nsew
rlabel metal1 s 26448 25820 26448 25820 4 vdd
port 513 nsew
rlabel metal1 s 25968 27109 25968 27109 4 vdd
port 513 nsew
rlabel metal1 s 26448 27400 26448 27400 4 vdd
port 513 nsew
rlabel metal1 s 25968 27400 25968 27400 4 vdd
port 513 nsew
rlabel metal1 s 26448 26319 26448 26319 4 vdd
port 513 nsew
rlabel metal1 s 27216 26319 27216 26319 4 vdd
port 513 nsew
rlabel metal1 s 25968 26319 25968 26319 4 vdd
port 513 nsew
rlabel metal1 s 26448 27109 26448 27109 4 vdd
port 513 nsew
rlabel metal1 s 27216 27400 27216 27400 4 vdd
port 513 nsew
rlabel metal1 s 25968 25529 25968 25529 4 vdd
port 513 nsew
rlabel metal1 s 25200 27109 25200 27109 4 vdd
port 513 nsew
rlabel metal1 s 25968 28190 25968 28190 4 vdd
port 513 nsew
rlabel metal1 s 27216 25820 27216 25820 4 vdd
port 513 nsew
rlabel metal1 s 25200 25820 25200 25820 4 vdd
port 513 nsew
rlabel metal1 s 27216 25529 27216 25529 4 vdd
port 513 nsew
rlabel metal1 s 26448 28190 26448 28190 4 vdd
port 513 nsew
rlabel metal1 s 27216 28190 27216 28190 4 vdd
port 513 nsew
rlabel metal1 s 25200 27400 25200 27400 4 vdd
port 513 nsew
rlabel metal1 s 27216 26610 27216 26610 4 vdd
port 513 nsew
rlabel metal1 s 26448 25529 26448 25529 4 vdd
port 513 nsew
rlabel metal1 s 25200 26319 25200 26319 4 vdd
port 513 nsew
rlabel metal1 s 25200 27899 25200 27899 4 vdd
port 513 nsew
rlabel metal1 s 25200 26610 25200 26610 4 vdd
port 513 nsew
rlabel metal1 s 25200 28190 25200 28190 4 vdd
port 513 nsew
rlabel metal1 s 27216 27109 27216 27109 4 vdd
port 513 nsew
rlabel metal1 s 26448 27899 26448 27899 4 vdd
port 513 nsew
rlabel metal1 s 27216 27899 27216 27899 4 vdd
port 513 nsew
rlabel metal1 s 25968 26610 25968 26610 4 vdd
port 513 nsew
rlabel metal1 s 25968 25820 25968 25820 4 vdd
port 513 nsew
rlabel metal1 s 25200 25529 25200 25529 4 vdd
port 513 nsew
rlabel metal1 s 25968 27899 25968 27899 4 vdd
port 513 nsew
rlabel metal1 s 26448 26610 26448 26610 4 vdd
port 513 nsew
rlabel metal1 s 28464 27400 28464 27400 4 vdd
port 513 nsew
rlabel metal1 s 28464 27109 28464 27109 4 vdd
port 513 nsew
rlabel metal1 s 27696 26319 27696 26319 4 vdd
port 513 nsew
rlabel metal1 s 27696 25820 27696 25820 4 vdd
port 513 nsew
rlabel metal1 s 28944 27109 28944 27109 4 vdd
port 513 nsew
rlabel metal1 s 28944 25529 28944 25529 4 vdd
port 513 nsew
rlabel metal1 s 29712 25820 29712 25820 4 vdd
port 513 nsew
rlabel metal1 s 27696 26610 27696 26610 4 vdd
port 513 nsew
rlabel metal1 s 28944 26610 28944 26610 4 vdd
port 513 nsew
rlabel metal1 s 27696 27109 27696 27109 4 vdd
port 513 nsew
rlabel metal1 s 29712 27899 29712 27899 4 vdd
port 513 nsew
rlabel metal1 s 29712 27109 29712 27109 4 vdd
port 513 nsew
rlabel metal1 s 28464 28190 28464 28190 4 vdd
port 513 nsew
rlabel metal1 s 29712 28190 29712 28190 4 vdd
port 513 nsew
rlabel metal1 s 27696 28190 27696 28190 4 vdd
port 513 nsew
rlabel metal1 s 29712 26319 29712 26319 4 vdd
port 513 nsew
rlabel metal1 s 28464 26319 28464 26319 4 vdd
port 513 nsew
rlabel metal1 s 28944 28190 28944 28190 4 vdd
port 513 nsew
rlabel metal1 s 29712 26610 29712 26610 4 vdd
port 513 nsew
rlabel metal1 s 28944 27899 28944 27899 4 vdd
port 513 nsew
rlabel metal1 s 29712 27400 29712 27400 4 vdd
port 513 nsew
rlabel metal1 s 27696 25529 27696 25529 4 vdd
port 513 nsew
rlabel metal1 s 28944 27400 28944 27400 4 vdd
port 513 nsew
rlabel metal1 s 28464 25820 28464 25820 4 vdd
port 513 nsew
rlabel metal1 s 29712 25529 29712 25529 4 vdd
port 513 nsew
rlabel metal1 s 27696 27400 27696 27400 4 vdd
port 513 nsew
rlabel metal1 s 28464 27899 28464 27899 4 vdd
port 513 nsew
rlabel metal1 s 28464 25529 28464 25529 4 vdd
port 513 nsew
rlabel metal1 s 27696 27899 27696 27899 4 vdd
port 513 nsew
rlabel metal1 s 28944 26319 28944 26319 4 vdd
port 513 nsew
rlabel metal1 s 28944 25820 28944 25820 4 vdd
port 513 nsew
rlabel metal1 s 28464 26610 28464 26610 4 vdd
port 513 nsew
rlabel metal1 s 38448 35799 38448 35799 4 vdd
port 513 nsew
rlabel metal1 s 38448 36880 38448 36880 4 vdd
port 513 nsew
rlabel metal1 s 38928 37379 38928 37379 4 vdd
port 513 nsew
rlabel metal1 s 38448 37379 38448 37379 4 vdd
port 513 nsew
rlabel metal1 s 37680 37670 37680 37670 4 vdd
port 513 nsew
rlabel metal1 s 39696 35799 39696 35799 4 vdd
port 513 nsew
rlabel metal1 s 37680 37379 37680 37379 4 vdd
port 513 nsew
rlabel metal1 s 38928 36589 38928 36589 4 vdd
port 513 nsew
rlabel metal1 s 39696 36880 39696 36880 4 vdd
port 513 nsew
rlabel metal1 s 38928 37670 38928 37670 4 vdd
port 513 nsew
rlabel metal1 s 38448 35300 38448 35300 4 vdd
port 513 nsew
rlabel metal1 s 37680 36589 37680 36589 4 vdd
port 513 nsew
rlabel metal1 s 38448 35009 38448 35009 4 vdd
port 513 nsew
rlabel metal1 s 39696 35009 39696 35009 4 vdd
port 513 nsew
rlabel metal1 s 39696 37379 39696 37379 4 vdd
port 513 nsew
rlabel metal1 s 39696 35300 39696 35300 4 vdd
port 513 nsew
rlabel metal1 s 38928 36090 38928 36090 4 vdd
port 513 nsew
rlabel metal1 s 38928 36880 38928 36880 4 vdd
port 513 nsew
rlabel metal1 s 37680 35799 37680 35799 4 vdd
port 513 nsew
rlabel metal1 s 39696 37670 39696 37670 4 vdd
port 513 nsew
rlabel metal1 s 38448 37670 38448 37670 4 vdd
port 513 nsew
rlabel metal1 s 38928 35799 38928 35799 4 vdd
port 513 nsew
rlabel metal1 s 38448 36589 38448 36589 4 vdd
port 513 nsew
rlabel metal1 s 39696 36090 39696 36090 4 vdd
port 513 nsew
rlabel metal1 s 38448 36090 38448 36090 4 vdd
port 513 nsew
rlabel metal1 s 37680 35009 37680 35009 4 vdd
port 513 nsew
rlabel metal1 s 37680 35300 37680 35300 4 vdd
port 513 nsew
rlabel metal1 s 38928 35009 38928 35009 4 vdd
port 513 nsew
rlabel metal1 s 38928 35300 38928 35300 4 vdd
port 513 nsew
rlabel metal1 s 37680 36880 37680 36880 4 vdd
port 513 nsew
rlabel metal1 s 39696 36589 39696 36589 4 vdd
port 513 nsew
rlabel metal1 s 37680 36090 37680 36090 4 vdd
port 513 nsew
rlabel metal1 s 35952 37670 35952 37670 4 vdd
port 513 nsew
rlabel metal1 s 36432 37670 36432 37670 4 vdd
port 513 nsew
rlabel metal1 s 36432 35009 36432 35009 4 vdd
port 513 nsew
rlabel metal1 s 35952 36880 35952 36880 4 vdd
port 513 nsew
rlabel metal1 s 37200 35799 37200 35799 4 vdd
port 513 nsew
rlabel metal1 s 37200 37670 37200 37670 4 vdd
port 513 nsew
rlabel metal1 s 35952 35799 35952 35799 4 vdd
port 513 nsew
rlabel metal1 s 35184 36090 35184 36090 4 vdd
port 513 nsew
rlabel metal1 s 37200 35009 37200 35009 4 vdd
port 513 nsew
rlabel metal1 s 37200 36880 37200 36880 4 vdd
port 513 nsew
rlabel metal1 s 35952 36090 35952 36090 4 vdd
port 513 nsew
rlabel metal1 s 36432 37379 36432 37379 4 vdd
port 513 nsew
rlabel metal1 s 36432 35300 36432 35300 4 vdd
port 513 nsew
rlabel metal1 s 35184 37670 35184 37670 4 vdd
port 513 nsew
rlabel metal1 s 35952 35009 35952 35009 4 vdd
port 513 nsew
rlabel metal1 s 35184 37379 35184 37379 4 vdd
port 513 nsew
rlabel metal1 s 36432 35799 36432 35799 4 vdd
port 513 nsew
rlabel metal1 s 35184 36880 35184 36880 4 vdd
port 513 nsew
rlabel metal1 s 37200 35300 37200 35300 4 vdd
port 513 nsew
rlabel metal1 s 36432 36880 36432 36880 4 vdd
port 513 nsew
rlabel metal1 s 36432 36090 36432 36090 4 vdd
port 513 nsew
rlabel metal1 s 36432 36589 36432 36589 4 vdd
port 513 nsew
rlabel metal1 s 35952 37379 35952 37379 4 vdd
port 513 nsew
rlabel metal1 s 37200 36589 37200 36589 4 vdd
port 513 nsew
rlabel metal1 s 37200 36090 37200 36090 4 vdd
port 513 nsew
rlabel metal1 s 35184 35009 35184 35009 4 vdd
port 513 nsew
rlabel metal1 s 35952 35300 35952 35300 4 vdd
port 513 nsew
rlabel metal1 s 35184 35300 35184 35300 4 vdd
port 513 nsew
rlabel metal1 s 35184 36589 35184 36589 4 vdd
port 513 nsew
rlabel metal1 s 37200 37379 37200 37379 4 vdd
port 513 nsew
rlabel metal1 s 35952 36589 35952 36589 4 vdd
port 513 nsew
rlabel metal1 s 35184 35799 35184 35799 4 vdd
port 513 nsew
rlabel metal1 s 35952 33429 35952 33429 4 vdd
port 513 nsew
rlabel metal1 s 35184 34510 35184 34510 4 vdd
port 513 nsew
rlabel metal1 s 35952 32639 35952 32639 4 vdd
port 513 nsew
rlabel metal1 s 36432 34510 36432 34510 4 vdd
port 513 nsew
rlabel metal1 s 36432 34219 36432 34219 4 vdd
port 513 nsew
rlabel metal1 s 35184 33720 35184 33720 4 vdd
port 513 nsew
rlabel metal1 s 36432 33429 36432 33429 4 vdd
port 513 nsew
rlabel metal1 s 35184 33429 35184 33429 4 vdd
port 513 nsew
rlabel metal1 s 35952 33720 35952 33720 4 vdd
port 513 nsew
rlabel metal1 s 37200 32140 37200 32140 4 vdd
port 513 nsew
rlabel metal1 s 35184 34219 35184 34219 4 vdd
port 513 nsew
rlabel metal1 s 35952 34219 35952 34219 4 vdd
port 513 nsew
rlabel metal1 s 35952 32930 35952 32930 4 vdd
port 513 nsew
rlabel metal1 s 36432 31849 36432 31849 4 vdd
port 513 nsew
rlabel metal1 s 37200 31849 37200 31849 4 vdd
port 513 nsew
rlabel metal1 s 35184 32140 35184 32140 4 vdd
port 513 nsew
rlabel metal1 s 35952 31849 35952 31849 4 vdd
port 513 nsew
rlabel metal1 s 35184 32930 35184 32930 4 vdd
port 513 nsew
rlabel metal1 s 37200 32930 37200 32930 4 vdd
port 513 nsew
rlabel metal1 s 36432 33720 36432 33720 4 vdd
port 513 nsew
rlabel metal1 s 35184 31849 35184 31849 4 vdd
port 513 nsew
rlabel metal1 s 36432 32930 36432 32930 4 vdd
port 513 nsew
rlabel metal1 s 37200 34219 37200 34219 4 vdd
port 513 nsew
rlabel metal1 s 36432 32639 36432 32639 4 vdd
port 513 nsew
rlabel metal1 s 37200 32639 37200 32639 4 vdd
port 513 nsew
rlabel metal1 s 37200 33720 37200 33720 4 vdd
port 513 nsew
rlabel metal1 s 35952 32140 35952 32140 4 vdd
port 513 nsew
rlabel metal1 s 36432 32140 36432 32140 4 vdd
port 513 nsew
rlabel metal1 s 37200 34510 37200 34510 4 vdd
port 513 nsew
rlabel metal1 s 35952 34510 35952 34510 4 vdd
port 513 nsew
rlabel metal1 s 35184 32639 35184 32639 4 vdd
port 513 nsew
rlabel metal1 s 37200 33429 37200 33429 4 vdd
port 513 nsew
rlabel metal1 s 37680 34219 37680 34219 4 vdd
port 513 nsew
rlabel metal1 s 39696 34510 39696 34510 4 vdd
port 513 nsew
rlabel metal1 s 37680 32930 37680 32930 4 vdd
port 513 nsew
rlabel metal1 s 37680 31849 37680 31849 4 vdd
port 513 nsew
rlabel metal1 s 39696 32639 39696 32639 4 vdd
port 513 nsew
rlabel metal1 s 38928 34219 38928 34219 4 vdd
port 513 nsew
rlabel metal1 s 38448 33429 38448 33429 4 vdd
port 513 nsew
rlabel metal1 s 38928 31849 38928 31849 4 vdd
port 513 nsew
rlabel metal1 s 38448 31849 38448 31849 4 vdd
port 513 nsew
rlabel metal1 s 38448 32140 38448 32140 4 vdd
port 513 nsew
rlabel metal1 s 38448 34219 38448 34219 4 vdd
port 513 nsew
rlabel metal1 s 37680 32140 37680 32140 4 vdd
port 513 nsew
rlabel metal1 s 39696 31849 39696 31849 4 vdd
port 513 nsew
rlabel metal1 s 38448 33720 38448 33720 4 vdd
port 513 nsew
rlabel metal1 s 37680 34510 37680 34510 4 vdd
port 513 nsew
rlabel metal1 s 39696 33720 39696 33720 4 vdd
port 513 nsew
rlabel metal1 s 39696 34219 39696 34219 4 vdd
port 513 nsew
rlabel metal1 s 37680 32639 37680 32639 4 vdd
port 513 nsew
rlabel metal1 s 38928 32930 38928 32930 4 vdd
port 513 nsew
rlabel metal1 s 39696 33429 39696 33429 4 vdd
port 513 nsew
rlabel metal1 s 39696 32930 39696 32930 4 vdd
port 513 nsew
rlabel metal1 s 38928 33720 38928 33720 4 vdd
port 513 nsew
rlabel metal1 s 37680 33429 37680 33429 4 vdd
port 513 nsew
rlabel metal1 s 38928 33429 38928 33429 4 vdd
port 513 nsew
rlabel metal1 s 37680 33720 37680 33720 4 vdd
port 513 nsew
rlabel metal1 s 38448 32930 38448 32930 4 vdd
port 513 nsew
rlabel metal1 s 38448 32639 38448 32639 4 vdd
port 513 nsew
rlabel metal1 s 38928 32639 38928 32639 4 vdd
port 513 nsew
rlabel metal1 s 38928 32140 38928 32140 4 vdd
port 513 nsew
rlabel metal1 s 38928 34510 38928 34510 4 vdd
port 513 nsew
rlabel metal1 s 38448 34510 38448 34510 4 vdd
port 513 nsew
rlabel metal1 s 39696 32140 39696 32140 4 vdd
port 513 nsew
rlabel metal1 s 32688 37379 32688 37379 4 vdd
port 513 nsew
rlabel metal1 s 34704 36589 34704 36589 4 vdd
port 513 nsew
rlabel metal1 s 33936 36589 33936 36589 4 vdd
port 513 nsew
rlabel metal1 s 33456 36880 33456 36880 4 vdd
port 513 nsew
rlabel metal1 s 33456 35300 33456 35300 4 vdd
port 513 nsew
rlabel metal1 s 33936 35300 33936 35300 4 vdd
port 513 nsew
rlabel metal1 s 33456 35799 33456 35799 4 vdd
port 513 nsew
rlabel metal1 s 34704 37379 34704 37379 4 vdd
port 513 nsew
rlabel metal1 s 32688 37670 32688 37670 4 vdd
port 513 nsew
rlabel metal1 s 32688 35009 32688 35009 4 vdd
port 513 nsew
rlabel metal1 s 34704 35799 34704 35799 4 vdd
port 513 nsew
rlabel metal1 s 32688 36090 32688 36090 4 vdd
port 513 nsew
rlabel metal1 s 33456 35009 33456 35009 4 vdd
port 513 nsew
rlabel metal1 s 34704 36090 34704 36090 4 vdd
port 513 nsew
rlabel metal1 s 34704 35300 34704 35300 4 vdd
port 513 nsew
rlabel metal1 s 33936 36880 33936 36880 4 vdd
port 513 nsew
rlabel metal1 s 34704 36880 34704 36880 4 vdd
port 513 nsew
rlabel metal1 s 34704 35009 34704 35009 4 vdd
port 513 nsew
rlabel metal1 s 34704 37670 34704 37670 4 vdd
port 513 nsew
rlabel metal1 s 32688 36880 32688 36880 4 vdd
port 513 nsew
rlabel metal1 s 33936 35799 33936 35799 4 vdd
port 513 nsew
rlabel metal1 s 33456 36589 33456 36589 4 vdd
port 513 nsew
rlabel metal1 s 33936 36090 33936 36090 4 vdd
port 513 nsew
rlabel metal1 s 32688 35300 32688 35300 4 vdd
port 513 nsew
rlabel metal1 s 33936 37670 33936 37670 4 vdd
port 513 nsew
rlabel metal1 s 32688 36589 32688 36589 4 vdd
port 513 nsew
rlabel metal1 s 33456 36090 33456 36090 4 vdd
port 513 nsew
rlabel metal1 s 33456 37670 33456 37670 4 vdd
port 513 nsew
rlabel metal1 s 32688 35799 32688 35799 4 vdd
port 513 nsew
rlabel metal1 s 33936 37379 33936 37379 4 vdd
port 513 nsew
rlabel metal1 s 33456 37379 33456 37379 4 vdd
port 513 nsew
rlabel metal1 s 33936 35009 33936 35009 4 vdd
port 513 nsew
rlabel metal1 s 31440 36589 31440 36589 4 vdd
port 513 nsew
rlabel metal1 s 30960 36589 30960 36589 4 vdd
port 513 nsew
rlabel metal1 s 30192 37379 30192 37379 4 vdd
port 513 nsew
rlabel metal1 s 31440 35300 31440 35300 4 vdd
port 513 nsew
rlabel metal1 s 30960 37379 30960 37379 4 vdd
port 513 nsew
rlabel metal1 s 32208 37670 32208 37670 4 vdd
port 513 nsew
rlabel metal1 s 31440 36880 31440 36880 4 vdd
port 513 nsew
rlabel metal1 s 30960 36880 30960 36880 4 vdd
port 513 nsew
rlabel metal1 s 30192 35799 30192 35799 4 vdd
port 513 nsew
rlabel metal1 s 30960 35009 30960 35009 4 vdd
port 513 nsew
rlabel metal1 s 32208 35300 32208 35300 4 vdd
port 513 nsew
rlabel metal1 s 31440 35009 31440 35009 4 vdd
port 513 nsew
rlabel metal1 s 32208 37379 32208 37379 4 vdd
port 513 nsew
rlabel metal1 s 30960 35300 30960 35300 4 vdd
port 513 nsew
rlabel metal1 s 30192 36589 30192 36589 4 vdd
port 513 nsew
rlabel metal1 s 32208 35009 32208 35009 4 vdd
port 513 nsew
rlabel metal1 s 32208 36589 32208 36589 4 vdd
port 513 nsew
rlabel metal1 s 30192 35009 30192 35009 4 vdd
port 513 nsew
rlabel metal1 s 31440 35799 31440 35799 4 vdd
port 513 nsew
rlabel metal1 s 32208 36090 32208 36090 4 vdd
port 513 nsew
rlabel metal1 s 30960 35799 30960 35799 4 vdd
port 513 nsew
rlabel metal1 s 30960 36090 30960 36090 4 vdd
port 513 nsew
rlabel metal1 s 30192 37670 30192 37670 4 vdd
port 513 nsew
rlabel metal1 s 30192 36880 30192 36880 4 vdd
port 513 nsew
rlabel metal1 s 32208 36880 32208 36880 4 vdd
port 513 nsew
rlabel metal1 s 31440 37670 31440 37670 4 vdd
port 513 nsew
rlabel metal1 s 31440 37379 31440 37379 4 vdd
port 513 nsew
rlabel metal1 s 30192 36090 30192 36090 4 vdd
port 513 nsew
rlabel metal1 s 31440 36090 31440 36090 4 vdd
port 513 nsew
rlabel metal1 s 32208 35799 32208 35799 4 vdd
port 513 nsew
rlabel metal1 s 30192 35300 30192 35300 4 vdd
port 513 nsew
rlabel metal1 s 30960 37670 30960 37670 4 vdd
port 513 nsew
rlabel metal1 s 31440 32930 31440 32930 4 vdd
port 513 nsew
rlabel metal1 s 32208 34510 32208 34510 4 vdd
port 513 nsew
rlabel metal1 s 30960 34219 30960 34219 4 vdd
port 513 nsew
rlabel metal1 s 31440 33720 31440 33720 4 vdd
port 513 nsew
rlabel metal1 s 30192 32639 30192 32639 4 vdd
port 513 nsew
rlabel metal1 s 30960 33720 30960 33720 4 vdd
port 513 nsew
rlabel metal1 s 30192 32930 30192 32930 4 vdd
port 513 nsew
rlabel metal1 s 30960 32930 30960 32930 4 vdd
port 513 nsew
rlabel metal1 s 31440 32140 31440 32140 4 vdd
port 513 nsew
rlabel metal1 s 32208 32930 32208 32930 4 vdd
port 513 nsew
rlabel metal1 s 30192 34219 30192 34219 4 vdd
port 513 nsew
rlabel metal1 s 32208 32140 32208 32140 4 vdd
port 513 nsew
rlabel metal1 s 31440 32639 31440 32639 4 vdd
port 513 nsew
rlabel metal1 s 30960 31849 30960 31849 4 vdd
port 513 nsew
rlabel metal1 s 30960 32639 30960 32639 4 vdd
port 513 nsew
rlabel metal1 s 30192 33429 30192 33429 4 vdd
port 513 nsew
rlabel metal1 s 30192 32140 30192 32140 4 vdd
port 513 nsew
rlabel metal1 s 31440 33429 31440 33429 4 vdd
port 513 nsew
rlabel metal1 s 31440 34510 31440 34510 4 vdd
port 513 nsew
rlabel metal1 s 31440 34219 31440 34219 4 vdd
port 513 nsew
rlabel metal1 s 31440 31849 31440 31849 4 vdd
port 513 nsew
rlabel metal1 s 32208 34219 32208 34219 4 vdd
port 513 nsew
rlabel metal1 s 32208 33720 32208 33720 4 vdd
port 513 nsew
rlabel metal1 s 30960 32140 30960 32140 4 vdd
port 513 nsew
rlabel metal1 s 32208 33429 32208 33429 4 vdd
port 513 nsew
rlabel metal1 s 30192 31849 30192 31849 4 vdd
port 513 nsew
rlabel metal1 s 30960 34510 30960 34510 4 vdd
port 513 nsew
rlabel metal1 s 32208 31849 32208 31849 4 vdd
port 513 nsew
rlabel metal1 s 30960 33429 30960 33429 4 vdd
port 513 nsew
rlabel metal1 s 30192 33720 30192 33720 4 vdd
port 513 nsew
rlabel metal1 s 30192 34510 30192 34510 4 vdd
port 513 nsew
rlabel metal1 s 32208 32639 32208 32639 4 vdd
port 513 nsew
rlabel metal1 s 33456 34510 33456 34510 4 vdd
port 513 nsew
rlabel metal1 s 33456 32930 33456 32930 4 vdd
port 513 nsew
rlabel metal1 s 34704 32639 34704 32639 4 vdd
port 513 nsew
rlabel metal1 s 33936 33720 33936 33720 4 vdd
port 513 nsew
rlabel metal1 s 32688 34219 32688 34219 4 vdd
port 513 nsew
rlabel metal1 s 33936 32930 33936 32930 4 vdd
port 513 nsew
rlabel metal1 s 34704 34510 34704 34510 4 vdd
port 513 nsew
rlabel metal1 s 33936 34510 33936 34510 4 vdd
port 513 nsew
rlabel metal1 s 32688 32140 32688 32140 4 vdd
port 513 nsew
rlabel metal1 s 33456 31849 33456 31849 4 vdd
port 513 nsew
rlabel metal1 s 34704 33720 34704 33720 4 vdd
port 513 nsew
rlabel metal1 s 34704 33429 34704 33429 4 vdd
port 513 nsew
rlabel metal1 s 33456 34219 33456 34219 4 vdd
port 513 nsew
rlabel metal1 s 34704 31849 34704 31849 4 vdd
port 513 nsew
rlabel metal1 s 32688 32930 32688 32930 4 vdd
port 513 nsew
rlabel metal1 s 32688 34510 32688 34510 4 vdd
port 513 nsew
rlabel metal1 s 33936 31849 33936 31849 4 vdd
port 513 nsew
rlabel metal1 s 32688 33720 32688 33720 4 vdd
port 513 nsew
rlabel metal1 s 33456 32639 33456 32639 4 vdd
port 513 nsew
rlabel metal1 s 32688 31849 32688 31849 4 vdd
port 513 nsew
rlabel metal1 s 33456 32140 33456 32140 4 vdd
port 513 nsew
rlabel metal1 s 33456 33720 33456 33720 4 vdd
port 513 nsew
rlabel metal1 s 33936 33429 33936 33429 4 vdd
port 513 nsew
rlabel metal1 s 34704 34219 34704 34219 4 vdd
port 513 nsew
rlabel metal1 s 34704 32140 34704 32140 4 vdd
port 513 nsew
rlabel metal1 s 32688 32639 32688 32639 4 vdd
port 513 nsew
rlabel metal1 s 33936 32140 33936 32140 4 vdd
port 513 nsew
rlabel metal1 s 33456 33429 33456 33429 4 vdd
port 513 nsew
rlabel metal1 s 32688 33429 32688 33429 4 vdd
port 513 nsew
rlabel metal1 s 34704 32930 34704 32930 4 vdd
port 513 nsew
rlabel metal1 s 33936 32639 33936 32639 4 vdd
port 513 nsew
rlabel metal1 s 33936 34219 33936 34219 4 vdd
port 513 nsew
rlabel metal1 s 32688 29770 32688 29770 4 vdd
port 513 nsew
rlabel metal1 s 33456 28980 33456 28980 4 vdd
port 513 nsew
rlabel metal1 s 33936 28980 33936 28980 4 vdd
port 513 nsew
rlabel metal1 s 33456 30269 33456 30269 4 vdd
port 513 nsew
rlabel metal1 s 33936 31059 33936 31059 4 vdd
port 513 nsew
rlabel metal1 s 33456 30560 33456 30560 4 vdd
port 513 nsew
rlabel metal1 s 34704 29479 34704 29479 4 vdd
port 513 nsew
rlabel metal1 s 34704 30560 34704 30560 4 vdd
port 513 nsew
rlabel metal1 s 34704 30269 34704 30269 4 vdd
port 513 nsew
rlabel metal1 s 34704 31059 34704 31059 4 vdd
port 513 nsew
rlabel metal1 s 33936 29770 33936 29770 4 vdd
port 513 nsew
rlabel metal1 s 33456 31350 33456 31350 4 vdd
port 513 nsew
rlabel metal1 s 32688 30269 32688 30269 4 vdd
port 513 nsew
rlabel metal1 s 33936 30560 33936 30560 4 vdd
port 513 nsew
rlabel metal1 s 34704 28689 34704 28689 4 vdd
port 513 nsew
rlabel metal1 s 32688 31059 32688 31059 4 vdd
port 513 nsew
rlabel metal1 s 33936 31350 33936 31350 4 vdd
port 513 nsew
rlabel metal1 s 32688 29479 32688 29479 4 vdd
port 513 nsew
rlabel metal1 s 32688 30560 32688 30560 4 vdd
port 513 nsew
rlabel metal1 s 33456 28689 33456 28689 4 vdd
port 513 nsew
rlabel metal1 s 33936 30269 33936 30269 4 vdd
port 513 nsew
rlabel metal1 s 33936 28689 33936 28689 4 vdd
port 513 nsew
rlabel metal1 s 32688 28980 32688 28980 4 vdd
port 513 nsew
rlabel metal1 s 32688 31350 32688 31350 4 vdd
port 513 nsew
rlabel metal1 s 33936 29479 33936 29479 4 vdd
port 513 nsew
rlabel metal1 s 33456 29479 33456 29479 4 vdd
port 513 nsew
rlabel metal1 s 34704 28980 34704 28980 4 vdd
port 513 nsew
rlabel metal1 s 32688 28689 32688 28689 4 vdd
port 513 nsew
rlabel metal1 s 33456 29770 33456 29770 4 vdd
port 513 nsew
rlabel metal1 s 33456 31059 33456 31059 4 vdd
port 513 nsew
rlabel metal1 s 34704 29770 34704 29770 4 vdd
port 513 nsew
rlabel metal1 s 34704 31350 34704 31350 4 vdd
port 513 nsew
rlabel metal1 s 32208 31350 32208 31350 4 vdd
port 513 nsew
rlabel metal1 s 30192 30269 30192 30269 4 vdd
port 513 nsew
rlabel metal1 s 32208 29770 32208 29770 4 vdd
port 513 nsew
rlabel metal1 s 30960 30560 30960 30560 4 vdd
port 513 nsew
rlabel metal1 s 32208 30269 32208 30269 4 vdd
port 513 nsew
rlabel metal1 s 32208 29479 32208 29479 4 vdd
port 513 nsew
rlabel metal1 s 31440 29770 31440 29770 4 vdd
port 513 nsew
rlabel metal1 s 30192 28689 30192 28689 4 vdd
port 513 nsew
rlabel metal1 s 31440 30560 31440 30560 4 vdd
port 513 nsew
rlabel metal1 s 31440 29479 31440 29479 4 vdd
port 513 nsew
rlabel metal1 s 30192 31059 30192 31059 4 vdd
port 513 nsew
rlabel metal1 s 32208 28980 32208 28980 4 vdd
port 513 nsew
rlabel metal1 s 30960 30269 30960 30269 4 vdd
port 513 nsew
rlabel metal1 s 30960 29479 30960 29479 4 vdd
port 513 nsew
rlabel metal1 s 31440 28980 31440 28980 4 vdd
port 513 nsew
rlabel metal1 s 31440 31059 31440 31059 4 vdd
port 513 nsew
rlabel metal1 s 31440 31350 31440 31350 4 vdd
port 513 nsew
rlabel metal1 s 30192 31350 30192 31350 4 vdd
port 513 nsew
rlabel metal1 s 30960 28689 30960 28689 4 vdd
port 513 nsew
rlabel metal1 s 30192 30560 30192 30560 4 vdd
port 513 nsew
rlabel metal1 s 32208 30560 32208 30560 4 vdd
port 513 nsew
rlabel metal1 s 30960 29770 30960 29770 4 vdd
port 513 nsew
rlabel metal1 s 31440 30269 31440 30269 4 vdd
port 513 nsew
rlabel metal1 s 30960 28980 30960 28980 4 vdd
port 513 nsew
rlabel metal1 s 30192 29479 30192 29479 4 vdd
port 513 nsew
rlabel metal1 s 32208 31059 32208 31059 4 vdd
port 513 nsew
rlabel metal1 s 32208 28689 32208 28689 4 vdd
port 513 nsew
rlabel metal1 s 30192 28980 30192 28980 4 vdd
port 513 nsew
rlabel metal1 s 31440 28689 31440 28689 4 vdd
port 513 nsew
rlabel metal1 s 30192 29770 30192 29770 4 vdd
port 513 nsew
rlabel metal1 s 30960 31059 30960 31059 4 vdd
port 513 nsew
rlabel metal1 s 30960 31350 30960 31350 4 vdd
port 513 nsew
rlabel metal1 s 30192 27109 30192 27109 4 vdd
port 513 nsew
rlabel metal1 s 30960 27400 30960 27400 4 vdd
port 513 nsew
rlabel metal1 s 30960 26319 30960 26319 4 vdd
port 513 nsew
rlabel metal1 s 30192 26319 30192 26319 4 vdd
port 513 nsew
rlabel metal1 s 31440 27400 31440 27400 4 vdd
port 513 nsew
rlabel metal1 s 31440 26610 31440 26610 4 vdd
port 513 nsew
rlabel metal1 s 30960 27899 30960 27899 4 vdd
port 513 nsew
rlabel metal1 s 30960 26610 30960 26610 4 vdd
port 513 nsew
rlabel metal1 s 30192 28190 30192 28190 4 vdd
port 513 nsew
rlabel metal1 s 32208 25820 32208 25820 4 vdd
port 513 nsew
rlabel metal1 s 30192 26610 30192 26610 4 vdd
port 513 nsew
rlabel metal1 s 31440 27899 31440 27899 4 vdd
port 513 nsew
rlabel metal1 s 30960 28190 30960 28190 4 vdd
port 513 nsew
rlabel metal1 s 30960 25820 30960 25820 4 vdd
port 513 nsew
rlabel metal1 s 30192 25820 30192 25820 4 vdd
port 513 nsew
rlabel metal1 s 32208 27109 32208 27109 4 vdd
port 513 nsew
rlabel metal1 s 31440 26319 31440 26319 4 vdd
port 513 nsew
rlabel metal1 s 31440 25820 31440 25820 4 vdd
port 513 nsew
rlabel metal1 s 30192 25529 30192 25529 4 vdd
port 513 nsew
rlabel metal1 s 31440 27109 31440 27109 4 vdd
port 513 nsew
rlabel metal1 s 30192 27899 30192 27899 4 vdd
port 513 nsew
rlabel metal1 s 30192 27400 30192 27400 4 vdd
port 513 nsew
rlabel metal1 s 31440 28190 31440 28190 4 vdd
port 513 nsew
rlabel metal1 s 31440 25529 31440 25529 4 vdd
port 513 nsew
rlabel metal1 s 32208 26319 32208 26319 4 vdd
port 513 nsew
rlabel metal1 s 32208 27400 32208 27400 4 vdd
port 513 nsew
rlabel metal1 s 30960 27109 30960 27109 4 vdd
port 513 nsew
rlabel metal1 s 30960 25529 30960 25529 4 vdd
port 513 nsew
rlabel metal1 s 32208 25529 32208 25529 4 vdd
port 513 nsew
rlabel metal1 s 32208 26610 32208 26610 4 vdd
port 513 nsew
rlabel metal1 s 32208 27899 32208 27899 4 vdd
port 513 nsew
rlabel metal1 s 32208 28190 32208 28190 4 vdd
port 513 nsew
rlabel metal1 s 34704 27109 34704 27109 4 vdd
port 513 nsew
rlabel metal1 s 33456 26319 33456 26319 4 vdd
port 513 nsew
rlabel metal1 s 33456 27899 33456 27899 4 vdd
port 513 nsew
rlabel metal1 s 34704 27400 34704 27400 4 vdd
port 513 nsew
rlabel metal1 s 33936 28190 33936 28190 4 vdd
port 513 nsew
rlabel metal1 s 33456 26610 33456 26610 4 vdd
port 513 nsew
rlabel metal1 s 33936 25529 33936 25529 4 vdd
port 513 nsew
rlabel metal1 s 32688 27899 32688 27899 4 vdd
port 513 nsew
rlabel metal1 s 33936 26610 33936 26610 4 vdd
port 513 nsew
rlabel metal1 s 33456 27400 33456 27400 4 vdd
port 513 nsew
rlabel metal1 s 33936 26319 33936 26319 4 vdd
port 513 nsew
rlabel metal1 s 33456 25820 33456 25820 4 vdd
port 513 nsew
rlabel metal1 s 33936 27400 33936 27400 4 vdd
port 513 nsew
rlabel metal1 s 33456 27109 33456 27109 4 vdd
port 513 nsew
rlabel metal1 s 33456 25529 33456 25529 4 vdd
port 513 nsew
rlabel metal1 s 32688 27109 32688 27109 4 vdd
port 513 nsew
rlabel metal1 s 34704 28190 34704 28190 4 vdd
port 513 nsew
rlabel metal1 s 33936 25820 33936 25820 4 vdd
port 513 nsew
rlabel metal1 s 34704 26319 34704 26319 4 vdd
port 513 nsew
rlabel metal1 s 34704 25820 34704 25820 4 vdd
port 513 nsew
rlabel metal1 s 34704 27899 34704 27899 4 vdd
port 513 nsew
rlabel metal1 s 33936 27899 33936 27899 4 vdd
port 513 nsew
rlabel metal1 s 32688 27400 32688 27400 4 vdd
port 513 nsew
rlabel metal1 s 32688 28190 32688 28190 4 vdd
port 513 nsew
rlabel metal1 s 33936 27109 33936 27109 4 vdd
port 513 nsew
rlabel metal1 s 32688 25529 32688 25529 4 vdd
port 513 nsew
rlabel metal1 s 32688 26610 32688 26610 4 vdd
port 513 nsew
rlabel metal1 s 32688 25820 32688 25820 4 vdd
port 513 nsew
rlabel metal1 s 33456 28190 33456 28190 4 vdd
port 513 nsew
rlabel metal1 s 32688 26319 32688 26319 4 vdd
port 513 nsew
rlabel metal1 s 34704 25529 34704 25529 4 vdd
port 513 nsew
rlabel metal1 s 34704 26610 34704 26610 4 vdd
port 513 nsew
rlabel metal1 s 39696 28980 39696 28980 4 vdd
port 513 nsew
rlabel metal1 s 38928 30560 38928 30560 4 vdd
port 513 nsew
rlabel metal1 s 38928 28980 38928 28980 4 vdd
port 513 nsew
rlabel metal1 s 37680 28689 37680 28689 4 vdd
port 513 nsew
rlabel metal1 s 38928 29770 38928 29770 4 vdd
port 513 nsew
rlabel metal1 s 38448 30269 38448 30269 4 vdd
port 513 nsew
rlabel metal1 s 37680 30269 37680 30269 4 vdd
port 513 nsew
rlabel metal1 s 39696 30269 39696 30269 4 vdd
port 513 nsew
rlabel metal1 s 39696 28689 39696 28689 4 vdd
port 513 nsew
rlabel metal1 s 37680 31059 37680 31059 4 vdd
port 513 nsew
rlabel metal1 s 38928 30269 38928 30269 4 vdd
port 513 nsew
rlabel metal1 s 38448 30560 38448 30560 4 vdd
port 513 nsew
rlabel metal1 s 39696 29770 39696 29770 4 vdd
port 513 nsew
rlabel metal1 s 38928 31350 38928 31350 4 vdd
port 513 nsew
rlabel metal1 s 39696 29479 39696 29479 4 vdd
port 513 nsew
rlabel metal1 s 38448 28980 38448 28980 4 vdd
port 513 nsew
rlabel metal1 s 38928 29479 38928 29479 4 vdd
port 513 nsew
rlabel metal1 s 38928 31059 38928 31059 4 vdd
port 513 nsew
rlabel metal1 s 38928 28689 38928 28689 4 vdd
port 513 nsew
rlabel metal1 s 39696 31350 39696 31350 4 vdd
port 513 nsew
rlabel metal1 s 39696 30560 39696 30560 4 vdd
port 513 nsew
rlabel metal1 s 38448 29770 38448 29770 4 vdd
port 513 nsew
rlabel metal1 s 38448 29479 38448 29479 4 vdd
port 513 nsew
rlabel metal1 s 38448 31350 38448 31350 4 vdd
port 513 nsew
rlabel metal1 s 37680 29770 37680 29770 4 vdd
port 513 nsew
rlabel metal1 s 37680 29479 37680 29479 4 vdd
port 513 nsew
rlabel metal1 s 38448 28689 38448 28689 4 vdd
port 513 nsew
rlabel metal1 s 38448 31059 38448 31059 4 vdd
port 513 nsew
rlabel metal1 s 37680 30560 37680 30560 4 vdd
port 513 nsew
rlabel metal1 s 39696 31059 39696 31059 4 vdd
port 513 nsew
rlabel metal1 s 37680 28980 37680 28980 4 vdd
port 513 nsew
rlabel metal1 s 37680 31350 37680 31350 4 vdd
port 513 nsew
rlabel metal1 s 36432 29479 36432 29479 4 vdd
port 513 nsew
rlabel metal1 s 37200 28689 37200 28689 4 vdd
port 513 nsew
rlabel metal1 s 36432 28980 36432 28980 4 vdd
port 513 nsew
rlabel metal1 s 35184 29770 35184 29770 4 vdd
port 513 nsew
rlabel metal1 s 35952 29770 35952 29770 4 vdd
port 513 nsew
rlabel metal1 s 35184 28689 35184 28689 4 vdd
port 513 nsew
rlabel metal1 s 37200 31059 37200 31059 4 vdd
port 513 nsew
rlabel metal1 s 36432 30269 36432 30269 4 vdd
port 513 nsew
rlabel metal1 s 35952 31350 35952 31350 4 vdd
port 513 nsew
rlabel metal1 s 37200 29770 37200 29770 4 vdd
port 513 nsew
rlabel metal1 s 35952 31059 35952 31059 4 vdd
port 513 nsew
rlabel metal1 s 35184 28980 35184 28980 4 vdd
port 513 nsew
rlabel metal1 s 35952 30269 35952 30269 4 vdd
port 513 nsew
rlabel metal1 s 35184 31350 35184 31350 4 vdd
port 513 nsew
rlabel metal1 s 36432 31350 36432 31350 4 vdd
port 513 nsew
rlabel metal1 s 36432 28689 36432 28689 4 vdd
port 513 nsew
rlabel metal1 s 35952 29479 35952 29479 4 vdd
port 513 nsew
rlabel metal1 s 36432 29770 36432 29770 4 vdd
port 513 nsew
rlabel metal1 s 36432 31059 36432 31059 4 vdd
port 513 nsew
rlabel metal1 s 36432 30560 36432 30560 4 vdd
port 513 nsew
rlabel metal1 s 35952 30560 35952 30560 4 vdd
port 513 nsew
rlabel metal1 s 35184 30269 35184 30269 4 vdd
port 513 nsew
rlabel metal1 s 35952 28980 35952 28980 4 vdd
port 513 nsew
rlabel metal1 s 37200 29479 37200 29479 4 vdd
port 513 nsew
rlabel metal1 s 37200 31350 37200 31350 4 vdd
port 513 nsew
rlabel metal1 s 35184 29479 35184 29479 4 vdd
port 513 nsew
rlabel metal1 s 37200 30560 37200 30560 4 vdd
port 513 nsew
rlabel metal1 s 35184 31059 35184 31059 4 vdd
port 513 nsew
rlabel metal1 s 35184 30560 35184 30560 4 vdd
port 513 nsew
rlabel metal1 s 37200 28980 37200 28980 4 vdd
port 513 nsew
rlabel metal1 s 37200 30269 37200 30269 4 vdd
port 513 nsew
rlabel metal1 s 35952 28689 35952 28689 4 vdd
port 513 nsew
rlabel metal1 s 37200 26610 37200 26610 4 vdd
port 513 nsew
rlabel metal1 s 37200 25529 37200 25529 4 vdd
port 513 nsew
rlabel metal1 s 37200 26319 37200 26319 4 vdd
port 513 nsew
rlabel metal1 s 35952 27899 35952 27899 4 vdd
port 513 nsew
rlabel metal1 s 35184 27400 35184 27400 4 vdd
port 513 nsew
rlabel metal1 s 37200 27109 37200 27109 4 vdd
port 513 nsew
rlabel metal1 s 36432 27899 36432 27899 4 vdd
port 513 nsew
rlabel metal1 s 37200 28190 37200 28190 4 vdd
port 513 nsew
rlabel metal1 s 37200 25820 37200 25820 4 vdd
port 513 nsew
rlabel metal1 s 36432 27400 36432 27400 4 vdd
port 513 nsew
rlabel metal1 s 35952 28190 35952 28190 4 vdd
port 513 nsew
rlabel metal1 s 35184 25820 35184 25820 4 vdd
port 513 nsew
rlabel metal1 s 35952 25529 35952 25529 4 vdd
port 513 nsew
rlabel metal1 s 36432 25529 36432 25529 4 vdd
port 513 nsew
rlabel metal1 s 36432 27109 36432 27109 4 vdd
port 513 nsew
rlabel metal1 s 35184 27109 35184 27109 4 vdd
port 513 nsew
rlabel metal1 s 35952 25820 35952 25820 4 vdd
port 513 nsew
rlabel metal1 s 37200 27400 37200 27400 4 vdd
port 513 nsew
rlabel metal1 s 35184 26610 35184 26610 4 vdd
port 513 nsew
rlabel metal1 s 35952 27400 35952 27400 4 vdd
port 513 nsew
rlabel metal1 s 35952 26319 35952 26319 4 vdd
port 513 nsew
rlabel metal1 s 36432 26610 36432 26610 4 vdd
port 513 nsew
rlabel metal1 s 37200 27899 37200 27899 4 vdd
port 513 nsew
rlabel metal1 s 35952 26610 35952 26610 4 vdd
port 513 nsew
rlabel metal1 s 36432 28190 36432 28190 4 vdd
port 513 nsew
rlabel metal1 s 36432 25820 36432 25820 4 vdd
port 513 nsew
rlabel metal1 s 35184 26319 35184 26319 4 vdd
port 513 nsew
rlabel metal1 s 36432 26319 36432 26319 4 vdd
port 513 nsew
rlabel metal1 s 35184 28190 35184 28190 4 vdd
port 513 nsew
rlabel metal1 s 35184 25529 35184 25529 4 vdd
port 513 nsew
rlabel metal1 s 35952 27109 35952 27109 4 vdd
port 513 nsew
rlabel metal1 s 35184 27899 35184 27899 4 vdd
port 513 nsew
rlabel metal1 s 37680 27109 37680 27109 4 vdd
port 513 nsew
rlabel metal1 s 39696 28190 39696 28190 4 vdd
port 513 nsew
rlabel metal1 s 37680 25820 37680 25820 4 vdd
port 513 nsew
rlabel metal1 s 38448 27899 38448 27899 4 vdd
port 513 nsew
rlabel metal1 s 38928 27400 38928 27400 4 vdd
port 513 nsew
rlabel metal1 s 37680 27899 37680 27899 4 vdd
port 513 nsew
rlabel metal1 s 39696 27899 39696 27899 4 vdd
port 513 nsew
rlabel metal1 s 39696 27400 39696 27400 4 vdd
port 513 nsew
rlabel metal1 s 39696 25820 39696 25820 4 vdd
port 513 nsew
rlabel metal1 s 37680 28190 37680 28190 4 vdd
port 513 nsew
rlabel metal1 s 38928 27109 38928 27109 4 vdd
port 513 nsew
rlabel metal1 s 37680 25529 37680 25529 4 vdd
port 513 nsew
rlabel metal1 s 38448 28190 38448 28190 4 vdd
port 513 nsew
rlabel metal1 s 38928 25529 38928 25529 4 vdd
port 513 nsew
rlabel metal1 s 38448 25820 38448 25820 4 vdd
port 513 nsew
rlabel metal1 s 39696 27109 39696 27109 4 vdd
port 513 nsew
rlabel metal1 s 38448 25529 38448 25529 4 vdd
port 513 nsew
rlabel metal1 s 39696 25529 39696 25529 4 vdd
port 513 nsew
rlabel metal1 s 38448 27109 38448 27109 4 vdd
port 513 nsew
rlabel metal1 s 38928 26319 38928 26319 4 vdd
port 513 nsew
rlabel metal1 s 37680 27400 37680 27400 4 vdd
port 513 nsew
rlabel metal1 s 37680 26319 37680 26319 4 vdd
port 513 nsew
rlabel metal1 s 38928 27899 38928 27899 4 vdd
port 513 nsew
rlabel metal1 s 38448 27400 38448 27400 4 vdd
port 513 nsew
rlabel metal1 s 39696 26610 39696 26610 4 vdd
port 513 nsew
rlabel metal1 s 38928 28190 38928 28190 4 vdd
port 513 nsew
rlabel metal1 s 38448 26319 38448 26319 4 vdd
port 513 nsew
rlabel metal1 s 39696 26319 39696 26319 4 vdd
port 513 nsew
rlabel metal1 s 38928 25820 38928 25820 4 vdd
port 513 nsew
rlabel metal1 s 38448 26610 38448 26610 4 vdd
port 513 nsew
rlabel metal1 s 37680 26610 37680 26610 4 vdd
port 513 nsew
rlabel metal1 s 38928 26610 38928 26610 4 vdd
port 513 nsew
rlabel metal1 s 18480 48730 18480 48730 4 vdd
port 513 nsew
rlabel metal1 s 19728 50019 19728 50019 4 vdd
port 513 nsew
rlabel metal1 s 18960 47649 18960 47649 4 vdd
port 513 nsew
rlabel metal1 s 17712 47649 17712 47649 4 vdd
port 513 nsew
rlabel metal1 s 18960 49520 18960 49520 4 vdd
port 513 nsew
rlabel metal1 s 17712 49229 17712 49229 4 vdd
port 513 nsew
rlabel metal1 s 17712 47940 17712 47940 4 vdd
port 513 nsew
rlabel metal1 s 18480 49520 18480 49520 4 vdd
port 513 nsew
rlabel metal1 s 18480 50019 18480 50019 4 vdd
port 513 nsew
rlabel metal1 s 19728 48730 19728 48730 4 vdd
port 513 nsew
rlabel metal1 s 17712 48439 17712 48439 4 vdd
port 513 nsew
rlabel metal1 s 18960 47940 18960 47940 4 vdd
port 513 nsew
rlabel metal1 s 19728 50310 19728 50310 4 vdd
port 513 nsew
rlabel metal1 s 17712 50310 17712 50310 4 vdd
port 513 nsew
rlabel metal1 s 19728 47649 19728 47649 4 vdd
port 513 nsew
rlabel metal1 s 17712 48730 17712 48730 4 vdd
port 513 nsew
rlabel metal1 s 18480 49229 18480 49229 4 vdd
port 513 nsew
rlabel metal1 s 18480 50310 18480 50310 4 vdd
port 513 nsew
rlabel metal1 s 19728 49229 19728 49229 4 vdd
port 513 nsew
rlabel metal1 s 18480 47940 18480 47940 4 vdd
port 513 nsew
rlabel metal1 s 18960 50019 18960 50019 4 vdd
port 513 nsew
rlabel metal1 s 18960 50310 18960 50310 4 vdd
port 513 nsew
rlabel metal1 s 19728 49520 19728 49520 4 vdd
port 513 nsew
rlabel metal1 s 18960 48439 18960 48439 4 vdd
port 513 nsew
rlabel metal1 s 18960 49229 18960 49229 4 vdd
port 513 nsew
rlabel metal1 s 19728 47940 19728 47940 4 vdd
port 513 nsew
rlabel metal1 s 18480 48439 18480 48439 4 vdd
port 513 nsew
rlabel metal1 s 17712 49520 17712 49520 4 vdd
port 513 nsew
rlabel metal1 s 18480 47649 18480 47649 4 vdd
port 513 nsew
rlabel metal1 s 19728 48439 19728 48439 4 vdd
port 513 nsew
rlabel metal1 s 18960 48730 18960 48730 4 vdd
port 513 nsew
rlabel metal1 s 17712 50019 17712 50019 4 vdd
port 513 nsew
rlabel metal1 s 17232 48439 17232 48439 4 vdd
port 513 nsew
rlabel metal1 s 15984 50310 15984 50310 4 vdd
port 513 nsew
rlabel metal1 s 15216 50019 15216 50019 4 vdd
port 513 nsew
rlabel metal1 s 17232 49520 17232 49520 4 vdd
port 513 nsew
rlabel metal1 s 15984 48439 15984 48439 4 vdd
port 513 nsew
rlabel metal1 s 15216 48439 15216 48439 4 vdd
port 513 nsew
rlabel metal1 s 15216 49229 15216 49229 4 vdd
port 513 nsew
rlabel metal1 s 16464 50310 16464 50310 4 vdd
port 513 nsew
rlabel metal1 s 15984 49229 15984 49229 4 vdd
port 513 nsew
rlabel metal1 s 15216 49520 15216 49520 4 vdd
port 513 nsew
rlabel metal1 s 16464 49520 16464 49520 4 vdd
port 513 nsew
rlabel metal1 s 15216 47940 15216 47940 4 vdd
port 513 nsew
rlabel metal1 s 15984 50019 15984 50019 4 vdd
port 513 nsew
rlabel metal1 s 16464 47940 16464 47940 4 vdd
port 513 nsew
rlabel metal1 s 17232 50310 17232 50310 4 vdd
port 513 nsew
rlabel metal1 s 15984 48730 15984 48730 4 vdd
port 513 nsew
rlabel metal1 s 16464 48730 16464 48730 4 vdd
port 513 nsew
rlabel metal1 s 17232 48730 17232 48730 4 vdd
port 513 nsew
rlabel metal1 s 15216 48730 15216 48730 4 vdd
port 513 nsew
rlabel metal1 s 17232 50019 17232 50019 4 vdd
port 513 nsew
rlabel metal1 s 16464 49229 16464 49229 4 vdd
port 513 nsew
rlabel metal1 s 15984 49520 15984 49520 4 vdd
port 513 nsew
rlabel metal1 s 15216 47649 15216 47649 4 vdd
port 513 nsew
rlabel metal1 s 16464 47649 16464 47649 4 vdd
port 513 nsew
rlabel metal1 s 17232 47649 17232 47649 4 vdd
port 513 nsew
rlabel metal1 s 15984 47649 15984 47649 4 vdd
port 513 nsew
rlabel metal1 s 17232 49229 17232 49229 4 vdd
port 513 nsew
rlabel metal1 s 16464 48439 16464 48439 4 vdd
port 513 nsew
rlabel metal1 s 15984 47940 15984 47940 4 vdd
port 513 nsew
rlabel metal1 s 17232 47940 17232 47940 4 vdd
port 513 nsew
rlabel metal1 s 16464 50019 16464 50019 4 vdd
port 513 nsew
rlabel metal1 s 15216 50310 15216 50310 4 vdd
port 513 nsew
rlabel metal1 s 16464 44489 16464 44489 4 vdd
port 513 nsew
rlabel metal1 s 15984 45279 15984 45279 4 vdd
port 513 nsew
rlabel metal1 s 15216 45570 15216 45570 4 vdd
port 513 nsew
rlabel metal1 s 17232 46360 17232 46360 4 vdd
port 513 nsew
rlabel metal1 s 17232 47150 17232 47150 4 vdd
port 513 nsew
rlabel metal1 s 15216 47150 15216 47150 4 vdd
port 513 nsew
rlabel metal1 s 17232 44780 17232 44780 4 vdd
port 513 nsew
rlabel metal1 s 15216 46069 15216 46069 4 vdd
port 513 nsew
rlabel metal1 s 16464 44780 16464 44780 4 vdd
port 513 nsew
rlabel metal1 s 15984 45570 15984 45570 4 vdd
port 513 nsew
rlabel metal1 s 16464 45279 16464 45279 4 vdd
port 513 nsew
rlabel metal1 s 15984 44780 15984 44780 4 vdd
port 513 nsew
rlabel metal1 s 15216 44780 15216 44780 4 vdd
port 513 nsew
rlabel metal1 s 15216 44489 15216 44489 4 vdd
port 513 nsew
rlabel metal1 s 15984 47150 15984 47150 4 vdd
port 513 nsew
rlabel metal1 s 17232 45570 17232 45570 4 vdd
port 513 nsew
rlabel metal1 s 17232 45279 17232 45279 4 vdd
port 513 nsew
rlabel metal1 s 16464 46360 16464 46360 4 vdd
port 513 nsew
rlabel metal1 s 15216 45279 15216 45279 4 vdd
port 513 nsew
rlabel metal1 s 16464 46069 16464 46069 4 vdd
port 513 nsew
rlabel metal1 s 17232 46069 17232 46069 4 vdd
port 513 nsew
rlabel metal1 s 17232 46859 17232 46859 4 vdd
port 513 nsew
rlabel metal1 s 15216 46360 15216 46360 4 vdd
port 513 nsew
rlabel metal1 s 15216 46859 15216 46859 4 vdd
port 513 nsew
rlabel metal1 s 17232 44489 17232 44489 4 vdd
port 513 nsew
rlabel metal1 s 16464 45570 16464 45570 4 vdd
port 513 nsew
rlabel metal1 s 15984 46859 15984 46859 4 vdd
port 513 nsew
rlabel metal1 s 15984 46360 15984 46360 4 vdd
port 513 nsew
rlabel metal1 s 16464 46859 16464 46859 4 vdd
port 513 nsew
rlabel metal1 s 16464 47150 16464 47150 4 vdd
port 513 nsew
rlabel metal1 s 15984 46069 15984 46069 4 vdd
port 513 nsew
rlabel metal1 s 15984 44489 15984 44489 4 vdd
port 513 nsew
rlabel metal1 s 17712 45570 17712 45570 4 vdd
port 513 nsew
rlabel metal1 s 19728 45570 19728 45570 4 vdd
port 513 nsew
rlabel metal1 s 19728 44780 19728 44780 4 vdd
port 513 nsew
rlabel metal1 s 18480 45570 18480 45570 4 vdd
port 513 nsew
rlabel metal1 s 18960 46069 18960 46069 4 vdd
port 513 nsew
rlabel metal1 s 18480 45279 18480 45279 4 vdd
port 513 nsew
rlabel metal1 s 19728 46360 19728 46360 4 vdd
port 513 nsew
rlabel metal1 s 17712 47150 17712 47150 4 vdd
port 513 nsew
rlabel metal1 s 18960 46360 18960 46360 4 vdd
port 513 nsew
rlabel metal1 s 17712 46859 17712 46859 4 vdd
port 513 nsew
rlabel metal1 s 17712 45279 17712 45279 4 vdd
port 513 nsew
rlabel metal1 s 19728 46859 19728 46859 4 vdd
port 513 nsew
rlabel metal1 s 18960 45570 18960 45570 4 vdd
port 513 nsew
rlabel metal1 s 18960 47150 18960 47150 4 vdd
port 513 nsew
rlabel metal1 s 18480 46069 18480 46069 4 vdd
port 513 nsew
rlabel metal1 s 17712 44489 17712 44489 4 vdd
port 513 nsew
rlabel metal1 s 18960 44489 18960 44489 4 vdd
port 513 nsew
rlabel metal1 s 18960 44780 18960 44780 4 vdd
port 513 nsew
rlabel metal1 s 19728 44489 19728 44489 4 vdd
port 513 nsew
rlabel metal1 s 18960 45279 18960 45279 4 vdd
port 513 nsew
rlabel metal1 s 18480 44489 18480 44489 4 vdd
port 513 nsew
rlabel metal1 s 17712 46360 17712 46360 4 vdd
port 513 nsew
rlabel metal1 s 18480 47150 18480 47150 4 vdd
port 513 nsew
rlabel metal1 s 17712 46069 17712 46069 4 vdd
port 513 nsew
rlabel metal1 s 19728 47150 19728 47150 4 vdd
port 513 nsew
rlabel metal1 s 18960 46859 18960 46859 4 vdd
port 513 nsew
rlabel metal1 s 19728 45279 19728 45279 4 vdd
port 513 nsew
rlabel metal1 s 18480 46360 18480 46360 4 vdd
port 513 nsew
rlabel metal1 s 18480 46859 18480 46859 4 vdd
port 513 nsew
rlabel metal1 s 18480 44780 18480 44780 4 vdd
port 513 nsew
rlabel metal1 s 17712 44780 17712 44780 4 vdd
port 513 nsew
rlabel metal1 s 19728 46069 19728 46069 4 vdd
port 513 nsew
rlabel metal1 s 12720 47649 12720 47649 4 vdd
port 513 nsew
rlabel metal1 s 12720 50019 12720 50019 4 vdd
port 513 nsew
rlabel metal1 s 12720 48730 12720 48730 4 vdd
port 513 nsew
rlabel metal1 s 13488 47649 13488 47649 4 vdd
port 513 nsew
rlabel metal1 s 14736 48439 14736 48439 4 vdd
port 513 nsew
rlabel metal1 s 13488 49520 13488 49520 4 vdd
port 513 nsew
rlabel metal1 s 14736 47940 14736 47940 4 vdd
port 513 nsew
rlabel metal1 s 14736 49229 14736 49229 4 vdd
port 513 nsew
rlabel metal1 s 12720 47940 12720 47940 4 vdd
port 513 nsew
rlabel metal1 s 13968 48730 13968 48730 4 vdd
port 513 nsew
rlabel metal1 s 14736 49520 14736 49520 4 vdd
port 513 nsew
rlabel metal1 s 13968 50019 13968 50019 4 vdd
port 513 nsew
rlabel metal1 s 14736 47649 14736 47649 4 vdd
port 513 nsew
rlabel metal1 s 13968 50310 13968 50310 4 vdd
port 513 nsew
rlabel metal1 s 12720 50310 12720 50310 4 vdd
port 513 nsew
rlabel metal1 s 12720 49520 12720 49520 4 vdd
port 513 nsew
rlabel metal1 s 13968 48439 13968 48439 4 vdd
port 513 nsew
rlabel metal1 s 12720 48439 12720 48439 4 vdd
port 513 nsew
rlabel metal1 s 13488 50310 13488 50310 4 vdd
port 513 nsew
rlabel metal1 s 13968 49520 13968 49520 4 vdd
port 513 nsew
rlabel metal1 s 13968 47649 13968 47649 4 vdd
port 513 nsew
rlabel metal1 s 14736 48730 14736 48730 4 vdd
port 513 nsew
rlabel metal1 s 13488 49229 13488 49229 4 vdd
port 513 nsew
rlabel metal1 s 12720 49229 12720 49229 4 vdd
port 513 nsew
rlabel metal1 s 13968 49229 13968 49229 4 vdd
port 513 nsew
rlabel metal1 s 13488 47940 13488 47940 4 vdd
port 513 nsew
rlabel metal1 s 14736 50019 14736 50019 4 vdd
port 513 nsew
rlabel metal1 s 13488 48730 13488 48730 4 vdd
port 513 nsew
rlabel metal1 s 13488 48439 13488 48439 4 vdd
port 513 nsew
rlabel metal1 s 14736 50310 14736 50310 4 vdd
port 513 nsew
rlabel metal1 s 13488 50019 13488 50019 4 vdd
port 513 nsew
rlabel metal1 s 13968 47940 13968 47940 4 vdd
port 513 nsew
rlabel metal1 s 12240 50310 12240 50310 4 vdd
port 513 nsew
rlabel metal1 s 10992 48439 10992 48439 4 vdd
port 513 nsew
rlabel metal1 s 11472 47940 11472 47940 4 vdd
port 513 nsew
rlabel metal1 s 11472 49520 11472 49520 4 vdd
port 513 nsew
rlabel metal1 s 10224 47940 10224 47940 4 vdd
port 513 nsew
rlabel metal1 s 12240 48439 12240 48439 4 vdd
port 513 nsew
rlabel metal1 s 12240 47649 12240 47649 4 vdd
port 513 nsew
rlabel metal1 s 12240 49229 12240 49229 4 vdd
port 513 nsew
rlabel metal1 s 10224 50310 10224 50310 4 vdd
port 513 nsew
rlabel metal1 s 10224 49520 10224 49520 4 vdd
port 513 nsew
rlabel metal1 s 11472 50019 11472 50019 4 vdd
port 513 nsew
rlabel metal1 s 11472 50310 11472 50310 4 vdd
port 513 nsew
rlabel metal1 s 12240 49520 12240 49520 4 vdd
port 513 nsew
rlabel metal1 s 11472 49229 11472 49229 4 vdd
port 513 nsew
rlabel metal1 s 10992 49520 10992 49520 4 vdd
port 513 nsew
rlabel metal1 s 10992 49229 10992 49229 4 vdd
port 513 nsew
rlabel metal1 s 10992 47649 10992 47649 4 vdd
port 513 nsew
rlabel metal1 s 10992 50310 10992 50310 4 vdd
port 513 nsew
rlabel metal1 s 11472 47649 11472 47649 4 vdd
port 513 nsew
rlabel metal1 s 10224 50019 10224 50019 4 vdd
port 513 nsew
rlabel metal1 s 11472 48730 11472 48730 4 vdd
port 513 nsew
rlabel metal1 s 10992 50019 10992 50019 4 vdd
port 513 nsew
rlabel metal1 s 10992 47940 10992 47940 4 vdd
port 513 nsew
rlabel metal1 s 10224 47649 10224 47649 4 vdd
port 513 nsew
rlabel metal1 s 12240 47940 12240 47940 4 vdd
port 513 nsew
rlabel metal1 s 12240 48730 12240 48730 4 vdd
port 513 nsew
rlabel metal1 s 10224 49229 10224 49229 4 vdd
port 513 nsew
rlabel metal1 s 10224 48730 10224 48730 4 vdd
port 513 nsew
rlabel metal1 s 10224 48439 10224 48439 4 vdd
port 513 nsew
rlabel metal1 s 12240 50019 12240 50019 4 vdd
port 513 nsew
rlabel metal1 s 10992 48730 10992 48730 4 vdd
port 513 nsew
rlabel metal1 s 11472 48439 11472 48439 4 vdd
port 513 nsew
rlabel metal1 s 12240 47150 12240 47150 4 vdd
port 513 nsew
rlabel metal1 s 10992 45570 10992 45570 4 vdd
port 513 nsew
rlabel metal1 s 10992 44489 10992 44489 4 vdd
port 513 nsew
rlabel metal1 s 12240 46360 12240 46360 4 vdd
port 513 nsew
rlabel metal1 s 10224 46360 10224 46360 4 vdd
port 513 nsew
rlabel metal1 s 10992 44780 10992 44780 4 vdd
port 513 nsew
rlabel metal1 s 11472 44780 11472 44780 4 vdd
port 513 nsew
rlabel metal1 s 10224 44489 10224 44489 4 vdd
port 513 nsew
rlabel metal1 s 12240 46069 12240 46069 4 vdd
port 513 nsew
rlabel metal1 s 11472 46069 11472 46069 4 vdd
port 513 nsew
rlabel metal1 s 12240 44489 12240 44489 4 vdd
port 513 nsew
rlabel metal1 s 11472 47150 11472 47150 4 vdd
port 513 nsew
rlabel metal1 s 11472 45279 11472 45279 4 vdd
port 513 nsew
rlabel metal1 s 10224 45570 10224 45570 4 vdd
port 513 nsew
rlabel metal1 s 10992 47150 10992 47150 4 vdd
port 513 nsew
rlabel metal1 s 12240 45570 12240 45570 4 vdd
port 513 nsew
rlabel metal1 s 11472 45570 11472 45570 4 vdd
port 513 nsew
rlabel metal1 s 10224 47150 10224 47150 4 vdd
port 513 nsew
rlabel metal1 s 11472 44489 11472 44489 4 vdd
port 513 nsew
rlabel metal1 s 10224 44780 10224 44780 4 vdd
port 513 nsew
rlabel metal1 s 11472 46360 11472 46360 4 vdd
port 513 nsew
rlabel metal1 s 10992 45279 10992 45279 4 vdd
port 513 nsew
rlabel metal1 s 10992 46859 10992 46859 4 vdd
port 513 nsew
rlabel metal1 s 12240 46859 12240 46859 4 vdd
port 513 nsew
rlabel metal1 s 12240 44780 12240 44780 4 vdd
port 513 nsew
rlabel metal1 s 12240 45279 12240 45279 4 vdd
port 513 nsew
rlabel metal1 s 10224 46859 10224 46859 4 vdd
port 513 nsew
rlabel metal1 s 10992 46360 10992 46360 4 vdd
port 513 nsew
rlabel metal1 s 10224 46069 10224 46069 4 vdd
port 513 nsew
rlabel metal1 s 11472 46859 11472 46859 4 vdd
port 513 nsew
rlabel metal1 s 10992 46069 10992 46069 4 vdd
port 513 nsew
rlabel metal1 s 10224 45279 10224 45279 4 vdd
port 513 nsew
rlabel metal1 s 13488 44489 13488 44489 4 vdd
port 513 nsew
rlabel metal1 s 13968 44780 13968 44780 4 vdd
port 513 nsew
rlabel metal1 s 13488 45570 13488 45570 4 vdd
port 513 nsew
rlabel metal1 s 13968 45279 13968 45279 4 vdd
port 513 nsew
rlabel metal1 s 14736 46360 14736 46360 4 vdd
port 513 nsew
rlabel metal1 s 12720 46859 12720 46859 4 vdd
port 513 nsew
rlabel metal1 s 13488 46859 13488 46859 4 vdd
port 513 nsew
rlabel metal1 s 13488 47150 13488 47150 4 vdd
port 513 nsew
rlabel metal1 s 14736 45279 14736 45279 4 vdd
port 513 nsew
rlabel metal1 s 13968 46360 13968 46360 4 vdd
port 513 nsew
rlabel metal1 s 14736 44780 14736 44780 4 vdd
port 513 nsew
rlabel metal1 s 12720 44780 12720 44780 4 vdd
port 513 nsew
rlabel metal1 s 13488 46360 13488 46360 4 vdd
port 513 nsew
rlabel metal1 s 12720 45279 12720 45279 4 vdd
port 513 nsew
rlabel metal1 s 13488 45279 13488 45279 4 vdd
port 513 nsew
rlabel metal1 s 14736 46069 14736 46069 4 vdd
port 513 nsew
rlabel metal1 s 13968 45570 13968 45570 4 vdd
port 513 nsew
rlabel metal1 s 13488 44780 13488 44780 4 vdd
port 513 nsew
rlabel metal1 s 12720 47150 12720 47150 4 vdd
port 513 nsew
rlabel metal1 s 12720 46069 12720 46069 4 vdd
port 513 nsew
rlabel metal1 s 13968 47150 13968 47150 4 vdd
port 513 nsew
rlabel metal1 s 12720 45570 12720 45570 4 vdd
port 513 nsew
rlabel metal1 s 13968 46859 13968 46859 4 vdd
port 513 nsew
rlabel metal1 s 12720 46360 12720 46360 4 vdd
port 513 nsew
rlabel metal1 s 13488 46069 13488 46069 4 vdd
port 513 nsew
rlabel metal1 s 12720 44489 12720 44489 4 vdd
port 513 nsew
rlabel metal1 s 13968 46069 13968 46069 4 vdd
port 513 nsew
rlabel metal1 s 13968 44489 13968 44489 4 vdd
port 513 nsew
rlabel metal1 s 14736 45570 14736 45570 4 vdd
port 513 nsew
rlabel metal1 s 14736 47150 14736 47150 4 vdd
port 513 nsew
rlabel metal1 s 14736 44489 14736 44489 4 vdd
port 513 nsew
rlabel metal1 s 14736 46859 14736 46859 4 vdd
port 513 nsew
rlabel metal1 s 13488 43699 13488 43699 4 vdd
port 513 nsew
rlabel metal1 s 12720 43200 12720 43200 4 vdd
port 513 nsew
rlabel metal1 s 13488 43200 13488 43200 4 vdd
port 513 nsew
rlabel metal1 s 13968 43200 13968 43200 4 vdd
port 513 nsew
rlabel metal1 s 14736 43200 14736 43200 4 vdd
port 513 nsew
rlabel metal1 s 13968 42410 13968 42410 4 vdd
port 513 nsew
rlabel metal1 s 13488 43990 13488 43990 4 vdd
port 513 nsew
rlabel metal1 s 12720 43699 12720 43699 4 vdd
port 513 nsew
rlabel metal1 s 12720 42909 12720 42909 4 vdd
port 513 nsew
rlabel metal1 s 14736 42410 14736 42410 4 vdd
port 513 nsew
rlabel metal1 s 12720 41329 12720 41329 4 vdd
port 513 nsew
rlabel metal1 s 13968 43990 13968 43990 4 vdd
port 513 nsew
rlabel metal1 s 13488 42909 13488 42909 4 vdd
port 513 nsew
rlabel metal1 s 13488 41329 13488 41329 4 vdd
port 513 nsew
rlabel metal1 s 12720 43990 12720 43990 4 vdd
port 513 nsew
rlabel metal1 s 12720 41620 12720 41620 4 vdd
port 513 nsew
rlabel metal1 s 14736 41620 14736 41620 4 vdd
port 513 nsew
rlabel metal1 s 13488 42410 13488 42410 4 vdd
port 513 nsew
rlabel metal1 s 14736 41329 14736 41329 4 vdd
port 513 nsew
rlabel metal1 s 14736 43990 14736 43990 4 vdd
port 513 nsew
rlabel metal1 s 13968 41329 13968 41329 4 vdd
port 513 nsew
rlabel metal1 s 12720 42119 12720 42119 4 vdd
port 513 nsew
rlabel metal1 s 14736 42119 14736 42119 4 vdd
port 513 nsew
rlabel metal1 s 14736 43699 14736 43699 4 vdd
port 513 nsew
rlabel metal1 s 13968 42909 13968 42909 4 vdd
port 513 nsew
rlabel metal1 s 12720 42410 12720 42410 4 vdd
port 513 nsew
rlabel metal1 s 13488 41620 13488 41620 4 vdd
port 513 nsew
rlabel metal1 s 13488 42119 13488 42119 4 vdd
port 513 nsew
rlabel metal1 s 14736 42909 14736 42909 4 vdd
port 513 nsew
rlabel metal1 s 13968 43699 13968 43699 4 vdd
port 513 nsew
rlabel metal1 s 13968 42119 13968 42119 4 vdd
port 513 nsew
rlabel metal1 s 13968 41620 13968 41620 4 vdd
port 513 nsew
rlabel metal1 s 10992 43699 10992 43699 4 vdd
port 513 nsew
rlabel metal1 s 11472 43699 11472 43699 4 vdd
port 513 nsew
rlabel metal1 s 11472 42410 11472 42410 4 vdd
port 513 nsew
rlabel metal1 s 12240 42909 12240 42909 4 vdd
port 513 nsew
rlabel metal1 s 10224 41620 10224 41620 4 vdd
port 513 nsew
rlabel metal1 s 12240 42119 12240 42119 4 vdd
port 513 nsew
rlabel metal1 s 11472 43990 11472 43990 4 vdd
port 513 nsew
rlabel metal1 s 10992 43990 10992 43990 4 vdd
port 513 nsew
rlabel metal1 s 12240 41620 12240 41620 4 vdd
port 513 nsew
rlabel metal1 s 10224 43990 10224 43990 4 vdd
port 513 nsew
rlabel metal1 s 10992 42909 10992 42909 4 vdd
port 513 nsew
rlabel metal1 s 10992 42119 10992 42119 4 vdd
port 513 nsew
rlabel metal1 s 12240 43200 12240 43200 4 vdd
port 513 nsew
rlabel metal1 s 10224 43200 10224 43200 4 vdd
port 513 nsew
rlabel metal1 s 10224 41329 10224 41329 4 vdd
port 513 nsew
rlabel metal1 s 12240 43699 12240 43699 4 vdd
port 513 nsew
rlabel metal1 s 10992 41329 10992 41329 4 vdd
port 513 nsew
rlabel metal1 s 10992 41620 10992 41620 4 vdd
port 513 nsew
rlabel metal1 s 10224 43699 10224 43699 4 vdd
port 513 nsew
rlabel metal1 s 10992 42410 10992 42410 4 vdd
port 513 nsew
rlabel metal1 s 11472 42909 11472 42909 4 vdd
port 513 nsew
rlabel metal1 s 12240 41329 12240 41329 4 vdd
port 513 nsew
rlabel metal1 s 12240 43990 12240 43990 4 vdd
port 513 nsew
rlabel metal1 s 10992 43200 10992 43200 4 vdd
port 513 nsew
rlabel metal1 s 10224 42119 10224 42119 4 vdd
port 513 nsew
rlabel metal1 s 12240 42410 12240 42410 4 vdd
port 513 nsew
rlabel metal1 s 11472 42119 11472 42119 4 vdd
port 513 nsew
rlabel metal1 s 11472 43200 11472 43200 4 vdd
port 513 nsew
rlabel metal1 s 11472 41329 11472 41329 4 vdd
port 513 nsew
rlabel metal1 s 10224 42909 10224 42909 4 vdd
port 513 nsew
rlabel metal1 s 10224 42410 10224 42410 4 vdd
port 513 nsew
rlabel metal1 s 11472 41620 11472 41620 4 vdd
port 513 nsew
rlabel metal1 s 10992 38169 10992 38169 4 vdd
port 513 nsew
rlabel metal1 s 12240 38460 12240 38460 4 vdd
port 513 nsew
rlabel metal1 s 10224 40830 10224 40830 4 vdd
port 513 nsew
rlabel metal1 s 11472 38460 11472 38460 4 vdd
port 513 nsew
rlabel metal1 s 10224 39749 10224 39749 4 vdd
port 513 nsew
rlabel metal1 s 12240 38169 12240 38169 4 vdd
port 513 nsew
rlabel metal1 s 10224 38169 10224 38169 4 vdd
port 513 nsew
rlabel metal1 s 10992 38959 10992 38959 4 vdd
port 513 nsew
rlabel metal1 s 11472 40539 11472 40539 4 vdd
port 513 nsew
rlabel metal1 s 11472 38959 11472 38959 4 vdd
port 513 nsew
rlabel metal1 s 12240 40539 12240 40539 4 vdd
port 513 nsew
rlabel metal1 s 12240 40830 12240 40830 4 vdd
port 513 nsew
rlabel metal1 s 12240 38959 12240 38959 4 vdd
port 513 nsew
rlabel metal1 s 10224 40539 10224 40539 4 vdd
port 513 nsew
rlabel metal1 s 10224 39250 10224 39250 4 vdd
port 513 nsew
rlabel metal1 s 11472 40040 11472 40040 4 vdd
port 513 nsew
rlabel metal1 s 12240 39749 12240 39749 4 vdd
port 513 nsew
rlabel metal1 s 10224 40040 10224 40040 4 vdd
port 513 nsew
rlabel metal1 s 10992 40539 10992 40539 4 vdd
port 513 nsew
rlabel metal1 s 11472 40830 11472 40830 4 vdd
port 513 nsew
rlabel metal1 s 10224 38460 10224 38460 4 vdd
port 513 nsew
rlabel metal1 s 12240 39250 12240 39250 4 vdd
port 513 nsew
rlabel metal1 s 10992 38460 10992 38460 4 vdd
port 513 nsew
rlabel metal1 s 12240 40040 12240 40040 4 vdd
port 513 nsew
rlabel metal1 s 10992 40040 10992 40040 4 vdd
port 513 nsew
rlabel metal1 s 10992 39749 10992 39749 4 vdd
port 513 nsew
rlabel metal1 s 11472 39250 11472 39250 4 vdd
port 513 nsew
rlabel metal1 s 10992 39250 10992 39250 4 vdd
port 513 nsew
rlabel metal1 s 10992 40830 10992 40830 4 vdd
port 513 nsew
rlabel metal1 s 11472 39749 11472 39749 4 vdd
port 513 nsew
rlabel metal1 s 11472 38169 11472 38169 4 vdd
port 513 nsew
rlabel metal1 s 10224 38959 10224 38959 4 vdd
port 513 nsew
rlabel metal1 s 14736 38169 14736 38169 4 vdd
port 513 nsew
rlabel metal1 s 14736 38460 14736 38460 4 vdd
port 513 nsew
rlabel metal1 s 12720 40040 12720 40040 4 vdd
port 513 nsew
rlabel metal1 s 13968 40040 13968 40040 4 vdd
port 513 nsew
rlabel metal1 s 12720 38460 12720 38460 4 vdd
port 513 nsew
rlabel metal1 s 14736 40040 14736 40040 4 vdd
port 513 nsew
rlabel metal1 s 13968 39250 13968 39250 4 vdd
port 513 nsew
rlabel metal1 s 13488 40040 13488 40040 4 vdd
port 513 nsew
rlabel metal1 s 13488 38460 13488 38460 4 vdd
port 513 nsew
rlabel metal1 s 13488 38959 13488 38959 4 vdd
port 513 nsew
rlabel metal1 s 14736 38959 14736 38959 4 vdd
port 513 nsew
rlabel metal1 s 14736 39250 14736 39250 4 vdd
port 513 nsew
rlabel metal1 s 12720 40539 12720 40539 4 vdd
port 513 nsew
rlabel metal1 s 13968 39749 13968 39749 4 vdd
port 513 nsew
rlabel metal1 s 13968 38460 13968 38460 4 vdd
port 513 nsew
rlabel metal1 s 13488 39749 13488 39749 4 vdd
port 513 nsew
rlabel metal1 s 13488 38169 13488 38169 4 vdd
port 513 nsew
rlabel metal1 s 13488 40830 13488 40830 4 vdd
port 513 nsew
rlabel metal1 s 12720 39749 12720 39749 4 vdd
port 513 nsew
rlabel metal1 s 13968 40539 13968 40539 4 vdd
port 513 nsew
rlabel metal1 s 12720 40830 12720 40830 4 vdd
port 513 nsew
rlabel metal1 s 13968 38169 13968 38169 4 vdd
port 513 nsew
rlabel metal1 s 13488 40539 13488 40539 4 vdd
port 513 nsew
rlabel metal1 s 14736 40539 14736 40539 4 vdd
port 513 nsew
rlabel metal1 s 14736 40830 14736 40830 4 vdd
port 513 nsew
rlabel metal1 s 12720 39250 12720 39250 4 vdd
port 513 nsew
rlabel metal1 s 13488 39250 13488 39250 4 vdd
port 513 nsew
rlabel metal1 s 13968 38959 13968 38959 4 vdd
port 513 nsew
rlabel metal1 s 14736 39749 14736 39749 4 vdd
port 513 nsew
rlabel metal1 s 13968 40830 13968 40830 4 vdd
port 513 nsew
rlabel metal1 s 12720 38169 12720 38169 4 vdd
port 513 nsew
rlabel metal1 s 12720 38959 12720 38959 4 vdd
port 513 nsew
rlabel metal1 s 18480 43990 18480 43990 4 vdd
port 513 nsew
rlabel metal1 s 17712 43990 17712 43990 4 vdd
port 513 nsew
rlabel metal1 s 18480 43200 18480 43200 4 vdd
port 513 nsew
rlabel metal1 s 18960 43990 18960 43990 4 vdd
port 513 nsew
rlabel metal1 s 18480 41620 18480 41620 4 vdd
port 513 nsew
rlabel metal1 s 18480 41329 18480 41329 4 vdd
port 513 nsew
rlabel metal1 s 18480 42119 18480 42119 4 vdd
port 513 nsew
rlabel metal1 s 17712 41620 17712 41620 4 vdd
port 513 nsew
rlabel metal1 s 19728 43699 19728 43699 4 vdd
port 513 nsew
rlabel metal1 s 17712 42410 17712 42410 4 vdd
port 513 nsew
rlabel metal1 s 18960 42410 18960 42410 4 vdd
port 513 nsew
rlabel metal1 s 19728 42119 19728 42119 4 vdd
port 513 nsew
rlabel metal1 s 19728 43200 19728 43200 4 vdd
port 513 nsew
rlabel metal1 s 17712 43200 17712 43200 4 vdd
port 513 nsew
rlabel metal1 s 19728 41620 19728 41620 4 vdd
port 513 nsew
rlabel metal1 s 18480 42410 18480 42410 4 vdd
port 513 nsew
rlabel metal1 s 18960 42909 18960 42909 4 vdd
port 513 nsew
rlabel metal1 s 19728 41329 19728 41329 4 vdd
port 513 nsew
rlabel metal1 s 17712 42909 17712 42909 4 vdd
port 513 nsew
rlabel metal1 s 18960 41620 18960 41620 4 vdd
port 513 nsew
rlabel metal1 s 17712 41329 17712 41329 4 vdd
port 513 nsew
rlabel metal1 s 18960 43200 18960 43200 4 vdd
port 513 nsew
rlabel metal1 s 18960 41329 18960 41329 4 vdd
port 513 nsew
rlabel metal1 s 19728 42909 19728 42909 4 vdd
port 513 nsew
rlabel metal1 s 19728 42410 19728 42410 4 vdd
port 513 nsew
rlabel metal1 s 17712 43699 17712 43699 4 vdd
port 513 nsew
rlabel metal1 s 18960 43699 18960 43699 4 vdd
port 513 nsew
rlabel metal1 s 18480 43699 18480 43699 4 vdd
port 513 nsew
rlabel metal1 s 19728 43990 19728 43990 4 vdd
port 513 nsew
rlabel metal1 s 17712 42119 17712 42119 4 vdd
port 513 nsew
rlabel metal1 s 18480 42909 18480 42909 4 vdd
port 513 nsew
rlabel metal1 s 18960 42119 18960 42119 4 vdd
port 513 nsew
rlabel metal1 s 15984 43200 15984 43200 4 vdd
port 513 nsew
rlabel metal1 s 16464 43699 16464 43699 4 vdd
port 513 nsew
rlabel metal1 s 16464 43200 16464 43200 4 vdd
port 513 nsew
rlabel metal1 s 15216 43200 15216 43200 4 vdd
port 513 nsew
rlabel metal1 s 15984 41329 15984 41329 4 vdd
port 513 nsew
rlabel metal1 s 15984 42410 15984 42410 4 vdd
port 513 nsew
rlabel metal1 s 15216 42909 15216 42909 4 vdd
port 513 nsew
rlabel metal1 s 17232 43990 17232 43990 4 vdd
port 513 nsew
rlabel metal1 s 17232 42410 17232 42410 4 vdd
port 513 nsew
rlabel metal1 s 17232 43200 17232 43200 4 vdd
port 513 nsew
rlabel metal1 s 15216 41620 15216 41620 4 vdd
port 513 nsew
rlabel metal1 s 17232 41620 17232 41620 4 vdd
port 513 nsew
rlabel metal1 s 15984 42119 15984 42119 4 vdd
port 513 nsew
rlabel metal1 s 15216 43990 15216 43990 4 vdd
port 513 nsew
rlabel metal1 s 15216 42410 15216 42410 4 vdd
port 513 nsew
rlabel metal1 s 17232 43699 17232 43699 4 vdd
port 513 nsew
rlabel metal1 s 15984 41620 15984 41620 4 vdd
port 513 nsew
rlabel metal1 s 15984 43699 15984 43699 4 vdd
port 513 nsew
rlabel metal1 s 17232 42909 17232 42909 4 vdd
port 513 nsew
rlabel metal1 s 15216 43699 15216 43699 4 vdd
port 513 nsew
rlabel metal1 s 15216 41329 15216 41329 4 vdd
port 513 nsew
rlabel metal1 s 17232 42119 17232 42119 4 vdd
port 513 nsew
rlabel metal1 s 16464 42909 16464 42909 4 vdd
port 513 nsew
rlabel metal1 s 15984 43990 15984 43990 4 vdd
port 513 nsew
rlabel metal1 s 16464 42410 16464 42410 4 vdd
port 513 nsew
rlabel metal1 s 17232 41329 17232 41329 4 vdd
port 513 nsew
rlabel metal1 s 16464 42119 16464 42119 4 vdd
port 513 nsew
rlabel metal1 s 16464 41620 16464 41620 4 vdd
port 513 nsew
rlabel metal1 s 15216 42119 15216 42119 4 vdd
port 513 nsew
rlabel metal1 s 15984 42909 15984 42909 4 vdd
port 513 nsew
rlabel metal1 s 16464 43990 16464 43990 4 vdd
port 513 nsew
rlabel metal1 s 16464 41329 16464 41329 4 vdd
port 513 nsew
rlabel metal1 s 15216 39250 15216 39250 4 vdd
port 513 nsew
rlabel metal1 s 16464 39749 16464 39749 4 vdd
port 513 nsew
rlabel metal1 s 15984 39749 15984 39749 4 vdd
port 513 nsew
rlabel metal1 s 15984 40539 15984 40539 4 vdd
port 513 nsew
rlabel metal1 s 15216 38959 15216 38959 4 vdd
port 513 nsew
rlabel metal1 s 16464 38169 16464 38169 4 vdd
port 513 nsew
rlabel metal1 s 15216 40539 15216 40539 4 vdd
port 513 nsew
rlabel metal1 s 17232 40830 17232 40830 4 vdd
port 513 nsew
rlabel metal1 s 17232 38460 17232 38460 4 vdd
port 513 nsew
rlabel metal1 s 15984 40830 15984 40830 4 vdd
port 513 nsew
rlabel metal1 s 15216 38460 15216 38460 4 vdd
port 513 nsew
rlabel metal1 s 16464 39250 16464 39250 4 vdd
port 513 nsew
rlabel metal1 s 15216 40040 15216 40040 4 vdd
port 513 nsew
rlabel metal1 s 16464 40539 16464 40539 4 vdd
port 513 nsew
rlabel metal1 s 17232 40539 17232 40539 4 vdd
port 513 nsew
rlabel metal1 s 15984 38959 15984 38959 4 vdd
port 513 nsew
rlabel metal1 s 16464 38460 16464 38460 4 vdd
port 513 nsew
rlabel metal1 s 17232 40040 17232 40040 4 vdd
port 513 nsew
rlabel metal1 s 15216 38169 15216 38169 4 vdd
port 513 nsew
rlabel metal1 s 17232 38169 17232 38169 4 vdd
port 513 nsew
rlabel metal1 s 17232 39749 17232 39749 4 vdd
port 513 nsew
rlabel metal1 s 15984 40040 15984 40040 4 vdd
port 513 nsew
rlabel metal1 s 15984 38460 15984 38460 4 vdd
port 513 nsew
rlabel metal1 s 16464 38959 16464 38959 4 vdd
port 513 nsew
rlabel metal1 s 16464 40040 16464 40040 4 vdd
port 513 nsew
rlabel metal1 s 15984 38169 15984 38169 4 vdd
port 513 nsew
rlabel metal1 s 15216 39749 15216 39749 4 vdd
port 513 nsew
rlabel metal1 s 17232 39250 17232 39250 4 vdd
port 513 nsew
rlabel metal1 s 15984 39250 15984 39250 4 vdd
port 513 nsew
rlabel metal1 s 15216 40830 15216 40830 4 vdd
port 513 nsew
rlabel metal1 s 16464 40830 16464 40830 4 vdd
port 513 nsew
rlabel metal1 s 17232 38959 17232 38959 4 vdd
port 513 nsew
rlabel metal1 s 19728 40539 19728 40539 4 vdd
port 513 nsew
rlabel metal1 s 18480 38959 18480 38959 4 vdd
port 513 nsew
rlabel metal1 s 17712 38169 17712 38169 4 vdd
port 513 nsew
rlabel metal1 s 17712 40830 17712 40830 4 vdd
port 513 nsew
rlabel metal1 s 19728 38169 19728 38169 4 vdd
port 513 nsew
rlabel metal1 s 18960 38460 18960 38460 4 vdd
port 513 nsew
rlabel metal1 s 19728 40040 19728 40040 4 vdd
port 513 nsew
rlabel metal1 s 19728 38959 19728 38959 4 vdd
port 513 nsew
rlabel metal1 s 17712 38460 17712 38460 4 vdd
port 513 nsew
rlabel metal1 s 18960 39749 18960 39749 4 vdd
port 513 nsew
rlabel metal1 s 18480 40830 18480 40830 4 vdd
port 513 nsew
rlabel metal1 s 18480 39250 18480 39250 4 vdd
port 513 nsew
rlabel metal1 s 17712 40040 17712 40040 4 vdd
port 513 nsew
rlabel metal1 s 19728 39749 19728 39749 4 vdd
port 513 nsew
rlabel metal1 s 17712 39250 17712 39250 4 vdd
port 513 nsew
rlabel metal1 s 17712 38959 17712 38959 4 vdd
port 513 nsew
rlabel metal1 s 18960 40830 18960 40830 4 vdd
port 513 nsew
rlabel metal1 s 18480 38169 18480 38169 4 vdd
port 513 nsew
rlabel metal1 s 19728 40830 19728 40830 4 vdd
port 513 nsew
rlabel metal1 s 19728 39250 19728 39250 4 vdd
port 513 nsew
rlabel metal1 s 18960 38959 18960 38959 4 vdd
port 513 nsew
rlabel metal1 s 18480 39749 18480 39749 4 vdd
port 513 nsew
rlabel metal1 s 18960 38169 18960 38169 4 vdd
port 513 nsew
rlabel metal1 s 18960 40040 18960 40040 4 vdd
port 513 nsew
rlabel metal1 s 18480 38460 18480 38460 4 vdd
port 513 nsew
rlabel metal1 s 17712 39749 17712 39749 4 vdd
port 513 nsew
rlabel metal1 s 18960 39250 18960 39250 4 vdd
port 513 nsew
rlabel metal1 s 18480 40539 18480 40539 4 vdd
port 513 nsew
rlabel metal1 s 18480 40040 18480 40040 4 vdd
port 513 nsew
rlabel metal1 s 17712 40539 17712 40539 4 vdd
port 513 nsew
rlabel metal1 s 19728 38460 19728 38460 4 vdd
port 513 nsew
rlabel metal1 s 18960 40539 18960 40539 4 vdd
port 513 nsew
rlabel metal1 s 8976 47649 8976 47649 4 vdd
port 513 nsew
rlabel metal1 s 7728 48730 7728 48730 4 vdd
port 513 nsew
rlabel metal1 s 9744 48439 9744 48439 4 vdd
port 513 nsew
rlabel metal1 s 8976 50019 8976 50019 4 vdd
port 513 nsew
rlabel metal1 s 8976 48730 8976 48730 4 vdd
port 513 nsew
rlabel metal1 s 9744 49520 9744 49520 4 vdd
port 513 nsew
rlabel metal1 s 8496 48439 8496 48439 4 vdd
port 513 nsew
rlabel metal1 s 8496 50310 8496 50310 4 vdd
port 513 nsew
rlabel metal1 s 7728 49229 7728 49229 4 vdd
port 513 nsew
rlabel metal1 s 8496 49229 8496 49229 4 vdd
port 513 nsew
rlabel metal1 s 8496 47649 8496 47649 4 vdd
port 513 nsew
rlabel metal1 s 8976 50310 8976 50310 4 vdd
port 513 nsew
rlabel metal1 s 7728 50019 7728 50019 4 vdd
port 513 nsew
rlabel metal1 s 7728 49520 7728 49520 4 vdd
port 513 nsew
rlabel metal1 s 7728 47940 7728 47940 4 vdd
port 513 nsew
rlabel metal1 s 8976 49229 8976 49229 4 vdd
port 513 nsew
rlabel metal1 s 8976 47940 8976 47940 4 vdd
port 513 nsew
rlabel metal1 s 9744 47940 9744 47940 4 vdd
port 513 nsew
rlabel metal1 s 7728 50310 7728 50310 4 vdd
port 513 nsew
rlabel metal1 s 9744 50310 9744 50310 4 vdd
port 513 nsew
rlabel metal1 s 9744 50019 9744 50019 4 vdd
port 513 nsew
rlabel metal1 s 9744 49229 9744 49229 4 vdd
port 513 nsew
rlabel metal1 s 8976 48439 8976 48439 4 vdd
port 513 nsew
rlabel metal1 s 8496 47940 8496 47940 4 vdd
port 513 nsew
rlabel metal1 s 9744 47649 9744 47649 4 vdd
port 513 nsew
rlabel metal1 s 8976 49520 8976 49520 4 vdd
port 513 nsew
rlabel metal1 s 7728 48439 7728 48439 4 vdd
port 513 nsew
rlabel metal1 s 7728 47649 7728 47649 4 vdd
port 513 nsew
rlabel metal1 s 9744 48730 9744 48730 4 vdd
port 513 nsew
rlabel metal1 s 8496 49520 8496 49520 4 vdd
port 513 nsew
rlabel metal1 s 8496 48730 8496 48730 4 vdd
port 513 nsew
rlabel metal1 s 8496 50019 8496 50019 4 vdd
port 513 nsew
rlabel metal1 s 5232 50019 5232 50019 4 vdd
port 513 nsew
rlabel metal1 s 6480 48730 6480 48730 4 vdd
port 513 nsew
rlabel metal1 s 5232 47649 5232 47649 4 vdd
port 513 nsew
rlabel metal1 s 5232 50310 5232 50310 4 vdd
port 513 nsew
rlabel metal1 s 6480 49229 6480 49229 4 vdd
port 513 nsew
rlabel metal1 s 6000 49520 6000 49520 4 vdd
port 513 nsew
rlabel metal1 s 5232 48730 5232 48730 4 vdd
port 513 nsew
rlabel metal1 s 7248 47649 7248 47649 4 vdd
port 513 nsew
rlabel metal1 s 6000 50019 6000 50019 4 vdd
port 513 nsew
rlabel metal1 s 7248 49520 7248 49520 4 vdd
port 513 nsew
rlabel metal1 s 5232 49229 5232 49229 4 vdd
port 513 nsew
rlabel metal1 s 6000 48730 6000 48730 4 vdd
port 513 nsew
rlabel metal1 s 7248 50019 7248 50019 4 vdd
port 513 nsew
rlabel metal1 s 6480 50310 6480 50310 4 vdd
port 513 nsew
rlabel metal1 s 5232 49520 5232 49520 4 vdd
port 513 nsew
rlabel metal1 s 6000 47649 6000 47649 4 vdd
port 513 nsew
rlabel metal1 s 6000 48439 6000 48439 4 vdd
port 513 nsew
rlabel metal1 s 6480 47649 6480 47649 4 vdd
port 513 nsew
rlabel metal1 s 5232 47940 5232 47940 4 vdd
port 513 nsew
rlabel metal1 s 6000 49229 6000 49229 4 vdd
port 513 nsew
rlabel metal1 s 6480 47940 6480 47940 4 vdd
port 513 nsew
rlabel metal1 s 7248 47940 7248 47940 4 vdd
port 513 nsew
rlabel metal1 s 5232 48439 5232 48439 4 vdd
port 513 nsew
rlabel metal1 s 7248 48730 7248 48730 4 vdd
port 513 nsew
rlabel metal1 s 7248 50310 7248 50310 4 vdd
port 513 nsew
rlabel metal1 s 6480 50019 6480 50019 4 vdd
port 513 nsew
rlabel metal1 s 6480 48439 6480 48439 4 vdd
port 513 nsew
rlabel metal1 s 7248 49229 7248 49229 4 vdd
port 513 nsew
rlabel metal1 s 6480 49520 6480 49520 4 vdd
port 513 nsew
rlabel metal1 s 6000 47940 6000 47940 4 vdd
port 513 nsew
rlabel metal1 s 6000 50310 6000 50310 4 vdd
port 513 nsew
rlabel metal1 s 7248 48439 7248 48439 4 vdd
port 513 nsew
rlabel metal1 s 6480 46360 6480 46360 4 vdd
port 513 nsew
rlabel metal1 s 5232 45279 5232 45279 4 vdd
port 513 nsew
rlabel metal1 s 5232 46360 5232 46360 4 vdd
port 513 nsew
rlabel metal1 s 7248 44489 7248 44489 4 vdd
port 513 nsew
rlabel metal1 s 7248 46069 7248 46069 4 vdd
port 513 nsew
rlabel metal1 s 5232 47150 5232 47150 4 vdd
port 513 nsew
rlabel metal1 s 7248 46360 7248 46360 4 vdd
port 513 nsew
rlabel metal1 s 5232 46069 5232 46069 4 vdd
port 513 nsew
rlabel metal1 s 6000 45570 6000 45570 4 vdd
port 513 nsew
rlabel metal1 s 6000 45279 6000 45279 4 vdd
port 513 nsew
rlabel metal1 s 7248 46859 7248 46859 4 vdd
port 513 nsew
rlabel metal1 s 6000 44780 6000 44780 4 vdd
port 513 nsew
rlabel metal1 s 6480 45279 6480 45279 4 vdd
port 513 nsew
rlabel metal1 s 6480 47150 6480 47150 4 vdd
port 513 nsew
rlabel metal1 s 5232 46859 5232 46859 4 vdd
port 513 nsew
rlabel metal1 s 6480 44780 6480 44780 4 vdd
port 513 nsew
rlabel metal1 s 5232 45570 5232 45570 4 vdd
port 513 nsew
rlabel metal1 s 6000 46069 6000 46069 4 vdd
port 513 nsew
rlabel metal1 s 6000 47150 6000 47150 4 vdd
port 513 nsew
rlabel metal1 s 6480 44489 6480 44489 4 vdd
port 513 nsew
rlabel metal1 s 6000 46859 6000 46859 4 vdd
port 513 nsew
rlabel metal1 s 6480 45570 6480 45570 4 vdd
port 513 nsew
rlabel metal1 s 5232 44489 5232 44489 4 vdd
port 513 nsew
rlabel metal1 s 6480 46859 6480 46859 4 vdd
port 513 nsew
rlabel metal1 s 6000 44489 6000 44489 4 vdd
port 513 nsew
rlabel metal1 s 6480 46069 6480 46069 4 vdd
port 513 nsew
rlabel metal1 s 5232 44780 5232 44780 4 vdd
port 513 nsew
rlabel metal1 s 7248 45279 7248 45279 4 vdd
port 513 nsew
rlabel metal1 s 6000 46360 6000 46360 4 vdd
port 513 nsew
rlabel metal1 s 7248 45570 7248 45570 4 vdd
port 513 nsew
rlabel metal1 s 7248 47150 7248 47150 4 vdd
port 513 nsew
rlabel metal1 s 7248 44780 7248 44780 4 vdd
port 513 nsew
rlabel metal1 s 8976 45279 8976 45279 4 vdd
port 513 nsew
rlabel metal1 s 8976 46069 8976 46069 4 vdd
port 513 nsew
rlabel metal1 s 8496 46859 8496 46859 4 vdd
port 513 nsew
rlabel metal1 s 8496 45570 8496 45570 4 vdd
port 513 nsew
rlabel metal1 s 8496 44780 8496 44780 4 vdd
port 513 nsew
rlabel metal1 s 8496 44489 8496 44489 4 vdd
port 513 nsew
rlabel metal1 s 8496 45279 8496 45279 4 vdd
port 513 nsew
rlabel metal1 s 7728 44780 7728 44780 4 vdd
port 513 nsew
rlabel metal1 s 7728 45570 7728 45570 4 vdd
port 513 nsew
rlabel metal1 s 8976 46859 8976 46859 4 vdd
port 513 nsew
rlabel metal1 s 7728 46360 7728 46360 4 vdd
port 513 nsew
rlabel metal1 s 8496 46360 8496 46360 4 vdd
port 513 nsew
rlabel metal1 s 9744 45570 9744 45570 4 vdd
port 513 nsew
rlabel metal1 s 9744 47150 9744 47150 4 vdd
port 513 nsew
rlabel metal1 s 8496 46069 8496 46069 4 vdd
port 513 nsew
rlabel metal1 s 8976 44489 8976 44489 4 vdd
port 513 nsew
rlabel metal1 s 9744 44489 9744 44489 4 vdd
port 513 nsew
rlabel metal1 s 7728 46859 7728 46859 4 vdd
port 513 nsew
rlabel metal1 s 9744 46859 9744 46859 4 vdd
port 513 nsew
rlabel metal1 s 7728 45279 7728 45279 4 vdd
port 513 nsew
rlabel metal1 s 9744 44780 9744 44780 4 vdd
port 513 nsew
rlabel metal1 s 7728 44489 7728 44489 4 vdd
port 513 nsew
rlabel metal1 s 7728 46069 7728 46069 4 vdd
port 513 nsew
rlabel metal1 s 8976 47150 8976 47150 4 vdd
port 513 nsew
rlabel metal1 s 8976 44780 8976 44780 4 vdd
port 513 nsew
rlabel metal1 s 8976 45570 8976 45570 4 vdd
port 513 nsew
rlabel metal1 s 8976 46360 8976 46360 4 vdd
port 513 nsew
rlabel metal1 s 8496 47150 8496 47150 4 vdd
port 513 nsew
rlabel metal1 s 9744 45279 9744 45279 4 vdd
port 513 nsew
rlabel metal1 s 9744 46360 9744 46360 4 vdd
port 513 nsew
rlabel metal1 s 9744 46069 9744 46069 4 vdd
port 513 nsew
rlabel metal1 s 7728 47150 7728 47150 4 vdd
port 513 nsew
rlabel metal1 s 3984 50310 3984 50310 4 vdd
port 513 nsew
rlabel metal1 s 3984 49229 3984 49229 4 vdd
port 513 nsew
rlabel metal1 s 3984 50019 3984 50019 4 vdd
port 513 nsew
rlabel metal1 s 2736 49520 2736 49520 4 vdd
port 513 nsew
rlabel metal1 s 4752 50310 4752 50310 4 vdd
port 513 nsew
rlabel metal1 s 4752 48730 4752 48730 4 vdd
port 513 nsew
rlabel metal1 s 2736 50310 2736 50310 4 vdd
port 513 nsew
rlabel metal1 s 3984 48439 3984 48439 4 vdd
port 513 nsew
rlabel metal1 s 3504 49229 3504 49229 4 vdd
port 513 nsew
rlabel metal1 s 4752 48439 4752 48439 4 vdd
port 513 nsew
rlabel metal1 s 3984 49520 3984 49520 4 vdd
port 513 nsew
rlabel metal1 s 3504 48439 3504 48439 4 vdd
port 513 nsew
rlabel metal1 s 4752 49520 4752 49520 4 vdd
port 513 nsew
rlabel metal1 s 2736 48730 2736 48730 4 vdd
port 513 nsew
rlabel metal1 s 4752 49229 4752 49229 4 vdd
port 513 nsew
rlabel metal1 s 4752 50019 4752 50019 4 vdd
port 513 nsew
rlabel metal1 s 3504 47940 3504 47940 4 vdd
port 513 nsew
rlabel metal1 s 2736 50019 2736 50019 4 vdd
port 513 nsew
rlabel metal1 s 3504 48730 3504 48730 4 vdd
port 513 nsew
rlabel metal1 s 3504 49520 3504 49520 4 vdd
port 513 nsew
rlabel metal1 s 3984 48730 3984 48730 4 vdd
port 513 nsew
rlabel metal1 s 3504 50310 3504 50310 4 vdd
port 513 nsew
rlabel metal1 s 3984 47940 3984 47940 4 vdd
port 513 nsew
rlabel metal1 s 2736 49229 2736 49229 4 vdd
port 513 nsew
rlabel metal1 s 2736 47649 2736 47649 4 vdd
port 513 nsew
rlabel metal1 s 3504 50019 3504 50019 4 vdd
port 513 nsew
rlabel metal1 s 3504 47649 3504 47649 4 vdd
port 513 nsew
rlabel metal1 s 4752 47940 4752 47940 4 vdd
port 513 nsew
rlabel metal1 s 3984 47649 3984 47649 4 vdd
port 513 nsew
rlabel metal1 s 4752 47649 4752 47649 4 vdd
port 513 nsew
rlabel metal1 s 2736 48439 2736 48439 4 vdd
port 513 nsew
rlabel metal1 s 2736 47940 2736 47940 4 vdd
port 513 nsew
rlabel metal1 s 1008 49520 1008 49520 4 vdd
port 513 nsew
rlabel metal1 s 1488 48439 1488 48439 4 vdd
port 513 nsew
rlabel metal1 s 2256 48730 2256 48730 4 vdd
port 513 nsew
rlabel metal1 s 1008 48439 1008 48439 4 vdd
port 513 nsew
rlabel metal1 s 1488 49520 1488 49520 4 vdd
port 513 nsew
rlabel metal1 s 240 49229 240 49229 4 vdd
port 513 nsew
rlabel metal1 s 1008 47649 1008 47649 4 vdd
port 513 nsew
rlabel metal1 s 240 49520 240 49520 4 vdd
port 513 nsew
rlabel metal1 s 1488 49229 1488 49229 4 vdd
port 513 nsew
rlabel metal1 s 2256 47940 2256 47940 4 vdd
port 513 nsew
rlabel metal1 s 1488 50310 1488 50310 4 vdd
port 513 nsew
rlabel metal1 s 1488 50019 1488 50019 4 vdd
port 513 nsew
rlabel metal1 s 1008 50019 1008 50019 4 vdd
port 513 nsew
rlabel metal1 s 2256 49520 2256 49520 4 vdd
port 513 nsew
rlabel metal1 s 1008 47940 1008 47940 4 vdd
port 513 nsew
rlabel metal1 s 240 47940 240 47940 4 vdd
port 513 nsew
rlabel metal1 s 240 50019 240 50019 4 vdd
port 513 nsew
rlabel metal1 s 240 47649 240 47649 4 vdd
port 513 nsew
rlabel metal1 s 1488 47940 1488 47940 4 vdd
port 513 nsew
rlabel metal1 s 240 48730 240 48730 4 vdd
port 513 nsew
rlabel metal1 s 1008 50310 1008 50310 4 vdd
port 513 nsew
rlabel metal1 s 1008 49229 1008 49229 4 vdd
port 513 nsew
rlabel metal1 s 2256 50310 2256 50310 4 vdd
port 513 nsew
rlabel metal1 s 1488 48730 1488 48730 4 vdd
port 513 nsew
rlabel metal1 s 2256 50019 2256 50019 4 vdd
port 513 nsew
rlabel metal1 s 240 48439 240 48439 4 vdd
port 513 nsew
rlabel metal1 s 1008 48730 1008 48730 4 vdd
port 513 nsew
rlabel metal1 s 2256 47649 2256 47649 4 vdd
port 513 nsew
rlabel metal1 s 1488 47649 1488 47649 4 vdd
port 513 nsew
rlabel metal1 s 240 50310 240 50310 4 vdd
port 513 nsew
rlabel metal1 s 2256 49229 2256 49229 4 vdd
port 513 nsew
rlabel metal1 s 2256 48439 2256 48439 4 vdd
port 513 nsew
rlabel metal1 s 1488 44489 1488 44489 4 vdd
port 513 nsew
rlabel metal1 s 1488 46360 1488 46360 4 vdd
port 513 nsew
rlabel metal1 s 1008 47150 1008 47150 4 vdd
port 513 nsew
rlabel metal1 s 240 44489 240 44489 4 vdd
port 513 nsew
rlabel metal1 s 1008 46069 1008 46069 4 vdd
port 513 nsew
rlabel metal1 s 2256 46069 2256 46069 4 vdd
port 513 nsew
rlabel metal1 s 1008 46360 1008 46360 4 vdd
port 513 nsew
rlabel metal1 s 1488 44780 1488 44780 4 vdd
port 513 nsew
rlabel metal1 s 1488 45279 1488 45279 4 vdd
port 513 nsew
rlabel metal1 s 1008 44489 1008 44489 4 vdd
port 513 nsew
rlabel metal1 s 240 44780 240 44780 4 vdd
port 513 nsew
rlabel metal1 s 2256 44489 2256 44489 4 vdd
port 513 nsew
rlabel metal1 s 240 47150 240 47150 4 vdd
port 513 nsew
rlabel metal1 s 2256 46859 2256 46859 4 vdd
port 513 nsew
rlabel metal1 s 2256 45279 2256 45279 4 vdd
port 513 nsew
rlabel metal1 s 1008 46859 1008 46859 4 vdd
port 513 nsew
rlabel metal1 s 1488 47150 1488 47150 4 vdd
port 513 nsew
rlabel metal1 s 240 45279 240 45279 4 vdd
port 513 nsew
rlabel metal1 s 2256 44780 2256 44780 4 vdd
port 513 nsew
rlabel metal1 s 2256 46360 2256 46360 4 vdd
port 513 nsew
rlabel metal1 s 240 46360 240 46360 4 vdd
port 513 nsew
rlabel metal1 s 1008 45279 1008 45279 4 vdd
port 513 nsew
rlabel metal1 s 1488 45570 1488 45570 4 vdd
port 513 nsew
rlabel metal1 s 2256 45570 2256 45570 4 vdd
port 513 nsew
rlabel metal1 s 240 46859 240 46859 4 vdd
port 513 nsew
rlabel metal1 s 240 45570 240 45570 4 vdd
port 513 nsew
rlabel metal1 s 1488 46859 1488 46859 4 vdd
port 513 nsew
rlabel metal1 s 1008 44780 1008 44780 4 vdd
port 513 nsew
rlabel metal1 s 240 46069 240 46069 4 vdd
port 513 nsew
rlabel metal1 s 1488 46069 1488 46069 4 vdd
port 513 nsew
rlabel metal1 s 2256 47150 2256 47150 4 vdd
port 513 nsew
rlabel metal1 s 1008 45570 1008 45570 4 vdd
port 513 nsew
rlabel metal1 s 3984 46069 3984 46069 4 vdd
port 513 nsew
rlabel metal1 s 3504 45279 3504 45279 4 vdd
port 513 nsew
rlabel metal1 s 4752 46069 4752 46069 4 vdd
port 513 nsew
rlabel metal1 s 2736 46859 2736 46859 4 vdd
port 513 nsew
rlabel metal1 s 4752 46859 4752 46859 4 vdd
port 513 nsew
rlabel metal1 s 3984 45570 3984 45570 4 vdd
port 513 nsew
rlabel metal1 s 3504 44489 3504 44489 4 vdd
port 513 nsew
rlabel metal1 s 4752 46360 4752 46360 4 vdd
port 513 nsew
rlabel metal1 s 3504 45570 3504 45570 4 vdd
port 513 nsew
rlabel metal1 s 3504 46360 3504 46360 4 vdd
port 513 nsew
rlabel metal1 s 2736 44489 2736 44489 4 vdd
port 513 nsew
rlabel metal1 s 2736 46069 2736 46069 4 vdd
port 513 nsew
rlabel metal1 s 3504 46859 3504 46859 4 vdd
port 513 nsew
rlabel metal1 s 2736 45279 2736 45279 4 vdd
port 513 nsew
rlabel metal1 s 4752 45570 4752 45570 4 vdd
port 513 nsew
rlabel metal1 s 3984 46859 3984 46859 4 vdd
port 513 nsew
rlabel metal1 s 4752 45279 4752 45279 4 vdd
port 513 nsew
rlabel metal1 s 3984 45279 3984 45279 4 vdd
port 513 nsew
rlabel metal1 s 3504 44780 3504 44780 4 vdd
port 513 nsew
rlabel metal1 s 4752 47150 4752 47150 4 vdd
port 513 nsew
rlabel metal1 s 2736 47150 2736 47150 4 vdd
port 513 nsew
rlabel metal1 s 3984 46360 3984 46360 4 vdd
port 513 nsew
rlabel metal1 s 3984 47150 3984 47150 4 vdd
port 513 nsew
rlabel metal1 s 3984 44489 3984 44489 4 vdd
port 513 nsew
rlabel metal1 s 3504 46069 3504 46069 4 vdd
port 513 nsew
rlabel metal1 s 2736 45570 2736 45570 4 vdd
port 513 nsew
rlabel metal1 s 3984 44780 3984 44780 4 vdd
port 513 nsew
rlabel metal1 s 2736 46360 2736 46360 4 vdd
port 513 nsew
rlabel metal1 s 2736 44780 2736 44780 4 vdd
port 513 nsew
rlabel metal1 s 4752 44780 4752 44780 4 vdd
port 513 nsew
rlabel metal1 s 4752 44489 4752 44489 4 vdd
port 513 nsew
rlabel metal1 s 3504 47150 3504 47150 4 vdd
port 513 nsew
rlabel metal1 s 4752 42119 4752 42119 4 vdd
port 513 nsew
rlabel metal1 s 3984 43990 3984 43990 4 vdd
port 513 nsew
rlabel metal1 s 3984 42909 3984 42909 4 vdd
port 513 nsew
rlabel metal1 s 4752 43990 4752 43990 4 vdd
port 513 nsew
rlabel metal1 s 2736 42410 2736 42410 4 vdd
port 513 nsew
rlabel metal1 s 2736 43200 2736 43200 4 vdd
port 513 nsew
rlabel metal1 s 2736 41620 2736 41620 4 vdd
port 513 nsew
rlabel metal1 s 4752 42410 4752 42410 4 vdd
port 513 nsew
rlabel metal1 s 3504 42909 3504 42909 4 vdd
port 513 nsew
rlabel metal1 s 3504 41620 3504 41620 4 vdd
port 513 nsew
rlabel metal1 s 3504 42119 3504 42119 4 vdd
port 513 nsew
rlabel metal1 s 4752 43200 4752 43200 4 vdd
port 513 nsew
rlabel metal1 s 4752 41329 4752 41329 4 vdd
port 513 nsew
rlabel metal1 s 3984 42410 3984 42410 4 vdd
port 513 nsew
rlabel metal1 s 3504 43699 3504 43699 4 vdd
port 513 nsew
rlabel metal1 s 3504 41329 3504 41329 4 vdd
port 513 nsew
rlabel metal1 s 2736 42119 2736 42119 4 vdd
port 513 nsew
rlabel metal1 s 4752 41620 4752 41620 4 vdd
port 513 nsew
rlabel metal1 s 4752 43699 4752 43699 4 vdd
port 513 nsew
rlabel metal1 s 2736 43699 2736 43699 4 vdd
port 513 nsew
rlabel metal1 s 4752 42909 4752 42909 4 vdd
port 513 nsew
rlabel metal1 s 3984 43200 3984 43200 4 vdd
port 513 nsew
rlabel metal1 s 3504 43200 3504 43200 4 vdd
port 513 nsew
rlabel metal1 s 3984 42119 3984 42119 4 vdd
port 513 nsew
rlabel metal1 s 3984 41329 3984 41329 4 vdd
port 513 nsew
rlabel metal1 s 2736 43990 2736 43990 4 vdd
port 513 nsew
rlabel metal1 s 3984 41620 3984 41620 4 vdd
port 513 nsew
rlabel metal1 s 3504 42410 3504 42410 4 vdd
port 513 nsew
rlabel metal1 s 2736 41329 2736 41329 4 vdd
port 513 nsew
rlabel metal1 s 2736 42909 2736 42909 4 vdd
port 513 nsew
rlabel metal1 s 3504 43990 3504 43990 4 vdd
port 513 nsew
rlabel metal1 s 3984 43699 3984 43699 4 vdd
port 513 nsew
rlabel metal1 s 240 43990 240 43990 4 vdd
port 513 nsew
rlabel metal1 s 240 43200 240 43200 4 vdd
port 513 nsew
rlabel metal1 s 1488 43699 1488 43699 4 vdd
port 513 nsew
rlabel metal1 s 240 42410 240 42410 4 vdd
port 513 nsew
rlabel metal1 s 2256 43990 2256 43990 4 vdd
port 513 nsew
rlabel metal1 s 1488 42119 1488 42119 4 vdd
port 513 nsew
rlabel metal1 s 1008 42119 1008 42119 4 vdd
port 513 nsew
rlabel metal1 s 240 42119 240 42119 4 vdd
port 513 nsew
rlabel metal1 s 2256 42410 2256 42410 4 vdd
port 513 nsew
rlabel metal1 s 2256 43200 2256 43200 4 vdd
port 513 nsew
rlabel metal1 s 1488 43990 1488 43990 4 vdd
port 513 nsew
rlabel metal1 s 1008 42410 1008 42410 4 vdd
port 513 nsew
rlabel metal1 s 2256 41329 2256 41329 4 vdd
port 513 nsew
rlabel metal1 s 240 43699 240 43699 4 vdd
port 513 nsew
rlabel metal1 s 2256 43699 2256 43699 4 vdd
port 513 nsew
rlabel metal1 s 1488 43200 1488 43200 4 vdd
port 513 nsew
rlabel metal1 s 1488 41329 1488 41329 4 vdd
port 513 nsew
rlabel metal1 s 1008 43990 1008 43990 4 vdd
port 513 nsew
rlabel metal1 s 240 42909 240 42909 4 vdd
port 513 nsew
rlabel metal1 s 1008 41329 1008 41329 4 vdd
port 513 nsew
rlabel metal1 s 2256 42119 2256 42119 4 vdd
port 513 nsew
rlabel metal1 s 2256 41620 2256 41620 4 vdd
port 513 nsew
rlabel metal1 s 240 41329 240 41329 4 vdd
port 513 nsew
rlabel metal1 s 2256 42909 2256 42909 4 vdd
port 513 nsew
rlabel metal1 s 1008 41620 1008 41620 4 vdd
port 513 nsew
rlabel metal1 s 240 41620 240 41620 4 vdd
port 513 nsew
rlabel metal1 s 1008 43200 1008 43200 4 vdd
port 513 nsew
rlabel metal1 s 1008 42909 1008 42909 4 vdd
port 513 nsew
rlabel metal1 s 1488 41620 1488 41620 4 vdd
port 513 nsew
rlabel metal1 s 1488 42909 1488 42909 4 vdd
port 513 nsew
rlabel metal1 s 1008 43699 1008 43699 4 vdd
port 513 nsew
rlabel metal1 s 1488 42410 1488 42410 4 vdd
port 513 nsew
rlabel metal1 s 240 38460 240 38460 4 vdd
port 513 nsew
rlabel metal1 s 2256 38460 2256 38460 4 vdd
port 513 nsew
rlabel metal1 s 1488 40539 1488 40539 4 vdd
port 513 nsew
rlabel metal1 s 2256 38169 2256 38169 4 vdd
port 513 nsew
rlabel metal1 s 1488 39749 1488 39749 4 vdd
port 513 nsew
rlabel metal1 s 1488 40830 1488 40830 4 vdd
port 513 nsew
rlabel metal1 s 1488 39250 1488 39250 4 vdd
port 513 nsew
rlabel metal1 s 1008 39749 1008 39749 4 vdd
port 513 nsew
rlabel metal1 s 240 40830 240 40830 4 vdd
port 513 nsew
rlabel metal1 s 240 39250 240 39250 4 vdd
port 513 nsew
rlabel metal1 s 2256 40040 2256 40040 4 vdd
port 513 nsew
rlabel metal1 s 1488 40040 1488 40040 4 vdd
port 513 nsew
rlabel metal1 s 1008 40830 1008 40830 4 vdd
port 513 nsew
rlabel metal1 s 2256 39749 2256 39749 4 vdd
port 513 nsew
rlabel metal1 s 240 40539 240 40539 4 vdd
port 513 nsew
rlabel metal1 s 240 38169 240 38169 4 vdd
port 513 nsew
rlabel metal1 s 240 38959 240 38959 4 vdd
port 513 nsew
rlabel metal1 s 1008 38169 1008 38169 4 vdd
port 513 nsew
rlabel metal1 s 1488 38460 1488 38460 4 vdd
port 513 nsew
rlabel metal1 s 1488 38169 1488 38169 4 vdd
port 513 nsew
rlabel metal1 s 1008 40539 1008 40539 4 vdd
port 513 nsew
rlabel metal1 s 1008 38959 1008 38959 4 vdd
port 513 nsew
rlabel metal1 s 2256 38959 2256 38959 4 vdd
port 513 nsew
rlabel metal1 s 240 39749 240 39749 4 vdd
port 513 nsew
rlabel metal1 s 2256 40539 2256 40539 4 vdd
port 513 nsew
rlabel metal1 s 2256 39250 2256 39250 4 vdd
port 513 nsew
rlabel metal1 s 2256 40830 2256 40830 4 vdd
port 513 nsew
rlabel metal1 s 1008 39250 1008 39250 4 vdd
port 513 nsew
rlabel metal1 s 240 40040 240 40040 4 vdd
port 513 nsew
rlabel metal1 s 1008 38460 1008 38460 4 vdd
port 513 nsew
rlabel metal1 s 1488 38959 1488 38959 4 vdd
port 513 nsew
rlabel metal1 s 1008 40040 1008 40040 4 vdd
port 513 nsew
rlabel metal1 s 3504 39749 3504 39749 4 vdd
port 513 nsew
rlabel metal1 s 2736 39250 2736 39250 4 vdd
port 513 nsew
rlabel metal1 s 3984 39749 3984 39749 4 vdd
port 513 nsew
rlabel metal1 s 3984 38460 3984 38460 4 vdd
port 513 nsew
rlabel metal1 s 2736 39749 2736 39749 4 vdd
port 513 nsew
rlabel metal1 s 3984 40040 3984 40040 4 vdd
port 513 nsew
rlabel metal1 s 3504 40040 3504 40040 4 vdd
port 513 nsew
rlabel metal1 s 2736 40830 2736 40830 4 vdd
port 513 nsew
rlabel metal1 s 4752 40040 4752 40040 4 vdd
port 513 nsew
rlabel metal1 s 3984 40830 3984 40830 4 vdd
port 513 nsew
rlabel metal1 s 2736 40539 2736 40539 4 vdd
port 513 nsew
rlabel metal1 s 2736 38460 2736 38460 4 vdd
port 513 nsew
rlabel metal1 s 2736 40040 2736 40040 4 vdd
port 513 nsew
rlabel metal1 s 4752 39749 4752 39749 4 vdd
port 513 nsew
rlabel metal1 s 4752 38460 4752 38460 4 vdd
port 513 nsew
rlabel metal1 s 4752 38169 4752 38169 4 vdd
port 513 nsew
rlabel metal1 s 3984 38959 3984 38959 4 vdd
port 513 nsew
rlabel metal1 s 2736 38169 2736 38169 4 vdd
port 513 nsew
rlabel metal1 s 3504 38460 3504 38460 4 vdd
port 513 nsew
rlabel metal1 s 3504 38169 3504 38169 4 vdd
port 513 nsew
rlabel metal1 s 3504 40830 3504 40830 4 vdd
port 513 nsew
rlabel metal1 s 3504 39250 3504 39250 4 vdd
port 513 nsew
rlabel metal1 s 3504 38959 3504 38959 4 vdd
port 513 nsew
rlabel metal1 s 4752 39250 4752 39250 4 vdd
port 513 nsew
rlabel metal1 s 3984 39250 3984 39250 4 vdd
port 513 nsew
rlabel metal1 s 4752 38959 4752 38959 4 vdd
port 513 nsew
rlabel metal1 s 3984 38169 3984 38169 4 vdd
port 513 nsew
rlabel metal1 s 4752 40830 4752 40830 4 vdd
port 513 nsew
rlabel metal1 s 3984 40539 3984 40539 4 vdd
port 513 nsew
rlabel metal1 s 3504 40539 3504 40539 4 vdd
port 513 nsew
rlabel metal1 s 4752 40539 4752 40539 4 vdd
port 513 nsew
rlabel metal1 s 2736 38959 2736 38959 4 vdd
port 513 nsew
rlabel metal1 s 8976 41329 8976 41329 4 vdd
port 513 nsew
rlabel metal1 s 8496 42119 8496 42119 4 vdd
port 513 nsew
rlabel metal1 s 8976 42909 8976 42909 4 vdd
port 513 nsew
rlabel metal1 s 8976 43990 8976 43990 4 vdd
port 513 nsew
rlabel metal1 s 9744 43200 9744 43200 4 vdd
port 513 nsew
rlabel metal1 s 8976 42410 8976 42410 4 vdd
port 513 nsew
rlabel metal1 s 9744 43990 9744 43990 4 vdd
port 513 nsew
rlabel metal1 s 8976 42119 8976 42119 4 vdd
port 513 nsew
rlabel metal1 s 8976 43699 8976 43699 4 vdd
port 513 nsew
rlabel metal1 s 8496 42909 8496 42909 4 vdd
port 513 nsew
rlabel metal1 s 8976 43200 8976 43200 4 vdd
port 513 nsew
rlabel metal1 s 8496 43990 8496 43990 4 vdd
port 513 nsew
rlabel metal1 s 7728 41329 7728 41329 4 vdd
port 513 nsew
rlabel metal1 s 8496 41620 8496 41620 4 vdd
port 513 nsew
rlabel metal1 s 9744 43699 9744 43699 4 vdd
port 513 nsew
rlabel metal1 s 9744 41620 9744 41620 4 vdd
port 513 nsew
rlabel metal1 s 8976 41620 8976 41620 4 vdd
port 513 nsew
rlabel metal1 s 9744 42909 9744 42909 4 vdd
port 513 nsew
rlabel metal1 s 7728 42909 7728 42909 4 vdd
port 513 nsew
rlabel metal1 s 7728 41620 7728 41620 4 vdd
port 513 nsew
rlabel metal1 s 8496 43699 8496 43699 4 vdd
port 513 nsew
rlabel metal1 s 8496 41329 8496 41329 4 vdd
port 513 nsew
rlabel metal1 s 7728 43990 7728 43990 4 vdd
port 513 nsew
rlabel metal1 s 8496 42410 8496 42410 4 vdd
port 513 nsew
rlabel metal1 s 9744 42410 9744 42410 4 vdd
port 513 nsew
rlabel metal1 s 7728 43200 7728 43200 4 vdd
port 513 nsew
rlabel metal1 s 9744 41329 9744 41329 4 vdd
port 513 nsew
rlabel metal1 s 7728 42410 7728 42410 4 vdd
port 513 nsew
rlabel metal1 s 7728 42119 7728 42119 4 vdd
port 513 nsew
rlabel metal1 s 9744 42119 9744 42119 4 vdd
port 513 nsew
rlabel metal1 s 7728 43699 7728 43699 4 vdd
port 513 nsew
rlabel metal1 s 8496 43200 8496 43200 4 vdd
port 513 nsew
rlabel metal1 s 5232 41329 5232 41329 4 vdd
port 513 nsew
rlabel metal1 s 5232 42909 5232 42909 4 vdd
port 513 nsew
rlabel metal1 s 6480 41620 6480 41620 4 vdd
port 513 nsew
rlabel metal1 s 7248 42119 7248 42119 4 vdd
port 513 nsew
rlabel metal1 s 7248 43699 7248 43699 4 vdd
port 513 nsew
rlabel metal1 s 6000 41620 6000 41620 4 vdd
port 513 nsew
rlabel metal1 s 7248 42909 7248 42909 4 vdd
port 513 nsew
rlabel metal1 s 6000 43990 6000 43990 4 vdd
port 513 nsew
rlabel metal1 s 6480 43990 6480 43990 4 vdd
port 513 nsew
rlabel metal1 s 5232 43200 5232 43200 4 vdd
port 513 nsew
rlabel metal1 s 7248 43990 7248 43990 4 vdd
port 513 nsew
rlabel metal1 s 5232 43699 5232 43699 4 vdd
port 513 nsew
rlabel metal1 s 5232 42119 5232 42119 4 vdd
port 513 nsew
rlabel metal1 s 6480 42410 6480 42410 4 vdd
port 513 nsew
rlabel metal1 s 6480 43699 6480 43699 4 vdd
port 513 nsew
rlabel metal1 s 5232 41620 5232 41620 4 vdd
port 513 nsew
rlabel metal1 s 6000 42410 6000 42410 4 vdd
port 513 nsew
rlabel metal1 s 7248 41620 7248 41620 4 vdd
port 513 nsew
rlabel metal1 s 7248 43200 7248 43200 4 vdd
port 513 nsew
rlabel metal1 s 5232 43990 5232 43990 4 vdd
port 513 nsew
rlabel metal1 s 6480 42119 6480 42119 4 vdd
port 513 nsew
rlabel metal1 s 6480 41329 6480 41329 4 vdd
port 513 nsew
rlabel metal1 s 6480 42909 6480 42909 4 vdd
port 513 nsew
rlabel metal1 s 6000 43200 6000 43200 4 vdd
port 513 nsew
rlabel metal1 s 6000 42119 6000 42119 4 vdd
port 513 nsew
rlabel metal1 s 6000 42909 6000 42909 4 vdd
port 513 nsew
rlabel metal1 s 6000 43699 6000 43699 4 vdd
port 513 nsew
rlabel metal1 s 6000 41329 6000 41329 4 vdd
port 513 nsew
rlabel metal1 s 5232 42410 5232 42410 4 vdd
port 513 nsew
rlabel metal1 s 6480 43200 6480 43200 4 vdd
port 513 nsew
rlabel metal1 s 7248 42410 7248 42410 4 vdd
port 513 nsew
rlabel metal1 s 7248 41329 7248 41329 4 vdd
port 513 nsew
rlabel metal1 s 5232 39749 5232 39749 4 vdd
port 513 nsew
rlabel metal1 s 6480 38169 6480 38169 4 vdd
port 513 nsew
rlabel metal1 s 6000 40040 6000 40040 4 vdd
port 513 nsew
rlabel metal1 s 6000 40539 6000 40539 4 vdd
port 513 nsew
rlabel metal1 s 7248 40539 7248 40539 4 vdd
port 513 nsew
rlabel metal1 s 6000 38460 6000 38460 4 vdd
port 513 nsew
rlabel metal1 s 7248 38460 7248 38460 4 vdd
port 513 nsew
rlabel metal1 s 5232 39250 5232 39250 4 vdd
port 513 nsew
rlabel metal1 s 6480 38460 6480 38460 4 vdd
port 513 nsew
rlabel metal1 s 6000 40830 6000 40830 4 vdd
port 513 nsew
rlabel metal1 s 5232 40539 5232 40539 4 vdd
port 513 nsew
rlabel metal1 s 6480 38959 6480 38959 4 vdd
port 513 nsew
rlabel metal1 s 6480 40830 6480 40830 4 vdd
port 513 nsew
rlabel metal1 s 6480 40539 6480 40539 4 vdd
port 513 nsew
rlabel metal1 s 6000 39749 6000 39749 4 vdd
port 513 nsew
rlabel metal1 s 5232 38169 5232 38169 4 vdd
port 513 nsew
rlabel metal1 s 7248 38169 7248 38169 4 vdd
port 513 nsew
rlabel metal1 s 6000 38169 6000 38169 4 vdd
port 513 nsew
rlabel metal1 s 7248 39749 7248 39749 4 vdd
port 513 nsew
rlabel metal1 s 7248 40830 7248 40830 4 vdd
port 513 nsew
rlabel metal1 s 6000 38959 6000 38959 4 vdd
port 513 nsew
rlabel metal1 s 5232 38460 5232 38460 4 vdd
port 513 nsew
rlabel metal1 s 7248 39250 7248 39250 4 vdd
port 513 nsew
rlabel metal1 s 6480 39250 6480 39250 4 vdd
port 513 nsew
rlabel metal1 s 5232 40830 5232 40830 4 vdd
port 513 nsew
rlabel metal1 s 5232 38959 5232 38959 4 vdd
port 513 nsew
rlabel metal1 s 7248 40040 7248 40040 4 vdd
port 513 nsew
rlabel metal1 s 6480 40040 6480 40040 4 vdd
port 513 nsew
rlabel metal1 s 7248 38959 7248 38959 4 vdd
port 513 nsew
rlabel metal1 s 6000 39250 6000 39250 4 vdd
port 513 nsew
rlabel metal1 s 5232 40040 5232 40040 4 vdd
port 513 nsew
rlabel metal1 s 6480 39749 6480 39749 4 vdd
port 513 nsew
rlabel metal1 s 7728 38959 7728 38959 4 vdd
port 513 nsew
rlabel metal1 s 8976 39749 8976 39749 4 vdd
port 513 nsew
rlabel metal1 s 7728 38169 7728 38169 4 vdd
port 513 nsew
rlabel metal1 s 8496 38169 8496 38169 4 vdd
port 513 nsew
rlabel metal1 s 8976 38959 8976 38959 4 vdd
port 513 nsew
rlabel metal1 s 8496 39250 8496 39250 4 vdd
port 513 nsew
rlabel metal1 s 8976 38460 8976 38460 4 vdd
port 513 nsew
rlabel metal1 s 9744 38959 9744 38959 4 vdd
port 513 nsew
rlabel metal1 s 7728 40539 7728 40539 4 vdd
port 513 nsew
rlabel metal1 s 8496 38460 8496 38460 4 vdd
port 513 nsew
rlabel metal1 s 7728 40830 7728 40830 4 vdd
port 513 nsew
rlabel metal1 s 7728 38460 7728 38460 4 vdd
port 513 nsew
rlabel metal1 s 9744 39749 9744 39749 4 vdd
port 513 nsew
rlabel metal1 s 8976 38169 8976 38169 4 vdd
port 513 nsew
rlabel metal1 s 8976 40539 8976 40539 4 vdd
port 513 nsew
rlabel metal1 s 8496 38959 8496 38959 4 vdd
port 513 nsew
rlabel metal1 s 7728 39749 7728 39749 4 vdd
port 513 nsew
rlabel metal1 s 8976 40830 8976 40830 4 vdd
port 513 nsew
rlabel metal1 s 9744 40830 9744 40830 4 vdd
port 513 nsew
rlabel metal1 s 8496 40830 8496 40830 4 vdd
port 513 nsew
rlabel metal1 s 8496 39749 8496 39749 4 vdd
port 513 nsew
rlabel metal1 s 7728 39250 7728 39250 4 vdd
port 513 nsew
rlabel metal1 s 7728 40040 7728 40040 4 vdd
port 513 nsew
rlabel metal1 s 8976 39250 8976 39250 4 vdd
port 513 nsew
rlabel metal1 s 9744 40040 9744 40040 4 vdd
port 513 nsew
rlabel metal1 s 8976 40040 8976 40040 4 vdd
port 513 nsew
rlabel metal1 s 8496 40539 8496 40539 4 vdd
port 513 nsew
rlabel metal1 s 9744 39250 9744 39250 4 vdd
port 513 nsew
rlabel metal1 s 9744 38169 9744 38169 4 vdd
port 513 nsew
rlabel metal1 s 9744 40539 9744 40539 4 vdd
port 513 nsew
rlabel metal1 s 9744 38460 9744 38460 4 vdd
port 513 nsew
rlabel metal1 s 8496 40040 8496 40040 4 vdd
port 513 nsew
rlabel metal1 s 7728 35009 7728 35009 4 vdd
port 513 nsew
rlabel metal1 s 9744 35799 9744 35799 4 vdd
port 513 nsew
rlabel metal1 s 9744 36589 9744 36589 4 vdd
port 513 nsew
rlabel metal1 s 8496 36090 8496 36090 4 vdd
port 513 nsew
rlabel metal1 s 9744 37379 9744 37379 4 vdd
port 513 nsew
rlabel metal1 s 7728 36880 7728 36880 4 vdd
port 513 nsew
rlabel metal1 s 8976 37670 8976 37670 4 vdd
port 513 nsew
rlabel metal1 s 7728 35799 7728 35799 4 vdd
port 513 nsew
rlabel metal1 s 8976 37379 8976 37379 4 vdd
port 513 nsew
rlabel metal1 s 9744 36090 9744 36090 4 vdd
port 513 nsew
rlabel metal1 s 8496 35799 8496 35799 4 vdd
port 513 nsew
rlabel metal1 s 7728 35300 7728 35300 4 vdd
port 513 nsew
rlabel metal1 s 8496 36880 8496 36880 4 vdd
port 513 nsew
rlabel metal1 s 7728 37379 7728 37379 4 vdd
port 513 nsew
rlabel metal1 s 8976 36880 8976 36880 4 vdd
port 513 nsew
rlabel metal1 s 8976 35009 8976 35009 4 vdd
port 513 nsew
rlabel metal1 s 8976 36090 8976 36090 4 vdd
port 513 nsew
rlabel metal1 s 7728 36090 7728 36090 4 vdd
port 513 nsew
rlabel metal1 s 8976 35300 8976 35300 4 vdd
port 513 nsew
rlabel metal1 s 9744 35009 9744 35009 4 vdd
port 513 nsew
rlabel metal1 s 7728 36589 7728 36589 4 vdd
port 513 nsew
rlabel metal1 s 8496 35009 8496 35009 4 vdd
port 513 nsew
rlabel metal1 s 9744 37670 9744 37670 4 vdd
port 513 nsew
rlabel metal1 s 8496 37379 8496 37379 4 vdd
port 513 nsew
rlabel metal1 s 8976 35799 8976 35799 4 vdd
port 513 nsew
rlabel metal1 s 9744 35300 9744 35300 4 vdd
port 513 nsew
rlabel metal1 s 8976 36589 8976 36589 4 vdd
port 513 nsew
rlabel metal1 s 7728 37670 7728 37670 4 vdd
port 513 nsew
rlabel metal1 s 8496 37670 8496 37670 4 vdd
port 513 nsew
rlabel metal1 s 8496 36589 8496 36589 4 vdd
port 513 nsew
rlabel metal1 s 9744 36880 9744 36880 4 vdd
port 513 nsew
rlabel metal1 s 8496 35300 8496 35300 4 vdd
port 513 nsew
rlabel metal1 s 5232 37670 5232 37670 4 vdd
port 513 nsew
rlabel metal1 s 6480 36589 6480 36589 4 vdd
port 513 nsew
rlabel metal1 s 6480 35009 6480 35009 4 vdd
port 513 nsew
rlabel metal1 s 6000 36880 6000 36880 4 vdd
port 513 nsew
rlabel metal1 s 5232 37379 5232 37379 4 vdd
port 513 nsew
rlabel metal1 s 6000 35300 6000 35300 4 vdd
port 513 nsew
rlabel metal1 s 7248 35300 7248 35300 4 vdd
port 513 nsew
rlabel metal1 s 6000 35009 6000 35009 4 vdd
port 513 nsew
rlabel metal1 s 6000 37379 6000 37379 4 vdd
port 513 nsew
rlabel metal1 s 6480 37379 6480 37379 4 vdd
port 513 nsew
rlabel metal1 s 6000 37670 6000 37670 4 vdd
port 513 nsew
rlabel metal1 s 6480 37670 6480 37670 4 vdd
port 513 nsew
rlabel metal1 s 6000 35799 6000 35799 4 vdd
port 513 nsew
rlabel metal1 s 7248 36589 7248 36589 4 vdd
port 513 nsew
rlabel metal1 s 7248 37379 7248 37379 4 vdd
port 513 nsew
rlabel metal1 s 7248 35799 7248 35799 4 vdd
port 513 nsew
rlabel metal1 s 5232 36090 5232 36090 4 vdd
port 513 nsew
rlabel metal1 s 7248 36090 7248 36090 4 vdd
port 513 nsew
rlabel metal1 s 7248 35009 7248 35009 4 vdd
port 513 nsew
rlabel metal1 s 5232 35009 5232 35009 4 vdd
port 513 nsew
rlabel metal1 s 6480 36090 6480 36090 4 vdd
port 513 nsew
rlabel metal1 s 5232 35799 5232 35799 4 vdd
port 513 nsew
rlabel metal1 s 5232 36589 5232 36589 4 vdd
port 513 nsew
rlabel metal1 s 6480 35799 6480 35799 4 vdd
port 513 nsew
rlabel metal1 s 5232 35300 5232 35300 4 vdd
port 513 nsew
rlabel metal1 s 5232 36880 5232 36880 4 vdd
port 513 nsew
rlabel metal1 s 6000 36589 6000 36589 4 vdd
port 513 nsew
rlabel metal1 s 7248 37670 7248 37670 4 vdd
port 513 nsew
rlabel metal1 s 6000 36090 6000 36090 4 vdd
port 513 nsew
rlabel metal1 s 7248 36880 7248 36880 4 vdd
port 513 nsew
rlabel metal1 s 6480 35300 6480 35300 4 vdd
port 513 nsew
rlabel metal1 s 6480 36880 6480 36880 4 vdd
port 513 nsew
rlabel metal1 s 7248 34510 7248 34510 4 vdd
port 513 nsew
rlabel metal1 s 6000 33720 6000 33720 4 vdd
port 513 nsew
rlabel metal1 s 7248 32140 7248 32140 4 vdd
port 513 nsew
rlabel metal1 s 6480 34219 6480 34219 4 vdd
port 513 nsew
rlabel metal1 s 6480 32930 6480 32930 4 vdd
port 513 nsew
rlabel metal1 s 6000 31849 6000 31849 4 vdd
port 513 nsew
rlabel metal1 s 7248 34219 7248 34219 4 vdd
port 513 nsew
rlabel metal1 s 5232 32930 5232 32930 4 vdd
port 513 nsew
rlabel metal1 s 6000 32639 6000 32639 4 vdd
port 513 nsew
rlabel metal1 s 7248 31849 7248 31849 4 vdd
port 513 nsew
rlabel metal1 s 7248 33429 7248 33429 4 vdd
port 513 nsew
rlabel metal1 s 5232 33720 5232 33720 4 vdd
port 513 nsew
rlabel metal1 s 6480 32140 6480 32140 4 vdd
port 513 nsew
rlabel metal1 s 5232 34510 5232 34510 4 vdd
port 513 nsew
rlabel metal1 s 5232 32140 5232 32140 4 vdd
port 513 nsew
rlabel metal1 s 6480 33720 6480 33720 4 vdd
port 513 nsew
rlabel metal1 s 6480 34510 6480 34510 4 vdd
port 513 nsew
rlabel metal1 s 7248 32930 7248 32930 4 vdd
port 513 nsew
rlabel metal1 s 6480 31849 6480 31849 4 vdd
port 513 nsew
rlabel metal1 s 5232 33429 5232 33429 4 vdd
port 513 nsew
rlabel metal1 s 5232 31849 5232 31849 4 vdd
port 513 nsew
rlabel metal1 s 5232 32639 5232 32639 4 vdd
port 513 nsew
rlabel metal1 s 6480 33429 6480 33429 4 vdd
port 513 nsew
rlabel metal1 s 6000 33429 6000 33429 4 vdd
port 513 nsew
rlabel metal1 s 7248 33720 7248 33720 4 vdd
port 513 nsew
rlabel metal1 s 6000 34510 6000 34510 4 vdd
port 513 nsew
rlabel metal1 s 6000 32140 6000 32140 4 vdd
port 513 nsew
rlabel metal1 s 6000 34219 6000 34219 4 vdd
port 513 nsew
rlabel metal1 s 7248 32639 7248 32639 4 vdd
port 513 nsew
rlabel metal1 s 5232 34219 5232 34219 4 vdd
port 513 nsew
rlabel metal1 s 6480 32639 6480 32639 4 vdd
port 513 nsew
rlabel metal1 s 6000 32930 6000 32930 4 vdd
port 513 nsew
rlabel metal1 s 8976 34219 8976 34219 4 vdd
port 513 nsew
rlabel metal1 s 9744 33720 9744 33720 4 vdd
port 513 nsew
rlabel metal1 s 8976 32639 8976 32639 4 vdd
port 513 nsew
rlabel metal1 s 8976 33720 8976 33720 4 vdd
port 513 nsew
rlabel metal1 s 8496 34510 8496 34510 4 vdd
port 513 nsew
rlabel metal1 s 7728 31849 7728 31849 4 vdd
port 513 nsew
rlabel metal1 s 7728 32930 7728 32930 4 vdd
port 513 nsew
rlabel metal1 s 8496 33429 8496 33429 4 vdd
port 513 nsew
rlabel metal1 s 7728 32140 7728 32140 4 vdd
port 513 nsew
rlabel metal1 s 8496 33720 8496 33720 4 vdd
port 513 nsew
rlabel metal1 s 7728 34219 7728 34219 4 vdd
port 513 nsew
rlabel metal1 s 8976 32930 8976 32930 4 vdd
port 513 nsew
rlabel metal1 s 9744 32140 9744 32140 4 vdd
port 513 nsew
rlabel metal1 s 9744 32639 9744 32639 4 vdd
port 513 nsew
rlabel metal1 s 8496 32140 8496 32140 4 vdd
port 513 nsew
rlabel metal1 s 7728 33429 7728 33429 4 vdd
port 513 nsew
rlabel metal1 s 9744 33429 9744 33429 4 vdd
port 513 nsew
rlabel metal1 s 8496 32930 8496 32930 4 vdd
port 513 nsew
rlabel metal1 s 7728 33720 7728 33720 4 vdd
port 513 nsew
rlabel metal1 s 8496 34219 8496 34219 4 vdd
port 513 nsew
rlabel metal1 s 9744 34219 9744 34219 4 vdd
port 513 nsew
rlabel metal1 s 8496 31849 8496 31849 4 vdd
port 513 nsew
rlabel metal1 s 7728 32639 7728 32639 4 vdd
port 513 nsew
rlabel metal1 s 8976 31849 8976 31849 4 vdd
port 513 nsew
rlabel metal1 s 9744 31849 9744 31849 4 vdd
port 513 nsew
rlabel metal1 s 8976 33429 8976 33429 4 vdd
port 513 nsew
rlabel metal1 s 9744 32930 9744 32930 4 vdd
port 513 nsew
rlabel metal1 s 7728 34510 7728 34510 4 vdd
port 513 nsew
rlabel metal1 s 8976 34510 8976 34510 4 vdd
port 513 nsew
rlabel metal1 s 8496 32639 8496 32639 4 vdd
port 513 nsew
rlabel metal1 s 9744 34510 9744 34510 4 vdd
port 513 nsew
rlabel metal1 s 8976 32140 8976 32140 4 vdd
port 513 nsew
rlabel metal1 s 3504 36090 3504 36090 4 vdd
port 513 nsew
rlabel metal1 s 2736 35799 2736 35799 4 vdd
port 513 nsew
rlabel metal1 s 3984 35799 3984 35799 4 vdd
port 513 nsew
rlabel metal1 s 2736 35300 2736 35300 4 vdd
port 513 nsew
rlabel metal1 s 4752 35300 4752 35300 4 vdd
port 513 nsew
rlabel metal1 s 4752 36589 4752 36589 4 vdd
port 513 nsew
rlabel metal1 s 2736 37670 2736 37670 4 vdd
port 513 nsew
rlabel metal1 s 2736 35009 2736 35009 4 vdd
port 513 nsew
rlabel metal1 s 3504 37379 3504 37379 4 vdd
port 513 nsew
rlabel metal1 s 3984 36589 3984 36589 4 vdd
port 513 nsew
rlabel metal1 s 2736 37379 2736 37379 4 vdd
port 513 nsew
rlabel metal1 s 3984 36880 3984 36880 4 vdd
port 513 nsew
rlabel metal1 s 2736 36589 2736 36589 4 vdd
port 513 nsew
rlabel metal1 s 3984 37379 3984 37379 4 vdd
port 513 nsew
rlabel metal1 s 3504 35799 3504 35799 4 vdd
port 513 nsew
rlabel metal1 s 3504 36880 3504 36880 4 vdd
port 513 nsew
rlabel metal1 s 3504 37670 3504 37670 4 vdd
port 513 nsew
rlabel metal1 s 3504 36589 3504 36589 4 vdd
port 513 nsew
rlabel metal1 s 3984 35300 3984 35300 4 vdd
port 513 nsew
rlabel metal1 s 3984 36090 3984 36090 4 vdd
port 513 nsew
rlabel metal1 s 3984 37670 3984 37670 4 vdd
port 513 nsew
rlabel metal1 s 3504 35009 3504 35009 4 vdd
port 513 nsew
rlabel metal1 s 4752 35799 4752 35799 4 vdd
port 513 nsew
rlabel metal1 s 4752 35009 4752 35009 4 vdd
port 513 nsew
rlabel metal1 s 3504 35300 3504 35300 4 vdd
port 513 nsew
rlabel metal1 s 3984 35009 3984 35009 4 vdd
port 513 nsew
rlabel metal1 s 4752 37670 4752 37670 4 vdd
port 513 nsew
rlabel metal1 s 4752 36090 4752 36090 4 vdd
port 513 nsew
rlabel metal1 s 2736 36880 2736 36880 4 vdd
port 513 nsew
rlabel metal1 s 2736 36090 2736 36090 4 vdd
port 513 nsew
rlabel metal1 s 4752 37379 4752 37379 4 vdd
port 513 nsew
rlabel metal1 s 4752 36880 4752 36880 4 vdd
port 513 nsew
rlabel metal1 s 240 35009 240 35009 4 vdd
port 513 nsew
rlabel metal1 s 2256 37670 2256 37670 4 vdd
port 513 nsew
rlabel metal1 s 1008 36589 1008 36589 4 vdd
port 513 nsew
rlabel metal1 s 2256 35300 2256 35300 4 vdd
port 513 nsew
rlabel metal1 s 1488 36880 1488 36880 4 vdd
port 513 nsew
rlabel metal1 s 240 36090 240 36090 4 vdd
port 513 nsew
rlabel metal1 s 1008 36880 1008 36880 4 vdd
port 513 nsew
rlabel metal1 s 240 37379 240 37379 4 vdd
port 513 nsew
rlabel metal1 s 2256 37379 2256 37379 4 vdd
port 513 nsew
rlabel metal1 s 1488 35009 1488 35009 4 vdd
port 513 nsew
rlabel metal1 s 1488 35799 1488 35799 4 vdd
port 513 nsew
rlabel metal1 s 1008 35799 1008 35799 4 vdd
port 513 nsew
rlabel metal1 s 1008 35300 1008 35300 4 vdd
port 513 nsew
rlabel metal1 s 240 36880 240 36880 4 vdd
port 513 nsew
rlabel metal1 s 240 36589 240 36589 4 vdd
port 513 nsew
rlabel metal1 s 240 35799 240 35799 4 vdd
port 513 nsew
rlabel metal1 s 2256 36090 2256 36090 4 vdd
port 513 nsew
rlabel metal1 s 2256 36880 2256 36880 4 vdd
port 513 nsew
rlabel metal1 s 240 37670 240 37670 4 vdd
port 513 nsew
rlabel metal1 s 1008 36090 1008 36090 4 vdd
port 513 nsew
rlabel metal1 s 2256 35799 2256 35799 4 vdd
port 513 nsew
rlabel metal1 s 1488 37379 1488 37379 4 vdd
port 513 nsew
rlabel metal1 s 1488 36589 1488 36589 4 vdd
port 513 nsew
rlabel metal1 s 1008 37379 1008 37379 4 vdd
port 513 nsew
rlabel metal1 s 1008 37670 1008 37670 4 vdd
port 513 nsew
rlabel metal1 s 1488 36090 1488 36090 4 vdd
port 513 nsew
rlabel metal1 s 2256 36589 2256 36589 4 vdd
port 513 nsew
rlabel metal1 s 1008 35009 1008 35009 4 vdd
port 513 nsew
rlabel metal1 s 2256 35009 2256 35009 4 vdd
port 513 nsew
rlabel metal1 s 240 35300 240 35300 4 vdd
port 513 nsew
rlabel metal1 s 1488 37670 1488 37670 4 vdd
port 513 nsew
rlabel metal1 s 1488 35300 1488 35300 4 vdd
port 513 nsew
rlabel metal1 s 240 33720 240 33720 4 vdd
port 513 nsew
rlabel metal1 s 2256 32639 2256 32639 4 vdd
port 513 nsew
rlabel metal1 s 1488 32639 1488 32639 4 vdd
port 513 nsew
rlabel metal1 s 1488 34219 1488 34219 4 vdd
port 513 nsew
rlabel metal1 s 2256 31849 2256 31849 4 vdd
port 513 nsew
rlabel metal1 s 2256 32930 2256 32930 4 vdd
port 513 nsew
rlabel metal1 s 1008 32930 1008 32930 4 vdd
port 513 nsew
rlabel metal1 s 2256 34510 2256 34510 4 vdd
port 513 nsew
rlabel metal1 s 1008 34219 1008 34219 4 vdd
port 513 nsew
rlabel metal1 s 2256 33720 2256 33720 4 vdd
port 513 nsew
rlabel metal1 s 2256 34219 2256 34219 4 vdd
port 513 nsew
rlabel metal1 s 2256 32140 2256 32140 4 vdd
port 513 nsew
rlabel metal1 s 1488 32140 1488 32140 4 vdd
port 513 nsew
rlabel metal1 s 240 34510 240 34510 4 vdd
port 513 nsew
rlabel metal1 s 1488 33429 1488 33429 4 vdd
port 513 nsew
rlabel metal1 s 1488 31849 1488 31849 4 vdd
port 513 nsew
rlabel metal1 s 1008 32140 1008 32140 4 vdd
port 513 nsew
rlabel metal1 s 1488 32930 1488 32930 4 vdd
port 513 nsew
rlabel metal1 s 240 34219 240 34219 4 vdd
port 513 nsew
rlabel metal1 s 1488 34510 1488 34510 4 vdd
port 513 nsew
rlabel metal1 s 1008 31849 1008 31849 4 vdd
port 513 nsew
rlabel metal1 s 240 31849 240 31849 4 vdd
port 513 nsew
rlabel metal1 s 1008 33429 1008 33429 4 vdd
port 513 nsew
rlabel metal1 s 1008 34510 1008 34510 4 vdd
port 513 nsew
rlabel metal1 s 240 33429 240 33429 4 vdd
port 513 nsew
rlabel metal1 s 1008 33720 1008 33720 4 vdd
port 513 nsew
rlabel metal1 s 2256 33429 2256 33429 4 vdd
port 513 nsew
rlabel metal1 s 240 32639 240 32639 4 vdd
port 513 nsew
rlabel metal1 s 1488 33720 1488 33720 4 vdd
port 513 nsew
rlabel metal1 s 240 32140 240 32140 4 vdd
port 513 nsew
rlabel metal1 s 1008 32639 1008 32639 4 vdd
port 513 nsew
rlabel metal1 s 240 32930 240 32930 4 vdd
port 513 nsew
rlabel metal1 s 4752 32930 4752 32930 4 vdd
port 513 nsew
rlabel metal1 s 3984 31849 3984 31849 4 vdd
port 513 nsew
rlabel metal1 s 4752 33429 4752 33429 4 vdd
port 513 nsew
rlabel metal1 s 4752 34219 4752 34219 4 vdd
port 513 nsew
rlabel metal1 s 4752 31849 4752 31849 4 vdd
port 513 nsew
rlabel metal1 s 3984 34510 3984 34510 4 vdd
port 513 nsew
rlabel metal1 s 2736 32639 2736 32639 4 vdd
port 513 nsew
rlabel metal1 s 3504 34219 3504 34219 4 vdd
port 513 nsew
rlabel metal1 s 2736 33720 2736 33720 4 vdd
port 513 nsew
rlabel metal1 s 3984 33720 3984 33720 4 vdd
port 513 nsew
rlabel metal1 s 3984 32140 3984 32140 4 vdd
port 513 nsew
rlabel metal1 s 3504 33720 3504 33720 4 vdd
port 513 nsew
rlabel metal1 s 3984 32639 3984 32639 4 vdd
port 513 nsew
rlabel metal1 s 4752 34510 4752 34510 4 vdd
port 513 nsew
rlabel metal1 s 2736 32930 2736 32930 4 vdd
port 513 nsew
rlabel metal1 s 2736 32140 2736 32140 4 vdd
port 513 nsew
rlabel metal1 s 2736 33429 2736 33429 4 vdd
port 513 nsew
rlabel metal1 s 3504 32639 3504 32639 4 vdd
port 513 nsew
rlabel metal1 s 4752 33720 4752 33720 4 vdd
port 513 nsew
rlabel metal1 s 3984 32930 3984 32930 4 vdd
port 513 nsew
rlabel metal1 s 3504 33429 3504 33429 4 vdd
port 513 nsew
rlabel metal1 s 3504 32930 3504 32930 4 vdd
port 513 nsew
rlabel metal1 s 4752 32140 4752 32140 4 vdd
port 513 nsew
rlabel metal1 s 3504 34510 3504 34510 4 vdd
port 513 nsew
rlabel metal1 s 2736 31849 2736 31849 4 vdd
port 513 nsew
rlabel metal1 s 2736 34219 2736 34219 4 vdd
port 513 nsew
rlabel metal1 s 3984 33429 3984 33429 4 vdd
port 513 nsew
rlabel metal1 s 3984 34219 3984 34219 4 vdd
port 513 nsew
rlabel metal1 s 3504 32140 3504 32140 4 vdd
port 513 nsew
rlabel metal1 s 2736 34510 2736 34510 4 vdd
port 513 nsew
rlabel metal1 s 3504 31849 3504 31849 4 vdd
port 513 nsew
rlabel metal1 s 4752 32639 4752 32639 4 vdd
port 513 nsew
rlabel metal1 s 3504 30560 3504 30560 4 vdd
port 513 nsew
rlabel metal1 s 3504 29770 3504 29770 4 vdd
port 513 nsew
rlabel metal1 s 4752 31059 4752 31059 4 vdd
port 513 nsew
rlabel metal1 s 4752 31350 4752 31350 4 vdd
port 513 nsew
rlabel metal1 s 3504 31059 3504 31059 4 vdd
port 513 nsew
rlabel metal1 s 2736 29770 2736 29770 4 vdd
port 513 nsew
rlabel metal1 s 4752 28980 4752 28980 4 vdd
port 513 nsew
rlabel metal1 s 2736 29479 2736 29479 4 vdd
port 513 nsew
rlabel metal1 s 4752 30269 4752 30269 4 vdd
port 513 nsew
rlabel metal1 s 3984 29479 3984 29479 4 vdd
port 513 nsew
rlabel metal1 s 4752 30560 4752 30560 4 vdd
port 513 nsew
rlabel metal1 s 2736 30269 2736 30269 4 vdd
port 513 nsew
rlabel metal1 s 2736 31059 2736 31059 4 vdd
port 513 nsew
rlabel metal1 s 3984 28689 3984 28689 4 vdd
port 513 nsew
rlabel metal1 s 3504 28980 3504 28980 4 vdd
port 513 nsew
rlabel metal1 s 3504 28689 3504 28689 4 vdd
port 513 nsew
rlabel metal1 s 4752 29479 4752 29479 4 vdd
port 513 nsew
rlabel metal1 s 2736 31350 2736 31350 4 vdd
port 513 nsew
rlabel metal1 s 4752 29770 4752 29770 4 vdd
port 513 nsew
rlabel metal1 s 3984 28980 3984 28980 4 vdd
port 513 nsew
rlabel metal1 s 4752 28689 4752 28689 4 vdd
port 513 nsew
rlabel metal1 s 2736 28980 2736 28980 4 vdd
port 513 nsew
rlabel metal1 s 3504 30269 3504 30269 4 vdd
port 513 nsew
rlabel metal1 s 3984 29770 3984 29770 4 vdd
port 513 nsew
rlabel metal1 s 2736 30560 2736 30560 4 vdd
port 513 nsew
rlabel metal1 s 3984 30560 3984 30560 4 vdd
port 513 nsew
rlabel metal1 s 3984 31059 3984 31059 4 vdd
port 513 nsew
rlabel metal1 s 3984 30269 3984 30269 4 vdd
port 513 nsew
rlabel metal1 s 3984 31350 3984 31350 4 vdd
port 513 nsew
rlabel metal1 s 3504 31350 3504 31350 4 vdd
port 513 nsew
rlabel metal1 s 2736 28689 2736 28689 4 vdd
port 513 nsew
rlabel metal1 s 3504 29479 3504 29479 4 vdd
port 513 nsew
rlabel metal1 s 1008 28980 1008 28980 4 vdd
port 513 nsew
rlabel metal1 s 240 30269 240 30269 4 vdd
port 513 nsew
rlabel metal1 s 1488 29479 1488 29479 4 vdd
port 513 nsew
rlabel metal1 s 240 29770 240 29770 4 vdd
port 513 nsew
rlabel metal1 s 2256 30269 2256 30269 4 vdd
port 513 nsew
rlabel metal1 s 1008 30560 1008 30560 4 vdd
port 513 nsew
rlabel metal1 s 240 31059 240 31059 4 vdd
port 513 nsew
rlabel metal1 s 1008 31059 1008 31059 4 vdd
port 513 nsew
rlabel metal1 s 2256 29479 2256 29479 4 vdd
port 513 nsew
rlabel metal1 s 1488 31350 1488 31350 4 vdd
port 513 nsew
rlabel metal1 s 240 28689 240 28689 4 vdd
port 513 nsew
rlabel metal1 s 2256 31059 2256 31059 4 vdd
port 513 nsew
rlabel metal1 s 1488 30560 1488 30560 4 vdd
port 513 nsew
rlabel metal1 s 240 31350 240 31350 4 vdd
port 513 nsew
rlabel metal1 s 1488 30269 1488 30269 4 vdd
port 513 nsew
rlabel metal1 s 1488 29770 1488 29770 4 vdd
port 513 nsew
rlabel metal1 s 1488 28980 1488 28980 4 vdd
port 513 nsew
rlabel metal1 s 1488 28689 1488 28689 4 vdd
port 513 nsew
rlabel metal1 s 1008 28689 1008 28689 4 vdd
port 513 nsew
rlabel metal1 s 1008 29770 1008 29770 4 vdd
port 513 nsew
rlabel metal1 s 2256 28980 2256 28980 4 vdd
port 513 nsew
rlabel metal1 s 1008 31350 1008 31350 4 vdd
port 513 nsew
rlabel metal1 s 2256 31350 2256 31350 4 vdd
port 513 nsew
rlabel metal1 s 2256 28689 2256 28689 4 vdd
port 513 nsew
rlabel metal1 s 1008 29479 1008 29479 4 vdd
port 513 nsew
rlabel metal1 s 240 30560 240 30560 4 vdd
port 513 nsew
rlabel metal1 s 1488 31059 1488 31059 4 vdd
port 513 nsew
rlabel metal1 s 2256 30560 2256 30560 4 vdd
port 513 nsew
rlabel metal1 s 240 29479 240 29479 4 vdd
port 513 nsew
rlabel metal1 s 1008 30269 1008 30269 4 vdd
port 513 nsew
rlabel metal1 s 2256 29770 2256 29770 4 vdd
port 513 nsew
rlabel metal1 s 240 28980 240 28980 4 vdd
port 513 nsew
rlabel metal1 s 240 26610 240 26610 4 vdd
port 513 nsew
rlabel metal1 s 2256 28190 2256 28190 4 vdd
port 513 nsew
rlabel metal1 s 240 28190 240 28190 4 vdd
port 513 nsew
rlabel metal1 s 2256 27109 2256 27109 4 vdd
port 513 nsew
rlabel metal1 s 240 25820 240 25820 4 vdd
port 513 nsew
rlabel metal1 s 1488 28190 1488 28190 4 vdd
port 513 nsew
rlabel metal1 s 240 27899 240 27899 4 vdd
port 513 nsew
rlabel metal1 s 1488 26610 1488 26610 4 vdd
port 513 nsew
rlabel metal1 s 1488 27400 1488 27400 4 vdd
port 513 nsew
rlabel metal1 s 240 27109 240 27109 4 vdd
port 513 nsew
rlabel metal1 s 2256 25820 2256 25820 4 vdd
port 513 nsew
rlabel metal1 s 1488 26319 1488 26319 4 vdd
port 513 nsew
rlabel metal1 s 1008 28190 1008 28190 4 vdd
port 513 nsew
rlabel metal1 s 2256 27400 2256 27400 4 vdd
port 513 nsew
rlabel metal1 s 2256 26610 2256 26610 4 vdd
port 513 nsew
rlabel metal1 s 1008 27109 1008 27109 4 vdd
port 513 nsew
rlabel metal1 s 1008 26610 1008 26610 4 vdd
port 513 nsew
rlabel metal1 s 1488 27899 1488 27899 4 vdd
port 513 nsew
rlabel metal1 s 1008 25529 1008 25529 4 vdd
port 513 nsew
rlabel metal1 s 2256 26319 2256 26319 4 vdd
port 513 nsew
rlabel metal1 s 1008 27400 1008 27400 4 vdd
port 513 nsew
rlabel metal1 s 2256 25529 2256 25529 4 vdd
port 513 nsew
rlabel metal1 s 1008 25820 1008 25820 4 vdd
port 513 nsew
rlabel metal1 s 1008 26319 1008 26319 4 vdd
port 513 nsew
rlabel metal1 s 240 27400 240 27400 4 vdd
port 513 nsew
rlabel metal1 s 240 25529 240 25529 4 vdd
port 513 nsew
rlabel metal1 s 1488 25820 1488 25820 4 vdd
port 513 nsew
rlabel metal1 s 2256 27899 2256 27899 4 vdd
port 513 nsew
rlabel metal1 s 1008 27899 1008 27899 4 vdd
port 513 nsew
rlabel metal1 s 240 26319 240 26319 4 vdd
port 513 nsew
rlabel metal1 s 1488 27109 1488 27109 4 vdd
port 513 nsew
rlabel metal1 s 1488 25529 1488 25529 4 vdd
port 513 nsew
rlabel metal1 s 3504 25820 3504 25820 4 vdd
port 513 nsew
rlabel metal1 s 2736 26610 2736 26610 4 vdd
port 513 nsew
rlabel metal1 s 2736 25820 2736 25820 4 vdd
port 513 nsew
rlabel metal1 s 3504 25529 3504 25529 4 vdd
port 513 nsew
rlabel metal1 s 2736 27400 2736 27400 4 vdd
port 513 nsew
rlabel metal1 s 3984 28190 3984 28190 4 vdd
port 513 nsew
rlabel metal1 s 4752 27400 4752 27400 4 vdd
port 513 nsew
rlabel metal1 s 4752 26610 4752 26610 4 vdd
port 513 nsew
rlabel metal1 s 3984 27400 3984 27400 4 vdd
port 513 nsew
rlabel metal1 s 4752 26319 4752 26319 4 vdd
port 513 nsew
rlabel metal1 s 3504 26319 3504 26319 4 vdd
port 513 nsew
rlabel metal1 s 4752 27899 4752 27899 4 vdd
port 513 nsew
rlabel metal1 s 3984 27109 3984 27109 4 vdd
port 513 nsew
rlabel metal1 s 4752 27109 4752 27109 4 vdd
port 513 nsew
rlabel metal1 s 3504 27899 3504 27899 4 vdd
port 513 nsew
rlabel metal1 s 3504 27109 3504 27109 4 vdd
port 513 nsew
rlabel metal1 s 2736 28190 2736 28190 4 vdd
port 513 nsew
rlabel metal1 s 3984 25529 3984 25529 4 vdd
port 513 nsew
rlabel metal1 s 3504 28190 3504 28190 4 vdd
port 513 nsew
rlabel metal1 s 2736 25529 2736 25529 4 vdd
port 513 nsew
rlabel metal1 s 3504 26610 3504 26610 4 vdd
port 513 nsew
rlabel metal1 s 4752 28190 4752 28190 4 vdd
port 513 nsew
rlabel metal1 s 4752 25820 4752 25820 4 vdd
port 513 nsew
rlabel metal1 s 3984 26610 3984 26610 4 vdd
port 513 nsew
rlabel metal1 s 3984 27899 3984 27899 4 vdd
port 513 nsew
rlabel metal1 s 2736 26319 2736 26319 4 vdd
port 513 nsew
rlabel metal1 s 4752 25529 4752 25529 4 vdd
port 513 nsew
rlabel metal1 s 2736 27899 2736 27899 4 vdd
port 513 nsew
rlabel metal1 s 3504 27400 3504 27400 4 vdd
port 513 nsew
rlabel metal1 s 2736 27109 2736 27109 4 vdd
port 513 nsew
rlabel metal1 s 3984 26319 3984 26319 4 vdd
port 513 nsew
rlabel metal1 s 3984 25820 3984 25820 4 vdd
port 513 nsew
rlabel metal1 s 7728 28689 7728 28689 4 vdd
port 513 nsew
rlabel metal1 s 8976 28980 8976 28980 4 vdd
port 513 nsew
rlabel metal1 s 8496 30269 8496 30269 4 vdd
port 513 nsew
rlabel metal1 s 7728 30560 7728 30560 4 vdd
port 513 nsew
rlabel metal1 s 9744 31059 9744 31059 4 vdd
port 513 nsew
rlabel metal1 s 7728 29479 7728 29479 4 vdd
port 513 nsew
rlabel metal1 s 8496 31350 8496 31350 4 vdd
port 513 nsew
rlabel metal1 s 8976 30560 8976 30560 4 vdd
port 513 nsew
rlabel metal1 s 8496 28689 8496 28689 4 vdd
port 513 nsew
rlabel metal1 s 7728 30269 7728 30269 4 vdd
port 513 nsew
rlabel metal1 s 8496 30560 8496 30560 4 vdd
port 513 nsew
rlabel metal1 s 9744 29770 9744 29770 4 vdd
port 513 nsew
rlabel metal1 s 9744 29479 9744 29479 4 vdd
port 513 nsew
rlabel metal1 s 9744 28980 9744 28980 4 vdd
port 513 nsew
rlabel metal1 s 8496 29479 8496 29479 4 vdd
port 513 nsew
rlabel metal1 s 8976 28689 8976 28689 4 vdd
port 513 nsew
rlabel metal1 s 8976 31059 8976 31059 4 vdd
port 513 nsew
rlabel metal1 s 7728 28980 7728 28980 4 vdd
port 513 nsew
rlabel metal1 s 8496 29770 8496 29770 4 vdd
port 513 nsew
rlabel metal1 s 8976 29770 8976 29770 4 vdd
port 513 nsew
rlabel metal1 s 8976 29479 8976 29479 4 vdd
port 513 nsew
rlabel metal1 s 8496 31059 8496 31059 4 vdd
port 513 nsew
rlabel metal1 s 8496 28980 8496 28980 4 vdd
port 513 nsew
rlabel metal1 s 8976 31350 8976 31350 4 vdd
port 513 nsew
rlabel metal1 s 7728 31059 7728 31059 4 vdd
port 513 nsew
rlabel metal1 s 9744 30269 9744 30269 4 vdd
port 513 nsew
rlabel metal1 s 7728 31350 7728 31350 4 vdd
port 513 nsew
rlabel metal1 s 9744 30560 9744 30560 4 vdd
port 513 nsew
rlabel metal1 s 9744 28689 9744 28689 4 vdd
port 513 nsew
rlabel metal1 s 9744 31350 9744 31350 4 vdd
port 513 nsew
rlabel metal1 s 8976 30269 8976 30269 4 vdd
port 513 nsew
rlabel metal1 s 7728 29770 7728 29770 4 vdd
port 513 nsew
rlabel metal1 s 6480 31350 6480 31350 4 vdd
port 513 nsew
rlabel metal1 s 5232 31350 5232 31350 4 vdd
port 513 nsew
rlabel metal1 s 6000 30269 6000 30269 4 vdd
port 513 nsew
rlabel metal1 s 7248 28980 7248 28980 4 vdd
port 513 nsew
rlabel metal1 s 7248 29770 7248 29770 4 vdd
port 513 nsew
rlabel metal1 s 5232 31059 5232 31059 4 vdd
port 513 nsew
rlabel metal1 s 6000 29479 6000 29479 4 vdd
port 513 nsew
rlabel metal1 s 5232 30560 5232 30560 4 vdd
port 513 nsew
rlabel metal1 s 6000 30560 6000 30560 4 vdd
port 513 nsew
rlabel metal1 s 5232 28689 5232 28689 4 vdd
port 513 nsew
rlabel metal1 s 6480 30560 6480 30560 4 vdd
port 513 nsew
rlabel metal1 s 6000 28689 6000 28689 4 vdd
port 513 nsew
rlabel metal1 s 6480 31059 6480 31059 4 vdd
port 513 nsew
rlabel metal1 s 7248 28689 7248 28689 4 vdd
port 513 nsew
rlabel metal1 s 6480 28980 6480 28980 4 vdd
port 513 nsew
rlabel metal1 s 6480 29479 6480 29479 4 vdd
port 513 nsew
rlabel metal1 s 6000 29770 6000 29770 4 vdd
port 513 nsew
rlabel metal1 s 6000 31350 6000 31350 4 vdd
port 513 nsew
rlabel metal1 s 6000 31059 6000 31059 4 vdd
port 513 nsew
rlabel metal1 s 5232 29479 5232 29479 4 vdd
port 513 nsew
rlabel metal1 s 6000 28980 6000 28980 4 vdd
port 513 nsew
rlabel metal1 s 7248 31350 7248 31350 4 vdd
port 513 nsew
rlabel metal1 s 6480 30269 6480 30269 4 vdd
port 513 nsew
rlabel metal1 s 7248 29479 7248 29479 4 vdd
port 513 nsew
rlabel metal1 s 5232 28980 5232 28980 4 vdd
port 513 nsew
rlabel metal1 s 5232 30269 5232 30269 4 vdd
port 513 nsew
rlabel metal1 s 7248 30269 7248 30269 4 vdd
port 513 nsew
rlabel metal1 s 7248 31059 7248 31059 4 vdd
port 513 nsew
rlabel metal1 s 6480 28689 6480 28689 4 vdd
port 513 nsew
rlabel metal1 s 5232 29770 5232 29770 4 vdd
port 513 nsew
rlabel metal1 s 6480 29770 6480 29770 4 vdd
port 513 nsew
rlabel metal1 s 7248 30560 7248 30560 4 vdd
port 513 nsew
rlabel metal1 s 7248 25529 7248 25529 4 vdd
port 513 nsew
rlabel metal1 s 7248 27109 7248 27109 4 vdd
port 513 nsew
rlabel metal1 s 6480 26610 6480 26610 4 vdd
port 513 nsew
rlabel metal1 s 5232 28190 5232 28190 4 vdd
port 513 nsew
rlabel metal1 s 6000 26610 6000 26610 4 vdd
port 513 nsew
rlabel metal1 s 7248 27899 7248 27899 4 vdd
port 513 nsew
rlabel metal1 s 6480 27109 6480 27109 4 vdd
port 513 nsew
rlabel metal1 s 5232 25820 5232 25820 4 vdd
port 513 nsew
rlabel metal1 s 7248 26610 7248 26610 4 vdd
port 513 nsew
rlabel metal1 s 7248 28190 7248 28190 4 vdd
port 513 nsew
rlabel metal1 s 6000 27899 6000 27899 4 vdd
port 513 nsew
rlabel metal1 s 5232 27400 5232 27400 4 vdd
port 513 nsew
rlabel metal1 s 6000 27400 6000 27400 4 vdd
port 513 nsew
rlabel metal1 s 6000 26319 6000 26319 4 vdd
port 513 nsew
rlabel metal1 s 6480 25820 6480 25820 4 vdd
port 513 nsew
rlabel metal1 s 6480 26319 6480 26319 4 vdd
port 513 nsew
rlabel metal1 s 7248 25820 7248 25820 4 vdd
port 513 nsew
rlabel metal1 s 6480 27899 6480 27899 4 vdd
port 513 nsew
rlabel metal1 s 5232 25529 5232 25529 4 vdd
port 513 nsew
rlabel metal1 s 5232 26319 5232 26319 4 vdd
port 513 nsew
rlabel metal1 s 6000 25529 6000 25529 4 vdd
port 513 nsew
rlabel metal1 s 5232 26610 5232 26610 4 vdd
port 513 nsew
rlabel metal1 s 6000 25820 6000 25820 4 vdd
port 513 nsew
rlabel metal1 s 5232 27109 5232 27109 4 vdd
port 513 nsew
rlabel metal1 s 6000 28190 6000 28190 4 vdd
port 513 nsew
rlabel metal1 s 6000 27109 6000 27109 4 vdd
port 513 nsew
rlabel metal1 s 5232 27899 5232 27899 4 vdd
port 513 nsew
rlabel metal1 s 6480 28190 6480 28190 4 vdd
port 513 nsew
rlabel metal1 s 6480 25529 6480 25529 4 vdd
port 513 nsew
rlabel metal1 s 7248 26319 7248 26319 4 vdd
port 513 nsew
rlabel metal1 s 6480 27400 6480 27400 4 vdd
port 513 nsew
rlabel metal1 s 7248 27400 7248 27400 4 vdd
port 513 nsew
rlabel metal1 s 8496 27109 8496 27109 4 vdd
port 513 nsew
rlabel metal1 s 9744 27899 9744 27899 4 vdd
port 513 nsew
rlabel metal1 s 9744 28190 9744 28190 4 vdd
port 513 nsew
rlabel metal1 s 8496 25820 8496 25820 4 vdd
port 513 nsew
rlabel metal1 s 8496 28190 8496 28190 4 vdd
port 513 nsew
rlabel metal1 s 9744 26319 9744 26319 4 vdd
port 513 nsew
rlabel metal1 s 8976 26319 8976 26319 4 vdd
port 513 nsew
rlabel metal1 s 7728 27899 7728 27899 4 vdd
port 513 nsew
rlabel metal1 s 8976 26610 8976 26610 4 vdd
port 513 nsew
rlabel metal1 s 8496 26319 8496 26319 4 vdd
port 513 nsew
rlabel metal1 s 9744 25529 9744 25529 4 vdd
port 513 nsew
rlabel metal1 s 8976 27400 8976 27400 4 vdd
port 513 nsew
rlabel metal1 s 9744 26610 9744 26610 4 vdd
port 513 nsew
rlabel metal1 s 7728 27109 7728 27109 4 vdd
port 513 nsew
rlabel metal1 s 9744 25820 9744 25820 4 vdd
port 513 nsew
rlabel metal1 s 7728 26319 7728 26319 4 vdd
port 513 nsew
rlabel metal1 s 7728 25820 7728 25820 4 vdd
port 513 nsew
rlabel metal1 s 8976 28190 8976 28190 4 vdd
port 513 nsew
rlabel metal1 s 8496 26610 8496 26610 4 vdd
port 513 nsew
rlabel metal1 s 8496 27400 8496 27400 4 vdd
port 513 nsew
rlabel metal1 s 9744 27400 9744 27400 4 vdd
port 513 nsew
rlabel metal1 s 8496 25529 8496 25529 4 vdd
port 513 nsew
rlabel metal1 s 7728 27400 7728 27400 4 vdd
port 513 nsew
rlabel metal1 s 8976 25529 8976 25529 4 vdd
port 513 nsew
rlabel metal1 s 8976 27899 8976 27899 4 vdd
port 513 nsew
rlabel metal1 s 7728 28190 7728 28190 4 vdd
port 513 nsew
rlabel metal1 s 7728 26610 7728 26610 4 vdd
port 513 nsew
rlabel metal1 s 8976 27109 8976 27109 4 vdd
port 513 nsew
rlabel metal1 s 8976 25820 8976 25820 4 vdd
port 513 nsew
rlabel metal1 s 8496 27899 8496 27899 4 vdd
port 513 nsew
rlabel metal1 s 9744 27109 9744 27109 4 vdd
port 513 nsew
rlabel metal1 s 7728 25529 7728 25529 4 vdd
port 513 nsew
rlabel metal1 s 17712 35300 17712 35300 4 vdd
port 513 nsew
rlabel metal1 s 18960 36880 18960 36880 4 vdd
port 513 nsew
rlabel metal1 s 19728 35300 19728 35300 4 vdd
port 513 nsew
rlabel metal1 s 19728 37670 19728 37670 4 vdd
port 513 nsew
rlabel metal1 s 18480 37670 18480 37670 4 vdd
port 513 nsew
rlabel metal1 s 17712 35009 17712 35009 4 vdd
port 513 nsew
rlabel metal1 s 19728 36090 19728 36090 4 vdd
port 513 nsew
rlabel metal1 s 17712 36589 17712 36589 4 vdd
port 513 nsew
rlabel metal1 s 17712 37379 17712 37379 4 vdd
port 513 nsew
rlabel metal1 s 19728 35799 19728 35799 4 vdd
port 513 nsew
rlabel metal1 s 18480 36880 18480 36880 4 vdd
port 513 nsew
rlabel metal1 s 18960 36090 18960 36090 4 vdd
port 513 nsew
rlabel metal1 s 18480 35799 18480 35799 4 vdd
port 513 nsew
rlabel metal1 s 18960 37379 18960 37379 4 vdd
port 513 nsew
rlabel metal1 s 18960 35799 18960 35799 4 vdd
port 513 nsew
rlabel metal1 s 18960 37670 18960 37670 4 vdd
port 513 nsew
rlabel metal1 s 18480 37379 18480 37379 4 vdd
port 513 nsew
rlabel metal1 s 18480 36589 18480 36589 4 vdd
port 513 nsew
rlabel metal1 s 18480 35300 18480 35300 4 vdd
port 513 nsew
rlabel metal1 s 19728 36589 19728 36589 4 vdd
port 513 nsew
rlabel metal1 s 17712 36880 17712 36880 4 vdd
port 513 nsew
rlabel metal1 s 19728 37379 19728 37379 4 vdd
port 513 nsew
rlabel metal1 s 18960 35009 18960 35009 4 vdd
port 513 nsew
rlabel metal1 s 18960 36589 18960 36589 4 vdd
port 513 nsew
rlabel metal1 s 18480 35009 18480 35009 4 vdd
port 513 nsew
rlabel metal1 s 17712 35799 17712 35799 4 vdd
port 513 nsew
rlabel metal1 s 18960 35300 18960 35300 4 vdd
port 513 nsew
rlabel metal1 s 17712 37670 17712 37670 4 vdd
port 513 nsew
rlabel metal1 s 19728 35009 19728 35009 4 vdd
port 513 nsew
rlabel metal1 s 17712 36090 17712 36090 4 vdd
port 513 nsew
rlabel metal1 s 18480 36090 18480 36090 4 vdd
port 513 nsew
rlabel metal1 s 19728 36880 19728 36880 4 vdd
port 513 nsew
rlabel metal1 s 17232 35799 17232 35799 4 vdd
port 513 nsew
rlabel metal1 s 15984 36589 15984 36589 4 vdd
port 513 nsew
rlabel metal1 s 16464 37670 16464 37670 4 vdd
port 513 nsew
rlabel metal1 s 16464 35300 16464 35300 4 vdd
port 513 nsew
rlabel metal1 s 15984 35009 15984 35009 4 vdd
port 513 nsew
rlabel metal1 s 15216 36880 15216 36880 4 vdd
port 513 nsew
rlabel metal1 s 15216 35300 15216 35300 4 vdd
port 513 nsew
rlabel metal1 s 17232 37379 17232 37379 4 vdd
port 513 nsew
rlabel metal1 s 15984 37670 15984 37670 4 vdd
port 513 nsew
rlabel metal1 s 17232 37670 17232 37670 4 vdd
port 513 nsew
rlabel metal1 s 15216 37670 15216 37670 4 vdd
port 513 nsew
rlabel metal1 s 15984 35300 15984 35300 4 vdd
port 513 nsew
rlabel metal1 s 15984 35799 15984 35799 4 vdd
port 513 nsew
rlabel metal1 s 17232 36589 17232 36589 4 vdd
port 513 nsew
rlabel metal1 s 15216 36090 15216 36090 4 vdd
port 513 nsew
rlabel metal1 s 16464 35799 16464 35799 4 vdd
port 513 nsew
rlabel metal1 s 17232 35300 17232 35300 4 vdd
port 513 nsew
rlabel metal1 s 16464 36090 16464 36090 4 vdd
port 513 nsew
rlabel metal1 s 15216 36589 15216 36589 4 vdd
port 513 nsew
rlabel metal1 s 15216 35799 15216 35799 4 vdd
port 513 nsew
rlabel metal1 s 17232 36090 17232 36090 4 vdd
port 513 nsew
rlabel metal1 s 15216 35009 15216 35009 4 vdd
port 513 nsew
rlabel metal1 s 15984 36090 15984 36090 4 vdd
port 513 nsew
rlabel metal1 s 17232 36880 17232 36880 4 vdd
port 513 nsew
rlabel metal1 s 16464 37379 16464 37379 4 vdd
port 513 nsew
rlabel metal1 s 16464 35009 16464 35009 4 vdd
port 513 nsew
rlabel metal1 s 15984 36880 15984 36880 4 vdd
port 513 nsew
rlabel metal1 s 16464 36880 16464 36880 4 vdd
port 513 nsew
rlabel metal1 s 17232 35009 17232 35009 4 vdd
port 513 nsew
rlabel metal1 s 15984 37379 15984 37379 4 vdd
port 513 nsew
rlabel metal1 s 15216 37379 15216 37379 4 vdd
port 513 nsew
rlabel metal1 s 16464 36589 16464 36589 4 vdd
port 513 nsew
rlabel metal1 s 16464 34510 16464 34510 4 vdd
port 513 nsew
rlabel metal1 s 15984 32930 15984 32930 4 vdd
port 513 nsew
rlabel metal1 s 17232 32140 17232 32140 4 vdd
port 513 nsew
rlabel metal1 s 17232 33429 17232 33429 4 vdd
port 513 nsew
rlabel metal1 s 15216 33720 15216 33720 4 vdd
port 513 nsew
rlabel metal1 s 15984 34510 15984 34510 4 vdd
port 513 nsew
rlabel metal1 s 15984 34219 15984 34219 4 vdd
port 513 nsew
rlabel metal1 s 15984 31849 15984 31849 4 vdd
port 513 nsew
rlabel metal1 s 15216 32140 15216 32140 4 vdd
port 513 nsew
rlabel metal1 s 17232 34510 17232 34510 4 vdd
port 513 nsew
rlabel metal1 s 17232 31849 17232 31849 4 vdd
port 513 nsew
rlabel metal1 s 16464 34219 16464 34219 4 vdd
port 513 nsew
rlabel metal1 s 16464 32930 16464 32930 4 vdd
port 513 nsew
rlabel metal1 s 15216 32639 15216 32639 4 vdd
port 513 nsew
rlabel metal1 s 17232 32930 17232 32930 4 vdd
port 513 nsew
rlabel metal1 s 15984 33429 15984 33429 4 vdd
port 513 nsew
rlabel metal1 s 16464 33720 16464 33720 4 vdd
port 513 nsew
rlabel metal1 s 16464 33429 16464 33429 4 vdd
port 513 nsew
rlabel metal1 s 17232 32639 17232 32639 4 vdd
port 513 nsew
rlabel metal1 s 15216 32930 15216 32930 4 vdd
port 513 nsew
rlabel metal1 s 15216 33429 15216 33429 4 vdd
port 513 nsew
rlabel metal1 s 17232 34219 17232 34219 4 vdd
port 513 nsew
rlabel metal1 s 16464 31849 16464 31849 4 vdd
port 513 nsew
rlabel metal1 s 15984 32140 15984 32140 4 vdd
port 513 nsew
rlabel metal1 s 15216 31849 15216 31849 4 vdd
port 513 nsew
rlabel metal1 s 16464 32639 16464 32639 4 vdd
port 513 nsew
rlabel metal1 s 16464 32140 16464 32140 4 vdd
port 513 nsew
rlabel metal1 s 15216 34219 15216 34219 4 vdd
port 513 nsew
rlabel metal1 s 15984 33720 15984 33720 4 vdd
port 513 nsew
rlabel metal1 s 17232 33720 17232 33720 4 vdd
port 513 nsew
rlabel metal1 s 15216 34510 15216 34510 4 vdd
port 513 nsew
rlabel metal1 s 15984 32639 15984 32639 4 vdd
port 513 nsew
rlabel metal1 s 19728 32639 19728 32639 4 vdd
port 513 nsew
rlabel metal1 s 18480 32639 18480 32639 4 vdd
port 513 nsew
rlabel metal1 s 18960 31849 18960 31849 4 vdd
port 513 nsew
rlabel metal1 s 17712 33429 17712 33429 4 vdd
port 513 nsew
rlabel metal1 s 19728 33720 19728 33720 4 vdd
port 513 nsew
rlabel metal1 s 17712 32639 17712 32639 4 vdd
port 513 nsew
rlabel metal1 s 18480 34510 18480 34510 4 vdd
port 513 nsew
rlabel metal1 s 19728 31849 19728 31849 4 vdd
port 513 nsew
rlabel metal1 s 17712 34510 17712 34510 4 vdd
port 513 nsew
rlabel metal1 s 17712 33720 17712 33720 4 vdd
port 513 nsew
rlabel metal1 s 18960 33429 18960 33429 4 vdd
port 513 nsew
rlabel metal1 s 17712 32930 17712 32930 4 vdd
port 513 nsew
rlabel metal1 s 19728 32140 19728 32140 4 vdd
port 513 nsew
rlabel metal1 s 17712 32140 17712 32140 4 vdd
port 513 nsew
rlabel metal1 s 18960 32639 18960 32639 4 vdd
port 513 nsew
rlabel metal1 s 19728 33429 19728 33429 4 vdd
port 513 nsew
rlabel metal1 s 17712 34219 17712 34219 4 vdd
port 513 nsew
rlabel metal1 s 18480 31849 18480 31849 4 vdd
port 513 nsew
rlabel metal1 s 18480 33720 18480 33720 4 vdd
port 513 nsew
rlabel metal1 s 18480 32930 18480 32930 4 vdd
port 513 nsew
rlabel metal1 s 18480 34219 18480 34219 4 vdd
port 513 nsew
rlabel metal1 s 18480 33429 18480 33429 4 vdd
port 513 nsew
rlabel metal1 s 18960 33720 18960 33720 4 vdd
port 513 nsew
rlabel metal1 s 18960 34219 18960 34219 4 vdd
port 513 nsew
rlabel metal1 s 18960 34510 18960 34510 4 vdd
port 513 nsew
rlabel metal1 s 18960 32140 18960 32140 4 vdd
port 513 nsew
rlabel metal1 s 18480 32140 18480 32140 4 vdd
port 513 nsew
rlabel metal1 s 19728 32930 19728 32930 4 vdd
port 513 nsew
rlabel metal1 s 18960 32930 18960 32930 4 vdd
port 513 nsew
rlabel metal1 s 19728 34510 19728 34510 4 vdd
port 513 nsew
rlabel metal1 s 17712 31849 17712 31849 4 vdd
port 513 nsew
rlabel metal1 s 19728 34219 19728 34219 4 vdd
port 513 nsew
rlabel metal1 s 14736 37670 14736 37670 4 vdd
port 513 nsew
rlabel metal1 s 12720 36090 12720 36090 4 vdd
port 513 nsew
rlabel metal1 s 13488 35009 13488 35009 4 vdd
port 513 nsew
rlabel metal1 s 14736 36880 14736 36880 4 vdd
port 513 nsew
rlabel metal1 s 12720 36880 12720 36880 4 vdd
port 513 nsew
rlabel metal1 s 13968 35009 13968 35009 4 vdd
port 513 nsew
rlabel metal1 s 12720 37379 12720 37379 4 vdd
port 513 nsew
rlabel metal1 s 14736 36589 14736 36589 4 vdd
port 513 nsew
rlabel metal1 s 13488 35300 13488 35300 4 vdd
port 513 nsew
rlabel metal1 s 13968 35300 13968 35300 4 vdd
port 513 nsew
rlabel metal1 s 13968 37379 13968 37379 4 vdd
port 513 nsew
rlabel metal1 s 12720 35300 12720 35300 4 vdd
port 513 nsew
rlabel metal1 s 12720 35799 12720 35799 4 vdd
port 513 nsew
rlabel metal1 s 12720 37670 12720 37670 4 vdd
port 513 nsew
rlabel metal1 s 14736 35300 14736 35300 4 vdd
port 513 nsew
rlabel metal1 s 13968 36589 13968 36589 4 vdd
port 513 nsew
rlabel metal1 s 13968 37670 13968 37670 4 vdd
port 513 nsew
rlabel metal1 s 12720 36589 12720 36589 4 vdd
port 513 nsew
rlabel metal1 s 14736 35009 14736 35009 4 vdd
port 513 nsew
rlabel metal1 s 13968 35799 13968 35799 4 vdd
port 513 nsew
rlabel metal1 s 13488 36880 13488 36880 4 vdd
port 513 nsew
rlabel metal1 s 12720 35009 12720 35009 4 vdd
port 513 nsew
rlabel metal1 s 13968 36090 13968 36090 4 vdd
port 513 nsew
rlabel metal1 s 13488 36589 13488 36589 4 vdd
port 513 nsew
rlabel metal1 s 14736 36090 14736 36090 4 vdd
port 513 nsew
rlabel metal1 s 13488 37670 13488 37670 4 vdd
port 513 nsew
rlabel metal1 s 14736 35799 14736 35799 4 vdd
port 513 nsew
rlabel metal1 s 13488 35799 13488 35799 4 vdd
port 513 nsew
rlabel metal1 s 14736 37379 14736 37379 4 vdd
port 513 nsew
rlabel metal1 s 13968 36880 13968 36880 4 vdd
port 513 nsew
rlabel metal1 s 13488 37379 13488 37379 4 vdd
port 513 nsew
rlabel metal1 s 13488 36090 13488 36090 4 vdd
port 513 nsew
rlabel metal1 s 10224 35300 10224 35300 4 vdd
port 513 nsew
rlabel metal1 s 10224 37670 10224 37670 4 vdd
port 513 nsew
rlabel metal1 s 11472 37379 11472 37379 4 vdd
port 513 nsew
rlabel metal1 s 10224 35799 10224 35799 4 vdd
port 513 nsew
rlabel metal1 s 12240 35799 12240 35799 4 vdd
port 513 nsew
rlabel metal1 s 10224 36589 10224 36589 4 vdd
port 513 nsew
rlabel metal1 s 10992 35009 10992 35009 4 vdd
port 513 nsew
rlabel metal1 s 12240 37670 12240 37670 4 vdd
port 513 nsew
rlabel metal1 s 10992 37670 10992 37670 4 vdd
port 513 nsew
rlabel metal1 s 12240 36880 12240 36880 4 vdd
port 513 nsew
rlabel metal1 s 11472 37670 11472 37670 4 vdd
port 513 nsew
rlabel metal1 s 10992 35300 10992 35300 4 vdd
port 513 nsew
rlabel metal1 s 12240 35300 12240 35300 4 vdd
port 513 nsew
rlabel metal1 s 10992 36880 10992 36880 4 vdd
port 513 nsew
rlabel metal1 s 10224 36880 10224 36880 4 vdd
port 513 nsew
rlabel metal1 s 12240 35009 12240 35009 4 vdd
port 513 nsew
rlabel metal1 s 10224 36090 10224 36090 4 vdd
port 513 nsew
rlabel metal1 s 10224 35009 10224 35009 4 vdd
port 513 nsew
rlabel metal1 s 10992 35799 10992 35799 4 vdd
port 513 nsew
rlabel metal1 s 10992 36589 10992 36589 4 vdd
port 513 nsew
rlabel metal1 s 12240 37379 12240 37379 4 vdd
port 513 nsew
rlabel metal1 s 11472 36589 11472 36589 4 vdd
port 513 nsew
rlabel metal1 s 11472 35009 11472 35009 4 vdd
port 513 nsew
rlabel metal1 s 11472 36090 11472 36090 4 vdd
port 513 nsew
rlabel metal1 s 11472 35799 11472 35799 4 vdd
port 513 nsew
rlabel metal1 s 10992 37379 10992 37379 4 vdd
port 513 nsew
rlabel metal1 s 12240 36090 12240 36090 4 vdd
port 513 nsew
rlabel metal1 s 10992 36090 10992 36090 4 vdd
port 513 nsew
rlabel metal1 s 11472 36880 11472 36880 4 vdd
port 513 nsew
rlabel metal1 s 11472 35300 11472 35300 4 vdd
port 513 nsew
rlabel metal1 s 10224 37379 10224 37379 4 vdd
port 513 nsew
rlabel metal1 s 12240 36589 12240 36589 4 vdd
port 513 nsew
rlabel metal1 s 11472 33429 11472 33429 4 vdd
port 513 nsew
rlabel metal1 s 10992 33720 10992 33720 4 vdd
port 513 nsew
rlabel metal1 s 10224 33720 10224 33720 4 vdd
port 513 nsew
rlabel metal1 s 11472 34219 11472 34219 4 vdd
port 513 nsew
rlabel metal1 s 11472 32930 11472 32930 4 vdd
port 513 nsew
rlabel metal1 s 12240 32639 12240 32639 4 vdd
port 513 nsew
rlabel metal1 s 10992 34219 10992 34219 4 vdd
port 513 nsew
rlabel metal1 s 11472 33720 11472 33720 4 vdd
port 513 nsew
rlabel metal1 s 11472 31849 11472 31849 4 vdd
port 513 nsew
rlabel metal1 s 10224 32930 10224 32930 4 vdd
port 513 nsew
rlabel metal1 s 12240 32930 12240 32930 4 vdd
port 513 nsew
rlabel metal1 s 10992 33429 10992 33429 4 vdd
port 513 nsew
rlabel metal1 s 10224 31849 10224 31849 4 vdd
port 513 nsew
rlabel metal1 s 10992 32140 10992 32140 4 vdd
port 513 nsew
rlabel metal1 s 10992 32930 10992 32930 4 vdd
port 513 nsew
rlabel metal1 s 11472 32140 11472 32140 4 vdd
port 513 nsew
rlabel metal1 s 10992 32639 10992 32639 4 vdd
port 513 nsew
rlabel metal1 s 10992 31849 10992 31849 4 vdd
port 513 nsew
rlabel metal1 s 10224 33429 10224 33429 4 vdd
port 513 nsew
rlabel metal1 s 12240 33720 12240 33720 4 vdd
port 513 nsew
rlabel metal1 s 12240 34219 12240 34219 4 vdd
port 513 nsew
rlabel metal1 s 10224 34510 10224 34510 4 vdd
port 513 nsew
rlabel metal1 s 10224 32140 10224 32140 4 vdd
port 513 nsew
rlabel metal1 s 10224 34219 10224 34219 4 vdd
port 513 nsew
rlabel metal1 s 12240 33429 12240 33429 4 vdd
port 513 nsew
rlabel metal1 s 10224 32639 10224 32639 4 vdd
port 513 nsew
rlabel metal1 s 12240 34510 12240 34510 4 vdd
port 513 nsew
rlabel metal1 s 11472 32639 11472 32639 4 vdd
port 513 nsew
rlabel metal1 s 10992 34510 10992 34510 4 vdd
port 513 nsew
rlabel metal1 s 12240 31849 12240 31849 4 vdd
port 513 nsew
rlabel metal1 s 12240 32140 12240 32140 4 vdd
port 513 nsew
rlabel metal1 s 11472 34510 11472 34510 4 vdd
port 513 nsew
rlabel metal1 s 12720 32639 12720 32639 4 vdd
port 513 nsew
rlabel metal1 s 12720 33429 12720 33429 4 vdd
port 513 nsew
rlabel metal1 s 14736 33720 14736 33720 4 vdd
port 513 nsew
rlabel metal1 s 13968 33429 13968 33429 4 vdd
port 513 nsew
rlabel metal1 s 13488 31849 13488 31849 4 vdd
port 513 nsew
rlabel metal1 s 14736 32639 14736 32639 4 vdd
port 513 nsew
rlabel metal1 s 13488 33429 13488 33429 4 vdd
port 513 nsew
rlabel metal1 s 12720 31849 12720 31849 4 vdd
port 513 nsew
rlabel metal1 s 13488 32930 13488 32930 4 vdd
port 513 nsew
rlabel metal1 s 13488 33720 13488 33720 4 vdd
port 513 nsew
rlabel metal1 s 13968 33720 13968 33720 4 vdd
port 513 nsew
rlabel metal1 s 13968 34510 13968 34510 4 vdd
port 513 nsew
rlabel metal1 s 13488 34219 13488 34219 4 vdd
port 513 nsew
rlabel metal1 s 14736 34510 14736 34510 4 vdd
port 513 nsew
rlabel metal1 s 13968 32140 13968 32140 4 vdd
port 513 nsew
rlabel metal1 s 13968 34219 13968 34219 4 vdd
port 513 nsew
rlabel metal1 s 14736 31849 14736 31849 4 vdd
port 513 nsew
rlabel metal1 s 13968 31849 13968 31849 4 vdd
port 513 nsew
rlabel metal1 s 12720 32930 12720 32930 4 vdd
port 513 nsew
rlabel metal1 s 12720 32140 12720 32140 4 vdd
port 513 nsew
rlabel metal1 s 14736 34219 14736 34219 4 vdd
port 513 nsew
rlabel metal1 s 12720 34510 12720 34510 4 vdd
port 513 nsew
rlabel metal1 s 12720 33720 12720 33720 4 vdd
port 513 nsew
rlabel metal1 s 13968 32930 13968 32930 4 vdd
port 513 nsew
rlabel metal1 s 13488 32639 13488 32639 4 vdd
port 513 nsew
rlabel metal1 s 13488 32140 13488 32140 4 vdd
port 513 nsew
rlabel metal1 s 12720 34219 12720 34219 4 vdd
port 513 nsew
rlabel metal1 s 13488 34510 13488 34510 4 vdd
port 513 nsew
rlabel metal1 s 14736 32930 14736 32930 4 vdd
port 513 nsew
rlabel metal1 s 14736 32140 14736 32140 4 vdd
port 513 nsew
rlabel metal1 s 13968 32639 13968 32639 4 vdd
port 513 nsew
rlabel metal1 s 14736 33429 14736 33429 4 vdd
port 513 nsew
rlabel metal1 s 13968 30560 13968 30560 4 vdd
port 513 nsew
rlabel metal1 s 13968 28689 13968 28689 4 vdd
port 513 nsew
rlabel metal1 s 13488 28689 13488 28689 4 vdd
port 513 nsew
rlabel metal1 s 14736 31350 14736 31350 4 vdd
port 513 nsew
rlabel metal1 s 13488 30560 13488 30560 4 vdd
port 513 nsew
rlabel metal1 s 13488 29770 13488 29770 4 vdd
port 513 nsew
rlabel metal1 s 12720 28689 12720 28689 4 vdd
port 513 nsew
rlabel metal1 s 13488 30269 13488 30269 4 vdd
port 513 nsew
rlabel metal1 s 12720 30269 12720 30269 4 vdd
port 513 nsew
rlabel metal1 s 14736 31059 14736 31059 4 vdd
port 513 nsew
rlabel metal1 s 13968 31059 13968 31059 4 vdd
port 513 nsew
rlabel metal1 s 13968 29479 13968 29479 4 vdd
port 513 nsew
rlabel metal1 s 13488 28980 13488 28980 4 vdd
port 513 nsew
rlabel metal1 s 13488 29479 13488 29479 4 vdd
port 513 nsew
rlabel metal1 s 12720 31059 12720 31059 4 vdd
port 513 nsew
rlabel metal1 s 14736 29479 14736 29479 4 vdd
port 513 nsew
rlabel metal1 s 12720 29479 12720 29479 4 vdd
port 513 nsew
rlabel metal1 s 13968 31350 13968 31350 4 vdd
port 513 nsew
rlabel metal1 s 14736 30560 14736 30560 4 vdd
port 513 nsew
rlabel metal1 s 14736 28689 14736 28689 4 vdd
port 513 nsew
rlabel metal1 s 13488 31350 13488 31350 4 vdd
port 513 nsew
rlabel metal1 s 12720 30560 12720 30560 4 vdd
port 513 nsew
rlabel metal1 s 13968 29770 13968 29770 4 vdd
port 513 nsew
rlabel metal1 s 14736 30269 14736 30269 4 vdd
port 513 nsew
rlabel metal1 s 13968 28980 13968 28980 4 vdd
port 513 nsew
rlabel metal1 s 13488 31059 13488 31059 4 vdd
port 513 nsew
rlabel metal1 s 14736 28980 14736 28980 4 vdd
port 513 nsew
rlabel metal1 s 13968 30269 13968 30269 4 vdd
port 513 nsew
rlabel metal1 s 12720 31350 12720 31350 4 vdd
port 513 nsew
rlabel metal1 s 14736 29770 14736 29770 4 vdd
port 513 nsew
rlabel metal1 s 12720 28980 12720 28980 4 vdd
port 513 nsew
rlabel metal1 s 12720 29770 12720 29770 4 vdd
port 513 nsew
rlabel metal1 s 10224 29479 10224 29479 4 vdd
port 513 nsew
rlabel metal1 s 10992 28980 10992 28980 4 vdd
port 513 nsew
rlabel metal1 s 11472 30560 11472 30560 4 vdd
port 513 nsew
rlabel metal1 s 10992 30269 10992 30269 4 vdd
port 513 nsew
rlabel metal1 s 12240 29770 12240 29770 4 vdd
port 513 nsew
rlabel metal1 s 12240 29479 12240 29479 4 vdd
port 513 nsew
rlabel metal1 s 10224 29770 10224 29770 4 vdd
port 513 nsew
rlabel metal1 s 10992 31350 10992 31350 4 vdd
port 513 nsew
rlabel metal1 s 11472 29770 11472 29770 4 vdd
port 513 nsew
rlabel metal1 s 10224 28980 10224 28980 4 vdd
port 513 nsew
rlabel metal1 s 10224 30269 10224 30269 4 vdd
port 513 nsew
rlabel metal1 s 10992 28689 10992 28689 4 vdd
port 513 nsew
rlabel metal1 s 11472 31350 11472 31350 4 vdd
port 513 nsew
rlabel metal1 s 11472 28689 11472 28689 4 vdd
port 513 nsew
rlabel metal1 s 12240 31059 12240 31059 4 vdd
port 513 nsew
rlabel metal1 s 10992 29770 10992 29770 4 vdd
port 513 nsew
rlabel metal1 s 10224 28689 10224 28689 4 vdd
port 513 nsew
rlabel metal1 s 12240 30560 12240 30560 4 vdd
port 513 nsew
rlabel metal1 s 12240 28980 12240 28980 4 vdd
port 513 nsew
rlabel metal1 s 10992 30560 10992 30560 4 vdd
port 513 nsew
rlabel metal1 s 11472 30269 11472 30269 4 vdd
port 513 nsew
rlabel metal1 s 11472 31059 11472 31059 4 vdd
port 513 nsew
rlabel metal1 s 10224 30560 10224 30560 4 vdd
port 513 nsew
rlabel metal1 s 12240 30269 12240 30269 4 vdd
port 513 nsew
rlabel metal1 s 10224 31350 10224 31350 4 vdd
port 513 nsew
rlabel metal1 s 11472 29479 11472 29479 4 vdd
port 513 nsew
rlabel metal1 s 12240 31350 12240 31350 4 vdd
port 513 nsew
rlabel metal1 s 10992 29479 10992 29479 4 vdd
port 513 nsew
rlabel metal1 s 11472 28980 11472 28980 4 vdd
port 513 nsew
rlabel metal1 s 12240 28689 12240 28689 4 vdd
port 513 nsew
rlabel metal1 s 10224 31059 10224 31059 4 vdd
port 513 nsew
rlabel metal1 s 10992 31059 10992 31059 4 vdd
port 513 nsew
rlabel metal1 s 12240 26610 12240 26610 4 vdd
port 513 nsew
rlabel metal1 s 10224 27109 10224 27109 4 vdd
port 513 nsew
rlabel metal1 s 10224 25820 10224 25820 4 vdd
port 513 nsew
rlabel metal1 s 11472 26319 11472 26319 4 vdd
port 513 nsew
rlabel metal1 s 11472 28190 11472 28190 4 vdd
port 513 nsew
rlabel metal1 s 11472 25820 11472 25820 4 vdd
port 513 nsew
rlabel metal1 s 10992 25529 10992 25529 4 vdd
port 513 nsew
rlabel metal1 s 10224 26319 10224 26319 4 vdd
port 513 nsew
rlabel metal1 s 10224 26610 10224 26610 4 vdd
port 513 nsew
rlabel metal1 s 10992 27400 10992 27400 4 vdd
port 513 nsew
rlabel metal1 s 11472 27400 11472 27400 4 vdd
port 513 nsew
rlabel metal1 s 11472 25529 11472 25529 4 vdd
port 513 nsew
rlabel metal1 s 10992 27109 10992 27109 4 vdd
port 513 nsew
rlabel metal1 s 10992 27899 10992 27899 4 vdd
port 513 nsew
rlabel metal1 s 10992 28190 10992 28190 4 vdd
port 513 nsew
rlabel metal1 s 12240 27109 12240 27109 4 vdd
port 513 nsew
rlabel metal1 s 10224 28190 10224 28190 4 vdd
port 513 nsew
rlabel metal1 s 10992 26319 10992 26319 4 vdd
port 513 nsew
rlabel metal1 s 12240 28190 12240 28190 4 vdd
port 513 nsew
rlabel metal1 s 12240 26319 12240 26319 4 vdd
port 513 nsew
rlabel metal1 s 11472 27899 11472 27899 4 vdd
port 513 nsew
rlabel metal1 s 11472 26610 11472 26610 4 vdd
port 513 nsew
rlabel metal1 s 10224 25529 10224 25529 4 vdd
port 513 nsew
rlabel metal1 s 10224 27400 10224 27400 4 vdd
port 513 nsew
rlabel metal1 s 12240 25529 12240 25529 4 vdd
port 513 nsew
rlabel metal1 s 11472 27109 11472 27109 4 vdd
port 513 nsew
rlabel metal1 s 10992 26610 10992 26610 4 vdd
port 513 nsew
rlabel metal1 s 12240 25820 12240 25820 4 vdd
port 513 nsew
rlabel metal1 s 10992 25820 10992 25820 4 vdd
port 513 nsew
rlabel metal1 s 12240 27400 12240 27400 4 vdd
port 513 nsew
rlabel metal1 s 10224 27899 10224 27899 4 vdd
port 513 nsew
rlabel metal1 s 12240 27899 12240 27899 4 vdd
port 513 nsew
rlabel metal1 s 13968 26319 13968 26319 4 vdd
port 513 nsew
rlabel metal1 s 13488 26610 13488 26610 4 vdd
port 513 nsew
rlabel metal1 s 14736 25529 14736 25529 4 vdd
port 513 nsew
rlabel metal1 s 12720 26610 12720 26610 4 vdd
port 513 nsew
rlabel metal1 s 14736 28190 14736 28190 4 vdd
port 513 nsew
rlabel metal1 s 13968 27109 13968 27109 4 vdd
port 513 nsew
rlabel metal1 s 13488 25820 13488 25820 4 vdd
port 513 nsew
rlabel metal1 s 12720 26319 12720 26319 4 vdd
port 513 nsew
rlabel metal1 s 13968 25820 13968 25820 4 vdd
port 513 nsew
rlabel metal1 s 13968 25529 13968 25529 4 vdd
port 513 nsew
rlabel metal1 s 14736 26610 14736 26610 4 vdd
port 513 nsew
rlabel metal1 s 12720 27109 12720 27109 4 vdd
port 513 nsew
rlabel metal1 s 13488 25529 13488 25529 4 vdd
port 513 nsew
rlabel metal1 s 13968 27899 13968 27899 4 vdd
port 513 nsew
rlabel metal1 s 13968 26610 13968 26610 4 vdd
port 513 nsew
rlabel metal1 s 14736 27109 14736 27109 4 vdd
port 513 nsew
rlabel metal1 s 12720 28190 12720 28190 4 vdd
port 513 nsew
rlabel metal1 s 12720 27899 12720 27899 4 vdd
port 513 nsew
rlabel metal1 s 13968 28190 13968 28190 4 vdd
port 513 nsew
rlabel metal1 s 14736 27400 14736 27400 4 vdd
port 513 nsew
rlabel metal1 s 14736 26319 14736 26319 4 vdd
port 513 nsew
rlabel metal1 s 14736 27899 14736 27899 4 vdd
port 513 nsew
rlabel metal1 s 13488 28190 13488 28190 4 vdd
port 513 nsew
rlabel metal1 s 12720 25529 12720 25529 4 vdd
port 513 nsew
rlabel metal1 s 14736 25820 14736 25820 4 vdd
port 513 nsew
rlabel metal1 s 13488 27400 13488 27400 4 vdd
port 513 nsew
rlabel metal1 s 13488 27109 13488 27109 4 vdd
port 513 nsew
rlabel metal1 s 12720 25820 12720 25820 4 vdd
port 513 nsew
rlabel metal1 s 13968 27400 13968 27400 4 vdd
port 513 nsew
rlabel metal1 s 12720 27400 12720 27400 4 vdd
port 513 nsew
rlabel metal1 s 13488 27899 13488 27899 4 vdd
port 513 nsew
rlabel metal1 s 13488 26319 13488 26319 4 vdd
port 513 nsew
rlabel metal1 s 19728 29770 19728 29770 4 vdd
port 513 nsew
rlabel metal1 s 19728 31350 19728 31350 4 vdd
port 513 nsew
rlabel metal1 s 18480 29770 18480 29770 4 vdd
port 513 nsew
rlabel metal1 s 18480 30269 18480 30269 4 vdd
port 513 nsew
rlabel metal1 s 19728 29479 19728 29479 4 vdd
port 513 nsew
rlabel metal1 s 18960 31350 18960 31350 4 vdd
port 513 nsew
rlabel metal1 s 18960 30560 18960 30560 4 vdd
port 513 nsew
rlabel metal1 s 19728 31059 19728 31059 4 vdd
port 513 nsew
rlabel metal1 s 17712 28980 17712 28980 4 vdd
port 513 nsew
rlabel metal1 s 18480 31059 18480 31059 4 vdd
port 513 nsew
rlabel metal1 s 17712 31059 17712 31059 4 vdd
port 513 nsew
rlabel metal1 s 18480 31350 18480 31350 4 vdd
port 513 nsew
rlabel metal1 s 18960 29770 18960 29770 4 vdd
port 513 nsew
rlabel metal1 s 19728 28980 19728 28980 4 vdd
port 513 nsew
rlabel metal1 s 17712 30269 17712 30269 4 vdd
port 513 nsew
rlabel metal1 s 18960 30269 18960 30269 4 vdd
port 513 nsew
rlabel metal1 s 19728 30269 19728 30269 4 vdd
port 513 nsew
rlabel metal1 s 17712 29770 17712 29770 4 vdd
port 513 nsew
rlabel metal1 s 19728 30560 19728 30560 4 vdd
port 513 nsew
rlabel metal1 s 18960 28980 18960 28980 4 vdd
port 513 nsew
rlabel metal1 s 18480 30560 18480 30560 4 vdd
port 513 nsew
rlabel metal1 s 17712 28689 17712 28689 4 vdd
port 513 nsew
rlabel metal1 s 18480 29479 18480 29479 4 vdd
port 513 nsew
rlabel metal1 s 17712 31350 17712 31350 4 vdd
port 513 nsew
rlabel metal1 s 18960 28689 18960 28689 4 vdd
port 513 nsew
rlabel metal1 s 18960 29479 18960 29479 4 vdd
port 513 nsew
rlabel metal1 s 18480 28980 18480 28980 4 vdd
port 513 nsew
rlabel metal1 s 18960 31059 18960 31059 4 vdd
port 513 nsew
rlabel metal1 s 17712 29479 17712 29479 4 vdd
port 513 nsew
rlabel metal1 s 19728 28689 19728 28689 4 vdd
port 513 nsew
rlabel metal1 s 17712 30560 17712 30560 4 vdd
port 513 nsew
rlabel metal1 s 18480 28689 18480 28689 4 vdd
port 513 nsew
rlabel metal1 s 16464 31350 16464 31350 4 vdd
port 513 nsew
rlabel metal1 s 16464 30560 16464 30560 4 vdd
port 513 nsew
rlabel metal1 s 16464 28980 16464 28980 4 vdd
port 513 nsew
rlabel metal1 s 17232 29479 17232 29479 4 vdd
port 513 nsew
rlabel metal1 s 17232 30560 17232 30560 4 vdd
port 513 nsew
rlabel metal1 s 15216 29770 15216 29770 4 vdd
port 513 nsew
rlabel metal1 s 15984 29479 15984 29479 4 vdd
port 513 nsew
rlabel metal1 s 16464 31059 16464 31059 4 vdd
port 513 nsew
rlabel metal1 s 15216 30560 15216 30560 4 vdd
port 513 nsew
rlabel metal1 s 16464 29770 16464 29770 4 vdd
port 513 nsew
rlabel metal1 s 15216 30269 15216 30269 4 vdd
port 513 nsew
rlabel metal1 s 15984 30269 15984 30269 4 vdd
port 513 nsew
rlabel metal1 s 15984 28980 15984 28980 4 vdd
port 513 nsew
rlabel metal1 s 16464 28689 16464 28689 4 vdd
port 513 nsew
rlabel metal1 s 15216 31059 15216 31059 4 vdd
port 513 nsew
rlabel metal1 s 17232 28689 17232 28689 4 vdd
port 513 nsew
rlabel metal1 s 15216 28980 15216 28980 4 vdd
port 513 nsew
rlabel metal1 s 15984 31350 15984 31350 4 vdd
port 513 nsew
rlabel metal1 s 15984 30560 15984 30560 4 vdd
port 513 nsew
rlabel metal1 s 15984 31059 15984 31059 4 vdd
port 513 nsew
rlabel metal1 s 15984 28689 15984 28689 4 vdd
port 513 nsew
rlabel metal1 s 15216 28689 15216 28689 4 vdd
port 513 nsew
rlabel metal1 s 15216 29479 15216 29479 4 vdd
port 513 nsew
rlabel metal1 s 15984 29770 15984 29770 4 vdd
port 513 nsew
rlabel metal1 s 16464 29479 16464 29479 4 vdd
port 513 nsew
rlabel metal1 s 17232 28980 17232 28980 4 vdd
port 513 nsew
rlabel metal1 s 17232 29770 17232 29770 4 vdd
port 513 nsew
rlabel metal1 s 17232 31059 17232 31059 4 vdd
port 513 nsew
rlabel metal1 s 17232 31350 17232 31350 4 vdd
port 513 nsew
rlabel metal1 s 17232 30269 17232 30269 4 vdd
port 513 nsew
rlabel metal1 s 16464 30269 16464 30269 4 vdd
port 513 nsew
rlabel metal1 s 15216 31350 15216 31350 4 vdd
port 513 nsew
rlabel metal1 s 16464 27899 16464 27899 4 vdd
port 513 nsew
rlabel metal1 s 15216 28190 15216 28190 4 vdd
port 513 nsew
rlabel metal1 s 17232 28190 17232 28190 4 vdd
port 513 nsew
rlabel metal1 s 15216 27899 15216 27899 4 vdd
port 513 nsew
rlabel metal1 s 15984 27400 15984 27400 4 vdd
port 513 nsew
rlabel metal1 s 15216 27109 15216 27109 4 vdd
port 513 nsew
rlabel metal1 s 16464 27400 16464 27400 4 vdd
port 513 nsew
rlabel metal1 s 15216 27400 15216 27400 4 vdd
port 513 nsew
rlabel metal1 s 15984 26610 15984 26610 4 vdd
port 513 nsew
rlabel metal1 s 17232 26610 17232 26610 4 vdd
port 513 nsew
rlabel metal1 s 15984 27899 15984 27899 4 vdd
port 513 nsew
rlabel metal1 s 15984 27109 15984 27109 4 vdd
port 513 nsew
rlabel metal1 s 16464 28190 16464 28190 4 vdd
port 513 nsew
rlabel metal1 s 16464 26319 16464 26319 4 vdd
port 513 nsew
rlabel metal1 s 17232 27109 17232 27109 4 vdd
port 513 nsew
rlabel metal1 s 17232 27400 17232 27400 4 vdd
port 513 nsew
rlabel metal1 s 15216 25820 15216 25820 4 vdd
port 513 nsew
rlabel metal1 s 15984 28190 15984 28190 4 vdd
port 513 nsew
rlabel metal1 s 15984 26319 15984 26319 4 vdd
port 513 nsew
rlabel metal1 s 17232 25820 17232 25820 4 vdd
port 513 nsew
rlabel metal1 s 17232 27899 17232 27899 4 vdd
port 513 nsew
rlabel metal1 s 16464 25820 16464 25820 4 vdd
port 513 nsew
rlabel metal1 s 16464 25529 16464 25529 4 vdd
port 513 nsew
rlabel metal1 s 15216 26319 15216 26319 4 vdd
port 513 nsew
rlabel metal1 s 15216 25529 15216 25529 4 vdd
port 513 nsew
rlabel metal1 s 16464 26610 16464 26610 4 vdd
port 513 nsew
rlabel metal1 s 16464 27109 16464 27109 4 vdd
port 513 nsew
rlabel metal1 s 17232 26319 17232 26319 4 vdd
port 513 nsew
rlabel metal1 s 15216 26610 15216 26610 4 vdd
port 513 nsew
rlabel metal1 s 17232 25529 17232 25529 4 vdd
port 513 nsew
rlabel metal1 s 15984 25820 15984 25820 4 vdd
port 513 nsew
rlabel metal1 s 15984 25529 15984 25529 4 vdd
port 513 nsew
rlabel metal1 s 17712 25529 17712 25529 4 vdd
port 513 nsew
rlabel metal1 s 18480 27899 18480 27899 4 vdd
port 513 nsew
rlabel metal1 s 19728 26319 19728 26319 4 vdd
port 513 nsew
rlabel metal1 s 18480 27400 18480 27400 4 vdd
port 513 nsew
rlabel metal1 s 18960 26610 18960 26610 4 vdd
port 513 nsew
rlabel metal1 s 18480 25820 18480 25820 4 vdd
port 513 nsew
rlabel metal1 s 19728 27400 19728 27400 4 vdd
port 513 nsew
rlabel metal1 s 17712 27899 17712 27899 4 vdd
port 513 nsew
rlabel metal1 s 18960 28190 18960 28190 4 vdd
port 513 nsew
rlabel metal1 s 19728 27109 19728 27109 4 vdd
port 513 nsew
rlabel metal1 s 18480 25529 18480 25529 4 vdd
port 513 nsew
rlabel metal1 s 19728 25820 19728 25820 4 vdd
port 513 nsew
rlabel metal1 s 18480 26319 18480 26319 4 vdd
port 513 nsew
rlabel metal1 s 18960 26319 18960 26319 4 vdd
port 513 nsew
rlabel metal1 s 18960 27400 18960 27400 4 vdd
port 513 nsew
rlabel metal1 s 18960 25820 18960 25820 4 vdd
port 513 nsew
rlabel metal1 s 18960 27899 18960 27899 4 vdd
port 513 nsew
rlabel metal1 s 19728 28190 19728 28190 4 vdd
port 513 nsew
rlabel metal1 s 17712 25820 17712 25820 4 vdd
port 513 nsew
rlabel metal1 s 18960 27109 18960 27109 4 vdd
port 513 nsew
rlabel metal1 s 18960 25529 18960 25529 4 vdd
port 513 nsew
rlabel metal1 s 18480 28190 18480 28190 4 vdd
port 513 nsew
rlabel metal1 s 17712 26610 17712 26610 4 vdd
port 513 nsew
rlabel metal1 s 19728 25529 19728 25529 4 vdd
port 513 nsew
rlabel metal1 s 18480 26610 18480 26610 4 vdd
port 513 nsew
rlabel metal1 s 17712 27400 17712 27400 4 vdd
port 513 nsew
rlabel metal1 s 19728 27899 19728 27899 4 vdd
port 513 nsew
rlabel metal1 s 19728 26610 19728 26610 4 vdd
port 513 nsew
rlabel metal1 s 18480 27109 18480 27109 4 vdd
port 513 nsew
rlabel metal1 s 17712 28190 17712 28190 4 vdd
port 513 nsew
rlabel metal1 s 17712 26319 17712 26319 4 vdd
port 513 nsew
rlabel metal1 s 17712 27109 17712 27109 4 vdd
port 513 nsew
rlabel metal1 s 18816 25280 18816 25280 4 bl0_30
port 121 nsew
rlabel metal1 s 19584 25280 19584 25280 4 br1_31
port 128 nsew
rlabel metal1 s 19728 23949 19728 23949 4 vdd
port 513 nsew
rlabel metal1 s 18624 25280 18624 25280 4 bl0_29
port 117 nsew
rlabel metal1 s 17712 24240 17712 24240 4 vdd
port 513 nsew
rlabel metal1 s 18960 24240 18960 24240 4 vdd
port 513 nsew
rlabel metal1 s 19800 25280 19800 25280 4 br0_31
port 126 nsew
rlabel metal1 s 18480 23949 18480 23949 4 vdd
port 513 nsew
rlabel metal1 s 18888 25280 18888 25280 4 br0_30
port 122 nsew
rlabel metal1 s 18480 24739 18480 24739 4 vdd
port 513 nsew
rlabel metal1 s 18336 25280 18336 25280 4 br1_29
port 120 nsew
rlabel metal1 s 17712 22369 17712 22369 4 vdd
port 513 nsew
rlabel metal1 s 19728 24240 19728 24240 4 vdd
port 513 nsew
rlabel metal1 s 18960 23159 18960 23159 4 vdd
port 513 nsew
rlabel metal1 s 19728 22369 19728 22369 4 vdd
port 513 nsew
rlabel metal1 s 19728 22660 19728 22660 4 vdd
port 513 nsew
rlabel metal1 s 18960 22660 18960 22660 4 vdd
port 513 nsew
rlabel metal1 s 18480 23450 18480 23450 4 vdd
port 513 nsew
rlabel metal1 s 17640 25280 17640 25280 4 br0_28
port 114 nsew
rlabel metal1 s 18960 24739 18960 24739 4 vdd
port 513 nsew
rlabel metal1 s 17712 24739 17712 24739 4 vdd
port 513 nsew
rlabel metal1 s 19728 24739 19728 24739 4 vdd
port 513 nsew
rlabel metal1 s 19656 25280 19656 25280 4 bl1_31
port 127 nsew
rlabel metal1 s 18480 23159 18480 23159 4 vdd
port 513 nsew
rlabel metal1 s 18480 22660 18480 22660 4 vdd
port 513 nsew
rlabel metal1 s 18960 22369 18960 22369 4 vdd
port 513 nsew
rlabel metal1 s 17712 23159 17712 23159 4 vdd
port 513 nsew
rlabel metal1 s 17856 25280 17856 25280 4 br1_28
port 116 nsew
rlabel metal1 s 19104 25280 19104 25280 4 br1_30
port 124 nsew
rlabel metal1 s 17712 23949 17712 23949 4 vdd
port 513 nsew
rlabel metal1 s 17712 23450 17712 23450 4 vdd
port 513 nsew
rlabel metal1 s 17712 25030 17712 25030 4 vdd
port 513 nsew
rlabel metal1 s 19032 25280 19032 25280 4 bl1_30
port 123 nsew
rlabel metal1 s 17712 22660 17712 22660 4 vdd
port 513 nsew
rlabel metal1 s 18960 25030 18960 25030 4 vdd
port 513 nsew
rlabel metal1 s 19728 25030 19728 25030 4 vdd
port 513 nsew
rlabel metal1 s 18960 23450 18960 23450 4 vdd
port 513 nsew
rlabel metal1 s 18480 24240 18480 24240 4 vdd
port 513 nsew
rlabel metal1 s 19728 23159 19728 23159 4 vdd
port 513 nsew
rlabel metal1 s 19872 25280 19872 25280 4 bl0_31
port 125 nsew
rlabel metal1 s 18960 23949 18960 23949 4 vdd
port 513 nsew
rlabel metal1 s 18480 25030 18480 25030 4 vdd
port 513 nsew
rlabel metal1 s 18480 22369 18480 22369 4 vdd
port 513 nsew
rlabel metal1 s 19728 23450 19728 23450 4 vdd
port 513 nsew
rlabel metal1 s 18408 25280 18408 25280 4 bl1_29
port 119 nsew
rlabel metal1 s 17784 25280 17784 25280 4 bl1_28
port 115 nsew
rlabel metal1 s 18552 25280 18552 25280 4 br0_29
port 118 nsew
rlabel metal1 s 17568 25280 17568 25280 4 bl0_28
port 113 nsew
rlabel metal1 s 16464 22369 16464 22369 4 vdd
port 513 nsew
rlabel metal1 s 17232 24240 17232 24240 4 vdd
port 513 nsew
rlabel metal1 s 15216 25030 15216 25030 4 vdd
port 513 nsew
rlabel metal1 s 17232 23949 17232 23949 4 vdd
port 513 nsew
rlabel metal1 s 17160 25280 17160 25280 4 bl1_27
port 111 nsew
rlabel metal1 s 16536 25280 16536 25280 4 bl1_26
port 107 nsew
rlabel metal1 s 15984 22369 15984 22369 4 vdd
port 513 nsew
rlabel metal1 s 16464 23159 16464 23159 4 vdd
port 513 nsew
rlabel metal1 s 17304 25280 17304 25280 4 br0_27
port 110 nsew
rlabel metal1 s 16464 23450 16464 23450 4 vdd
port 513 nsew
rlabel metal1 s 16392 25280 16392 25280 4 br0_26
port 106 nsew
rlabel metal1 s 17232 22369 17232 22369 4 vdd
port 513 nsew
rlabel metal1 s 16056 25280 16056 25280 4 br0_25
port 102 nsew
rlabel metal1 s 15984 22660 15984 22660 4 vdd
port 513 nsew
rlabel metal1 s 17232 22660 17232 22660 4 vdd
port 513 nsew
rlabel metal1 s 15840 25280 15840 25280 4 br1_25
port 104 nsew
rlabel metal1 s 15144 25280 15144 25280 4 br0_24
port 98 nsew
rlabel metal1 s 15216 24240 15216 24240 4 vdd
port 513 nsew
rlabel metal1 s 15072 25280 15072 25280 4 bl0_24
port 97 nsew
rlabel metal1 s 15984 23949 15984 23949 4 vdd
port 513 nsew
rlabel metal1 s 17232 24739 17232 24739 4 vdd
port 513 nsew
rlabel metal1 s 16464 24240 16464 24240 4 vdd
port 513 nsew
rlabel metal1 s 17232 23450 17232 23450 4 vdd
port 513 nsew
rlabel metal1 s 17376 25280 17376 25280 4 bl0_27
port 109 nsew
rlabel metal1 s 17232 25030 17232 25030 4 vdd
port 513 nsew
rlabel metal1 s 16464 22660 16464 22660 4 vdd
port 513 nsew
rlabel metal1 s 15984 24240 15984 24240 4 vdd
port 513 nsew
rlabel metal1 s 16464 25030 16464 25030 4 vdd
port 513 nsew
rlabel metal1 s 15360 25280 15360 25280 4 br1_24
port 100 nsew
rlabel metal1 s 17232 23159 17232 23159 4 vdd
port 513 nsew
rlabel metal1 s 15216 23450 15216 23450 4 vdd
port 513 nsew
rlabel metal1 s 15216 22660 15216 22660 4 vdd
port 513 nsew
rlabel metal1 s 15216 24739 15216 24739 4 vdd
port 513 nsew
rlabel metal1 s 16128 25280 16128 25280 4 bl0_25
port 101 nsew
rlabel metal1 s 15984 25030 15984 25030 4 vdd
port 513 nsew
rlabel metal1 s 15216 23159 15216 23159 4 vdd
port 513 nsew
rlabel metal1 s 15288 25280 15288 25280 4 bl1_24
port 99 nsew
rlabel metal1 s 16464 24739 16464 24739 4 vdd
port 513 nsew
rlabel metal1 s 16320 25280 16320 25280 4 bl0_26
port 105 nsew
rlabel metal1 s 15984 23450 15984 23450 4 vdd
port 513 nsew
rlabel metal1 s 15984 24739 15984 24739 4 vdd
port 513 nsew
rlabel metal1 s 16464 23949 16464 23949 4 vdd
port 513 nsew
rlabel metal1 s 15984 23159 15984 23159 4 vdd
port 513 nsew
rlabel metal1 s 17088 25280 17088 25280 4 br1_27
port 112 nsew
rlabel metal1 s 16608 25280 16608 25280 4 br1_26
port 108 nsew
rlabel metal1 s 15216 22369 15216 22369 4 vdd
port 513 nsew
rlabel metal1 s 15912 25280 15912 25280 4 bl1_25
port 103 nsew
rlabel metal1 s 15216 23949 15216 23949 4 vdd
port 513 nsew
rlabel metal1 s 17232 19209 17232 19209 4 vdd
port 513 nsew
rlabel metal1 s 16464 21870 16464 21870 4 vdd
port 513 nsew
rlabel metal1 s 15984 20789 15984 20789 4 vdd
port 513 nsew
rlabel metal1 s 15984 20290 15984 20290 4 vdd
port 513 nsew
rlabel metal1 s 17232 20290 17232 20290 4 vdd
port 513 nsew
rlabel metal1 s 15984 19500 15984 19500 4 vdd
port 513 nsew
rlabel metal1 s 15984 19999 15984 19999 4 vdd
port 513 nsew
rlabel metal1 s 17232 21579 17232 21579 4 vdd
port 513 nsew
rlabel metal1 s 15984 21579 15984 21579 4 vdd
port 513 nsew
rlabel metal1 s 17232 19999 17232 19999 4 vdd
port 513 nsew
rlabel metal1 s 17232 20789 17232 20789 4 vdd
port 513 nsew
rlabel metal1 s 15216 21870 15216 21870 4 vdd
port 513 nsew
rlabel metal1 s 17232 19500 17232 19500 4 vdd
port 513 nsew
rlabel metal1 s 15984 21870 15984 21870 4 vdd
port 513 nsew
rlabel metal1 s 16464 20789 16464 20789 4 vdd
port 513 nsew
rlabel metal1 s 17232 21080 17232 21080 4 vdd
port 513 nsew
rlabel metal1 s 16464 20290 16464 20290 4 vdd
port 513 nsew
rlabel metal1 s 16464 21080 16464 21080 4 vdd
port 513 nsew
rlabel metal1 s 15984 21080 15984 21080 4 vdd
port 513 nsew
rlabel metal1 s 17232 21870 17232 21870 4 vdd
port 513 nsew
rlabel metal1 s 16464 19209 16464 19209 4 vdd
port 513 nsew
rlabel metal1 s 15216 21080 15216 21080 4 vdd
port 513 nsew
rlabel metal1 s 15216 21579 15216 21579 4 vdd
port 513 nsew
rlabel metal1 s 15984 19209 15984 19209 4 vdd
port 513 nsew
rlabel metal1 s 15216 20290 15216 20290 4 vdd
port 513 nsew
rlabel metal1 s 15216 19500 15216 19500 4 vdd
port 513 nsew
rlabel metal1 s 15216 19999 15216 19999 4 vdd
port 513 nsew
rlabel metal1 s 16464 21579 16464 21579 4 vdd
port 513 nsew
rlabel metal1 s 16464 19500 16464 19500 4 vdd
port 513 nsew
rlabel metal1 s 16464 19999 16464 19999 4 vdd
port 513 nsew
rlabel metal1 s 15216 20789 15216 20789 4 vdd
port 513 nsew
rlabel metal1 s 15216 19209 15216 19209 4 vdd
port 513 nsew
rlabel metal1 s 18960 21870 18960 21870 4 vdd
port 513 nsew
rlabel metal1 s 18960 21579 18960 21579 4 vdd
port 513 nsew
rlabel metal1 s 19728 20290 19728 20290 4 vdd
port 513 nsew
rlabel metal1 s 17712 19209 17712 19209 4 vdd
port 513 nsew
rlabel metal1 s 17712 19999 17712 19999 4 vdd
port 513 nsew
rlabel metal1 s 18480 21080 18480 21080 4 vdd
port 513 nsew
rlabel metal1 s 18960 19500 18960 19500 4 vdd
port 513 nsew
rlabel metal1 s 17712 21579 17712 21579 4 vdd
port 513 nsew
rlabel metal1 s 18960 20789 18960 20789 4 vdd
port 513 nsew
rlabel metal1 s 19728 21080 19728 21080 4 vdd
port 513 nsew
rlabel metal1 s 17712 21870 17712 21870 4 vdd
port 513 nsew
rlabel metal1 s 18960 21080 18960 21080 4 vdd
port 513 nsew
rlabel metal1 s 18960 19999 18960 19999 4 vdd
port 513 nsew
rlabel metal1 s 17712 19500 17712 19500 4 vdd
port 513 nsew
rlabel metal1 s 19728 19500 19728 19500 4 vdd
port 513 nsew
rlabel metal1 s 18480 21579 18480 21579 4 vdd
port 513 nsew
rlabel metal1 s 19728 20789 19728 20789 4 vdd
port 513 nsew
rlabel metal1 s 18480 21870 18480 21870 4 vdd
port 513 nsew
rlabel metal1 s 18480 19999 18480 19999 4 vdd
port 513 nsew
rlabel metal1 s 18960 19209 18960 19209 4 vdd
port 513 nsew
rlabel metal1 s 17712 20290 17712 20290 4 vdd
port 513 nsew
rlabel metal1 s 19728 21579 19728 21579 4 vdd
port 513 nsew
rlabel metal1 s 19728 19209 19728 19209 4 vdd
port 513 nsew
rlabel metal1 s 18960 20290 18960 20290 4 vdd
port 513 nsew
rlabel metal1 s 18480 20789 18480 20789 4 vdd
port 513 nsew
rlabel metal1 s 17712 20789 17712 20789 4 vdd
port 513 nsew
rlabel metal1 s 19728 19999 19728 19999 4 vdd
port 513 nsew
rlabel metal1 s 18480 20290 18480 20290 4 vdd
port 513 nsew
rlabel metal1 s 17712 21080 17712 21080 4 vdd
port 513 nsew
rlabel metal1 s 19728 21870 19728 21870 4 vdd
port 513 nsew
rlabel metal1 s 18480 19209 18480 19209 4 vdd
port 513 nsew
rlabel metal1 s 18480 19500 18480 19500 4 vdd
port 513 nsew
rlabel metal1 s 13968 23159 13968 23159 4 vdd
port 513 nsew
rlabel metal1 s 13968 23949 13968 23949 4 vdd
port 513 nsew
rlabel metal1 s 13488 22369 13488 22369 4 vdd
port 513 nsew
rlabel metal1 s 14736 23159 14736 23159 4 vdd
port 513 nsew
rlabel metal1 s 12720 23949 12720 23949 4 vdd
port 513 nsew
rlabel metal1 s 13968 25030 13968 25030 4 vdd
port 513 nsew
rlabel metal1 s 14040 25280 14040 25280 4 bl1_22
port 91 nsew
rlabel metal1 s 14736 22660 14736 22660 4 vdd
port 513 nsew
rlabel metal1 s 14736 23450 14736 23450 4 vdd
port 513 nsew
rlabel metal1 s 12720 22660 12720 22660 4 vdd
port 513 nsew
rlabel metal1 s 13344 25280 13344 25280 4 br1_21
port 88 nsew
rlabel metal1 s 14736 22369 14736 22369 4 vdd
port 513 nsew
rlabel metal1 s 14736 23949 14736 23949 4 vdd
port 513 nsew
rlabel metal1 s 13560 25280 13560 25280 4 br0_21
port 86 nsew
rlabel metal1 s 13968 24739 13968 24739 4 vdd
port 513 nsew
rlabel metal1 s 13896 25280 13896 25280 4 br0_22
port 90 nsew
rlabel metal1 s 13488 23450 13488 23450 4 vdd
port 513 nsew
rlabel metal1 s 13488 23159 13488 23159 4 vdd
port 513 nsew
rlabel metal1 s 12648 25280 12648 25280 4 br0_20
port 82 nsew
rlabel metal1 s 13488 25030 13488 25030 4 vdd
port 513 nsew
rlabel metal1 s 13416 25280 13416 25280 4 bl1_21
port 87 nsew
rlabel metal1 s 14736 25030 14736 25030 4 vdd
port 513 nsew
rlabel metal1 s 14112 25280 14112 25280 4 br1_22
port 92 nsew
rlabel metal1 s 13968 22369 13968 22369 4 vdd
port 513 nsew
rlabel metal1 s 12720 22369 12720 22369 4 vdd
port 513 nsew
rlabel metal1 s 14592 25280 14592 25280 4 br1_23
port 96 nsew
rlabel metal1 s 13488 22660 13488 22660 4 vdd
port 513 nsew
rlabel metal1 s 13968 23450 13968 23450 4 vdd
port 513 nsew
rlabel metal1 s 13488 24739 13488 24739 4 vdd
port 513 nsew
rlabel metal1 s 13968 24240 13968 24240 4 vdd
port 513 nsew
rlabel metal1 s 14736 24240 14736 24240 4 vdd
port 513 nsew
rlabel metal1 s 13488 24240 13488 24240 4 vdd
port 513 nsew
rlabel metal1 s 12720 23450 12720 23450 4 vdd
port 513 nsew
rlabel metal1 s 12720 25030 12720 25030 4 vdd
port 513 nsew
rlabel metal1 s 12720 24739 12720 24739 4 vdd
port 513 nsew
rlabel metal1 s 13632 25280 13632 25280 4 bl0_21
port 85 nsew
rlabel metal1 s 14880 25280 14880 25280 4 bl0_23
port 93 nsew
rlabel metal1 s 12792 25280 12792 25280 4 bl1_20
port 83 nsew
rlabel metal1 s 12720 24240 12720 24240 4 vdd
port 513 nsew
rlabel metal1 s 14736 24739 14736 24739 4 vdd
port 513 nsew
rlabel metal1 s 12720 23159 12720 23159 4 vdd
port 513 nsew
rlabel metal1 s 13488 23949 13488 23949 4 vdd
port 513 nsew
rlabel metal1 s 14664 25280 14664 25280 4 bl1_23
port 95 nsew
rlabel metal1 s 14808 25280 14808 25280 4 br0_23
port 94 nsew
rlabel metal1 s 12576 25280 12576 25280 4 bl0_20
port 81 nsew
rlabel metal1 s 13968 22660 13968 22660 4 vdd
port 513 nsew
rlabel metal1 s 13824 25280 13824 25280 4 bl0_22
port 89 nsew
rlabel metal1 s 12864 25280 12864 25280 4 br1_20
port 84 nsew
rlabel metal1 s 10992 25030 10992 25030 4 vdd
port 513 nsew
rlabel metal1 s 11472 23450 11472 23450 4 vdd
port 513 nsew
rlabel metal1 s 10296 25280 10296 25280 4 bl1_16
port 67 nsew
rlabel metal1 s 12240 23450 12240 23450 4 vdd
port 513 nsew
rlabel metal1 s 12240 22660 12240 22660 4 vdd
port 513 nsew
rlabel metal1 s 10224 24739 10224 24739 4 vdd
port 513 nsew
rlabel metal1 s 12240 23949 12240 23949 4 vdd
port 513 nsew
rlabel metal1 s 12240 25030 12240 25030 4 vdd
port 513 nsew
rlabel metal1 s 10224 22660 10224 22660 4 vdd
port 513 nsew
rlabel metal1 s 10224 23949 10224 23949 4 vdd
port 513 nsew
rlabel metal1 s 11472 23949 11472 23949 4 vdd
port 513 nsew
rlabel metal1 s 10224 23450 10224 23450 4 vdd
port 513 nsew
rlabel metal1 s 11472 22369 11472 22369 4 vdd
port 513 nsew
rlabel metal1 s 11472 23159 11472 23159 4 vdd
port 513 nsew
rlabel metal1 s 11472 24739 11472 24739 4 vdd
port 513 nsew
rlabel metal1 s 10992 22369 10992 22369 4 vdd
port 513 nsew
rlabel metal1 s 12168 25280 12168 25280 4 bl1_19
port 79 nsew
rlabel metal1 s 11400 25280 11400 25280 4 br0_18
port 74 nsew
rlabel metal1 s 12240 24739 12240 24739 4 vdd
port 513 nsew
rlabel metal1 s 11064 25280 11064 25280 4 br0_17
port 70 nsew
rlabel metal1 s 11136 25280 11136 25280 4 bl0_17
port 69 nsew
rlabel metal1 s 12240 22369 12240 22369 4 vdd
port 513 nsew
rlabel metal1 s 10152 25280 10152 25280 4 br0_16
port 66 nsew
rlabel metal1 s 11472 24240 11472 24240 4 vdd
port 513 nsew
rlabel metal1 s 10848 25280 10848 25280 4 br1_17
port 72 nsew
rlabel metal1 s 10080 25280 10080 25280 4 bl0_16
port 65 nsew
rlabel metal1 s 11472 25030 11472 25030 4 vdd
port 513 nsew
rlabel metal1 s 12312 25280 12312 25280 4 br0_19
port 78 nsew
rlabel metal1 s 10920 25280 10920 25280 4 bl1_17
port 71 nsew
rlabel metal1 s 10224 25030 10224 25030 4 vdd
port 513 nsew
rlabel metal1 s 11616 25280 11616 25280 4 br1_18
port 76 nsew
rlabel metal1 s 12384 25280 12384 25280 4 bl0_19
port 77 nsew
rlabel metal1 s 10992 22660 10992 22660 4 vdd
port 513 nsew
rlabel metal1 s 10224 24240 10224 24240 4 vdd
port 513 nsew
rlabel metal1 s 12240 24240 12240 24240 4 vdd
port 513 nsew
rlabel metal1 s 10992 23159 10992 23159 4 vdd
port 513 nsew
rlabel metal1 s 10992 24240 10992 24240 4 vdd
port 513 nsew
rlabel metal1 s 12240 23159 12240 23159 4 vdd
port 513 nsew
rlabel metal1 s 10368 25280 10368 25280 4 br1_16
port 68 nsew
rlabel metal1 s 10992 23949 10992 23949 4 vdd
port 513 nsew
rlabel metal1 s 11544 25280 11544 25280 4 bl1_18
port 75 nsew
rlabel metal1 s 10224 23159 10224 23159 4 vdd
port 513 nsew
rlabel metal1 s 11472 22660 11472 22660 4 vdd
port 513 nsew
rlabel metal1 s 10992 23450 10992 23450 4 vdd
port 513 nsew
rlabel metal1 s 11328 25280 11328 25280 4 bl0_18
port 73 nsew
rlabel metal1 s 10992 24739 10992 24739 4 vdd
port 513 nsew
rlabel metal1 s 12096 25280 12096 25280 4 br1_19
port 80 nsew
rlabel metal1 s 10224 22369 10224 22369 4 vdd
port 513 nsew
rlabel metal1 s 12240 20789 12240 20789 4 vdd
port 513 nsew
rlabel metal1 s 11472 19500 11472 19500 4 vdd
port 513 nsew
rlabel metal1 s 10224 19500 10224 19500 4 vdd
port 513 nsew
rlabel metal1 s 10224 20290 10224 20290 4 vdd
port 513 nsew
rlabel metal1 s 11472 21870 11472 21870 4 vdd
port 513 nsew
rlabel metal1 s 11472 20290 11472 20290 4 vdd
port 513 nsew
rlabel metal1 s 10992 19209 10992 19209 4 vdd
port 513 nsew
rlabel metal1 s 12240 20290 12240 20290 4 vdd
port 513 nsew
rlabel metal1 s 12240 21080 12240 21080 4 vdd
port 513 nsew
rlabel metal1 s 11472 19209 11472 19209 4 vdd
port 513 nsew
rlabel metal1 s 10992 21870 10992 21870 4 vdd
port 513 nsew
rlabel metal1 s 12240 21870 12240 21870 4 vdd
port 513 nsew
rlabel metal1 s 12240 19500 12240 19500 4 vdd
port 513 nsew
rlabel metal1 s 10224 19209 10224 19209 4 vdd
port 513 nsew
rlabel metal1 s 11472 19999 11472 19999 4 vdd
port 513 nsew
rlabel metal1 s 10992 19500 10992 19500 4 vdd
port 513 nsew
rlabel metal1 s 10224 19999 10224 19999 4 vdd
port 513 nsew
rlabel metal1 s 10992 21080 10992 21080 4 vdd
port 513 nsew
rlabel metal1 s 11472 21579 11472 21579 4 vdd
port 513 nsew
rlabel metal1 s 12240 19999 12240 19999 4 vdd
port 513 nsew
rlabel metal1 s 10992 21579 10992 21579 4 vdd
port 513 nsew
rlabel metal1 s 12240 21579 12240 21579 4 vdd
port 513 nsew
rlabel metal1 s 10992 19999 10992 19999 4 vdd
port 513 nsew
rlabel metal1 s 10224 21080 10224 21080 4 vdd
port 513 nsew
rlabel metal1 s 10992 20789 10992 20789 4 vdd
port 513 nsew
rlabel metal1 s 11472 20789 11472 20789 4 vdd
port 513 nsew
rlabel metal1 s 10224 21870 10224 21870 4 vdd
port 513 nsew
rlabel metal1 s 12240 19209 12240 19209 4 vdd
port 513 nsew
rlabel metal1 s 10224 21579 10224 21579 4 vdd
port 513 nsew
rlabel metal1 s 11472 21080 11472 21080 4 vdd
port 513 nsew
rlabel metal1 s 10992 20290 10992 20290 4 vdd
port 513 nsew
rlabel metal1 s 10224 20789 10224 20789 4 vdd
port 513 nsew
rlabel metal1 s 14736 20290 14736 20290 4 vdd
port 513 nsew
rlabel metal1 s 13968 21579 13968 21579 4 vdd
port 513 nsew
rlabel metal1 s 12720 21579 12720 21579 4 vdd
port 513 nsew
rlabel metal1 s 12720 19209 12720 19209 4 vdd
port 513 nsew
rlabel metal1 s 13488 20290 13488 20290 4 vdd
port 513 nsew
rlabel metal1 s 12720 19500 12720 19500 4 vdd
port 513 nsew
rlabel metal1 s 13968 21080 13968 21080 4 vdd
port 513 nsew
rlabel metal1 s 14736 21870 14736 21870 4 vdd
port 513 nsew
rlabel metal1 s 13968 19999 13968 19999 4 vdd
port 513 nsew
rlabel metal1 s 14736 20789 14736 20789 4 vdd
port 513 nsew
rlabel metal1 s 12720 21870 12720 21870 4 vdd
port 513 nsew
rlabel metal1 s 13488 21579 13488 21579 4 vdd
port 513 nsew
rlabel metal1 s 13968 21870 13968 21870 4 vdd
port 513 nsew
rlabel metal1 s 12720 20290 12720 20290 4 vdd
port 513 nsew
rlabel metal1 s 13968 19500 13968 19500 4 vdd
port 513 nsew
rlabel metal1 s 14736 19209 14736 19209 4 vdd
port 513 nsew
rlabel metal1 s 13488 20789 13488 20789 4 vdd
port 513 nsew
rlabel metal1 s 13488 19999 13488 19999 4 vdd
port 513 nsew
rlabel metal1 s 13968 20789 13968 20789 4 vdd
port 513 nsew
rlabel metal1 s 13488 19500 13488 19500 4 vdd
port 513 nsew
rlabel metal1 s 13488 19209 13488 19209 4 vdd
port 513 nsew
rlabel metal1 s 14736 21579 14736 21579 4 vdd
port 513 nsew
rlabel metal1 s 13968 20290 13968 20290 4 vdd
port 513 nsew
rlabel metal1 s 14736 19999 14736 19999 4 vdd
port 513 nsew
rlabel metal1 s 14736 21080 14736 21080 4 vdd
port 513 nsew
rlabel metal1 s 12720 21080 12720 21080 4 vdd
port 513 nsew
rlabel metal1 s 13488 21870 13488 21870 4 vdd
port 513 nsew
rlabel metal1 s 12720 19999 12720 19999 4 vdd
port 513 nsew
rlabel metal1 s 12720 20789 12720 20789 4 vdd
port 513 nsew
rlabel metal1 s 13488 21080 13488 21080 4 vdd
port 513 nsew
rlabel metal1 s 13968 19209 13968 19209 4 vdd
port 513 nsew
rlabel metal1 s 14736 19500 14736 19500 4 vdd
port 513 nsew
rlabel metal1 s 13968 18710 13968 18710 4 vdd
port 513 nsew
rlabel metal1 s 12720 17629 12720 17629 4 vdd
port 513 nsew
rlabel metal1 s 12720 16839 12720 16839 4 vdd
port 513 nsew
rlabel metal1 s 13488 16839 13488 16839 4 vdd
port 513 nsew
rlabel metal1 s 13488 18419 13488 18419 4 vdd
port 513 nsew
rlabel metal1 s 13488 18710 13488 18710 4 vdd
port 513 nsew
rlabel metal1 s 12720 16049 12720 16049 4 vdd
port 513 nsew
rlabel metal1 s 13488 17130 13488 17130 4 vdd
port 513 nsew
rlabel metal1 s 13968 18419 13968 18419 4 vdd
port 513 nsew
rlabel metal1 s 13488 17629 13488 17629 4 vdd
port 513 nsew
rlabel metal1 s 13968 16839 13968 16839 4 vdd
port 513 nsew
rlabel metal1 s 14736 17130 14736 17130 4 vdd
port 513 nsew
rlabel metal1 s 13488 16049 13488 16049 4 vdd
port 513 nsew
rlabel metal1 s 12720 16340 12720 16340 4 vdd
port 513 nsew
rlabel metal1 s 12720 18419 12720 18419 4 vdd
port 513 nsew
rlabel metal1 s 13968 16049 13968 16049 4 vdd
port 513 nsew
rlabel metal1 s 14736 17629 14736 17629 4 vdd
port 513 nsew
rlabel metal1 s 12720 17920 12720 17920 4 vdd
port 513 nsew
rlabel metal1 s 13488 16340 13488 16340 4 vdd
port 513 nsew
rlabel metal1 s 14736 16340 14736 16340 4 vdd
port 513 nsew
rlabel metal1 s 14736 16839 14736 16839 4 vdd
port 513 nsew
rlabel metal1 s 13968 17920 13968 17920 4 vdd
port 513 nsew
rlabel metal1 s 14736 18710 14736 18710 4 vdd
port 513 nsew
rlabel metal1 s 13488 17920 13488 17920 4 vdd
port 513 nsew
rlabel metal1 s 13968 17629 13968 17629 4 vdd
port 513 nsew
rlabel metal1 s 14736 16049 14736 16049 4 vdd
port 513 nsew
rlabel metal1 s 12720 18710 12720 18710 4 vdd
port 513 nsew
rlabel metal1 s 13968 16340 13968 16340 4 vdd
port 513 nsew
rlabel metal1 s 14736 17920 14736 17920 4 vdd
port 513 nsew
rlabel metal1 s 12720 17130 12720 17130 4 vdd
port 513 nsew
rlabel metal1 s 14736 18419 14736 18419 4 vdd
port 513 nsew
rlabel metal1 s 13968 17130 13968 17130 4 vdd
port 513 nsew
rlabel metal1 s 10224 18419 10224 18419 4 vdd
port 513 nsew
rlabel metal1 s 10992 17130 10992 17130 4 vdd
port 513 nsew
rlabel metal1 s 11472 17629 11472 17629 4 vdd
port 513 nsew
rlabel metal1 s 10992 17629 10992 17629 4 vdd
port 513 nsew
rlabel metal1 s 10224 17629 10224 17629 4 vdd
port 513 nsew
rlabel metal1 s 12240 16340 12240 16340 4 vdd
port 513 nsew
rlabel metal1 s 11472 18710 11472 18710 4 vdd
port 513 nsew
rlabel metal1 s 12240 17920 12240 17920 4 vdd
port 513 nsew
rlabel metal1 s 11472 17920 11472 17920 4 vdd
port 513 nsew
rlabel metal1 s 12240 17130 12240 17130 4 vdd
port 513 nsew
rlabel metal1 s 11472 16340 11472 16340 4 vdd
port 513 nsew
rlabel metal1 s 10224 17130 10224 17130 4 vdd
port 513 nsew
rlabel metal1 s 12240 16839 12240 16839 4 vdd
port 513 nsew
rlabel metal1 s 10224 16340 10224 16340 4 vdd
port 513 nsew
rlabel metal1 s 10224 18710 10224 18710 4 vdd
port 513 nsew
rlabel metal1 s 10992 16049 10992 16049 4 vdd
port 513 nsew
rlabel metal1 s 11472 16049 11472 16049 4 vdd
port 513 nsew
rlabel metal1 s 10992 18419 10992 18419 4 vdd
port 513 nsew
rlabel metal1 s 11472 17130 11472 17130 4 vdd
port 513 nsew
rlabel metal1 s 10224 16049 10224 16049 4 vdd
port 513 nsew
rlabel metal1 s 10992 16839 10992 16839 4 vdd
port 513 nsew
rlabel metal1 s 11472 16839 11472 16839 4 vdd
port 513 nsew
rlabel metal1 s 12240 18419 12240 18419 4 vdd
port 513 nsew
rlabel metal1 s 10224 17920 10224 17920 4 vdd
port 513 nsew
rlabel metal1 s 10992 17920 10992 17920 4 vdd
port 513 nsew
rlabel metal1 s 10992 16340 10992 16340 4 vdd
port 513 nsew
rlabel metal1 s 12240 16049 12240 16049 4 vdd
port 513 nsew
rlabel metal1 s 12240 18710 12240 18710 4 vdd
port 513 nsew
rlabel metal1 s 10992 18710 10992 18710 4 vdd
port 513 nsew
rlabel metal1 s 10224 16839 10224 16839 4 vdd
port 513 nsew
rlabel metal1 s 11472 18419 11472 18419 4 vdd
port 513 nsew
rlabel metal1 s 12240 17629 12240 17629 4 vdd
port 513 nsew
rlabel metal1 s 10224 13679 10224 13679 4 vdd
port 513 nsew
rlabel metal1 s 10224 15259 10224 15259 4 vdd
port 513 nsew
rlabel metal1 s 11472 13679 11472 13679 4 vdd
port 513 nsew
rlabel metal1 s 12240 13180 12240 13180 4 vdd
port 513 nsew
rlabel metal1 s 10992 14469 10992 14469 4 vdd
port 513 nsew
rlabel metal1 s 12240 14760 12240 14760 4 vdd
port 513 nsew
rlabel metal1 s 10224 13970 10224 13970 4 vdd
port 513 nsew
rlabel metal1 s 12240 15259 12240 15259 4 vdd
port 513 nsew
rlabel metal1 s 12240 13970 12240 13970 4 vdd
port 513 nsew
rlabel metal1 s 11472 13970 11472 13970 4 vdd
port 513 nsew
rlabel metal1 s 10992 12889 10992 12889 4 vdd
port 513 nsew
rlabel metal1 s 10992 13970 10992 13970 4 vdd
port 513 nsew
rlabel metal1 s 11472 15550 11472 15550 4 vdd
port 513 nsew
rlabel metal1 s 12240 13679 12240 13679 4 vdd
port 513 nsew
rlabel metal1 s 10224 12889 10224 12889 4 vdd
port 513 nsew
rlabel metal1 s 12240 12889 12240 12889 4 vdd
port 513 nsew
rlabel metal1 s 10992 13180 10992 13180 4 vdd
port 513 nsew
rlabel metal1 s 10224 14469 10224 14469 4 vdd
port 513 nsew
rlabel metal1 s 12240 15550 12240 15550 4 vdd
port 513 nsew
rlabel metal1 s 11472 14760 11472 14760 4 vdd
port 513 nsew
rlabel metal1 s 12240 14469 12240 14469 4 vdd
port 513 nsew
rlabel metal1 s 10992 13679 10992 13679 4 vdd
port 513 nsew
rlabel metal1 s 10992 15550 10992 15550 4 vdd
port 513 nsew
rlabel metal1 s 10224 14760 10224 14760 4 vdd
port 513 nsew
rlabel metal1 s 11472 13180 11472 13180 4 vdd
port 513 nsew
rlabel metal1 s 11472 14469 11472 14469 4 vdd
port 513 nsew
rlabel metal1 s 11472 12889 11472 12889 4 vdd
port 513 nsew
rlabel metal1 s 10992 15259 10992 15259 4 vdd
port 513 nsew
rlabel metal1 s 11472 15259 11472 15259 4 vdd
port 513 nsew
rlabel metal1 s 10992 14760 10992 14760 4 vdd
port 513 nsew
rlabel metal1 s 10224 13180 10224 13180 4 vdd
port 513 nsew
rlabel metal1 s 10224 15550 10224 15550 4 vdd
port 513 nsew
rlabel metal1 s 14736 13970 14736 13970 4 vdd
port 513 nsew
rlabel metal1 s 14736 15550 14736 15550 4 vdd
port 513 nsew
rlabel metal1 s 13488 15259 13488 15259 4 vdd
port 513 nsew
rlabel metal1 s 14736 14469 14736 14469 4 vdd
port 513 nsew
rlabel metal1 s 14736 12889 14736 12889 4 vdd
port 513 nsew
rlabel metal1 s 12720 13970 12720 13970 4 vdd
port 513 nsew
rlabel metal1 s 13968 13679 13968 13679 4 vdd
port 513 nsew
rlabel metal1 s 12720 13180 12720 13180 4 vdd
port 513 nsew
rlabel metal1 s 13968 13970 13968 13970 4 vdd
port 513 nsew
rlabel metal1 s 14736 13679 14736 13679 4 vdd
port 513 nsew
rlabel metal1 s 13968 14760 13968 14760 4 vdd
port 513 nsew
rlabel metal1 s 13488 12889 13488 12889 4 vdd
port 513 nsew
rlabel metal1 s 13968 15550 13968 15550 4 vdd
port 513 nsew
rlabel metal1 s 12720 13679 12720 13679 4 vdd
port 513 nsew
rlabel metal1 s 13488 13180 13488 13180 4 vdd
port 513 nsew
rlabel metal1 s 13488 13970 13488 13970 4 vdd
port 513 nsew
rlabel metal1 s 12720 12889 12720 12889 4 vdd
port 513 nsew
rlabel metal1 s 13488 13679 13488 13679 4 vdd
port 513 nsew
rlabel metal1 s 12720 14469 12720 14469 4 vdd
port 513 nsew
rlabel metal1 s 14736 14760 14736 14760 4 vdd
port 513 nsew
rlabel metal1 s 13488 14469 13488 14469 4 vdd
port 513 nsew
rlabel metal1 s 12720 15550 12720 15550 4 vdd
port 513 nsew
rlabel metal1 s 13968 15259 13968 15259 4 vdd
port 513 nsew
rlabel metal1 s 14736 15259 14736 15259 4 vdd
port 513 nsew
rlabel metal1 s 13968 13180 13968 13180 4 vdd
port 513 nsew
rlabel metal1 s 12720 14760 12720 14760 4 vdd
port 513 nsew
rlabel metal1 s 14736 13180 14736 13180 4 vdd
port 513 nsew
rlabel metal1 s 13968 12889 13968 12889 4 vdd
port 513 nsew
rlabel metal1 s 13488 14760 13488 14760 4 vdd
port 513 nsew
rlabel metal1 s 12720 15259 12720 15259 4 vdd
port 513 nsew
rlabel metal1 s 13488 15550 13488 15550 4 vdd
port 513 nsew
rlabel metal1 s 13968 14469 13968 14469 4 vdd
port 513 nsew
rlabel metal1 s 18480 17130 18480 17130 4 vdd
port 513 nsew
rlabel metal1 s 19728 16340 19728 16340 4 vdd
port 513 nsew
rlabel metal1 s 18480 16340 18480 16340 4 vdd
port 513 nsew
rlabel metal1 s 18960 16340 18960 16340 4 vdd
port 513 nsew
rlabel metal1 s 18480 16049 18480 16049 4 vdd
port 513 nsew
rlabel metal1 s 17712 18710 17712 18710 4 vdd
port 513 nsew
rlabel metal1 s 18960 18419 18960 18419 4 vdd
port 513 nsew
rlabel metal1 s 18960 17920 18960 17920 4 vdd
port 513 nsew
rlabel metal1 s 17712 18419 17712 18419 4 vdd
port 513 nsew
rlabel metal1 s 19728 17629 19728 17629 4 vdd
port 513 nsew
rlabel metal1 s 18480 18419 18480 18419 4 vdd
port 513 nsew
rlabel metal1 s 19728 18419 19728 18419 4 vdd
port 513 nsew
rlabel metal1 s 17712 17920 17712 17920 4 vdd
port 513 nsew
rlabel metal1 s 18960 16049 18960 16049 4 vdd
port 513 nsew
rlabel metal1 s 17712 16340 17712 16340 4 vdd
port 513 nsew
rlabel metal1 s 17712 17629 17712 17629 4 vdd
port 513 nsew
rlabel metal1 s 18480 18710 18480 18710 4 vdd
port 513 nsew
rlabel metal1 s 18960 17130 18960 17130 4 vdd
port 513 nsew
rlabel metal1 s 18480 16839 18480 16839 4 vdd
port 513 nsew
rlabel metal1 s 18960 16839 18960 16839 4 vdd
port 513 nsew
rlabel metal1 s 17712 17130 17712 17130 4 vdd
port 513 nsew
rlabel metal1 s 19728 17920 19728 17920 4 vdd
port 513 nsew
rlabel metal1 s 19728 16049 19728 16049 4 vdd
port 513 nsew
rlabel metal1 s 19728 17130 19728 17130 4 vdd
port 513 nsew
rlabel metal1 s 18480 17920 18480 17920 4 vdd
port 513 nsew
rlabel metal1 s 18960 18710 18960 18710 4 vdd
port 513 nsew
rlabel metal1 s 17712 16049 17712 16049 4 vdd
port 513 nsew
rlabel metal1 s 18480 17629 18480 17629 4 vdd
port 513 nsew
rlabel metal1 s 18960 17629 18960 17629 4 vdd
port 513 nsew
rlabel metal1 s 17712 16839 17712 16839 4 vdd
port 513 nsew
rlabel metal1 s 19728 18710 19728 18710 4 vdd
port 513 nsew
rlabel metal1 s 19728 16839 19728 16839 4 vdd
port 513 nsew
rlabel metal1 s 15216 18710 15216 18710 4 vdd
port 513 nsew
rlabel metal1 s 17232 18710 17232 18710 4 vdd
port 513 nsew
rlabel metal1 s 16464 16839 16464 16839 4 vdd
port 513 nsew
rlabel metal1 s 17232 16839 17232 16839 4 vdd
port 513 nsew
rlabel metal1 s 17232 17629 17232 17629 4 vdd
port 513 nsew
rlabel metal1 s 17232 17920 17232 17920 4 vdd
port 513 nsew
rlabel metal1 s 15216 17130 15216 17130 4 vdd
port 513 nsew
rlabel metal1 s 16464 18419 16464 18419 4 vdd
port 513 nsew
rlabel metal1 s 16464 16049 16464 16049 4 vdd
port 513 nsew
rlabel metal1 s 17232 16340 17232 16340 4 vdd
port 513 nsew
rlabel metal1 s 15984 17130 15984 17130 4 vdd
port 513 nsew
rlabel metal1 s 17232 18419 17232 18419 4 vdd
port 513 nsew
rlabel metal1 s 15984 16839 15984 16839 4 vdd
port 513 nsew
rlabel metal1 s 15216 17629 15216 17629 4 vdd
port 513 nsew
rlabel metal1 s 16464 17130 16464 17130 4 vdd
port 513 nsew
rlabel metal1 s 15216 16049 15216 16049 4 vdd
port 513 nsew
rlabel metal1 s 15984 18710 15984 18710 4 vdd
port 513 nsew
rlabel metal1 s 15216 16340 15216 16340 4 vdd
port 513 nsew
rlabel metal1 s 17232 16049 17232 16049 4 vdd
port 513 nsew
rlabel metal1 s 15984 16049 15984 16049 4 vdd
port 513 nsew
rlabel metal1 s 16464 16340 16464 16340 4 vdd
port 513 nsew
rlabel metal1 s 15216 16839 15216 16839 4 vdd
port 513 nsew
rlabel metal1 s 15984 17920 15984 17920 4 vdd
port 513 nsew
rlabel metal1 s 15984 18419 15984 18419 4 vdd
port 513 nsew
rlabel metal1 s 15216 18419 15216 18419 4 vdd
port 513 nsew
rlabel metal1 s 16464 17920 16464 17920 4 vdd
port 513 nsew
rlabel metal1 s 17232 17130 17232 17130 4 vdd
port 513 nsew
rlabel metal1 s 15216 17920 15216 17920 4 vdd
port 513 nsew
rlabel metal1 s 15984 16340 15984 16340 4 vdd
port 513 nsew
rlabel metal1 s 16464 18710 16464 18710 4 vdd
port 513 nsew
rlabel metal1 s 16464 17629 16464 17629 4 vdd
port 513 nsew
rlabel metal1 s 15984 17629 15984 17629 4 vdd
port 513 nsew
rlabel metal1 s 16464 13970 16464 13970 4 vdd
port 513 nsew
rlabel metal1 s 15984 13970 15984 13970 4 vdd
port 513 nsew
rlabel metal1 s 17232 12889 17232 12889 4 vdd
port 513 nsew
rlabel metal1 s 15984 13679 15984 13679 4 vdd
port 513 nsew
rlabel metal1 s 16464 12889 16464 12889 4 vdd
port 513 nsew
rlabel metal1 s 15216 15550 15216 15550 4 vdd
port 513 nsew
rlabel metal1 s 15984 15550 15984 15550 4 vdd
port 513 nsew
rlabel metal1 s 15216 14469 15216 14469 4 vdd
port 513 nsew
rlabel metal1 s 16464 14469 16464 14469 4 vdd
port 513 nsew
rlabel metal1 s 15984 14469 15984 14469 4 vdd
port 513 nsew
rlabel metal1 s 17232 14469 17232 14469 4 vdd
port 513 nsew
rlabel metal1 s 15984 15259 15984 15259 4 vdd
port 513 nsew
rlabel metal1 s 16464 14760 16464 14760 4 vdd
port 513 nsew
rlabel metal1 s 16464 13679 16464 13679 4 vdd
port 513 nsew
rlabel metal1 s 15216 13679 15216 13679 4 vdd
port 513 nsew
rlabel metal1 s 16464 13180 16464 13180 4 vdd
port 513 nsew
rlabel metal1 s 17232 15259 17232 15259 4 vdd
port 513 nsew
rlabel metal1 s 17232 15550 17232 15550 4 vdd
port 513 nsew
rlabel metal1 s 17232 13679 17232 13679 4 vdd
port 513 nsew
rlabel metal1 s 15216 13180 15216 13180 4 vdd
port 513 nsew
rlabel metal1 s 17232 14760 17232 14760 4 vdd
port 513 nsew
rlabel metal1 s 17232 13970 17232 13970 4 vdd
port 513 nsew
rlabel metal1 s 15216 15259 15216 15259 4 vdd
port 513 nsew
rlabel metal1 s 16464 15259 16464 15259 4 vdd
port 513 nsew
rlabel metal1 s 15984 13180 15984 13180 4 vdd
port 513 nsew
rlabel metal1 s 15984 12889 15984 12889 4 vdd
port 513 nsew
rlabel metal1 s 15216 13970 15216 13970 4 vdd
port 513 nsew
rlabel metal1 s 17232 13180 17232 13180 4 vdd
port 513 nsew
rlabel metal1 s 15984 14760 15984 14760 4 vdd
port 513 nsew
rlabel metal1 s 15216 12889 15216 12889 4 vdd
port 513 nsew
rlabel metal1 s 15216 14760 15216 14760 4 vdd
port 513 nsew
rlabel metal1 s 16464 15550 16464 15550 4 vdd
port 513 nsew
rlabel metal1 s 19728 14469 19728 14469 4 vdd
port 513 nsew
rlabel metal1 s 18480 15550 18480 15550 4 vdd
port 513 nsew
rlabel metal1 s 18960 14760 18960 14760 4 vdd
port 513 nsew
rlabel metal1 s 17712 13970 17712 13970 4 vdd
port 513 nsew
rlabel metal1 s 18480 12889 18480 12889 4 vdd
port 513 nsew
rlabel metal1 s 18960 15550 18960 15550 4 vdd
port 513 nsew
rlabel metal1 s 19728 12889 19728 12889 4 vdd
port 513 nsew
rlabel metal1 s 18480 14760 18480 14760 4 vdd
port 513 nsew
rlabel metal1 s 18480 14469 18480 14469 4 vdd
port 513 nsew
rlabel metal1 s 17712 13180 17712 13180 4 vdd
port 513 nsew
rlabel metal1 s 17712 13679 17712 13679 4 vdd
port 513 nsew
rlabel metal1 s 19728 13679 19728 13679 4 vdd
port 513 nsew
rlabel metal1 s 17712 12889 17712 12889 4 vdd
port 513 nsew
rlabel metal1 s 19728 13180 19728 13180 4 vdd
port 513 nsew
rlabel metal1 s 18960 12889 18960 12889 4 vdd
port 513 nsew
rlabel metal1 s 18480 13970 18480 13970 4 vdd
port 513 nsew
rlabel metal1 s 19728 15550 19728 15550 4 vdd
port 513 nsew
rlabel metal1 s 18960 13180 18960 13180 4 vdd
port 513 nsew
rlabel metal1 s 18480 15259 18480 15259 4 vdd
port 513 nsew
rlabel metal1 s 18960 13970 18960 13970 4 vdd
port 513 nsew
rlabel metal1 s 17712 15259 17712 15259 4 vdd
port 513 nsew
rlabel metal1 s 18960 15259 18960 15259 4 vdd
port 513 nsew
rlabel metal1 s 18960 14469 18960 14469 4 vdd
port 513 nsew
rlabel metal1 s 19728 13970 19728 13970 4 vdd
port 513 nsew
rlabel metal1 s 19728 15259 19728 15259 4 vdd
port 513 nsew
rlabel metal1 s 19728 14760 19728 14760 4 vdd
port 513 nsew
rlabel metal1 s 17712 15550 17712 15550 4 vdd
port 513 nsew
rlabel metal1 s 17712 14760 17712 14760 4 vdd
port 513 nsew
rlabel metal1 s 18480 13679 18480 13679 4 vdd
port 513 nsew
rlabel metal1 s 17712 14469 17712 14469 4 vdd
port 513 nsew
rlabel metal1 s 18480 13180 18480 13180 4 vdd
port 513 nsew
rlabel metal1 s 18960 13679 18960 13679 4 vdd
port 513 nsew
rlabel metal1 s 8496 25030 8496 25030 4 vdd
port 513 nsew
rlabel metal1 s 7872 25280 7872 25280 4 br1_12
port 52 nsew
rlabel metal1 s 9744 22660 9744 22660 4 vdd
port 513 nsew
rlabel metal1 s 8496 22369 8496 22369 4 vdd
port 513 nsew
rlabel metal1 s 7728 24739 7728 24739 4 vdd
port 513 nsew
rlabel metal1 s 8496 24739 8496 24739 4 vdd
port 513 nsew
rlabel metal1 s 9744 25030 9744 25030 4 vdd
port 513 nsew
rlabel metal1 s 7800 25280 7800 25280 4 bl1_12
port 51 nsew
rlabel metal1 s 7656 25280 7656 25280 4 br0_12
port 50 nsew
rlabel metal1 s 9600 25280 9600 25280 4 br1_15
port 64 nsew
rlabel metal1 s 8496 22660 8496 22660 4 vdd
port 513 nsew
rlabel metal1 s 9744 23159 9744 23159 4 vdd
port 513 nsew
rlabel metal1 s 8496 24240 8496 24240 4 vdd
port 513 nsew
rlabel metal1 s 9744 22369 9744 22369 4 vdd
port 513 nsew
rlabel metal1 s 8976 22660 8976 22660 4 vdd
port 513 nsew
rlabel metal1 s 8976 22369 8976 22369 4 vdd
port 513 nsew
rlabel metal1 s 8496 23949 8496 23949 4 vdd
port 513 nsew
rlabel metal1 s 8976 23159 8976 23159 4 vdd
port 513 nsew
rlabel metal1 s 8496 23159 8496 23159 4 vdd
port 513 nsew
rlabel metal1 s 8568 25280 8568 25280 4 br0_13
port 54 nsew
rlabel metal1 s 8640 25280 8640 25280 4 bl0_13
port 53 nsew
rlabel metal1 s 7728 23949 7728 23949 4 vdd
port 513 nsew
rlabel metal1 s 8976 24240 8976 24240 4 vdd
port 513 nsew
rlabel metal1 s 7728 23450 7728 23450 4 vdd
port 513 nsew
rlabel metal1 s 9744 23949 9744 23949 4 vdd
port 513 nsew
rlabel metal1 s 7728 22369 7728 22369 4 vdd
port 513 nsew
rlabel metal1 s 7728 24240 7728 24240 4 vdd
port 513 nsew
rlabel metal1 s 7728 23159 7728 23159 4 vdd
port 513 nsew
rlabel metal1 s 9744 23450 9744 23450 4 vdd
port 513 nsew
rlabel metal1 s 8976 25030 8976 25030 4 vdd
port 513 nsew
rlabel metal1 s 8904 25280 8904 25280 4 br0_14
port 58 nsew
rlabel metal1 s 9744 24739 9744 24739 4 vdd
port 513 nsew
rlabel metal1 s 8496 23450 8496 23450 4 vdd
port 513 nsew
rlabel metal1 s 7728 22660 7728 22660 4 vdd
port 513 nsew
rlabel metal1 s 9672 25280 9672 25280 4 bl1_15
port 63 nsew
rlabel metal1 s 7728 25030 7728 25030 4 vdd
port 513 nsew
rlabel metal1 s 8976 23949 8976 23949 4 vdd
port 513 nsew
rlabel metal1 s 9888 25280 9888 25280 4 bl0_15
port 61 nsew
rlabel metal1 s 8976 23450 8976 23450 4 vdd
port 513 nsew
rlabel metal1 s 8832 25280 8832 25280 4 bl0_14
port 57 nsew
rlabel metal1 s 9048 25280 9048 25280 4 bl1_14
port 59 nsew
rlabel metal1 s 9120 25280 9120 25280 4 br1_14
port 60 nsew
rlabel metal1 s 8424 25280 8424 25280 4 bl1_13
port 55 nsew
rlabel metal1 s 9744 24240 9744 24240 4 vdd
port 513 nsew
rlabel metal1 s 8352 25280 8352 25280 4 br1_13
port 56 nsew
rlabel metal1 s 9816 25280 9816 25280 4 br0_15
port 62 nsew
rlabel metal1 s 7584 25280 7584 25280 4 bl0_12
port 49 nsew
rlabel metal1 s 8976 24739 8976 24739 4 vdd
port 513 nsew
rlabel metal1 s 7392 25280 7392 25280 4 bl0_11
port 45 nsew
rlabel metal1 s 6408 25280 6408 25280 4 br0_10
port 42 nsew
rlabel metal1 s 5160 25280 5160 25280 4 br0_8
port 34 nsew
rlabel metal1 s 5304 25280 5304 25280 4 bl1_8
port 35 nsew
rlabel metal1 s 6000 24739 6000 24739 4 vdd
port 513 nsew
rlabel metal1 s 5232 24739 5232 24739 4 vdd
port 513 nsew
rlabel metal1 s 6480 24240 6480 24240 4 vdd
port 513 nsew
rlabel metal1 s 7248 24739 7248 24739 4 vdd
port 513 nsew
rlabel metal1 s 7248 22660 7248 22660 4 vdd
port 513 nsew
rlabel metal1 s 6000 23949 6000 23949 4 vdd
port 513 nsew
rlabel metal1 s 6000 22660 6000 22660 4 vdd
port 513 nsew
rlabel metal1 s 7248 23159 7248 23159 4 vdd
port 513 nsew
rlabel metal1 s 6000 23159 6000 23159 4 vdd
port 513 nsew
rlabel metal1 s 7248 24240 7248 24240 4 vdd
port 513 nsew
rlabel metal1 s 5088 25280 5088 25280 4 bl0_8
port 33 nsew
rlabel metal1 s 7248 22369 7248 22369 4 vdd
port 513 nsew
rlabel metal1 s 5856 25280 5856 25280 4 br1_9
port 40 nsew
rlabel metal1 s 5232 22369 5232 22369 4 vdd
port 513 nsew
rlabel metal1 s 6480 24739 6480 24739 4 vdd
port 513 nsew
rlabel metal1 s 6480 25030 6480 25030 4 vdd
port 513 nsew
rlabel metal1 s 6624 25280 6624 25280 4 br1_10
port 44 nsew
rlabel metal1 s 6480 23949 6480 23949 4 vdd
port 513 nsew
rlabel metal1 s 7176 25280 7176 25280 4 bl1_11
port 47 nsew
rlabel metal1 s 7248 25030 7248 25030 4 vdd
port 513 nsew
rlabel metal1 s 5232 24240 5232 24240 4 vdd
port 513 nsew
rlabel metal1 s 6144 25280 6144 25280 4 bl0_9
port 37 nsew
rlabel metal1 s 5232 23949 5232 23949 4 vdd
port 513 nsew
rlabel metal1 s 5232 22660 5232 22660 4 vdd
port 513 nsew
rlabel metal1 s 6000 24240 6000 24240 4 vdd
port 513 nsew
rlabel metal1 s 5232 23450 5232 23450 4 vdd
port 513 nsew
rlabel metal1 s 7248 23949 7248 23949 4 vdd
port 513 nsew
rlabel metal1 s 6480 22369 6480 22369 4 vdd
port 513 nsew
rlabel metal1 s 7320 25280 7320 25280 4 br0_11
port 46 nsew
rlabel metal1 s 6000 23450 6000 23450 4 vdd
port 513 nsew
rlabel metal1 s 6336 25280 6336 25280 4 bl0_10
port 41 nsew
rlabel metal1 s 5232 25030 5232 25030 4 vdd
port 513 nsew
rlabel metal1 s 6480 23450 6480 23450 4 vdd
port 513 nsew
rlabel metal1 s 6000 22369 6000 22369 4 vdd
port 513 nsew
rlabel metal1 s 7104 25280 7104 25280 4 br1_11
port 48 nsew
rlabel metal1 s 6552 25280 6552 25280 4 bl1_10
port 43 nsew
rlabel metal1 s 5928 25280 5928 25280 4 bl1_9
port 39 nsew
rlabel metal1 s 6000 25030 6000 25030 4 vdd
port 513 nsew
rlabel metal1 s 6072 25280 6072 25280 4 br0_9
port 38 nsew
rlabel metal1 s 5376 25280 5376 25280 4 br1_8
port 36 nsew
rlabel metal1 s 6480 23159 6480 23159 4 vdd
port 513 nsew
rlabel metal1 s 5232 23159 5232 23159 4 vdd
port 513 nsew
rlabel metal1 s 6480 22660 6480 22660 4 vdd
port 513 nsew
rlabel metal1 s 7248 23450 7248 23450 4 vdd
port 513 nsew
rlabel metal1 s 6480 20789 6480 20789 4 vdd
port 513 nsew
rlabel metal1 s 5232 20789 5232 20789 4 vdd
port 513 nsew
rlabel metal1 s 7248 21080 7248 21080 4 vdd
port 513 nsew
rlabel metal1 s 6480 21579 6480 21579 4 vdd
port 513 nsew
rlabel metal1 s 5232 21870 5232 21870 4 vdd
port 513 nsew
rlabel metal1 s 6000 20789 6000 20789 4 vdd
port 513 nsew
rlabel metal1 s 7248 19500 7248 19500 4 vdd
port 513 nsew
rlabel metal1 s 5232 19500 5232 19500 4 vdd
port 513 nsew
rlabel metal1 s 6480 21080 6480 21080 4 vdd
port 513 nsew
rlabel metal1 s 7248 20290 7248 20290 4 vdd
port 513 nsew
rlabel metal1 s 7248 21870 7248 21870 4 vdd
port 513 nsew
rlabel metal1 s 7248 19999 7248 19999 4 vdd
port 513 nsew
rlabel metal1 s 6000 21080 6000 21080 4 vdd
port 513 nsew
rlabel metal1 s 6000 21579 6000 21579 4 vdd
port 513 nsew
rlabel metal1 s 5232 19209 5232 19209 4 vdd
port 513 nsew
rlabel metal1 s 5232 20290 5232 20290 4 vdd
port 513 nsew
rlabel metal1 s 6000 19999 6000 19999 4 vdd
port 513 nsew
rlabel metal1 s 6480 19999 6480 19999 4 vdd
port 513 nsew
rlabel metal1 s 6480 21870 6480 21870 4 vdd
port 513 nsew
rlabel metal1 s 6000 19500 6000 19500 4 vdd
port 513 nsew
rlabel metal1 s 5232 21579 5232 21579 4 vdd
port 513 nsew
rlabel metal1 s 6480 19500 6480 19500 4 vdd
port 513 nsew
rlabel metal1 s 7248 21579 7248 21579 4 vdd
port 513 nsew
rlabel metal1 s 6000 20290 6000 20290 4 vdd
port 513 nsew
rlabel metal1 s 7248 20789 7248 20789 4 vdd
port 513 nsew
rlabel metal1 s 7248 19209 7248 19209 4 vdd
port 513 nsew
rlabel metal1 s 6480 20290 6480 20290 4 vdd
port 513 nsew
rlabel metal1 s 6000 19209 6000 19209 4 vdd
port 513 nsew
rlabel metal1 s 6000 21870 6000 21870 4 vdd
port 513 nsew
rlabel metal1 s 5232 19999 5232 19999 4 vdd
port 513 nsew
rlabel metal1 s 5232 21080 5232 21080 4 vdd
port 513 nsew
rlabel metal1 s 6480 19209 6480 19209 4 vdd
port 513 nsew
rlabel metal1 s 8976 19999 8976 19999 4 vdd
port 513 nsew
rlabel metal1 s 8976 20290 8976 20290 4 vdd
port 513 nsew
rlabel metal1 s 8976 19500 8976 19500 4 vdd
port 513 nsew
rlabel metal1 s 8976 21579 8976 21579 4 vdd
port 513 nsew
rlabel metal1 s 9744 21870 9744 21870 4 vdd
port 513 nsew
rlabel metal1 s 8976 20789 8976 20789 4 vdd
port 513 nsew
rlabel metal1 s 7728 20290 7728 20290 4 vdd
port 513 nsew
rlabel metal1 s 8496 19999 8496 19999 4 vdd
port 513 nsew
rlabel metal1 s 9744 19209 9744 19209 4 vdd
port 513 nsew
rlabel metal1 s 7728 21579 7728 21579 4 vdd
port 513 nsew
rlabel metal1 s 7728 19999 7728 19999 4 vdd
port 513 nsew
rlabel metal1 s 7728 20789 7728 20789 4 vdd
port 513 nsew
rlabel metal1 s 9744 20789 9744 20789 4 vdd
port 513 nsew
rlabel metal1 s 8496 20290 8496 20290 4 vdd
port 513 nsew
rlabel metal1 s 8496 21870 8496 21870 4 vdd
port 513 nsew
rlabel metal1 s 7728 21870 7728 21870 4 vdd
port 513 nsew
rlabel metal1 s 8976 19209 8976 19209 4 vdd
port 513 nsew
rlabel metal1 s 9744 19999 9744 19999 4 vdd
port 513 nsew
rlabel metal1 s 7728 19500 7728 19500 4 vdd
port 513 nsew
rlabel metal1 s 8976 21870 8976 21870 4 vdd
port 513 nsew
rlabel metal1 s 8496 21579 8496 21579 4 vdd
port 513 nsew
rlabel metal1 s 9744 21579 9744 21579 4 vdd
port 513 nsew
rlabel metal1 s 8496 21080 8496 21080 4 vdd
port 513 nsew
rlabel metal1 s 8496 19209 8496 19209 4 vdd
port 513 nsew
rlabel metal1 s 8976 21080 8976 21080 4 vdd
port 513 nsew
rlabel metal1 s 7728 21080 7728 21080 4 vdd
port 513 nsew
rlabel metal1 s 7728 19209 7728 19209 4 vdd
port 513 nsew
rlabel metal1 s 9744 20290 9744 20290 4 vdd
port 513 nsew
rlabel metal1 s 8496 19500 8496 19500 4 vdd
port 513 nsew
rlabel metal1 s 8496 20789 8496 20789 4 vdd
port 513 nsew
rlabel metal1 s 9744 19500 9744 19500 4 vdd
port 513 nsew
rlabel metal1 s 9744 21080 9744 21080 4 vdd
port 513 nsew
rlabel metal1 s 4752 23949 4752 23949 4 vdd
port 513 nsew
rlabel metal1 s 4752 24240 4752 24240 4 vdd
port 513 nsew
rlabel metal1 s 4752 24739 4752 24739 4 vdd
port 513 nsew
rlabel metal1 s 2736 23949 2736 23949 4 vdd
port 513 nsew
rlabel metal1 s 2736 22369 2736 22369 4 vdd
port 513 nsew
rlabel metal1 s 3984 23949 3984 23949 4 vdd
port 513 nsew
rlabel metal1 s 2736 24240 2736 24240 4 vdd
port 513 nsew
rlabel metal1 s 3504 23159 3504 23159 4 vdd
port 513 nsew
rlabel metal1 s 3432 25280 3432 25280 4 bl1_5
port 23 nsew
rlabel metal1 s 3984 22369 3984 22369 4 vdd
port 513 nsew
rlabel metal1 s 3504 24739 3504 24739 4 vdd
port 513 nsew
rlabel metal1 s 4752 23159 4752 23159 4 vdd
port 513 nsew
rlabel metal1 s 3984 24240 3984 24240 4 vdd
port 513 nsew
rlabel metal1 s 3984 22660 3984 22660 4 vdd
port 513 nsew
rlabel metal1 s 2736 24739 2736 24739 4 vdd
port 513 nsew
rlabel metal1 s 4608 25280 4608 25280 4 br1_7
port 32 nsew
rlabel metal1 s 2736 25030 2736 25030 4 vdd
port 513 nsew
rlabel metal1 s 4752 22369 4752 22369 4 vdd
port 513 nsew
rlabel metal1 s 2808 25280 2808 25280 4 bl1_4
port 19 nsew
rlabel metal1 s 3504 23450 3504 23450 4 vdd
port 513 nsew
rlabel metal1 s 4752 25030 4752 25030 4 vdd
port 513 nsew
rlabel metal1 s 3984 25030 3984 25030 4 vdd
port 513 nsew
rlabel metal1 s 4752 22660 4752 22660 4 vdd
port 513 nsew
rlabel metal1 s 3360 25280 3360 25280 4 br1_5
port 24 nsew
rlabel metal1 s 2736 23450 2736 23450 4 vdd
port 513 nsew
rlabel metal1 s 3504 24240 3504 24240 4 vdd
port 513 nsew
rlabel metal1 s 3504 22369 3504 22369 4 vdd
port 513 nsew
rlabel metal1 s 2592 25280 2592 25280 4 bl0_4
port 17 nsew
rlabel metal1 s 3504 23949 3504 23949 4 vdd
port 513 nsew
rlabel metal1 s 3984 24739 3984 24739 4 vdd
port 513 nsew
rlabel metal1 s 3504 22660 3504 22660 4 vdd
port 513 nsew
rlabel metal1 s 3648 25280 3648 25280 4 bl0_5
port 21 nsew
rlabel metal1 s 2736 23159 2736 23159 4 vdd
port 513 nsew
rlabel metal1 s 4752 23450 4752 23450 4 vdd
port 513 nsew
rlabel metal1 s 3504 25030 3504 25030 4 vdd
port 513 nsew
rlabel metal1 s 2736 22660 2736 22660 4 vdd
port 513 nsew
rlabel metal1 s 3984 23159 3984 23159 4 vdd
port 513 nsew
rlabel metal1 s 4896 25280 4896 25280 4 bl0_7
port 29 nsew
rlabel metal1 s 3840 25280 3840 25280 4 bl0_6
port 25 nsew
rlabel metal1 s 4680 25280 4680 25280 4 bl1_7
port 31 nsew
rlabel metal1 s 4056 25280 4056 25280 4 bl1_6
port 27 nsew
rlabel metal1 s 3576 25280 3576 25280 4 br0_5
port 22 nsew
rlabel metal1 s 4128 25280 4128 25280 4 br1_6
port 28 nsew
rlabel metal1 s 3912 25280 3912 25280 4 br0_6
port 26 nsew
rlabel metal1 s 3984 23450 3984 23450 4 vdd
port 513 nsew
rlabel metal1 s 2880 25280 2880 25280 4 br1_4
port 20 nsew
rlabel metal1 s 2664 25280 2664 25280 4 br0_4
port 18 nsew
rlabel metal1 s 4824 25280 4824 25280 4 br0_7
port 30 nsew
rlabel metal1 s 2256 23450 2256 23450 4 vdd
port 513 nsew
rlabel metal1 s 2256 23949 2256 23949 4 vdd
port 513 nsew
rlabel metal1 s 1488 24739 1488 24739 4 vdd
port 513 nsew
rlabel metal1 s 1008 23949 1008 23949 4 vdd
port 513 nsew
rlabel metal1 s 1488 24240 1488 24240 4 vdd
port 513 nsew
rlabel metal1 s 1344 25280 1344 25280 4 bl0_2
port 9 nsew
rlabel metal1 s 2256 24739 2256 24739 4 vdd
port 513 nsew
rlabel metal1 s 2256 25030 2256 25030 4 vdd
port 513 nsew
rlabel metal1 s 2400 25280 2400 25280 4 bl0_3
port 13 nsew
rlabel metal1 s 2256 22369 2256 22369 4 vdd
port 513 nsew
rlabel metal1 s 1416 25280 1416 25280 4 br0_2
port 10 nsew
rlabel metal1 s 1008 22369 1008 22369 4 vdd
port 513 nsew
rlabel metal1 s 240 24739 240 24739 4 vdd
port 513 nsew
rlabel metal1 s 864 25280 864 25280 4 br1_1
port 8 nsew
rlabel metal1 s 1008 25030 1008 25030 4 vdd
port 513 nsew
rlabel metal1 s 240 22660 240 22660 4 vdd
port 513 nsew
rlabel metal1 s 1488 25030 1488 25030 4 vdd
port 513 nsew
rlabel metal1 s 312 25280 312 25280 4 bl1_0
port 3 nsew
rlabel metal1 s 1008 23450 1008 23450 4 vdd
port 513 nsew
rlabel metal1 s 2256 24240 2256 24240 4 vdd
port 513 nsew
rlabel metal1 s 1632 25280 1632 25280 4 br1_2
port 12 nsew
rlabel metal1 s 2256 22660 2256 22660 4 vdd
port 513 nsew
rlabel metal1 s 1152 25280 1152 25280 4 bl0_1
port 5 nsew
rlabel metal1 s 240 23949 240 23949 4 vdd
port 513 nsew
rlabel metal1 s 384 25280 384 25280 4 br1_0
port 4 nsew
rlabel metal1 s 240 25030 240 25030 4 vdd
port 513 nsew
rlabel metal1 s 1008 22660 1008 22660 4 vdd
port 513 nsew
rlabel metal1 s 240 23159 240 23159 4 vdd
port 513 nsew
rlabel metal1 s 936 25280 936 25280 4 bl1_1
port 7 nsew
rlabel metal1 s 1008 24739 1008 24739 4 vdd
port 513 nsew
rlabel metal1 s 2112 25280 2112 25280 4 br1_3
port 16 nsew
rlabel metal1 s 240 23450 240 23450 4 vdd
port 513 nsew
rlabel metal1 s 168 25280 168 25280 4 br0_0
port 2 nsew
rlabel metal1 s 1488 22369 1488 22369 4 vdd
port 513 nsew
rlabel metal1 s 240 24240 240 24240 4 vdd
port 513 nsew
rlabel metal1 s 2328 25280 2328 25280 4 br0_3
port 14 nsew
rlabel metal1 s 96 25280 96 25280 4 bl0_0
port 1 nsew
rlabel metal1 s 1008 23159 1008 23159 4 vdd
port 513 nsew
rlabel metal1 s 1080 25280 1080 25280 4 br0_1
port 6 nsew
rlabel metal1 s 2184 25280 2184 25280 4 bl1_3
port 15 nsew
rlabel metal1 s 2256 23159 2256 23159 4 vdd
port 513 nsew
rlabel metal1 s 240 22369 240 22369 4 vdd
port 513 nsew
rlabel metal1 s 1488 23159 1488 23159 4 vdd
port 513 nsew
rlabel metal1 s 1560 25280 1560 25280 4 bl1_2
port 11 nsew
rlabel metal1 s 1488 23949 1488 23949 4 vdd
port 513 nsew
rlabel metal1 s 1008 24240 1008 24240 4 vdd
port 513 nsew
rlabel metal1 s 1488 23450 1488 23450 4 vdd
port 513 nsew
rlabel metal1 s 1488 22660 1488 22660 4 vdd
port 513 nsew
rlabel metal1 s 240 21870 240 21870 4 vdd
port 513 nsew
rlabel metal1 s 1488 19999 1488 19999 4 vdd
port 513 nsew
rlabel metal1 s 240 21080 240 21080 4 vdd
port 513 nsew
rlabel metal1 s 1488 21579 1488 21579 4 vdd
port 513 nsew
rlabel metal1 s 240 19500 240 19500 4 vdd
port 513 nsew
rlabel metal1 s 1488 20789 1488 20789 4 vdd
port 513 nsew
rlabel metal1 s 1008 19500 1008 19500 4 vdd
port 513 nsew
rlabel metal1 s 2256 21080 2256 21080 4 vdd
port 513 nsew
rlabel metal1 s 240 20789 240 20789 4 vdd
port 513 nsew
rlabel metal1 s 1488 21080 1488 21080 4 vdd
port 513 nsew
rlabel metal1 s 1008 19999 1008 19999 4 vdd
port 513 nsew
rlabel metal1 s 2256 21870 2256 21870 4 vdd
port 513 nsew
rlabel metal1 s 1008 20789 1008 20789 4 vdd
port 513 nsew
rlabel metal1 s 1488 21870 1488 21870 4 vdd
port 513 nsew
rlabel metal1 s 1488 19500 1488 19500 4 vdd
port 513 nsew
rlabel metal1 s 240 20290 240 20290 4 vdd
port 513 nsew
rlabel metal1 s 1488 19209 1488 19209 4 vdd
port 513 nsew
rlabel metal1 s 1008 19209 1008 19209 4 vdd
port 513 nsew
rlabel metal1 s 240 21579 240 21579 4 vdd
port 513 nsew
rlabel metal1 s 240 19209 240 19209 4 vdd
port 513 nsew
rlabel metal1 s 2256 19999 2256 19999 4 vdd
port 513 nsew
rlabel metal1 s 1008 21870 1008 21870 4 vdd
port 513 nsew
rlabel metal1 s 1008 20290 1008 20290 4 vdd
port 513 nsew
rlabel metal1 s 1008 21080 1008 21080 4 vdd
port 513 nsew
rlabel metal1 s 2256 19500 2256 19500 4 vdd
port 513 nsew
rlabel metal1 s 2256 20290 2256 20290 4 vdd
port 513 nsew
rlabel metal1 s 2256 21579 2256 21579 4 vdd
port 513 nsew
rlabel metal1 s 2256 19209 2256 19209 4 vdd
port 513 nsew
rlabel metal1 s 2256 20789 2256 20789 4 vdd
port 513 nsew
rlabel metal1 s 240 19999 240 19999 4 vdd
port 513 nsew
rlabel metal1 s 1488 20290 1488 20290 4 vdd
port 513 nsew
rlabel metal1 s 1008 21579 1008 21579 4 vdd
port 513 nsew
rlabel metal1 s 4752 19209 4752 19209 4 vdd
port 513 nsew
rlabel metal1 s 3984 21080 3984 21080 4 vdd
port 513 nsew
rlabel metal1 s 4752 19999 4752 19999 4 vdd
port 513 nsew
rlabel metal1 s 3984 21579 3984 21579 4 vdd
port 513 nsew
rlabel metal1 s 3504 21870 3504 21870 4 vdd
port 513 nsew
rlabel metal1 s 3984 20789 3984 20789 4 vdd
port 513 nsew
rlabel metal1 s 3984 19999 3984 19999 4 vdd
port 513 nsew
rlabel metal1 s 2736 20290 2736 20290 4 vdd
port 513 nsew
rlabel metal1 s 2736 21870 2736 21870 4 vdd
port 513 nsew
rlabel metal1 s 2736 21080 2736 21080 4 vdd
port 513 nsew
rlabel metal1 s 3984 19500 3984 19500 4 vdd
port 513 nsew
rlabel metal1 s 3504 20290 3504 20290 4 vdd
port 513 nsew
rlabel metal1 s 2736 19500 2736 19500 4 vdd
port 513 nsew
rlabel metal1 s 3504 20789 3504 20789 4 vdd
port 513 nsew
rlabel metal1 s 3984 19209 3984 19209 4 vdd
port 513 nsew
rlabel metal1 s 2736 20789 2736 20789 4 vdd
port 513 nsew
rlabel metal1 s 4752 21080 4752 21080 4 vdd
port 513 nsew
rlabel metal1 s 4752 20789 4752 20789 4 vdd
port 513 nsew
rlabel metal1 s 3504 19500 3504 19500 4 vdd
port 513 nsew
rlabel metal1 s 4752 21579 4752 21579 4 vdd
port 513 nsew
rlabel metal1 s 2736 21579 2736 21579 4 vdd
port 513 nsew
rlabel metal1 s 4752 19500 4752 19500 4 vdd
port 513 nsew
rlabel metal1 s 4752 20290 4752 20290 4 vdd
port 513 nsew
rlabel metal1 s 3984 21870 3984 21870 4 vdd
port 513 nsew
rlabel metal1 s 2736 19209 2736 19209 4 vdd
port 513 nsew
rlabel metal1 s 4752 21870 4752 21870 4 vdd
port 513 nsew
rlabel metal1 s 3504 19209 3504 19209 4 vdd
port 513 nsew
rlabel metal1 s 2736 19999 2736 19999 4 vdd
port 513 nsew
rlabel metal1 s 3504 21080 3504 21080 4 vdd
port 513 nsew
rlabel metal1 s 3984 20290 3984 20290 4 vdd
port 513 nsew
rlabel metal1 s 3504 21579 3504 21579 4 vdd
port 513 nsew
rlabel metal1 s 3504 19999 3504 19999 4 vdd
port 513 nsew
rlabel metal1 s 3504 18710 3504 18710 4 vdd
port 513 nsew
rlabel metal1 s 3504 16049 3504 16049 4 vdd
port 513 nsew
rlabel metal1 s 3504 17920 3504 17920 4 vdd
port 513 nsew
rlabel metal1 s 2736 18710 2736 18710 4 vdd
port 513 nsew
rlabel metal1 s 4752 17629 4752 17629 4 vdd
port 513 nsew
rlabel metal1 s 2736 16839 2736 16839 4 vdd
port 513 nsew
rlabel metal1 s 3984 16049 3984 16049 4 vdd
port 513 nsew
rlabel metal1 s 3504 17130 3504 17130 4 vdd
port 513 nsew
rlabel metal1 s 3504 16340 3504 16340 4 vdd
port 513 nsew
rlabel metal1 s 4752 16340 4752 16340 4 vdd
port 513 nsew
rlabel metal1 s 3504 17629 3504 17629 4 vdd
port 513 nsew
rlabel metal1 s 2736 16049 2736 16049 4 vdd
port 513 nsew
rlabel metal1 s 3984 16839 3984 16839 4 vdd
port 513 nsew
rlabel metal1 s 2736 18419 2736 18419 4 vdd
port 513 nsew
rlabel metal1 s 3984 17629 3984 17629 4 vdd
port 513 nsew
rlabel metal1 s 3504 16839 3504 16839 4 vdd
port 513 nsew
rlabel metal1 s 4752 17130 4752 17130 4 vdd
port 513 nsew
rlabel metal1 s 2736 17130 2736 17130 4 vdd
port 513 nsew
rlabel metal1 s 3984 18710 3984 18710 4 vdd
port 513 nsew
rlabel metal1 s 2736 16340 2736 16340 4 vdd
port 513 nsew
rlabel metal1 s 3984 17920 3984 17920 4 vdd
port 513 nsew
rlabel metal1 s 3984 16340 3984 16340 4 vdd
port 513 nsew
rlabel metal1 s 2736 17920 2736 17920 4 vdd
port 513 nsew
rlabel metal1 s 4752 16839 4752 16839 4 vdd
port 513 nsew
rlabel metal1 s 3504 18419 3504 18419 4 vdd
port 513 nsew
rlabel metal1 s 4752 18710 4752 18710 4 vdd
port 513 nsew
rlabel metal1 s 4752 16049 4752 16049 4 vdd
port 513 nsew
rlabel metal1 s 4752 17920 4752 17920 4 vdd
port 513 nsew
rlabel metal1 s 4752 18419 4752 18419 4 vdd
port 513 nsew
rlabel metal1 s 3984 18419 3984 18419 4 vdd
port 513 nsew
rlabel metal1 s 3984 17130 3984 17130 4 vdd
port 513 nsew
rlabel metal1 s 2736 17629 2736 17629 4 vdd
port 513 nsew
rlabel metal1 s 1488 17629 1488 17629 4 vdd
port 513 nsew
rlabel metal1 s 1488 16340 1488 16340 4 vdd
port 513 nsew
rlabel metal1 s 240 16049 240 16049 4 vdd
port 513 nsew
rlabel metal1 s 240 16340 240 16340 4 vdd
port 513 nsew
rlabel metal1 s 1488 16049 1488 16049 4 vdd
port 513 nsew
rlabel metal1 s 1488 18419 1488 18419 4 vdd
port 513 nsew
rlabel metal1 s 2256 18419 2256 18419 4 vdd
port 513 nsew
rlabel metal1 s 240 16839 240 16839 4 vdd
port 513 nsew
rlabel metal1 s 240 17130 240 17130 4 vdd
port 513 nsew
rlabel metal1 s 1488 16839 1488 16839 4 vdd
port 513 nsew
rlabel metal1 s 2256 17920 2256 17920 4 vdd
port 513 nsew
rlabel metal1 s 240 17629 240 17629 4 vdd
port 513 nsew
rlabel metal1 s 1008 17920 1008 17920 4 vdd
port 513 nsew
rlabel metal1 s 1008 16340 1008 16340 4 vdd
port 513 nsew
rlabel metal1 s 1488 17920 1488 17920 4 vdd
port 513 nsew
rlabel metal1 s 2256 16340 2256 16340 4 vdd
port 513 nsew
rlabel metal1 s 2256 17130 2256 17130 4 vdd
port 513 nsew
rlabel metal1 s 1008 17629 1008 17629 4 vdd
port 513 nsew
rlabel metal1 s 1008 17130 1008 17130 4 vdd
port 513 nsew
rlabel metal1 s 1008 16839 1008 16839 4 vdd
port 513 nsew
rlabel metal1 s 1008 18710 1008 18710 4 vdd
port 513 nsew
rlabel metal1 s 2256 16049 2256 16049 4 vdd
port 513 nsew
rlabel metal1 s 1488 17130 1488 17130 4 vdd
port 513 nsew
rlabel metal1 s 240 18710 240 18710 4 vdd
port 513 nsew
rlabel metal1 s 240 18419 240 18419 4 vdd
port 513 nsew
rlabel metal1 s 2256 18710 2256 18710 4 vdd
port 513 nsew
rlabel metal1 s 2256 17629 2256 17629 4 vdd
port 513 nsew
rlabel metal1 s 1008 16049 1008 16049 4 vdd
port 513 nsew
rlabel metal1 s 240 17920 240 17920 4 vdd
port 513 nsew
rlabel metal1 s 1488 18710 1488 18710 4 vdd
port 513 nsew
rlabel metal1 s 1008 18419 1008 18419 4 vdd
port 513 nsew
rlabel metal1 s 2256 16839 2256 16839 4 vdd
port 513 nsew
rlabel metal1 s 1008 13970 1008 13970 4 vdd
port 513 nsew
rlabel metal1 s 2256 14469 2256 14469 4 vdd
port 513 nsew
rlabel metal1 s 240 13970 240 13970 4 vdd
port 513 nsew
rlabel metal1 s 2256 15259 2256 15259 4 vdd
port 513 nsew
rlabel metal1 s 2256 12889 2256 12889 4 vdd
port 513 nsew
rlabel metal1 s 2256 13180 2256 13180 4 vdd
port 513 nsew
rlabel metal1 s 1488 12889 1488 12889 4 vdd
port 513 nsew
rlabel metal1 s 2256 14760 2256 14760 4 vdd
port 513 nsew
rlabel metal1 s 1008 12889 1008 12889 4 vdd
port 513 nsew
rlabel metal1 s 1488 15550 1488 15550 4 vdd
port 513 nsew
rlabel metal1 s 240 15550 240 15550 4 vdd
port 513 nsew
rlabel metal1 s 1488 13679 1488 13679 4 vdd
port 513 nsew
rlabel metal1 s 240 14760 240 14760 4 vdd
port 513 nsew
rlabel metal1 s 1008 13679 1008 13679 4 vdd
port 513 nsew
rlabel metal1 s 1488 15259 1488 15259 4 vdd
port 513 nsew
rlabel metal1 s 2256 13970 2256 13970 4 vdd
port 513 nsew
rlabel metal1 s 1008 15259 1008 15259 4 vdd
port 513 nsew
rlabel metal1 s 2256 15550 2256 15550 4 vdd
port 513 nsew
rlabel metal1 s 240 15259 240 15259 4 vdd
port 513 nsew
rlabel metal1 s 1488 13180 1488 13180 4 vdd
port 513 nsew
rlabel metal1 s 2256 13679 2256 13679 4 vdd
port 513 nsew
rlabel metal1 s 1008 14760 1008 14760 4 vdd
port 513 nsew
rlabel metal1 s 240 13180 240 13180 4 vdd
port 513 nsew
rlabel metal1 s 240 12889 240 12889 4 vdd
port 513 nsew
rlabel metal1 s 240 13679 240 13679 4 vdd
port 513 nsew
rlabel metal1 s 1008 14469 1008 14469 4 vdd
port 513 nsew
rlabel metal1 s 1488 14469 1488 14469 4 vdd
port 513 nsew
rlabel metal1 s 1488 13970 1488 13970 4 vdd
port 513 nsew
rlabel metal1 s 1008 15550 1008 15550 4 vdd
port 513 nsew
rlabel metal1 s 1488 14760 1488 14760 4 vdd
port 513 nsew
rlabel metal1 s 240 14469 240 14469 4 vdd
port 513 nsew
rlabel metal1 s 1008 13180 1008 13180 4 vdd
port 513 nsew
rlabel metal1 s 3984 13180 3984 13180 4 vdd
port 513 nsew
rlabel metal1 s 4752 14469 4752 14469 4 vdd
port 513 nsew
rlabel metal1 s 2736 13679 2736 13679 4 vdd
port 513 nsew
rlabel metal1 s 2736 14760 2736 14760 4 vdd
port 513 nsew
rlabel metal1 s 3504 13180 3504 13180 4 vdd
port 513 nsew
rlabel metal1 s 3504 15550 3504 15550 4 vdd
port 513 nsew
rlabel metal1 s 2736 13180 2736 13180 4 vdd
port 513 nsew
rlabel metal1 s 3984 14469 3984 14469 4 vdd
port 513 nsew
rlabel metal1 s 2736 14469 2736 14469 4 vdd
port 513 nsew
rlabel metal1 s 4752 12889 4752 12889 4 vdd
port 513 nsew
rlabel metal1 s 3984 12889 3984 12889 4 vdd
port 513 nsew
rlabel metal1 s 3504 15259 3504 15259 4 vdd
port 513 nsew
rlabel metal1 s 3984 15550 3984 15550 4 vdd
port 513 nsew
rlabel metal1 s 4752 15550 4752 15550 4 vdd
port 513 nsew
rlabel metal1 s 3504 14469 3504 14469 4 vdd
port 513 nsew
rlabel metal1 s 3504 13679 3504 13679 4 vdd
port 513 nsew
rlabel metal1 s 2736 12889 2736 12889 4 vdd
port 513 nsew
rlabel metal1 s 3504 13970 3504 13970 4 vdd
port 513 nsew
rlabel metal1 s 2736 15259 2736 15259 4 vdd
port 513 nsew
rlabel metal1 s 2736 15550 2736 15550 4 vdd
port 513 nsew
rlabel metal1 s 4752 13970 4752 13970 4 vdd
port 513 nsew
rlabel metal1 s 3504 12889 3504 12889 4 vdd
port 513 nsew
rlabel metal1 s 4752 15259 4752 15259 4 vdd
port 513 nsew
rlabel metal1 s 2736 13970 2736 13970 4 vdd
port 513 nsew
rlabel metal1 s 3984 14760 3984 14760 4 vdd
port 513 nsew
rlabel metal1 s 4752 14760 4752 14760 4 vdd
port 513 nsew
rlabel metal1 s 4752 13679 4752 13679 4 vdd
port 513 nsew
rlabel metal1 s 3984 13970 3984 13970 4 vdd
port 513 nsew
rlabel metal1 s 3984 15259 3984 15259 4 vdd
port 513 nsew
rlabel metal1 s 3984 13679 3984 13679 4 vdd
port 513 nsew
rlabel metal1 s 3504 14760 3504 14760 4 vdd
port 513 nsew
rlabel metal1 s 4752 13180 4752 13180 4 vdd
port 513 nsew
rlabel metal1 s 7728 17130 7728 17130 4 vdd
port 513 nsew
rlabel metal1 s 8976 17920 8976 17920 4 vdd
port 513 nsew
rlabel metal1 s 8976 17130 8976 17130 4 vdd
port 513 nsew
rlabel metal1 s 9744 18710 9744 18710 4 vdd
port 513 nsew
rlabel metal1 s 7728 18710 7728 18710 4 vdd
port 513 nsew
rlabel metal1 s 8496 17920 8496 17920 4 vdd
port 513 nsew
rlabel metal1 s 9744 17629 9744 17629 4 vdd
port 513 nsew
rlabel metal1 s 7728 17629 7728 17629 4 vdd
port 513 nsew
rlabel metal1 s 8496 16340 8496 16340 4 vdd
port 513 nsew
rlabel metal1 s 8496 16049 8496 16049 4 vdd
port 513 nsew
rlabel metal1 s 9744 18419 9744 18419 4 vdd
port 513 nsew
rlabel metal1 s 8496 17130 8496 17130 4 vdd
port 513 nsew
rlabel metal1 s 7728 16049 7728 16049 4 vdd
port 513 nsew
rlabel metal1 s 8976 16340 8976 16340 4 vdd
port 513 nsew
rlabel metal1 s 8976 16049 8976 16049 4 vdd
port 513 nsew
rlabel metal1 s 9744 16340 9744 16340 4 vdd
port 513 nsew
rlabel metal1 s 8496 17629 8496 17629 4 vdd
port 513 nsew
rlabel metal1 s 8496 18419 8496 18419 4 vdd
port 513 nsew
rlabel metal1 s 8976 18710 8976 18710 4 vdd
port 513 nsew
rlabel metal1 s 7728 18419 7728 18419 4 vdd
port 513 nsew
rlabel metal1 s 7728 17920 7728 17920 4 vdd
port 513 nsew
rlabel metal1 s 7728 16839 7728 16839 4 vdd
port 513 nsew
rlabel metal1 s 8976 18419 8976 18419 4 vdd
port 513 nsew
rlabel metal1 s 9744 16049 9744 16049 4 vdd
port 513 nsew
rlabel metal1 s 9744 17920 9744 17920 4 vdd
port 513 nsew
rlabel metal1 s 9744 17130 9744 17130 4 vdd
port 513 nsew
rlabel metal1 s 8976 17629 8976 17629 4 vdd
port 513 nsew
rlabel metal1 s 8496 16839 8496 16839 4 vdd
port 513 nsew
rlabel metal1 s 7728 16340 7728 16340 4 vdd
port 513 nsew
rlabel metal1 s 8496 18710 8496 18710 4 vdd
port 513 nsew
rlabel metal1 s 9744 16839 9744 16839 4 vdd
port 513 nsew
rlabel metal1 s 8976 16839 8976 16839 4 vdd
port 513 nsew
rlabel metal1 s 6000 18710 6000 18710 4 vdd
port 513 nsew
rlabel metal1 s 6000 16049 6000 16049 4 vdd
port 513 nsew
rlabel metal1 s 5232 16049 5232 16049 4 vdd
port 513 nsew
rlabel metal1 s 5232 17130 5232 17130 4 vdd
port 513 nsew
rlabel metal1 s 6000 16839 6000 16839 4 vdd
port 513 nsew
rlabel metal1 s 7248 17629 7248 17629 4 vdd
port 513 nsew
rlabel metal1 s 6000 17130 6000 17130 4 vdd
port 513 nsew
rlabel metal1 s 6000 16340 6000 16340 4 vdd
port 513 nsew
rlabel metal1 s 5232 16839 5232 16839 4 vdd
port 513 nsew
rlabel metal1 s 6480 16839 6480 16839 4 vdd
port 513 nsew
rlabel metal1 s 6000 17629 6000 17629 4 vdd
port 513 nsew
rlabel metal1 s 5232 17920 5232 17920 4 vdd
port 513 nsew
rlabel metal1 s 7248 17130 7248 17130 4 vdd
port 513 nsew
rlabel metal1 s 5232 18710 5232 18710 4 vdd
port 513 nsew
rlabel metal1 s 7248 16340 7248 16340 4 vdd
port 513 nsew
rlabel metal1 s 5232 18419 5232 18419 4 vdd
port 513 nsew
rlabel metal1 s 6480 17629 6480 17629 4 vdd
port 513 nsew
rlabel metal1 s 7248 16839 7248 16839 4 vdd
port 513 nsew
rlabel metal1 s 5232 16340 5232 16340 4 vdd
port 513 nsew
rlabel metal1 s 6480 18710 6480 18710 4 vdd
port 513 nsew
rlabel metal1 s 6480 16049 6480 16049 4 vdd
port 513 nsew
rlabel metal1 s 7248 18419 7248 18419 4 vdd
port 513 nsew
rlabel metal1 s 6480 17920 6480 17920 4 vdd
port 513 nsew
rlabel metal1 s 6000 18419 6000 18419 4 vdd
port 513 nsew
rlabel metal1 s 5232 17629 5232 17629 4 vdd
port 513 nsew
rlabel metal1 s 7248 18710 7248 18710 4 vdd
port 513 nsew
rlabel metal1 s 7248 17920 7248 17920 4 vdd
port 513 nsew
rlabel metal1 s 7248 16049 7248 16049 4 vdd
port 513 nsew
rlabel metal1 s 6480 17130 6480 17130 4 vdd
port 513 nsew
rlabel metal1 s 6480 18419 6480 18419 4 vdd
port 513 nsew
rlabel metal1 s 6480 16340 6480 16340 4 vdd
port 513 nsew
rlabel metal1 s 6000 17920 6000 17920 4 vdd
port 513 nsew
rlabel metal1 s 6480 14469 6480 14469 4 vdd
port 513 nsew
rlabel metal1 s 5232 13970 5232 13970 4 vdd
port 513 nsew
rlabel metal1 s 6000 13180 6000 13180 4 vdd
port 513 nsew
rlabel metal1 s 6000 15259 6000 15259 4 vdd
port 513 nsew
rlabel metal1 s 5232 15550 5232 15550 4 vdd
port 513 nsew
rlabel metal1 s 5232 15259 5232 15259 4 vdd
port 513 nsew
rlabel metal1 s 7248 15550 7248 15550 4 vdd
port 513 nsew
rlabel metal1 s 5232 13180 5232 13180 4 vdd
port 513 nsew
rlabel metal1 s 6480 14760 6480 14760 4 vdd
port 513 nsew
rlabel metal1 s 5232 13679 5232 13679 4 vdd
port 513 nsew
rlabel metal1 s 5232 14469 5232 14469 4 vdd
port 513 nsew
rlabel metal1 s 7248 12889 7248 12889 4 vdd
port 513 nsew
rlabel metal1 s 6000 15550 6000 15550 4 vdd
port 513 nsew
rlabel metal1 s 6000 13679 6000 13679 4 vdd
port 513 nsew
rlabel metal1 s 7248 13679 7248 13679 4 vdd
port 513 nsew
rlabel metal1 s 7248 14469 7248 14469 4 vdd
port 513 nsew
rlabel metal1 s 7248 14760 7248 14760 4 vdd
port 513 nsew
rlabel metal1 s 6480 12889 6480 12889 4 vdd
port 513 nsew
rlabel metal1 s 6480 15259 6480 15259 4 vdd
port 513 nsew
rlabel metal1 s 7248 15259 7248 15259 4 vdd
port 513 nsew
rlabel metal1 s 6480 13679 6480 13679 4 vdd
port 513 nsew
rlabel metal1 s 6480 13970 6480 13970 4 vdd
port 513 nsew
rlabel metal1 s 7248 13180 7248 13180 4 vdd
port 513 nsew
rlabel metal1 s 5232 14760 5232 14760 4 vdd
port 513 nsew
rlabel metal1 s 6480 13180 6480 13180 4 vdd
port 513 nsew
rlabel metal1 s 6000 14469 6000 14469 4 vdd
port 513 nsew
rlabel metal1 s 6000 13970 6000 13970 4 vdd
port 513 nsew
rlabel metal1 s 6000 12889 6000 12889 4 vdd
port 513 nsew
rlabel metal1 s 6480 15550 6480 15550 4 vdd
port 513 nsew
rlabel metal1 s 6000 14760 6000 14760 4 vdd
port 513 nsew
rlabel metal1 s 5232 12889 5232 12889 4 vdd
port 513 nsew
rlabel metal1 s 7248 13970 7248 13970 4 vdd
port 513 nsew
rlabel metal1 s 8496 13180 8496 13180 4 vdd
port 513 nsew
rlabel metal1 s 8496 15259 8496 15259 4 vdd
port 513 nsew
rlabel metal1 s 7728 14760 7728 14760 4 vdd
port 513 nsew
rlabel metal1 s 8976 13970 8976 13970 4 vdd
port 513 nsew
rlabel metal1 s 7728 13180 7728 13180 4 vdd
port 513 nsew
rlabel metal1 s 7728 13970 7728 13970 4 vdd
port 513 nsew
rlabel metal1 s 8976 15259 8976 15259 4 vdd
port 513 nsew
rlabel metal1 s 7728 15550 7728 15550 4 vdd
port 513 nsew
rlabel metal1 s 8976 13679 8976 13679 4 vdd
port 513 nsew
rlabel metal1 s 8976 12889 8976 12889 4 vdd
port 513 nsew
rlabel metal1 s 7728 13679 7728 13679 4 vdd
port 513 nsew
rlabel metal1 s 8496 13970 8496 13970 4 vdd
port 513 nsew
rlabel metal1 s 8496 12889 8496 12889 4 vdd
port 513 nsew
rlabel metal1 s 9744 13679 9744 13679 4 vdd
port 513 nsew
rlabel metal1 s 7728 15259 7728 15259 4 vdd
port 513 nsew
rlabel metal1 s 8976 14760 8976 14760 4 vdd
port 513 nsew
rlabel metal1 s 7728 14469 7728 14469 4 vdd
port 513 nsew
rlabel metal1 s 9744 15259 9744 15259 4 vdd
port 513 nsew
rlabel metal1 s 8976 14469 8976 14469 4 vdd
port 513 nsew
rlabel metal1 s 8496 14760 8496 14760 4 vdd
port 513 nsew
rlabel metal1 s 8976 15550 8976 15550 4 vdd
port 513 nsew
rlabel metal1 s 8496 13679 8496 13679 4 vdd
port 513 nsew
rlabel metal1 s 7728 12889 7728 12889 4 vdd
port 513 nsew
rlabel metal1 s 9744 13970 9744 13970 4 vdd
port 513 nsew
rlabel metal1 s 9744 15550 9744 15550 4 vdd
port 513 nsew
rlabel metal1 s 9744 14469 9744 14469 4 vdd
port 513 nsew
rlabel metal1 s 8496 14469 8496 14469 4 vdd
port 513 nsew
rlabel metal1 s 9744 14760 9744 14760 4 vdd
port 513 nsew
rlabel metal1 s 9744 12889 9744 12889 4 vdd
port 513 nsew
rlabel metal1 s 8976 13180 8976 13180 4 vdd
port 513 nsew
rlabel metal1 s 9744 13180 9744 13180 4 vdd
port 513 nsew
rlabel metal1 s 8496 15550 8496 15550 4 vdd
port 513 nsew
rlabel metal1 s 7728 9729 7728 9729 4 vdd
port 513 nsew
rlabel metal1 s 7728 11309 7728 11309 4 vdd
port 513 nsew
rlabel metal1 s 9744 10020 9744 10020 4 vdd
port 513 nsew
rlabel metal1 s 9744 11309 9744 11309 4 vdd
port 513 nsew
rlabel metal1 s 8496 10020 8496 10020 4 vdd
port 513 nsew
rlabel metal1 s 9744 12390 9744 12390 4 vdd
port 513 nsew
rlabel metal1 s 8976 10519 8976 10519 4 vdd
port 513 nsew
rlabel metal1 s 9744 10519 9744 10519 4 vdd
port 513 nsew
rlabel metal1 s 9744 12099 9744 12099 4 vdd
port 513 nsew
rlabel metal1 s 8496 11600 8496 11600 4 vdd
port 513 nsew
rlabel metal1 s 7728 12099 7728 12099 4 vdd
port 513 nsew
rlabel metal1 s 7728 10810 7728 10810 4 vdd
port 513 nsew
rlabel metal1 s 8496 12390 8496 12390 4 vdd
port 513 nsew
rlabel metal1 s 9744 11600 9744 11600 4 vdd
port 513 nsew
rlabel metal1 s 7728 12390 7728 12390 4 vdd
port 513 nsew
rlabel metal1 s 8496 10810 8496 10810 4 vdd
port 513 nsew
rlabel metal1 s 8976 11309 8976 11309 4 vdd
port 513 nsew
rlabel metal1 s 8976 12099 8976 12099 4 vdd
port 513 nsew
rlabel metal1 s 8496 11309 8496 11309 4 vdd
port 513 nsew
rlabel metal1 s 8496 9729 8496 9729 4 vdd
port 513 nsew
rlabel metal1 s 8976 11600 8976 11600 4 vdd
port 513 nsew
rlabel metal1 s 8976 10810 8976 10810 4 vdd
port 513 nsew
rlabel metal1 s 8496 10519 8496 10519 4 vdd
port 513 nsew
rlabel metal1 s 7728 10020 7728 10020 4 vdd
port 513 nsew
rlabel metal1 s 9744 10810 9744 10810 4 vdd
port 513 nsew
rlabel metal1 s 7728 11600 7728 11600 4 vdd
port 513 nsew
rlabel metal1 s 8976 12390 8976 12390 4 vdd
port 513 nsew
rlabel metal1 s 8496 12099 8496 12099 4 vdd
port 513 nsew
rlabel metal1 s 8976 10020 8976 10020 4 vdd
port 513 nsew
rlabel metal1 s 9744 9729 9744 9729 4 vdd
port 513 nsew
rlabel metal1 s 7728 10519 7728 10519 4 vdd
port 513 nsew
rlabel metal1 s 8976 9729 8976 9729 4 vdd
port 513 nsew
rlabel metal1 s 6000 12390 6000 12390 4 vdd
port 513 nsew
rlabel metal1 s 6480 12390 6480 12390 4 vdd
port 513 nsew
rlabel metal1 s 6480 10020 6480 10020 4 vdd
port 513 nsew
rlabel metal1 s 5232 11309 5232 11309 4 vdd
port 513 nsew
rlabel metal1 s 7248 12099 7248 12099 4 vdd
port 513 nsew
rlabel metal1 s 6480 11309 6480 11309 4 vdd
port 513 nsew
rlabel metal1 s 7248 10810 7248 10810 4 vdd
port 513 nsew
rlabel metal1 s 6000 10020 6000 10020 4 vdd
port 513 nsew
rlabel metal1 s 6480 11600 6480 11600 4 vdd
port 513 nsew
rlabel metal1 s 7248 10519 7248 10519 4 vdd
port 513 nsew
rlabel metal1 s 5232 11600 5232 11600 4 vdd
port 513 nsew
rlabel metal1 s 5232 9729 5232 9729 4 vdd
port 513 nsew
rlabel metal1 s 6000 10810 6000 10810 4 vdd
port 513 nsew
rlabel metal1 s 6480 9729 6480 9729 4 vdd
port 513 nsew
rlabel metal1 s 6480 12099 6480 12099 4 vdd
port 513 nsew
rlabel metal1 s 5232 10519 5232 10519 4 vdd
port 513 nsew
rlabel metal1 s 6000 10519 6000 10519 4 vdd
port 513 nsew
rlabel metal1 s 7248 12390 7248 12390 4 vdd
port 513 nsew
rlabel metal1 s 7248 10020 7248 10020 4 vdd
port 513 nsew
rlabel metal1 s 6480 10810 6480 10810 4 vdd
port 513 nsew
rlabel metal1 s 7248 11309 7248 11309 4 vdd
port 513 nsew
rlabel metal1 s 6000 11309 6000 11309 4 vdd
port 513 nsew
rlabel metal1 s 6000 11600 6000 11600 4 vdd
port 513 nsew
rlabel metal1 s 5232 10810 5232 10810 4 vdd
port 513 nsew
rlabel metal1 s 5232 10020 5232 10020 4 vdd
port 513 nsew
rlabel metal1 s 6480 10519 6480 10519 4 vdd
port 513 nsew
rlabel metal1 s 6000 9729 6000 9729 4 vdd
port 513 nsew
rlabel metal1 s 5232 12390 5232 12390 4 vdd
port 513 nsew
rlabel metal1 s 7248 9729 7248 9729 4 vdd
port 513 nsew
rlabel metal1 s 7248 11600 7248 11600 4 vdd
port 513 nsew
rlabel metal1 s 5232 12099 5232 12099 4 vdd
port 513 nsew
rlabel metal1 s 6000 12099 6000 12099 4 vdd
port 513 nsew
rlabel metal1 s 5232 7650 5232 7650 4 vdd
port 513 nsew
rlabel metal1 s 6000 6569 6000 6569 4 vdd
port 513 nsew
rlabel metal1 s 7248 6860 7248 6860 4 vdd
port 513 nsew
rlabel metal1 s 5232 6860 5232 6860 4 vdd
port 513 nsew
rlabel metal1 s 6480 7650 6480 7650 4 vdd
port 513 nsew
rlabel metal1 s 6480 7359 6480 7359 4 vdd
port 513 nsew
rlabel metal1 s 5232 8440 5232 8440 4 vdd
port 513 nsew
rlabel metal1 s 7248 7359 7248 7359 4 vdd
port 513 nsew
rlabel metal1 s 5232 8149 5232 8149 4 vdd
port 513 nsew
rlabel metal1 s 5232 7359 5232 7359 4 vdd
port 513 nsew
rlabel metal1 s 7248 9230 7248 9230 4 vdd
port 513 nsew
rlabel metal1 s 6480 6569 6480 6569 4 vdd
port 513 nsew
rlabel metal1 s 7248 8440 7248 8440 4 vdd
port 513 nsew
rlabel metal1 s 5232 9230 5232 9230 4 vdd
port 513 nsew
rlabel metal1 s 7248 6569 7248 6569 4 vdd
port 513 nsew
rlabel metal1 s 6000 8939 6000 8939 4 vdd
port 513 nsew
rlabel metal1 s 6000 6860 6000 6860 4 vdd
port 513 nsew
rlabel metal1 s 6480 8440 6480 8440 4 vdd
port 513 nsew
rlabel metal1 s 6000 7650 6000 7650 4 vdd
port 513 nsew
rlabel metal1 s 6000 8440 6000 8440 4 vdd
port 513 nsew
rlabel metal1 s 7248 8149 7248 8149 4 vdd
port 513 nsew
rlabel metal1 s 5232 8939 5232 8939 4 vdd
port 513 nsew
rlabel metal1 s 6480 8149 6480 8149 4 vdd
port 513 nsew
rlabel metal1 s 7248 7650 7248 7650 4 vdd
port 513 nsew
rlabel metal1 s 6000 9230 6000 9230 4 vdd
port 513 nsew
rlabel metal1 s 6000 7359 6000 7359 4 vdd
port 513 nsew
rlabel metal1 s 7248 8939 7248 8939 4 vdd
port 513 nsew
rlabel metal1 s 5232 6569 5232 6569 4 vdd
port 513 nsew
rlabel metal1 s 6000 8149 6000 8149 4 vdd
port 513 nsew
rlabel metal1 s 6480 6860 6480 6860 4 vdd
port 513 nsew
rlabel metal1 s 6480 8939 6480 8939 4 vdd
port 513 nsew
rlabel metal1 s 6480 9230 6480 9230 4 vdd
port 513 nsew
rlabel metal1 s 8496 9230 8496 9230 4 vdd
port 513 nsew
rlabel metal1 s 8976 6569 8976 6569 4 vdd
port 513 nsew
rlabel metal1 s 8496 8149 8496 8149 4 vdd
port 513 nsew
rlabel metal1 s 7728 7650 7728 7650 4 vdd
port 513 nsew
rlabel metal1 s 8976 6860 8976 6860 4 vdd
port 513 nsew
rlabel metal1 s 8976 8149 8976 8149 4 vdd
port 513 nsew
rlabel metal1 s 8976 7650 8976 7650 4 vdd
port 513 nsew
rlabel metal1 s 9744 6569 9744 6569 4 vdd
port 513 nsew
rlabel metal1 s 8976 8939 8976 8939 4 vdd
port 513 nsew
rlabel metal1 s 9744 8939 9744 8939 4 vdd
port 513 nsew
rlabel metal1 s 8976 8440 8976 8440 4 vdd
port 513 nsew
rlabel metal1 s 7728 6569 7728 6569 4 vdd
port 513 nsew
rlabel metal1 s 8496 8939 8496 8939 4 vdd
port 513 nsew
rlabel metal1 s 7728 8149 7728 8149 4 vdd
port 513 nsew
rlabel metal1 s 9744 9230 9744 9230 4 vdd
port 513 nsew
rlabel metal1 s 7728 8939 7728 8939 4 vdd
port 513 nsew
rlabel metal1 s 9744 8440 9744 8440 4 vdd
port 513 nsew
rlabel metal1 s 8496 6569 8496 6569 4 vdd
port 513 nsew
rlabel metal1 s 8496 7359 8496 7359 4 vdd
port 513 nsew
rlabel metal1 s 9744 8149 9744 8149 4 vdd
port 513 nsew
rlabel metal1 s 8496 7650 8496 7650 4 vdd
port 513 nsew
rlabel metal1 s 8496 8440 8496 8440 4 vdd
port 513 nsew
rlabel metal1 s 7728 8440 7728 8440 4 vdd
port 513 nsew
rlabel metal1 s 9744 7650 9744 7650 4 vdd
port 513 nsew
rlabel metal1 s 8496 6860 8496 6860 4 vdd
port 513 nsew
rlabel metal1 s 9744 7359 9744 7359 4 vdd
port 513 nsew
rlabel metal1 s 7728 7359 7728 7359 4 vdd
port 513 nsew
rlabel metal1 s 9744 6860 9744 6860 4 vdd
port 513 nsew
rlabel metal1 s 7728 6860 7728 6860 4 vdd
port 513 nsew
rlabel metal1 s 7728 9230 7728 9230 4 vdd
port 513 nsew
rlabel metal1 s 8976 9230 8976 9230 4 vdd
port 513 nsew
rlabel metal1 s 8976 7359 8976 7359 4 vdd
port 513 nsew
rlabel metal1 s 3504 12390 3504 12390 4 vdd
port 513 nsew
rlabel metal1 s 3984 10810 3984 10810 4 vdd
port 513 nsew
rlabel metal1 s 4752 12390 4752 12390 4 vdd
port 513 nsew
rlabel metal1 s 3504 10519 3504 10519 4 vdd
port 513 nsew
rlabel metal1 s 3984 10020 3984 10020 4 vdd
port 513 nsew
rlabel metal1 s 4752 10020 4752 10020 4 vdd
port 513 nsew
rlabel metal1 s 3504 10020 3504 10020 4 vdd
port 513 nsew
rlabel metal1 s 4752 11600 4752 11600 4 vdd
port 513 nsew
rlabel metal1 s 3984 12099 3984 12099 4 vdd
port 513 nsew
rlabel metal1 s 2736 10020 2736 10020 4 vdd
port 513 nsew
rlabel metal1 s 3984 12390 3984 12390 4 vdd
port 513 nsew
rlabel metal1 s 2736 11600 2736 11600 4 vdd
port 513 nsew
rlabel metal1 s 3504 12099 3504 12099 4 vdd
port 513 nsew
rlabel metal1 s 4752 11309 4752 11309 4 vdd
port 513 nsew
rlabel metal1 s 4752 10519 4752 10519 4 vdd
port 513 nsew
rlabel metal1 s 3504 10810 3504 10810 4 vdd
port 513 nsew
rlabel metal1 s 2736 9729 2736 9729 4 vdd
port 513 nsew
rlabel metal1 s 4752 12099 4752 12099 4 vdd
port 513 nsew
rlabel metal1 s 2736 12099 2736 12099 4 vdd
port 513 nsew
rlabel metal1 s 3504 11309 3504 11309 4 vdd
port 513 nsew
rlabel metal1 s 3984 11600 3984 11600 4 vdd
port 513 nsew
rlabel metal1 s 2736 12390 2736 12390 4 vdd
port 513 nsew
rlabel metal1 s 2736 10519 2736 10519 4 vdd
port 513 nsew
rlabel metal1 s 2736 11309 2736 11309 4 vdd
port 513 nsew
rlabel metal1 s 2736 10810 2736 10810 4 vdd
port 513 nsew
rlabel metal1 s 3984 11309 3984 11309 4 vdd
port 513 nsew
rlabel metal1 s 3984 9729 3984 9729 4 vdd
port 513 nsew
rlabel metal1 s 4752 10810 4752 10810 4 vdd
port 513 nsew
rlabel metal1 s 3504 9729 3504 9729 4 vdd
port 513 nsew
rlabel metal1 s 3504 11600 3504 11600 4 vdd
port 513 nsew
rlabel metal1 s 4752 9729 4752 9729 4 vdd
port 513 nsew
rlabel metal1 s 3984 10519 3984 10519 4 vdd
port 513 nsew
rlabel metal1 s 2256 10020 2256 10020 4 vdd
port 513 nsew
rlabel metal1 s 2256 12390 2256 12390 4 vdd
port 513 nsew
rlabel metal1 s 240 10810 240 10810 4 vdd
port 513 nsew
rlabel metal1 s 1008 10810 1008 10810 4 vdd
port 513 nsew
rlabel metal1 s 1488 11600 1488 11600 4 vdd
port 513 nsew
rlabel metal1 s 240 10020 240 10020 4 vdd
port 513 nsew
rlabel metal1 s 2256 9729 2256 9729 4 vdd
port 513 nsew
rlabel metal1 s 1488 9729 1488 9729 4 vdd
port 513 nsew
rlabel metal1 s 240 10519 240 10519 4 vdd
port 513 nsew
rlabel metal1 s 1008 9729 1008 9729 4 vdd
port 513 nsew
rlabel metal1 s 240 11600 240 11600 4 vdd
port 513 nsew
rlabel metal1 s 1008 10519 1008 10519 4 vdd
port 513 nsew
rlabel metal1 s 240 11309 240 11309 4 vdd
port 513 nsew
rlabel metal1 s 2256 10810 2256 10810 4 vdd
port 513 nsew
rlabel metal1 s 2256 12099 2256 12099 4 vdd
port 513 nsew
rlabel metal1 s 1488 10810 1488 10810 4 vdd
port 513 nsew
rlabel metal1 s 1008 10020 1008 10020 4 vdd
port 513 nsew
rlabel metal1 s 1008 11600 1008 11600 4 vdd
port 513 nsew
rlabel metal1 s 2256 11600 2256 11600 4 vdd
port 513 nsew
rlabel metal1 s 2256 11309 2256 11309 4 vdd
port 513 nsew
rlabel metal1 s 1488 11309 1488 11309 4 vdd
port 513 nsew
rlabel metal1 s 1008 12390 1008 12390 4 vdd
port 513 nsew
rlabel metal1 s 1488 10519 1488 10519 4 vdd
port 513 nsew
rlabel metal1 s 2256 10519 2256 10519 4 vdd
port 513 nsew
rlabel metal1 s 1008 12099 1008 12099 4 vdd
port 513 nsew
rlabel metal1 s 240 12099 240 12099 4 vdd
port 513 nsew
rlabel metal1 s 240 9729 240 9729 4 vdd
port 513 nsew
rlabel metal1 s 240 12390 240 12390 4 vdd
port 513 nsew
rlabel metal1 s 1008 11309 1008 11309 4 vdd
port 513 nsew
rlabel metal1 s 1488 12099 1488 12099 4 vdd
port 513 nsew
rlabel metal1 s 1488 10020 1488 10020 4 vdd
port 513 nsew
rlabel metal1 s 1488 12390 1488 12390 4 vdd
port 513 nsew
rlabel metal1 s 2256 8149 2256 8149 4 vdd
port 513 nsew
rlabel metal1 s 1008 8939 1008 8939 4 vdd
port 513 nsew
rlabel metal1 s 1488 8440 1488 8440 4 vdd
port 513 nsew
rlabel metal1 s 1488 6569 1488 6569 4 vdd
port 513 nsew
rlabel metal1 s 2256 7359 2256 7359 4 vdd
port 513 nsew
rlabel metal1 s 240 8440 240 8440 4 vdd
port 513 nsew
rlabel metal1 s 2256 6860 2256 6860 4 vdd
port 513 nsew
rlabel metal1 s 1488 7359 1488 7359 4 vdd
port 513 nsew
rlabel metal1 s 1488 9230 1488 9230 4 vdd
port 513 nsew
rlabel metal1 s 1008 6569 1008 6569 4 vdd
port 513 nsew
rlabel metal1 s 1488 8149 1488 8149 4 vdd
port 513 nsew
rlabel metal1 s 1488 7650 1488 7650 4 vdd
port 513 nsew
rlabel metal1 s 1008 8149 1008 8149 4 vdd
port 513 nsew
rlabel metal1 s 240 9230 240 9230 4 vdd
port 513 nsew
rlabel metal1 s 240 8939 240 8939 4 vdd
port 513 nsew
rlabel metal1 s 2256 6569 2256 6569 4 vdd
port 513 nsew
rlabel metal1 s 1488 6860 1488 6860 4 vdd
port 513 nsew
rlabel metal1 s 1008 6860 1008 6860 4 vdd
port 513 nsew
rlabel metal1 s 240 8149 240 8149 4 vdd
port 513 nsew
rlabel metal1 s 2256 9230 2256 9230 4 vdd
port 513 nsew
rlabel metal1 s 1008 8440 1008 8440 4 vdd
port 513 nsew
rlabel metal1 s 1008 7650 1008 7650 4 vdd
port 513 nsew
rlabel metal1 s 240 7359 240 7359 4 vdd
port 513 nsew
rlabel metal1 s 2256 7650 2256 7650 4 vdd
port 513 nsew
rlabel metal1 s 2256 8939 2256 8939 4 vdd
port 513 nsew
rlabel metal1 s 240 7650 240 7650 4 vdd
port 513 nsew
rlabel metal1 s 1008 7359 1008 7359 4 vdd
port 513 nsew
rlabel metal1 s 240 6569 240 6569 4 vdd
port 513 nsew
rlabel metal1 s 1008 9230 1008 9230 4 vdd
port 513 nsew
rlabel metal1 s 2256 8440 2256 8440 4 vdd
port 513 nsew
rlabel metal1 s 240 6860 240 6860 4 vdd
port 513 nsew
rlabel metal1 s 1488 8939 1488 8939 4 vdd
port 513 nsew
rlabel metal1 s 3504 7650 3504 7650 4 vdd
port 513 nsew
rlabel metal1 s 3504 6860 3504 6860 4 vdd
port 513 nsew
rlabel metal1 s 2736 6860 2736 6860 4 vdd
port 513 nsew
rlabel metal1 s 4752 6860 4752 6860 4 vdd
port 513 nsew
rlabel metal1 s 2736 6569 2736 6569 4 vdd
port 513 nsew
rlabel metal1 s 3504 9230 3504 9230 4 vdd
port 513 nsew
rlabel metal1 s 3504 6569 3504 6569 4 vdd
port 513 nsew
rlabel metal1 s 4752 7359 4752 7359 4 vdd
port 513 nsew
rlabel metal1 s 3504 7359 3504 7359 4 vdd
port 513 nsew
rlabel metal1 s 2736 9230 2736 9230 4 vdd
port 513 nsew
rlabel metal1 s 3984 9230 3984 9230 4 vdd
port 513 nsew
rlabel metal1 s 3984 6569 3984 6569 4 vdd
port 513 nsew
rlabel metal1 s 4752 8440 4752 8440 4 vdd
port 513 nsew
rlabel metal1 s 3504 8149 3504 8149 4 vdd
port 513 nsew
rlabel metal1 s 3504 8939 3504 8939 4 vdd
port 513 nsew
rlabel metal1 s 3504 8440 3504 8440 4 vdd
port 513 nsew
rlabel metal1 s 2736 7359 2736 7359 4 vdd
port 513 nsew
rlabel metal1 s 2736 8939 2736 8939 4 vdd
port 513 nsew
rlabel metal1 s 3984 7359 3984 7359 4 vdd
port 513 nsew
rlabel metal1 s 3984 8149 3984 8149 4 vdd
port 513 nsew
rlabel metal1 s 2736 8149 2736 8149 4 vdd
port 513 nsew
rlabel metal1 s 4752 6569 4752 6569 4 vdd
port 513 nsew
rlabel metal1 s 3984 8440 3984 8440 4 vdd
port 513 nsew
rlabel metal1 s 3984 8939 3984 8939 4 vdd
port 513 nsew
rlabel metal1 s 3984 6860 3984 6860 4 vdd
port 513 nsew
rlabel metal1 s 4752 9230 4752 9230 4 vdd
port 513 nsew
rlabel metal1 s 4752 7650 4752 7650 4 vdd
port 513 nsew
rlabel metal1 s 2736 7650 2736 7650 4 vdd
port 513 nsew
rlabel metal1 s 2736 8440 2736 8440 4 vdd
port 513 nsew
rlabel metal1 s 4752 8939 4752 8939 4 vdd
port 513 nsew
rlabel metal1 s 3984 7650 3984 7650 4 vdd
port 513 nsew
rlabel metal1 s 4752 8149 4752 8149 4 vdd
port 513 nsew
rlabel metal1 s 3984 6070 3984 6070 4 vdd
port 513 nsew
rlabel metal1 s 3984 4199 3984 4199 4 vdd
port 513 nsew
rlabel metal1 s 4752 3409 4752 3409 4 vdd
port 513 nsew
rlabel metal1 s 3504 5280 3504 5280 4 vdd
port 513 nsew
rlabel metal1 s 3504 6070 3504 6070 4 vdd
port 513 nsew
rlabel metal1 s 3984 4490 3984 4490 4 vdd
port 513 nsew
rlabel metal1 s 4752 5779 4752 5779 4 vdd
port 513 nsew
rlabel metal1 s 4752 5280 4752 5280 4 vdd
port 513 nsew
rlabel metal1 s 3984 3700 3984 3700 4 vdd
port 513 nsew
rlabel metal1 s 4752 4199 4752 4199 4 vdd
port 513 nsew
rlabel metal1 s 3504 4490 3504 4490 4 vdd
port 513 nsew
rlabel metal1 s 3504 4199 3504 4199 4 vdd
port 513 nsew
rlabel metal1 s 3984 5280 3984 5280 4 vdd
port 513 nsew
rlabel metal1 s 2736 4490 2736 4490 4 vdd
port 513 nsew
rlabel metal1 s 3504 4989 3504 4989 4 vdd
port 513 nsew
rlabel metal1 s 4752 6070 4752 6070 4 vdd
port 513 nsew
rlabel metal1 s 2736 6070 2736 6070 4 vdd
port 513 nsew
rlabel metal1 s 4752 3700 4752 3700 4 vdd
port 513 nsew
rlabel metal1 s 4752 4989 4752 4989 4 vdd
port 513 nsew
rlabel metal1 s 3504 5779 3504 5779 4 vdd
port 513 nsew
rlabel metal1 s 3984 3409 3984 3409 4 vdd
port 513 nsew
rlabel metal1 s 2736 3700 2736 3700 4 vdd
port 513 nsew
rlabel metal1 s 2736 5779 2736 5779 4 vdd
port 513 nsew
rlabel metal1 s 3984 4989 3984 4989 4 vdd
port 513 nsew
rlabel metal1 s 4752 4490 4752 4490 4 vdd
port 513 nsew
rlabel metal1 s 2736 5280 2736 5280 4 vdd
port 513 nsew
rlabel metal1 s 2736 4199 2736 4199 4 vdd
port 513 nsew
rlabel metal1 s 3504 3409 3504 3409 4 vdd
port 513 nsew
rlabel metal1 s 3504 3700 3504 3700 4 vdd
port 513 nsew
rlabel metal1 s 3984 5779 3984 5779 4 vdd
port 513 nsew
rlabel metal1 s 2736 4989 2736 4989 4 vdd
port 513 nsew
rlabel metal1 s 2736 3409 2736 3409 4 vdd
port 513 nsew
rlabel metal1 s 2256 3700 2256 3700 4 vdd
port 513 nsew
rlabel metal1 s 1008 5280 1008 5280 4 vdd
port 513 nsew
rlabel metal1 s 1008 4199 1008 4199 4 vdd
port 513 nsew
rlabel metal1 s 240 3409 240 3409 4 vdd
port 513 nsew
rlabel metal1 s 2256 4989 2256 4989 4 vdd
port 513 nsew
rlabel metal1 s 2256 5779 2256 5779 4 vdd
port 513 nsew
rlabel metal1 s 240 5779 240 5779 4 vdd
port 513 nsew
rlabel metal1 s 2256 4199 2256 4199 4 vdd
port 513 nsew
rlabel metal1 s 1488 4989 1488 4989 4 vdd
port 513 nsew
rlabel metal1 s 1488 5280 1488 5280 4 vdd
port 513 nsew
rlabel metal1 s 2256 6070 2256 6070 4 vdd
port 513 nsew
rlabel metal1 s 2256 5280 2256 5280 4 vdd
port 513 nsew
rlabel metal1 s 1008 5779 1008 5779 4 vdd
port 513 nsew
rlabel metal1 s 240 4199 240 4199 4 vdd
port 513 nsew
rlabel metal1 s 2256 3409 2256 3409 4 vdd
port 513 nsew
rlabel metal1 s 1488 4199 1488 4199 4 vdd
port 513 nsew
rlabel metal1 s 1488 3700 1488 3700 4 vdd
port 513 nsew
rlabel metal1 s 1488 6070 1488 6070 4 vdd
port 513 nsew
rlabel metal1 s 1488 3409 1488 3409 4 vdd
port 513 nsew
rlabel metal1 s 1488 5779 1488 5779 4 vdd
port 513 nsew
rlabel metal1 s 240 4989 240 4989 4 vdd
port 513 nsew
rlabel metal1 s 240 6070 240 6070 4 vdd
port 513 nsew
rlabel metal1 s 240 3700 240 3700 4 vdd
port 513 nsew
rlabel metal1 s 240 4490 240 4490 4 vdd
port 513 nsew
rlabel metal1 s 1488 4490 1488 4490 4 vdd
port 513 nsew
rlabel metal1 s 1008 4490 1008 4490 4 vdd
port 513 nsew
rlabel metal1 s 240 5280 240 5280 4 vdd
port 513 nsew
rlabel metal1 s 1008 6070 1008 6070 4 vdd
port 513 nsew
rlabel metal1 s 1008 3700 1008 3700 4 vdd
port 513 nsew
rlabel metal1 s 2256 4490 2256 4490 4 vdd
port 513 nsew
rlabel metal1 s 1008 3409 1008 3409 4 vdd
port 513 nsew
rlabel metal1 s 1008 4989 1008 4989 4 vdd
port 513 nsew
rlabel metal1 s 2256 1330 2256 1330 4 vdd
port 513 nsew
rlabel metal1 s 1008 2120 1008 2120 4 vdd
port 513 nsew
rlabel metal1 s 240 1039 240 1039 4 vdd
port 513 nsew
rlabel metal1 s 240 1829 240 1829 4 vdd
port 513 nsew
rlabel metal1 s 1488 2120 1488 2120 4 vdd
port 513 nsew
rlabel metal1 s 1008 1330 1008 1330 4 vdd
port 513 nsew
rlabel metal1 s 240 2120 240 2120 4 vdd
port 513 nsew
rlabel metal1 s 1008 1829 1008 1829 4 vdd
port 513 nsew
rlabel metal1 s 1488 1330 1488 1330 4 vdd
port 513 nsew
rlabel metal1 s 1488 1039 1488 1039 4 vdd
port 513 nsew
rlabel metal1 s 240 2619 240 2619 4 vdd
port 513 nsew
rlabel metal1 s 240 540 240 540 4 vdd
port 513 nsew
rlabel metal1 s 2256 2120 2256 2120 4 vdd
port 513 nsew
rlabel metal1 s 240 249 240 249 4 vdd
port 513 nsew
rlabel metal1 s 2256 1829 2256 1829 4 vdd
port 513 nsew
rlabel metal1 s 1008 2910 1008 2910 4 vdd
port 513 nsew
rlabel metal1 s 1488 2619 1488 2619 4 vdd
port 513 nsew
rlabel metal1 s 2256 249 2256 249 4 vdd
port 513 nsew
rlabel metal1 s 1488 540 1488 540 4 vdd
port 513 nsew
rlabel metal1 s 1008 249 1008 249 4 vdd
port 513 nsew
rlabel metal1 s 1008 1039 1008 1039 4 vdd
port 513 nsew
rlabel metal1 s 1488 249 1488 249 4 vdd
port 513 nsew
rlabel metal1 s 1008 540 1008 540 4 vdd
port 513 nsew
rlabel metal1 s 1488 1829 1488 1829 4 vdd
port 513 nsew
rlabel metal1 s 2256 1039 2256 1039 4 vdd
port 513 nsew
rlabel metal1 s 240 2910 240 2910 4 vdd
port 513 nsew
rlabel metal1 s 240 1330 240 1330 4 vdd
port 513 nsew
rlabel metal1 s 1008 2619 1008 2619 4 vdd
port 513 nsew
rlabel metal1 s 2256 540 2256 540 4 vdd
port 513 nsew
rlabel metal1 s 1488 2910 1488 2910 4 vdd
port 513 nsew
rlabel metal1 s 2256 2910 2256 2910 4 vdd
port 513 nsew
rlabel metal1 s 2256 2619 2256 2619 4 vdd
port 513 nsew
rlabel metal1 s 4752 1039 4752 1039 4 vdd
port 513 nsew
rlabel metal1 s 3504 540 3504 540 4 vdd
port 513 nsew
rlabel metal1 s 3984 249 3984 249 4 vdd
port 513 nsew
rlabel metal1 s 4752 2619 4752 2619 4 vdd
port 513 nsew
rlabel metal1 s 3504 2120 3504 2120 4 vdd
port 513 nsew
rlabel metal1 s 3984 540 3984 540 4 vdd
port 513 nsew
rlabel metal1 s 4752 540 4752 540 4 vdd
port 513 nsew
rlabel metal1 s 3984 1829 3984 1829 4 vdd
port 513 nsew
rlabel metal1 s 4752 1829 4752 1829 4 vdd
port 513 nsew
rlabel metal1 s 3984 1039 3984 1039 4 vdd
port 513 nsew
rlabel metal1 s 4752 2120 4752 2120 4 vdd
port 513 nsew
rlabel metal1 s 2736 1330 2736 1330 4 vdd
port 513 nsew
rlabel metal1 s 3984 1330 3984 1330 4 vdd
port 513 nsew
rlabel metal1 s 2736 2120 2736 2120 4 vdd
port 513 nsew
rlabel metal1 s 3504 249 3504 249 4 vdd
port 513 nsew
rlabel metal1 s 4752 2910 4752 2910 4 vdd
port 513 nsew
rlabel metal1 s 2736 1829 2736 1829 4 vdd
port 513 nsew
rlabel metal1 s 3984 2910 3984 2910 4 vdd
port 513 nsew
rlabel metal1 s 3984 2120 3984 2120 4 vdd
port 513 nsew
rlabel metal1 s 2736 1039 2736 1039 4 vdd
port 513 nsew
rlabel metal1 s 4752 1330 4752 1330 4 vdd
port 513 nsew
rlabel metal1 s 2736 540 2736 540 4 vdd
port 513 nsew
rlabel metal1 s 2736 249 2736 249 4 vdd
port 513 nsew
rlabel metal1 s 3984 2619 3984 2619 4 vdd
port 513 nsew
rlabel metal1 s 2736 2619 2736 2619 4 vdd
port 513 nsew
rlabel metal1 s 3504 2910 3504 2910 4 vdd
port 513 nsew
rlabel metal1 s 2736 2910 2736 2910 4 vdd
port 513 nsew
rlabel metal1 s 3504 2619 3504 2619 4 vdd
port 513 nsew
rlabel metal1 s 3504 1330 3504 1330 4 vdd
port 513 nsew
rlabel metal1 s 3504 1039 3504 1039 4 vdd
port 513 nsew
rlabel metal1 s 3504 1829 3504 1829 4 vdd
port 513 nsew
rlabel metal1 s 4752 249 4752 249 4 vdd
port 513 nsew
rlabel metal1 s 9744 4989 9744 4989 4 vdd
port 513 nsew
rlabel metal1 s 7728 3700 7728 3700 4 vdd
port 513 nsew
rlabel metal1 s 8976 4490 8976 4490 4 vdd
port 513 nsew
rlabel metal1 s 8976 5280 8976 5280 4 vdd
port 513 nsew
rlabel metal1 s 8496 5779 8496 5779 4 vdd
port 513 nsew
rlabel metal1 s 7728 4490 7728 4490 4 vdd
port 513 nsew
rlabel metal1 s 8496 3409 8496 3409 4 vdd
port 513 nsew
rlabel metal1 s 8496 6070 8496 6070 4 vdd
port 513 nsew
rlabel metal1 s 8496 4989 8496 4989 4 vdd
port 513 nsew
rlabel metal1 s 9744 4490 9744 4490 4 vdd
port 513 nsew
rlabel metal1 s 8496 3700 8496 3700 4 vdd
port 513 nsew
rlabel metal1 s 8976 4989 8976 4989 4 vdd
port 513 nsew
rlabel metal1 s 8496 4199 8496 4199 4 vdd
port 513 nsew
rlabel metal1 s 7728 4989 7728 4989 4 vdd
port 513 nsew
rlabel metal1 s 8976 3409 8976 3409 4 vdd
port 513 nsew
rlabel metal1 s 9744 3409 9744 3409 4 vdd
port 513 nsew
rlabel metal1 s 8976 3700 8976 3700 4 vdd
port 513 nsew
rlabel metal1 s 7728 6070 7728 6070 4 vdd
port 513 nsew
rlabel metal1 s 8976 4199 8976 4199 4 vdd
port 513 nsew
rlabel metal1 s 7728 3409 7728 3409 4 vdd
port 513 nsew
rlabel metal1 s 8976 6070 8976 6070 4 vdd
port 513 nsew
rlabel metal1 s 7728 5280 7728 5280 4 vdd
port 513 nsew
rlabel metal1 s 9744 4199 9744 4199 4 vdd
port 513 nsew
rlabel metal1 s 8976 5779 8976 5779 4 vdd
port 513 nsew
rlabel metal1 s 9744 5779 9744 5779 4 vdd
port 513 nsew
rlabel metal1 s 7728 4199 7728 4199 4 vdd
port 513 nsew
rlabel metal1 s 8496 5280 8496 5280 4 vdd
port 513 nsew
rlabel metal1 s 7728 5779 7728 5779 4 vdd
port 513 nsew
rlabel metal1 s 9744 5280 9744 5280 4 vdd
port 513 nsew
rlabel metal1 s 8496 4490 8496 4490 4 vdd
port 513 nsew
rlabel metal1 s 9744 3700 9744 3700 4 vdd
port 513 nsew
rlabel metal1 s 9744 6070 9744 6070 4 vdd
port 513 nsew
rlabel metal1 s 5232 6070 5232 6070 4 vdd
port 513 nsew
rlabel metal1 s 6000 4490 6000 4490 4 vdd
port 513 nsew
rlabel metal1 s 6480 4199 6480 4199 4 vdd
port 513 nsew
rlabel metal1 s 6000 5280 6000 5280 4 vdd
port 513 nsew
rlabel metal1 s 6480 4989 6480 4989 4 vdd
port 513 nsew
rlabel metal1 s 6000 4199 6000 4199 4 vdd
port 513 nsew
rlabel metal1 s 6000 3700 6000 3700 4 vdd
port 513 nsew
rlabel metal1 s 7248 6070 7248 6070 4 vdd
port 513 nsew
rlabel metal1 s 5232 5280 5232 5280 4 vdd
port 513 nsew
rlabel metal1 s 6480 4490 6480 4490 4 vdd
port 513 nsew
rlabel metal1 s 7248 4199 7248 4199 4 vdd
port 513 nsew
rlabel metal1 s 6480 3700 6480 3700 4 vdd
port 513 nsew
rlabel metal1 s 5232 3700 5232 3700 4 vdd
port 513 nsew
rlabel metal1 s 5232 4490 5232 4490 4 vdd
port 513 nsew
rlabel metal1 s 7248 4490 7248 4490 4 vdd
port 513 nsew
rlabel metal1 s 6480 3409 6480 3409 4 vdd
port 513 nsew
rlabel metal1 s 5232 4989 5232 4989 4 vdd
port 513 nsew
rlabel metal1 s 5232 3409 5232 3409 4 vdd
port 513 nsew
rlabel metal1 s 7248 5280 7248 5280 4 vdd
port 513 nsew
rlabel metal1 s 7248 3409 7248 3409 4 vdd
port 513 nsew
rlabel metal1 s 7248 3700 7248 3700 4 vdd
port 513 nsew
rlabel metal1 s 6000 3409 6000 3409 4 vdd
port 513 nsew
rlabel metal1 s 6000 4989 6000 4989 4 vdd
port 513 nsew
rlabel metal1 s 6000 5779 6000 5779 4 vdd
port 513 nsew
rlabel metal1 s 7248 5779 7248 5779 4 vdd
port 513 nsew
rlabel metal1 s 6480 6070 6480 6070 4 vdd
port 513 nsew
rlabel metal1 s 5232 4199 5232 4199 4 vdd
port 513 nsew
rlabel metal1 s 7248 4989 7248 4989 4 vdd
port 513 nsew
rlabel metal1 s 6000 6070 6000 6070 4 vdd
port 513 nsew
rlabel metal1 s 5232 5779 5232 5779 4 vdd
port 513 nsew
rlabel metal1 s 6480 5779 6480 5779 4 vdd
port 513 nsew
rlabel metal1 s 6480 5280 6480 5280 4 vdd
port 513 nsew
rlabel metal1 s 5232 2619 5232 2619 4 vdd
port 513 nsew
rlabel metal1 s 6000 540 6000 540 4 vdd
port 513 nsew
rlabel metal1 s 7248 2619 7248 2619 4 vdd
port 513 nsew
rlabel metal1 s 6480 1829 6480 1829 4 vdd
port 513 nsew
rlabel metal1 s 6480 2619 6480 2619 4 vdd
port 513 nsew
rlabel metal1 s 5232 1829 5232 1829 4 vdd
port 513 nsew
rlabel metal1 s 7248 1330 7248 1330 4 vdd
port 513 nsew
rlabel metal1 s 6480 1039 6480 1039 4 vdd
port 513 nsew
rlabel metal1 s 6480 1330 6480 1330 4 vdd
port 513 nsew
rlabel metal1 s 5232 249 5232 249 4 vdd
port 513 nsew
rlabel metal1 s 7248 1039 7248 1039 4 vdd
port 513 nsew
rlabel metal1 s 6000 1829 6000 1829 4 vdd
port 513 nsew
rlabel metal1 s 7248 249 7248 249 4 vdd
port 513 nsew
rlabel metal1 s 6000 2120 6000 2120 4 vdd
port 513 nsew
rlabel metal1 s 6000 1039 6000 1039 4 vdd
port 513 nsew
rlabel metal1 s 6000 2619 6000 2619 4 vdd
port 513 nsew
rlabel metal1 s 7248 540 7248 540 4 vdd
port 513 nsew
rlabel metal1 s 6480 540 6480 540 4 vdd
port 513 nsew
rlabel metal1 s 6480 2910 6480 2910 4 vdd
port 513 nsew
rlabel metal1 s 5232 1039 5232 1039 4 vdd
port 513 nsew
rlabel metal1 s 6480 2120 6480 2120 4 vdd
port 513 nsew
rlabel metal1 s 5232 540 5232 540 4 vdd
port 513 nsew
rlabel metal1 s 6000 249 6000 249 4 vdd
port 513 nsew
rlabel metal1 s 5232 2120 5232 2120 4 vdd
port 513 nsew
rlabel metal1 s 5232 1330 5232 1330 4 vdd
port 513 nsew
rlabel metal1 s 6480 249 6480 249 4 vdd
port 513 nsew
rlabel metal1 s 5232 2910 5232 2910 4 vdd
port 513 nsew
rlabel metal1 s 6000 2910 6000 2910 4 vdd
port 513 nsew
rlabel metal1 s 7248 1829 7248 1829 4 vdd
port 513 nsew
rlabel metal1 s 7248 2910 7248 2910 4 vdd
port 513 nsew
rlabel metal1 s 7248 2120 7248 2120 4 vdd
port 513 nsew
rlabel metal1 s 6000 1330 6000 1330 4 vdd
port 513 nsew
rlabel metal1 s 8976 1039 8976 1039 4 vdd
port 513 nsew
rlabel metal1 s 8496 1330 8496 1330 4 vdd
port 513 nsew
rlabel metal1 s 9744 249 9744 249 4 vdd
port 513 nsew
rlabel metal1 s 8496 249 8496 249 4 vdd
port 513 nsew
rlabel metal1 s 8496 2910 8496 2910 4 vdd
port 513 nsew
rlabel metal1 s 8496 540 8496 540 4 vdd
port 513 nsew
rlabel metal1 s 8496 2120 8496 2120 4 vdd
port 513 nsew
rlabel metal1 s 7728 1039 7728 1039 4 vdd
port 513 nsew
rlabel metal1 s 8976 2619 8976 2619 4 vdd
port 513 nsew
rlabel metal1 s 9744 2120 9744 2120 4 vdd
port 513 nsew
rlabel metal1 s 9744 540 9744 540 4 vdd
port 513 nsew
rlabel metal1 s 8976 1829 8976 1829 4 vdd
port 513 nsew
rlabel metal1 s 8496 2619 8496 2619 4 vdd
port 513 nsew
rlabel metal1 s 7728 1330 7728 1330 4 vdd
port 513 nsew
rlabel metal1 s 8976 540 8976 540 4 vdd
port 513 nsew
rlabel metal1 s 9744 2619 9744 2619 4 vdd
port 513 nsew
rlabel metal1 s 8496 1039 8496 1039 4 vdd
port 513 nsew
rlabel metal1 s 8976 1330 8976 1330 4 vdd
port 513 nsew
rlabel metal1 s 9744 1829 9744 1829 4 vdd
port 513 nsew
rlabel metal1 s 8976 2910 8976 2910 4 vdd
port 513 nsew
rlabel metal1 s 9744 2910 9744 2910 4 vdd
port 513 nsew
rlabel metal1 s 7728 2120 7728 2120 4 vdd
port 513 nsew
rlabel metal1 s 8976 2120 8976 2120 4 vdd
port 513 nsew
rlabel metal1 s 7728 540 7728 540 4 vdd
port 513 nsew
rlabel metal1 s 9744 1039 9744 1039 4 vdd
port 513 nsew
rlabel metal1 s 7728 2910 7728 2910 4 vdd
port 513 nsew
rlabel metal1 s 8976 249 8976 249 4 vdd
port 513 nsew
rlabel metal1 s 7728 2619 7728 2619 4 vdd
port 513 nsew
rlabel metal1 s 8496 1829 8496 1829 4 vdd
port 513 nsew
rlabel metal1 s 7728 249 7728 249 4 vdd
port 513 nsew
rlabel metal1 s 7728 1829 7728 1829 4 vdd
port 513 nsew
rlabel metal1 s 9744 1330 9744 1330 4 vdd
port 513 nsew
rlabel metal1 s 18480 11309 18480 11309 4 vdd
port 513 nsew
rlabel metal1 s 19728 12099 19728 12099 4 vdd
port 513 nsew
rlabel metal1 s 18960 10020 18960 10020 4 vdd
port 513 nsew
rlabel metal1 s 17712 9729 17712 9729 4 vdd
port 513 nsew
rlabel metal1 s 19728 11600 19728 11600 4 vdd
port 513 nsew
rlabel metal1 s 17712 10810 17712 10810 4 vdd
port 513 nsew
rlabel metal1 s 18480 10519 18480 10519 4 vdd
port 513 nsew
rlabel metal1 s 19728 12390 19728 12390 4 vdd
port 513 nsew
rlabel metal1 s 18960 12390 18960 12390 4 vdd
port 513 nsew
rlabel metal1 s 18480 9729 18480 9729 4 vdd
port 513 nsew
rlabel metal1 s 18960 11600 18960 11600 4 vdd
port 513 nsew
rlabel metal1 s 18960 12099 18960 12099 4 vdd
port 513 nsew
rlabel metal1 s 19728 10810 19728 10810 4 vdd
port 513 nsew
rlabel metal1 s 17712 12390 17712 12390 4 vdd
port 513 nsew
rlabel metal1 s 18960 9729 18960 9729 4 vdd
port 513 nsew
rlabel metal1 s 17712 11600 17712 11600 4 vdd
port 513 nsew
rlabel metal1 s 17712 11309 17712 11309 4 vdd
port 513 nsew
rlabel metal1 s 19728 10020 19728 10020 4 vdd
port 513 nsew
rlabel metal1 s 18960 11309 18960 11309 4 vdd
port 513 nsew
rlabel metal1 s 19728 10519 19728 10519 4 vdd
port 513 nsew
rlabel metal1 s 18960 10810 18960 10810 4 vdd
port 513 nsew
rlabel metal1 s 18480 10020 18480 10020 4 vdd
port 513 nsew
rlabel metal1 s 18480 11600 18480 11600 4 vdd
port 513 nsew
rlabel metal1 s 18480 12390 18480 12390 4 vdd
port 513 nsew
rlabel metal1 s 17712 10020 17712 10020 4 vdd
port 513 nsew
rlabel metal1 s 18960 10519 18960 10519 4 vdd
port 513 nsew
rlabel metal1 s 19728 11309 19728 11309 4 vdd
port 513 nsew
rlabel metal1 s 19728 9729 19728 9729 4 vdd
port 513 nsew
rlabel metal1 s 18480 10810 18480 10810 4 vdd
port 513 nsew
rlabel metal1 s 17712 12099 17712 12099 4 vdd
port 513 nsew
rlabel metal1 s 18480 12099 18480 12099 4 vdd
port 513 nsew
rlabel metal1 s 17712 10519 17712 10519 4 vdd
port 513 nsew
rlabel metal1 s 15216 10810 15216 10810 4 vdd
port 513 nsew
rlabel metal1 s 17232 10519 17232 10519 4 vdd
port 513 nsew
rlabel metal1 s 15216 10519 15216 10519 4 vdd
port 513 nsew
rlabel metal1 s 16464 10519 16464 10519 4 vdd
port 513 nsew
rlabel metal1 s 15216 12099 15216 12099 4 vdd
port 513 nsew
rlabel metal1 s 15984 10519 15984 10519 4 vdd
port 513 nsew
rlabel metal1 s 15216 11600 15216 11600 4 vdd
port 513 nsew
rlabel metal1 s 15216 11309 15216 11309 4 vdd
port 513 nsew
rlabel metal1 s 15984 12390 15984 12390 4 vdd
port 513 nsew
rlabel metal1 s 15216 12390 15216 12390 4 vdd
port 513 nsew
rlabel metal1 s 15984 12099 15984 12099 4 vdd
port 513 nsew
rlabel metal1 s 15216 10020 15216 10020 4 vdd
port 513 nsew
rlabel metal1 s 16464 11309 16464 11309 4 vdd
port 513 nsew
rlabel metal1 s 15984 10020 15984 10020 4 vdd
port 513 nsew
rlabel metal1 s 15984 9729 15984 9729 4 vdd
port 513 nsew
rlabel metal1 s 17232 9729 17232 9729 4 vdd
port 513 nsew
rlabel metal1 s 17232 12390 17232 12390 4 vdd
port 513 nsew
rlabel metal1 s 15984 11600 15984 11600 4 vdd
port 513 nsew
rlabel metal1 s 16464 12099 16464 12099 4 vdd
port 513 nsew
rlabel metal1 s 17232 11600 17232 11600 4 vdd
port 513 nsew
rlabel metal1 s 16464 9729 16464 9729 4 vdd
port 513 nsew
rlabel metal1 s 17232 12099 17232 12099 4 vdd
port 513 nsew
rlabel metal1 s 17232 10020 17232 10020 4 vdd
port 513 nsew
rlabel metal1 s 15216 9729 15216 9729 4 vdd
port 513 nsew
rlabel metal1 s 15984 11309 15984 11309 4 vdd
port 513 nsew
rlabel metal1 s 16464 10810 16464 10810 4 vdd
port 513 nsew
rlabel metal1 s 16464 11600 16464 11600 4 vdd
port 513 nsew
rlabel metal1 s 17232 11309 17232 11309 4 vdd
port 513 nsew
rlabel metal1 s 17232 10810 17232 10810 4 vdd
port 513 nsew
rlabel metal1 s 16464 10020 16464 10020 4 vdd
port 513 nsew
rlabel metal1 s 15984 10810 15984 10810 4 vdd
port 513 nsew
rlabel metal1 s 16464 12390 16464 12390 4 vdd
port 513 nsew
rlabel metal1 s 16464 6569 16464 6569 4 vdd
port 513 nsew
rlabel metal1 s 16464 8939 16464 8939 4 vdd
port 513 nsew
rlabel metal1 s 15216 6860 15216 6860 4 vdd
port 513 nsew
rlabel metal1 s 17232 8939 17232 8939 4 vdd
port 513 nsew
rlabel metal1 s 15216 8149 15216 8149 4 vdd
port 513 nsew
rlabel metal1 s 15984 6569 15984 6569 4 vdd
port 513 nsew
rlabel metal1 s 15984 8149 15984 8149 4 vdd
port 513 nsew
rlabel metal1 s 17232 8440 17232 8440 4 vdd
port 513 nsew
rlabel metal1 s 15216 8440 15216 8440 4 vdd
port 513 nsew
rlabel metal1 s 15216 6569 15216 6569 4 vdd
port 513 nsew
rlabel metal1 s 15216 9230 15216 9230 4 vdd
port 513 nsew
rlabel metal1 s 17232 6860 17232 6860 4 vdd
port 513 nsew
rlabel metal1 s 17232 9230 17232 9230 4 vdd
port 513 nsew
rlabel metal1 s 15216 8939 15216 8939 4 vdd
port 513 nsew
rlabel metal1 s 15984 8939 15984 8939 4 vdd
port 513 nsew
rlabel metal1 s 15216 7650 15216 7650 4 vdd
port 513 nsew
rlabel metal1 s 15984 7359 15984 7359 4 vdd
port 513 nsew
rlabel metal1 s 15216 7359 15216 7359 4 vdd
port 513 nsew
rlabel metal1 s 17232 7650 17232 7650 4 vdd
port 513 nsew
rlabel metal1 s 15984 8440 15984 8440 4 vdd
port 513 nsew
rlabel metal1 s 17232 7359 17232 7359 4 vdd
port 513 nsew
rlabel metal1 s 16464 7359 16464 7359 4 vdd
port 513 nsew
rlabel metal1 s 16464 6860 16464 6860 4 vdd
port 513 nsew
rlabel metal1 s 16464 8149 16464 8149 4 vdd
port 513 nsew
rlabel metal1 s 17232 8149 17232 8149 4 vdd
port 513 nsew
rlabel metal1 s 16464 7650 16464 7650 4 vdd
port 513 nsew
rlabel metal1 s 15984 6860 15984 6860 4 vdd
port 513 nsew
rlabel metal1 s 17232 6569 17232 6569 4 vdd
port 513 nsew
rlabel metal1 s 16464 9230 16464 9230 4 vdd
port 513 nsew
rlabel metal1 s 15984 9230 15984 9230 4 vdd
port 513 nsew
rlabel metal1 s 15984 7650 15984 7650 4 vdd
port 513 nsew
rlabel metal1 s 16464 8440 16464 8440 4 vdd
port 513 nsew
rlabel metal1 s 19728 7650 19728 7650 4 vdd
port 513 nsew
rlabel metal1 s 17712 9230 17712 9230 4 vdd
port 513 nsew
rlabel metal1 s 17712 6860 17712 6860 4 vdd
port 513 nsew
rlabel metal1 s 18960 6569 18960 6569 4 vdd
port 513 nsew
rlabel metal1 s 18960 8440 18960 8440 4 vdd
port 513 nsew
rlabel metal1 s 17712 8440 17712 8440 4 vdd
port 513 nsew
rlabel metal1 s 19728 6569 19728 6569 4 vdd
port 513 nsew
rlabel metal1 s 17712 7650 17712 7650 4 vdd
port 513 nsew
rlabel metal1 s 18480 9230 18480 9230 4 vdd
port 513 nsew
rlabel metal1 s 18960 9230 18960 9230 4 vdd
port 513 nsew
rlabel metal1 s 18480 6569 18480 6569 4 vdd
port 513 nsew
rlabel metal1 s 18960 7359 18960 7359 4 vdd
port 513 nsew
rlabel metal1 s 18480 6860 18480 6860 4 vdd
port 513 nsew
rlabel metal1 s 19728 8440 19728 8440 4 vdd
port 513 nsew
rlabel metal1 s 17712 7359 17712 7359 4 vdd
port 513 nsew
rlabel metal1 s 19728 9230 19728 9230 4 vdd
port 513 nsew
rlabel metal1 s 19728 6860 19728 6860 4 vdd
port 513 nsew
rlabel metal1 s 18960 8149 18960 8149 4 vdd
port 513 nsew
rlabel metal1 s 17712 8939 17712 8939 4 vdd
port 513 nsew
rlabel metal1 s 19728 7359 19728 7359 4 vdd
port 513 nsew
rlabel metal1 s 18480 7359 18480 7359 4 vdd
port 513 nsew
rlabel metal1 s 18960 6860 18960 6860 4 vdd
port 513 nsew
rlabel metal1 s 17712 6569 17712 6569 4 vdd
port 513 nsew
rlabel metal1 s 19728 8149 19728 8149 4 vdd
port 513 nsew
rlabel metal1 s 18480 8149 18480 8149 4 vdd
port 513 nsew
rlabel metal1 s 18960 8939 18960 8939 4 vdd
port 513 nsew
rlabel metal1 s 17712 8149 17712 8149 4 vdd
port 513 nsew
rlabel metal1 s 18960 7650 18960 7650 4 vdd
port 513 nsew
rlabel metal1 s 19728 8939 19728 8939 4 vdd
port 513 nsew
rlabel metal1 s 18480 8440 18480 8440 4 vdd
port 513 nsew
rlabel metal1 s 18480 7650 18480 7650 4 vdd
port 513 nsew
rlabel metal1 s 18480 8939 18480 8939 4 vdd
port 513 nsew
rlabel metal1 s 14736 11309 14736 11309 4 vdd
port 513 nsew
rlabel metal1 s 13488 11600 13488 11600 4 vdd
port 513 nsew
rlabel metal1 s 14736 11600 14736 11600 4 vdd
port 513 nsew
rlabel metal1 s 14736 12099 14736 12099 4 vdd
port 513 nsew
rlabel metal1 s 13968 9729 13968 9729 4 vdd
port 513 nsew
rlabel metal1 s 12720 9729 12720 9729 4 vdd
port 513 nsew
rlabel metal1 s 12720 12390 12720 12390 4 vdd
port 513 nsew
rlabel metal1 s 13968 11600 13968 11600 4 vdd
port 513 nsew
rlabel metal1 s 13968 11309 13968 11309 4 vdd
port 513 nsew
rlabel metal1 s 13968 10810 13968 10810 4 vdd
port 513 nsew
rlabel metal1 s 14736 10810 14736 10810 4 vdd
port 513 nsew
rlabel metal1 s 12720 11600 12720 11600 4 vdd
port 513 nsew
rlabel metal1 s 13488 12099 13488 12099 4 vdd
port 513 nsew
rlabel metal1 s 13488 10020 13488 10020 4 vdd
port 513 nsew
rlabel metal1 s 12720 10020 12720 10020 4 vdd
port 513 nsew
rlabel metal1 s 13968 12390 13968 12390 4 vdd
port 513 nsew
rlabel metal1 s 12720 12099 12720 12099 4 vdd
port 513 nsew
rlabel metal1 s 13968 10020 13968 10020 4 vdd
port 513 nsew
rlabel metal1 s 12720 10519 12720 10519 4 vdd
port 513 nsew
rlabel metal1 s 12720 10810 12720 10810 4 vdd
port 513 nsew
rlabel metal1 s 14736 12390 14736 12390 4 vdd
port 513 nsew
rlabel metal1 s 13488 12390 13488 12390 4 vdd
port 513 nsew
rlabel metal1 s 14736 9729 14736 9729 4 vdd
port 513 nsew
rlabel metal1 s 13488 11309 13488 11309 4 vdd
port 513 nsew
rlabel metal1 s 14736 10519 14736 10519 4 vdd
port 513 nsew
rlabel metal1 s 13968 12099 13968 12099 4 vdd
port 513 nsew
rlabel metal1 s 13968 10519 13968 10519 4 vdd
port 513 nsew
rlabel metal1 s 14736 10020 14736 10020 4 vdd
port 513 nsew
rlabel metal1 s 13488 10519 13488 10519 4 vdd
port 513 nsew
rlabel metal1 s 12720 11309 12720 11309 4 vdd
port 513 nsew
rlabel metal1 s 13488 9729 13488 9729 4 vdd
port 513 nsew
rlabel metal1 s 13488 10810 13488 10810 4 vdd
port 513 nsew
rlabel metal1 s 12240 12390 12240 12390 4 vdd
port 513 nsew
rlabel metal1 s 11472 10810 11472 10810 4 vdd
port 513 nsew
rlabel metal1 s 10992 10810 10992 10810 4 vdd
port 513 nsew
rlabel metal1 s 12240 12099 12240 12099 4 vdd
port 513 nsew
rlabel metal1 s 10992 12390 10992 12390 4 vdd
port 513 nsew
rlabel metal1 s 11472 12390 11472 12390 4 vdd
port 513 nsew
rlabel metal1 s 10224 12390 10224 12390 4 vdd
port 513 nsew
rlabel metal1 s 11472 10020 11472 10020 4 vdd
port 513 nsew
rlabel metal1 s 12240 10519 12240 10519 4 vdd
port 513 nsew
rlabel metal1 s 12240 10810 12240 10810 4 vdd
port 513 nsew
rlabel metal1 s 11472 10519 11472 10519 4 vdd
port 513 nsew
rlabel metal1 s 10992 11600 10992 11600 4 vdd
port 513 nsew
rlabel metal1 s 10224 10810 10224 10810 4 vdd
port 513 nsew
rlabel metal1 s 12240 10020 12240 10020 4 vdd
port 513 nsew
rlabel metal1 s 11472 9729 11472 9729 4 vdd
port 513 nsew
rlabel metal1 s 10224 9729 10224 9729 4 vdd
port 513 nsew
rlabel metal1 s 12240 11309 12240 11309 4 vdd
port 513 nsew
rlabel metal1 s 10992 10519 10992 10519 4 vdd
port 513 nsew
rlabel metal1 s 10992 11309 10992 11309 4 vdd
port 513 nsew
rlabel metal1 s 10224 12099 10224 12099 4 vdd
port 513 nsew
rlabel metal1 s 10992 10020 10992 10020 4 vdd
port 513 nsew
rlabel metal1 s 11472 11309 11472 11309 4 vdd
port 513 nsew
rlabel metal1 s 10992 12099 10992 12099 4 vdd
port 513 nsew
rlabel metal1 s 12240 9729 12240 9729 4 vdd
port 513 nsew
rlabel metal1 s 10224 11600 10224 11600 4 vdd
port 513 nsew
rlabel metal1 s 10224 11309 10224 11309 4 vdd
port 513 nsew
rlabel metal1 s 11472 11600 11472 11600 4 vdd
port 513 nsew
rlabel metal1 s 10992 9729 10992 9729 4 vdd
port 513 nsew
rlabel metal1 s 10224 10519 10224 10519 4 vdd
port 513 nsew
rlabel metal1 s 10224 10020 10224 10020 4 vdd
port 513 nsew
rlabel metal1 s 11472 12099 11472 12099 4 vdd
port 513 nsew
rlabel metal1 s 12240 11600 12240 11600 4 vdd
port 513 nsew
rlabel metal1 s 11472 6569 11472 6569 4 vdd
port 513 nsew
rlabel metal1 s 10224 9230 10224 9230 4 vdd
port 513 nsew
rlabel metal1 s 10224 6860 10224 6860 4 vdd
port 513 nsew
rlabel metal1 s 11472 8440 11472 8440 4 vdd
port 513 nsew
rlabel metal1 s 12240 7650 12240 7650 4 vdd
port 513 nsew
rlabel metal1 s 10992 8440 10992 8440 4 vdd
port 513 nsew
rlabel metal1 s 10224 8939 10224 8939 4 vdd
port 513 nsew
rlabel metal1 s 11472 8149 11472 8149 4 vdd
port 513 nsew
rlabel metal1 s 10992 7359 10992 7359 4 vdd
port 513 nsew
rlabel metal1 s 10992 6569 10992 6569 4 vdd
port 513 nsew
rlabel metal1 s 12240 6569 12240 6569 4 vdd
port 513 nsew
rlabel metal1 s 12240 8939 12240 8939 4 vdd
port 513 nsew
rlabel metal1 s 10992 9230 10992 9230 4 vdd
port 513 nsew
rlabel metal1 s 10224 8149 10224 8149 4 vdd
port 513 nsew
rlabel metal1 s 10992 6860 10992 6860 4 vdd
port 513 nsew
rlabel metal1 s 10224 7359 10224 7359 4 vdd
port 513 nsew
rlabel metal1 s 10224 7650 10224 7650 4 vdd
port 513 nsew
rlabel metal1 s 11472 8939 11472 8939 4 vdd
port 513 nsew
rlabel metal1 s 12240 8149 12240 8149 4 vdd
port 513 nsew
rlabel metal1 s 10224 6569 10224 6569 4 vdd
port 513 nsew
rlabel metal1 s 12240 7359 12240 7359 4 vdd
port 513 nsew
rlabel metal1 s 12240 6860 12240 6860 4 vdd
port 513 nsew
rlabel metal1 s 10992 8149 10992 8149 4 vdd
port 513 nsew
rlabel metal1 s 10992 7650 10992 7650 4 vdd
port 513 nsew
rlabel metal1 s 11472 7359 11472 7359 4 vdd
port 513 nsew
rlabel metal1 s 11472 9230 11472 9230 4 vdd
port 513 nsew
rlabel metal1 s 11472 6860 11472 6860 4 vdd
port 513 nsew
rlabel metal1 s 11472 7650 11472 7650 4 vdd
port 513 nsew
rlabel metal1 s 10992 8939 10992 8939 4 vdd
port 513 nsew
rlabel metal1 s 12240 8440 12240 8440 4 vdd
port 513 nsew
rlabel metal1 s 10224 8440 10224 8440 4 vdd
port 513 nsew
rlabel metal1 s 12240 9230 12240 9230 4 vdd
port 513 nsew
rlabel metal1 s 13488 6569 13488 6569 4 vdd
port 513 nsew
rlabel metal1 s 13488 8149 13488 8149 4 vdd
port 513 nsew
rlabel metal1 s 13968 8440 13968 8440 4 vdd
port 513 nsew
rlabel metal1 s 13968 7359 13968 7359 4 vdd
port 513 nsew
rlabel metal1 s 13488 8440 13488 8440 4 vdd
port 513 nsew
rlabel metal1 s 13488 9230 13488 9230 4 vdd
port 513 nsew
rlabel metal1 s 13488 6860 13488 6860 4 vdd
port 513 nsew
rlabel metal1 s 12720 8939 12720 8939 4 vdd
port 513 nsew
rlabel metal1 s 12720 6569 12720 6569 4 vdd
port 513 nsew
rlabel metal1 s 12720 7650 12720 7650 4 vdd
port 513 nsew
rlabel metal1 s 13488 8939 13488 8939 4 vdd
port 513 nsew
rlabel metal1 s 14736 9230 14736 9230 4 vdd
port 513 nsew
rlabel metal1 s 14736 6860 14736 6860 4 vdd
port 513 nsew
rlabel metal1 s 13488 7359 13488 7359 4 vdd
port 513 nsew
rlabel metal1 s 13968 6860 13968 6860 4 vdd
port 513 nsew
rlabel metal1 s 12720 9230 12720 9230 4 vdd
port 513 nsew
rlabel metal1 s 12720 8149 12720 8149 4 vdd
port 513 nsew
rlabel metal1 s 12720 7359 12720 7359 4 vdd
port 513 nsew
rlabel metal1 s 14736 7650 14736 7650 4 vdd
port 513 nsew
rlabel metal1 s 13968 9230 13968 9230 4 vdd
port 513 nsew
rlabel metal1 s 14736 6569 14736 6569 4 vdd
port 513 nsew
rlabel metal1 s 14736 8939 14736 8939 4 vdd
port 513 nsew
rlabel metal1 s 13488 7650 13488 7650 4 vdd
port 513 nsew
rlabel metal1 s 14736 8440 14736 8440 4 vdd
port 513 nsew
rlabel metal1 s 13968 8939 13968 8939 4 vdd
port 513 nsew
rlabel metal1 s 14736 7359 14736 7359 4 vdd
port 513 nsew
rlabel metal1 s 14736 8149 14736 8149 4 vdd
port 513 nsew
rlabel metal1 s 13968 6569 13968 6569 4 vdd
port 513 nsew
rlabel metal1 s 13968 7650 13968 7650 4 vdd
port 513 nsew
rlabel metal1 s 12720 8440 12720 8440 4 vdd
port 513 nsew
rlabel metal1 s 13968 8149 13968 8149 4 vdd
port 513 nsew
rlabel metal1 s 12720 6860 12720 6860 4 vdd
port 513 nsew
rlabel metal1 s 13488 4989 13488 4989 4 vdd
port 513 nsew
rlabel metal1 s 13968 5280 13968 5280 4 vdd
port 513 nsew
rlabel metal1 s 14736 4989 14736 4989 4 vdd
port 513 nsew
rlabel metal1 s 12720 4989 12720 4989 4 vdd
port 513 nsew
rlabel metal1 s 13968 3700 13968 3700 4 vdd
port 513 nsew
rlabel metal1 s 14736 5779 14736 5779 4 vdd
port 513 nsew
rlabel metal1 s 12720 3700 12720 3700 4 vdd
port 513 nsew
rlabel metal1 s 12720 5280 12720 5280 4 vdd
port 513 nsew
rlabel metal1 s 12720 4490 12720 4490 4 vdd
port 513 nsew
rlabel metal1 s 13488 5779 13488 5779 4 vdd
port 513 nsew
rlabel metal1 s 14736 6070 14736 6070 4 vdd
port 513 nsew
rlabel metal1 s 14736 3700 14736 3700 4 vdd
port 513 nsew
rlabel metal1 s 12720 5779 12720 5779 4 vdd
port 513 nsew
rlabel metal1 s 13488 4490 13488 4490 4 vdd
port 513 nsew
rlabel metal1 s 13488 4199 13488 4199 4 vdd
port 513 nsew
rlabel metal1 s 13968 4989 13968 4989 4 vdd
port 513 nsew
rlabel metal1 s 12720 3409 12720 3409 4 vdd
port 513 nsew
rlabel metal1 s 14736 4199 14736 4199 4 vdd
port 513 nsew
rlabel metal1 s 13488 5280 13488 5280 4 vdd
port 513 nsew
rlabel metal1 s 13968 6070 13968 6070 4 vdd
port 513 nsew
rlabel metal1 s 12720 4199 12720 4199 4 vdd
port 513 nsew
rlabel metal1 s 13488 6070 13488 6070 4 vdd
port 513 nsew
rlabel metal1 s 14736 3409 14736 3409 4 vdd
port 513 nsew
rlabel metal1 s 13968 4490 13968 4490 4 vdd
port 513 nsew
rlabel metal1 s 14736 5280 14736 5280 4 vdd
port 513 nsew
rlabel metal1 s 13968 4199 13968 4199 4 vdd
port 513 nsew
rlabel metal1 s 13488 3409 13488 3409 4 vdd
port 513 nsew
rlabel metal1 s 13968 3409 13968 3409 4 vdd
port 513 nsew
rlabel metal1 s 14736 4490 14736 4490 4 vdd
port 513 nsew
rlabel metal1 s 13968 5779 13968 5779 4 vdd
port 513 nsew
rlabel metal1 s 12720 6070 12720 6070 4 vdd
port 513 nsew
rlabel metal1 s 13488 3700 13488 3700 4 vdd
port 513 nsew
rlabel metal1 s 10224 6070 10224 6070 4 vdd
port 513 nsew
rlabel metal1 s 10224 5280 10224 5280 4 vdd
port 513 nsew
rlabel metal1 s 11472 6070 11472 6070 4 vdd
port 513 nsew
rlabel metal1 s 12240 5779 12240 5779 4 vdd
port 513 nsew
rlabel metal1 s 10224 4490 10224 4490 4 vdd
port 513 nsew
rlabel metal1 s 12240 3700 12240 3700 4 vdd
port 513 nsew
rlabel metal1 s 12240 3409 12240 3409 4 vdd
port 513 nsew
rlabel metal1 s 11472 5779 11472 5779 4 vdd
port 513 nsew
rlabel metal1 s 10992 4199 10992 4199 4 vdd
port 513 nsew
rlabel metal1 s 10992 4490 10992 4490 4 vdd
port 513 nsew
rlabel metal1 s 10224 4199 10224 4199 4 vdd
port 513 nsew
rlabel metal1 s 12240 4989 12240 4989 4 vdd
port 513 nsew
rlabel metal1 s 11472 3700 11472 3700 4 vdd
port 513 nsew
rlabel metal1 s 12240 6070 12240 6070 4 vdd
port 513 nsew
rlabel metal1 s 10992 5280 10992 5280 4 vdd
port 513 nsew
rlabel metal1 s 11472 4199 11472 4199 4 vdd
port 513 nsew
rlabel metal1 s 10224 5779 10224 5779 4 vdd
port 513 nsew
rlabel metal1 s 10224 3409 10224 3409 4 vdd
port 513 nsew
rlabel metal1 s 12240 4490 12240 4490 4 vdd
port 513 nsew
rlabel metal1 s 10224 3700 10224 3700 4 vdd
port 513 nsew
rlabel metal1 s 10992 3409 10992 3409 4 vdd
port 513 nsew
rlabel metal1 s 10224 4989 10224 4989 4 vdd
port 513 nsew
rlabel metal1 s 11472 3409 11472 3409 4 vdd
port 513 nsew
rlabel metal1 s 11472 5280 11472 5280 4 vdd
port 513 nsew
rlabel metal1 s 10992 3700 10992 3700 4 vdd
port 513 nsew
rlabel metal1 s 10992 6070 10992 6070 4 vdd
port 513 nsew
rlabel metal1 s 10992 5779 10992 5779 4 vdd
port 513 nsew
rlabel metal1 s 12240 5280 12240 5280 4 vdd
port 513 nsew
rlabel metal1 s 10992 4989 10992 4989 4 vdd
port 513 nsew
rlabel metal1 s 11472 4490 11472 4490 4 vdd
port 513 nsew
rlabel metal1 s 11472 4989 11472 4989 4 vdd
port 513 nsew
rlabel metal1 s 12240 4199 12240 4199 4 vdd
port 513 nsew
rlabel metal1 s 10224 1829 10224 1829 4 vdd
port 513 nsew
rlabel metal1 s 11472 2910 11472 2910 4 vdd
port 513 nsew
rlabel metal1 s 11472 1829 11472 1829 4 vdd
port 513 nsew
rlabel metal1 s 11472 2120 11472 2120 4 vdd
port 513 nsew
rlabel metal1 s 10224 1330 10224 1330 4 vdd
port 513 nsew
rlabel metal1 s 10992 249 10992 249 4 vdd
port 513 nsew
rlabel metal1 s 11472 1330 11472 1330 4 vdd
port 513 nsew
rlabel metal1 s 10992 1039 10992 1039 4 vdd
port 513 nsew
rlabel metal1 s 10992 540 10992 540 4 vdd
port 513 nsew
rlabel metal1 s 10224 249 10224 249 4 vdd
port 513 nsew
rlabel metal1 s 11472 540 11472 540 4 vdd
port 513 nsew
rlabel metal1 s 10224 1039 10224 1039 4 vdd
port 513 nsew
rlabel metal1 s 12240 1330 12240 1330 4 vdd
port 513 nsew
rlabel metal1 s 10224 540 10224 540 4 vdd
port 513 nsew
rlabel metal1 s 12240 540 12240 540 4 vdd
port 513 nsew
rlabel metal1 s 10992 2120 10992 2120 4 vdd
port 513 nsew
rlabel metal1 s 10992 2619 10992 2619 4 vdd
port 513 nsew
rlabel metal1 s 11472 249 11472 249 4 vdd
port 513 nsew
rlabel metal1 s 12240 1039 12240 1039 4 vdd
port 513 nsew
rlabel metal1 s 10992 1829 10992 1829 4 vdd
port 513 nsew
rlabel metal1 s 12240 2619 12240 2619 4 vdd
port 513 nsew
rlabel metal1 s 12240 2120 12240 2120 4 vdd
port 513 nsew
rlabel metal1 s 12240 249 12240 249 4 vdd
port 513 nsew
rlabel metal1 s 10992 2910 10992 2910 4 vdd
port 513 nsew
rlabel metal1 s 12240 2910 12240 2910 4 vdd
port 513 nsew
rlabel metal1 s 11472 2619 11472 2619 4 vdd
port 513 nsew
rlabel metal1 s 10224 2619 10224 2619 4 vdd
port 513 nsew
rlabel metal1 s 10224 2120 10224 2120 4 vdd
port 513 nsew
rlabel metal1 s 10224 2910 10224 2910 4 vdd
port 513 nsew
rlabel metal1 s 10992 1330 10992 1330 4 vdd
port 513 nsew
rlabel metal1 s 12240 1829 12240 1829 4 vdd
port 513 nsew
rlabel metal1 s 11472 1039 11472 1039 4 vdd
port 513 nsew
rlabel metal1 s 13968 2619 13968 2619 4 vdd
port 513 nsew
rlabel metal1 s 13488 1330 13488 1330 4 vdd
port 513 nsew
rlabel metal1 s 13968 2120 13968 2120 4 vdd
port 513 nsew
rlabel metal1 s 13488 540 13488 540 4 vdd
port 513 nsew
rlabel metal1 s 13488 2910 13488 2910 4 vdd
port 513 nsew
rlabel metal1 s 13488 1829 13488 1829 4 vdd
port 513 nsew
rlabel metal1 s 12720 2910 12720 2910 4 vdd
port 513 nsew
rlabel metal1 s 13968 540 13968 540 4 vdd
port 513 nsew
rlabel metal1 s 14736 249 14736 249 4 vdd
port 513 nsew
rlabel metal1 s 13968 249 13968 249 4 vdd
port 513 nsew
rlabel metal1 s 13968 2910 13968 2910 4 vdd
port 513 nsew
rlabel metal1 s 12720 1039 12720 1039 4 vdd
port 513 nsew
rlabel metal1 s 12720 2619 12720 2619 4 vdd
port 513 nsew
rlabel metal1 s 13488 1039 13488 1039 4 vdd
port 513 nsew
rlabel metal1 s 14736 1039 14736 1039 4 vdd
port 513 nsew
rlabel metal1 s 14736 540 14736 540 4 vdd
port 513 nsew
rlabel metal1 s 14736 1330 14736 1330 4 vdd
port 513 nsew
rlabel metal1 s 13488 2619 13488 2619 4 vdd
port 513 nsew
rlabel metal1 s 13968 1330 13968 1330 4 vdd
port 513 nsew
rlabel metal1 s 13968 1039 13968 1039 4 vdd
port 513 nsew
rlabel metal1 s 12720 1829 12720 1829 4 vdd
port 513 nsew
rlabel metal1 s 12720 540 12720 540 4 vdd
port 513 nsew
rlabel metal1 s 14736 2120 14736 2120 4 vdd
port 513 nsew
rlabel metal1 s 12720 249 12720 249 4 vdd
port 513 nsew
rlabel metal1 s 12720 1330 12720 1330 4 vdd
port 513 nsew
rlabel metal1 s 12720 2120 12720 2120 4 vdd
port 513 nsew
rlabel metal1 s 13968 1829 13968 1829 4 vdd
port 513 nsew
rlabel metal1 s 13488 249 13488 249 4 vdd
port 513 nsew
rlabel metal1 s 14736 1829 14736 1829 4 vdd
port 513 nsew
rlabel metal1 s 14736 2910 14736 2910 4 vdd
port 513 nsew
rlabel metal1 s 14736 2619 14736 2619 4 vdd
port 513 nsew
rlabel metal1 s 13488 2120 13488 2120 4 vdd
port 513 nsew
rlabel metal1 s 18480 4490 18480 4490 4 vdd
port 513 nsew
rlabel metal1 s 19728 4989 19728 4989 4 vdd
port 513 nsew
rlabel metal1 s 17712 3409 17712 3409 4 vdd
port 513 nsew
rlabel metal1 s 18480 5280 18480 5280 4 vdd
port 513 nsew
rlabel metal1 s 18480 5779 18480 5779 4 vdd
port 513 nsew
rlabel metal1 s 19728 3700 19728 3700 4 vdd
port 513 nsew
rlabel metal1 s 18960 5779 18960 5779 4 vdd
port 513 nsew
rlabel metal1 s 19728 5779 19728 5779 4 vdd
port 513 nsew
rlabel metal1 s 19728 4490 19728 4490 4 vdd
port 513 nsew
rlabel metal1 s 19728 5280 19728 5280 4 vdd
port 513 nsew
rlabel metal1 s 18480 3409 18480 3409 4 vdd
port 513 nsew
rlabel metal1 s 18960 3700 18960 3700 4 vdd
port 513 nsew
rlabel metal1 s 18480 3700 18480 3700 4 vdd
port 513 nsew
rlabel metal1 s 17712 4490 17712 4490 4 vdd
port 513 nsew
rlabel metal1 s 19728 4199 19728 4199 4 vdd
port 513 nsew
rlabel metal1 s 17712 3700 17712 3700 4 vdd
port 513 nsew
rlabel metal1 s 18960 3409 18960 3409 4 vdd
port 513 nsew
rlabel metal1 s 18960 6070 18960 6070 4 vdd
port 513 nsew
rlabel metal1 s 18480 4989 18480 4989 4 vdd
port 513 nsew
rlabel metal1 s 18480 6070 18480 6070 4 vdd
port 513 nsew
rlabel metal1 s 19728 6070 19728 6070 4 vdd
port 513 nsew
rlabel metal1 s 18480 4199 18480 4199 4 vdd
port 513 nsew
rlabel metal1 s 18960 4199 18960 4199 4 vdd
port 513 nsew
rlabel metal1 s 18960 4989 18960 4989 4 vdd
port 513 nsew
rlabel metal1 s 17712 5779 17712 5779 4 vdd
port 513 nsew
rlabel metal1 s 17712 4989 17712 4989 4 vdd
port 513 nsew
rlabel metal1 s 18960 4490 18960 4490 4 vdd
port 513 nsew
rlabel metal1 s 17712 4199 17712 4199 4 vdd
port 513 nsew
rlabel metal1 s 17712 5280 17712 5280 4 vdd
port 513 nsew
rlabel metal1 s 18960 5280 18960 5280 4 vdd
port 513 nsew
rlabel metal1 s 17712 6070 17712 6070 4 vdd
port 513 nsew
rlabel metal1 s 19728 3409 19728 3409 4 vdd
port 513 nsew
rlabel metal1 s 15984 3700 15984 3700 4 vdd
port 513 nsew
rlabel metal1 s 15984 5280 15984 5280 4 vdd
port 513 nsew
rlabel metal1 s 17232 3409 17232 3409 4 vdd
port 513 nsew
rlabel metal1 s 16464 5280 16464 5280 4 vdd
port 513 nsew
rlabel metal1 s 15984 5779 15984 5779 4 vdd
port 513 nsew
rlabel metal1 s 15216 3700 15216 3700 4 vdd
port 513 nsew
rlabel metal1 s 15216 5280 15216 5280 4 vdd
port 513 nsew
rlabel metal1 s 16464 6070 16464 6070 4 vdd
port 513 nsew
rlabel metal1 s 16464 3700 16464 3700 4 vdd
port 513 nsew
rlabel metal1 s 15216 6070 15216 6070 4 vdd
port 513 nsew
rlabel metal1 s 15984 6070 15984 6070 4 vdd
port 513 nsew
rlabel metal1 s 16464 5779 16464 5779 4 vdd
port 513 nsew
rlabel metal1 s 15216 3409 15216 3409 4 vdd
port 513 nsew
rlabel metal1 s 16464 3409 16464 3409 4 vdd
port 513 nsew
rlabel metal1 s 15984 4989 15984 4989 4 vdd
port 513 nsew
rlabel metal1 s 17232 5280 17232 5280 4 vdd
port 513 nsew
rlabel metal1 s 17232 4490 17232 4490 4 vdd
port 513 nsew
rlabel metal1 s 15216 5779 15216 5779 4 vdd
port 513 nsew
rlabel metal1 s 16464 4989 16464 4989 4 vdd
port 513 nsew
rlabel metal1 s 15216 4199 15216 4199 4 vdd
port 513 nsew
rlabel metal1 s 17232 4989 17232 4989 4 vdd
port 513 nsew
rlabel metal1 s 17232 4199 17232 4199 4 vdd
port 513 nsew
rlabel metal1 s 16464 4490 16464 4490 4 vdd
port 513 nsew
rlabel metal1 s 17232 6070 17232 6070 4 vdd
port 513 nsew
rlabel metal1 s 15984 4199 15984 4199 4 vdd
port 513 nsew
rlabel metal1 s 16464 4199 16464 4199 4 vdd
port 513 nsew
rlabel metal1 s 17232 5779 17232 5779 4 vdd
port 513 nsew
rlabel metal1 s 15216 4989 15216 4989 4 vdd
port 513 nsew
rlabel metal1 s 15216 4490 15216 4490 4 vdd
port 513 nsew
rlabel metal1 s 17232 3700 17232 3700 4 vdd
port 513 nsew
rlabel metal1 s 15984 4490 15984 4490 4 vdd
port 513 nsew
rlabel metal1 s 15984 3409 15984 3409 4 vdd
port 513 nsew
rlabel metal1 s 16464 2910 16464 2910 4 vdd
port 513 nsew
rlabel metal1 s 15216 1330 15216 1330 4 vdd
port 513 nsew
rlabel metal1 s 15984 2619 15984 2619 4 vdd
port 513 nsew
rlabel metal1 s 15216 540 15216 540 4 vdd
port 513 nsew
rlabel metal1 s 17232 2619 17232 2619 4 vdd
port 513 nsew
rlabel metal1 s 17232 1039 17232 1039 4 vdd
port 513 nsew
rlabel metal1 s 15984 1039 15984 1039 4 vdd
port 513 nsew
rlabel metal1 s 15984 2120 15984 2120 4 vdd
port 513 nsew
rlabel metal1 s 15216 1829 15216 1829 4 vdd
port 513 nsew
rlabel metal1 s 17232 2910 17232 2910 4 vdd
port 513 nsew
rlabel metal1 s 16464 249 16464 249 4 vdd
port 513 nsew
rlabel metal1 s 16464 1039 16464 1039 4 vdd
port 513 nsew
rlabel metal1 s 15216 2619 15216 2619 4 vdd
port 513 nsew
rlabel metal1 s 15984 249 15984 249 4 vdd
port 513 nsew
rlabel metal1 s 15984 1330 15984 1330 4 vdd
port 513 nsew
rlabel metal1 s 15984 1829 15984 1829 4 vdd
port 513 nsew
rlabel metal1 s 15984 2910 15984 2910 4 vdd
port 513 nsew
rlabel metal1 s 15216 2910 15216 2910 4 vdd
port 513 nsew
rlabel metal1 s 17232 1829 17232 1829 4 vdd
port 513 nsew
rlabel metal1 s 16464 2619 16464 2619 4 vdd
port 513 nsew
rlabel metal1 s 16464 1330 16464 1330 4 vdd
port 513 nsew
rlabel metal1 s 17232 540 17232 540 4 vdd
port 513 nsew
rlabel metal1 s 15216 249 15216 249 4 vdd
port 513 nsew
rlabel metal1 s 15216 2120 15216 2120 4 vdd
port 513 nsew
rlabel metal1 s 16464 540 16464 540 4 vdd
port 513 nsew
rlabel metal1 s 16464 2120 16464 2120 4 vdd
port 513 nsew
rlabel metal1 s 15216 1039 15216 1039 4 vdd
port 513 nsew
rlabel metal1 s 16464 1829 16464 1829 4 vdd
port 513 nsew
rlabel metal1 s 17232 1330 17232 1330 4 vdd
port 513 nsew
rlabel metal1 s 17232 2120 17232 2120 4 vdd
port 513 nsew
rlabel metal1 s 17232 249 17232 249 4 vdd
port 513 nsew
rlabel metal1 s 15984 540 15984 540 4 vdd
port 513 nsew
rlabel metal1 s 19728 2619 19728 2619 4 vdd
port 513 nsew
rlabel metal1 s 19728 2120 19728 2120 4 vdd
port 513 nsew
rlabel metal1 s 18960 249 18960 249 4 vdd
port 513 nsew
rlabel metal1 s 18960 1039 18960 1039 4 vdd
port 513 nsew
rlabel metal1 s 17712 2120 17712 2120 4 vdd
port 513 nsew
rlabel metal1 s 19728 1039 19728 1039 4 vdd
port 513 nsew
rlabel metal1 s 18960 2619 18960 2619 4 vdd
port 513 nsew
rlabel metal1 s 18960 2120 18960 2120 4 vdd
port 513 nsew
rlabel metal1 s 17712 1039 17712 1039 4 vdd
port 513 nsew
rlabel metal1 s 17712 2910 17712 2910 4 vdd
port 513 nsew
rlabel metal1 s 17712 249 17712 249 4 vdd
port 513 nsew
rlabel metal1 s 18480 249 18480 249 4 vdd
port 513 nsew
rlabel metal1 s 18480 2910 18480 2910 4 vdd
port 513 nsew
rlabel metal1 s 18960 2910 18960 2910 4 vdd
port 513 nsew
rlabel metal1 s 18960 1330 18960 1330 4 vdd
port 513 nsew
rlabel metal1 s 17712 540 17712 540 4 vdd
port 513 nsew
rlabel metal1 s 18480 2619 18480 2619 4 vdd
port 513 nsew
rlabel metal1 s 19728 1330 19728 1330 4 vdd
port 513 nsew
rlabel metal1 s 17712 1829 17712 1829 4 vdd
port 513 nsew
rlabel metal1 s 19728 540 19728 540 4 vdd
port 513 nsew
rlabel metal1 s 18480 2120 18480 2120 4 vdd
port 513 nsew
rlabel metal1 s 19728 249 19728 249 4 vdd
port 513 nsew
rlabel metal1 s 18480 1829 18480 1829 4 vdd
port 513 nsew
rlabel metal1 s 19728 1829 19728 1829 4 vdd
port 513 nsew
rlabel metal1 s 17712 1330 17712 1330 4 vdd
port 513 nsew
rlabel metal1 s 19728 2910 19728 2910 4 vdd
port 513 nsew
rlabel metal1 s 18480 1330 18480 1330 4 vdd
port 513 nsew
rlabel metal1 s 18960 540 18960 540 4 vdd
port 513 nsew
rlabel metal1 s 17712 2619 17712 2619 4 vdd
port 513 nsew
rlabel metal1 s 18480 540 18480 540 4 vdd
port 513 nsew
rlabel metal1 s 18960 1829 18960 1829 4 vdd
port 513 nsew
rlabel metal1 s 18480 1039 18480 1039 4 vdd
port 513 nsew
rlabel metal1 s 39552 25280 39552 25280 4 br1_63
port 256 nsew
rlabel metal1 s 38928 25030 38928 25030 4 vdd
port 513 nsew
rlabel metal1 s 38448 23949 38448 23949 4 vdd
port 513 nsew
rlabel metal1 s 39696 22369 39696 22369 4 vdd
port 513 nsew
rlabel metal1 s 38928 23949 38928 23949 4 vdd
port 513 nsew
rlabel metal1 s 38928 22369 38928 22369 4 vdd
port 513 nsew
rlabel metal1 s 37680 23159 37680 23159 4 vdd
port 513 nsew
rlabel metal1 s 37680 24739 37680 24739 4 vdd
port 513 nsew
rlabel metal1 s 38304 25280 38304 25280 4 br1_61
port 248 nsew
rlabel metal1 s 37680 23949 37680 23949 4 vdd
port 513 nsew
rlabel metal1 s 38448 24739 38448 24739 4 vdd
port 513 nsew
rlabel metal1 s 38448 24240 38448 24240 4 vdd
port 513 nsew
rlabel metal1 s 39696 23949 39696 23949 4 vdd
port 513 nsew
rlabel metal1 s 38592 25280 38592 25280 4 bl0_61
port 245 nsew
rlabel metal1 s 38928 24240 38928 24240 4 vdd
port 513 nsew
rlabel metal1 s 38928 23450 38928 23450 4 vdd
port 513 nsew
rlabel metal1 s 39696 25030 39696 25030 4 vdd
port 513 nsew
rlabel metal1 s 39696 24739 39696 24739 4 vdd
port 513 nsew
rlabel metal1 s 37680 23450 37680 23450 4 vdd
port 513 nsew
rlabel metal1 s 39696 23159 39696 23159 4 vdd
port 513 nsew
rlabel metal1 s 37680 22660 37680 22660 4 vdd
port 513 nsew
rlabel metal1 s 38448 23159 38448 23159 4 vdd
port 513 nsew
rlabel metal1 s 39840 25280 39840 25280 4 bl0_63
port 253 nsew
rlabel metal1 s 37680 25030 37680 25030 4 vdd
port 513 nsew
rlabel metal1 s 38448 22660 38448 22660 4 vdd
port 513 nsew
rlabel metal1 s 39696 23450 39696 23450 4 vdd
port 513 nsew
rlabel metal1 s 38448 22369 38448 22369 4 vdd
port 513 nsew
rlabel metal1 s 37680 22369 37680 22369 4 vdd
port 513 nsew
rlabel metal1 s 38448 25030 38448 25030 4 vdd
port 513 nsew
rlabel metal1 s 39768 25280 39768 25280 4 br0_63
port 254 nsew
rlabel metal1 s 38928 22660 38928 22660 4 vdd
port 513 nsew
rlabel metal1 s 37680 24240 37680 24240 4 vdd
port 513 nsew
rlabel metal1 s 37824 25280 37824 25280 4 br1_60
port 244 nsew
rlabel metal1 s 39696 22660 39696 22660 4 vdd
port 513 nsew
rlabel metal1 s 39696 24240 39696 24240 4 vdd
port 513 nsew
rlabel metal1 s 38928 24739 38928 24739 4 vdd
port 513 nsew
rlabel metal1 s 38784 25280 38784 25280 4 bl0_62
port 249 nsew
rlabel metal1 s 38928 23159 38928 23159 4 vdd
port 513 nsew
rlabel metal1 s 38448 23450 38448 23450 4 vdd
port 513 nsew
rlabel metal1 s 39072 25280 39072 25280 4 br1_62
port 252 nsew
rlabel metal1 s 39624 25280 39624 25280 4 bl1_63
port 255 nsew
rlabel metal1 s 37752 25280 37752 25280 4 bl1_60
port 243 nsew
rlabel metal1 s 37536 25280 37536 25280 4 bl0_60
port 241 nsew
rlabel metal1 s 39000 25280 39000 25280 4 bl1_62
port 251 nsew
rlabel metal1 s 38376 25280 38376 25280 4 bl1_61
port 247 nsew
rlabel metal1 s 37608 25280 37608 25280 4 br0_60
port 242 nsew
rlabel metal1 s 38856 25280 38856 25280 4 br0_62
port 250 nsew
rlabel metal1 s 38520 25280 38520 25280 4 br0_61
port 246 nsew
rlabel metal1 s 37200 23159 37200 23159 4 vdd
port 513 nsew
rlabel metal1 s 36432 23450 36432 23450 4 vdd
port 513 nsew
rlabel metal1 s 35184 22369 35184 22369 4 vdd
port 513 nsew
rlabel metal1 s 35952 23949 35952 23949 4 vdd
port 513 nsew
rlabel metal1 s 35952 24739 35952 24739 4 vdd
port 513 nsew
rlabel metal1 s 35952 23159 35952 23159 4 vdd
port 513 nsew
rlabel metal1 s 37056 25280 37056 25280 4 br1_59
port 240 nsew
rlabel metal1 s 36432 22660 36432 22660 4 vdd
port 513 nsew
rlabel metal1 s 36360 25280 36360 25280 4 br0_58
port 234 nsew
rlabel metal1 s 36432 24240 36432 24240 4 vdd
port 513 nsew
rlabel metal1 s 36432 24739 36432 24739 4 vdd
port 513 nsew
rlabel metal1 s 35184 24240 35184 24240 4 vdd
port 513 nsew
rlabel metal1 s 35184 23949 35184 23949 4 vdd
port 513 nsew
rlabel metal1 s 37200 24739 37200 24739 4 vdd
port 513 nsew
rlabel metal1 s 35184 25030 35184 25030 4 vdd
port 513 nsew
rlabel metal1 s 36432 23159 36432 23159 4 vdd
port 513 nsew
rlabel metal1 s 35184 24739 35184 24739 4 vdd
port 513 nsew
rlabel metal1 s 37200 23949 37200 23949 4 vdd
port 513 nsew
rlabel metal1 s 35952 22660 35952 22660 4 vdd
port 513 nsew
rlabel metal1 s 37200 22660 37200 22660 4 vdd
port 513 nsew
rlabel metal1 s 37344 25280 37344 25280 4 bl0_59
port 237 nsew
rlabel metal1 s 35952 25030 35952 25030 4 vdd
port 513 nsew
rlabel metal1 s 36432 25030 36432 25030 4 vdd
port 513 nsew
rlabel metal1 s 37200 22369 37200 22369 4 vdd
port 513 nsew
rlabel metal1 s 35952 24240 35952 24240 4 vdd
port 513 nsew
rlabel metal1 s 36288 25280 36288 25280 4 bl0_58
port 233 nsew
rlabel metal1 s 36432 22369 36432 22369 4 vdd
port 513 nsew
rlabel metal1 s 36504 25280 36504 25280 4 bl1_58
port 235 nsew
rlabel metal1 s 36096 25280 36096 25280 4 bl0_57
port 229 nsew
rlabel metal1 s 37200 23450 37200 23450 4 vdd
port 513 nsew
rlabel metal1 s 35040 25280 35040 25280 4 bl0_56
port 225 nsew
rlabel metal1 s 35184 23450 35184 23450 4 vdd
port 513 nsew
rlabel metal1 s 35952 22369 35952 22369 4 vdd
port 513 nsew
rlabel metal1 s 35256 25280 35256 25280 4 bl1_56
port 227 nsew
rlabel metal1 s 35328 25280 35328 25280 4 br1_56
port 228 nsew
rlabel metal1 s 37200 24240 37200 24240 4 vdd
port 513 nsew
rlabel metal1 s 36024 25280 36024 25280 4 br0_57
port 230 nsew
rlabel metal1 s 35184 23159 35184 23159 4 vdd
port 513 nsew
rlabel metal1 s 36432 23949 36432 23949 4 vdd
port 513 nsew
rlabel metal1 s 35952 23450 35952 23450 4 vdd
port 513 nsew
rlabel metal1 s 37200 25030 37200 25030 4 vdd
port 513 nsew
rlabel metal1 s 35880 25280 35880 25280 4 bl1_57
port 231 nsew
rlabel metal1 s 35112 25280 35112 25280 4 br0_56
port 226 nsew
rlabel metal1 s 37128 25280 37128 25280 4 bl1_59
port 239 nsew
rlabel metal1 s 36576 25280 36576 25280 4 br1_58
port 236 nsew
rlabel metal1 s 35184 22660 35184 22660 4 vdd
port 513 nsew
rlabel metal1 s 35808 25280 35808 25280 4 br1_57
port 232 nsew
rlabel metal1 s 37272 25280 37272 25280 4 br0_59
port 238 nsew
rlabel metal1 s 35952 21579 35952 21579 4 vdd
port 513 nsew
rlabel metal1 s 35184 21870 35184 21870 4 vdd
port 513 nsew
rlabel metal1 s 36432 20789 36432 20789 4 vdd
port 513 nsew
rlabel metal1 s 36432 20290 36432 20290 4 vdd
port 513 nsew
rlabel metal1 s 35184 19999 35184 19999 4 vdd
port 513 nsew
rlabel metal1 s 37200 19999 37200 19999 4 vdd
port 513 nsew
rlabel metal1 s 36432 19500 36432 19500 4 vdd
port 513 nsew
rlabel metal1 s 37200 20290 37200 20290 4 vdd
port 513 nsew
rlabel metal1 s 37200 21870 37200 21870 4 vdd
port 513 nsew
rlabel metal1 s 35184 19209 35184 19209 4 vdd
port 513 nsew
rlabel metal1 s 35952 21870 35952 21870 4 vdd
port 513 nsew
rlabel metal1 s 35952 20789 35952 20789 4 vdd
port 513 nsew
rlabel metal1 s 35952 19209 35952 19209 4 vdd
port 513 nsew
rlabel metal1 s 35184 19500 35184 19500 4 vdd
port 513 nsew
rlabel metal1 s 37200 19209 37200 19209 4 vdd
port 513 nsew
rlabel metal1 s 35952 19999 35952 19999 4 vdd
port 513 nsew
rlabel metal1 s 37200 21579 37200 21579 4 vdd
port 513 nsew
rlabel metal1 s 36432 21870 36432 21870 4 vdd
port 513 nsew
rlabel metal1 s 36432 19209 36432 19209 4 vdd
port 513 nsew
rlabel metal1 s 35952 20290 35952 20290 4 vdd
port 513 nsew
rlabel metal1 s 35952 19500 35952 19500 4 vdd
port 513 nsew
rlabel metal1 s 36432 19999 36432 19999 4 vdd
port 513 nsew
rlabel metal1 s 35184 21080 35184 21080 4 vdd
port 513 nsew
rlabel metal1 s 36432 21579 36432 21579 4 vdd
port 513 nsew
rlabel metal1 s 37200 20789 37200 20789 4 vdd
port 513 nsew
rlabel metal1 s 35952 21080 35952 21080 4 vdd
port 513 nsew
rlabel metal1 s 35184 20789 35184 20789 4 vdd
port 513 nsew
rlabel metal1 s 37200 21080 37200 21080 4 vdd
port 513 nsew
rlabel metal1 s 35184 21579 35184 21579 4 vdd
port 513 nsew
rlabel metal1 s 35184 20290 35184 20290 4 vdd
port 513 nsew
rlabel metal1 s 36432 21080 36432 21080 4 vdd
port 513 nsew
rlabel metal1 s 37200 19500 37200 19500 4 vdd
port 513 nsew
rlabel metal1 s 37680 19209 37680 19209 4 vdd
port 513 nsew
rlabel metal1 s 38928 21870 38928 21870 4 vdd
port 513 nsew
rlabel metal1 s 38448 21579 38448 21579 4 vdd
port 513 nsew
rlabel metal1 s 37680 20290 37680 20290 4 vdd
port 513 nsew
rlabel metal1 s 39696 21579 39696 21579 4 vdd
port 513 nsew
rlabel metal1 s 38448 19500 38448 19500 4 vdd
port 513 nsew
rlabel metal1 s 38448 20290 38448 20290 4 vdd
port 513 nsew
rlabel metal1 s 38448 21080 38448 21080 4 vdd
port 513 nsew
rlabel metal1 s 38928 20789 38928 20789 4 vdd
port 513 nsew
rlabel metal1 s 37680 21870 37680 21870 4 vdd
port 513 nsew
rlabel metal1 s 38448 19999 38448 19999 4 vdd
port 513 nsew
rlabel metal1 s 38928 19999 38928 19999 4 vdd
port 513 nsew
rlabel metal1 s 39696 19999 39696 19999 4 vdd
port 513 nsew
rlabel metal1 s 37680 21579 37680 21579 4 vdd
port 513 nsew
rlabel metal1 s 39696 21870 39696 21870 4 vdd
port 513 nsew
rlabel metal1 s 39696 20789 39696 20789 4 vdd
port 513 nsew
rlabel metal1 s 38928 21080 38928 21080 4 vdd
port 513 nsew
rlabel metal1 s 39696 19209 39696 19209 4 vdd
port 513 nsew
rlabel metal1 s 38928 19209 38928 19209 4 vdd
port 513 nsew
rlabel metal1 s 37680 21080 37680 21080 4 vdd
port 513 nsew
rlabel metal1 s 38448 20789 38448 20789 4 vdd
port 513 nsew
rlabel metal1 s 38928 20290 38928 20290 4 vdd
port 513 nsew
rlabel metal1 s 39696 20290 39696 20290 4 vdd
port 513 nsew
rlabel metal1 s 37680 20789 37680 20789 4 vdd
port 513 nsew
rlabel metal1 s 38448 21870 38448 21870 4 vdd
port 513 nsew
rlabel metal1 s 38448 19209 38448 19209 4 vdd
port 513 nsew
rlabel metal1 s 39696 21080 39696 21080 4 vdd
port 513 nsew
rlabel metal1 s 38928 21579 38928 21579 4 vdd
port 513 nsew
rlabel metal1 s 39696 19500 39696 19500 4 vdd
port 513 nsew
rlabel metal1 s 37680 19500 37680 19500 4 vdd
port 513 nsew
rlabel metal1 s 37680 19999 37680 19999 4 vdd
port 513 nsew
rlabel metal1 s 38928 19500 38928 19500 4 vdd
port 513 nsew
rlabel metal1 s 33936 24739 33936 24739 4 vdd
port 513 nsew
rlabel metal1 s 32688 24240 32688 24240 4 vdd
port 513 nsew
rlabel metal1 s 33864 25280 33864 25280 4 br0_54
port 218 nsew
rlabel metal1 s 33936 24240 33936 24240 4 vdd
port 513 nsew
rlabel metal1 s 32688 25030 32688 25030 4 vdd
port 513 nsew
rlabel metal1 s 34704 25030 34704 25030 4 vdd
port 513 nsew
rlabel metal1 s 32688 23949 32688 23949 4 vdd
port 513 nsew
rlabel metal1 s 33456 25030 33456 25030 4 vdd
port 513 nsew
rlabel metal1 s 34704 23949 34704 23949 4 vdd
port 513 nsew
rlabel metal1 s 32688 22369 32688 22369 4 vdd
port 513 nsew
rlabel metal1 s 33936 23159 33936 23159 4 vdd
port 513 nsew
rlabel metal1 s 33456 23949 33456 23949 4 vdd
port 513 nsew
rlabel metal1 s 34704 23450 34704 23450 4 vdd
port 513 nsew
rlabel metal1 s 32688 23450 32688 23450 4 vdd
port 513 nsew
rlabel metal1 s 34704 23159 34704 23159 4 vdd
port 513 nsew
rlabel metal1 s 33456 23159 33456 23159 4 vdd
port 513 nsew
rlabel metal1 s 34848 25280 34848 25280 4 bl0_55
port 221 nsew
rlabel metal1 s 32832 25280 32832 25280 4 br1_52
port 212 nsew
rlabel metal1 s 34704 24240 34704 24240 4 vdd
port 513 nsew
rlabel metal1 s 33936 25030 33936 25030 4 vdd
port 513 nsew
rlabel metal1 s 33936 23450 33936 23450 4 vdd
port 513 nsew
rlabel metal1 s 34776 25280 34776 25280 4 br0_55
port 222 nsew
rlabel metal1 s 34560 25280 34560 25280 4 br1_55
port 224 nsew
rlabel metal1 s 32688 23159 32688 23159 4 vdd
port 513 nsew
rlabel metal1 s 34632 25280 34632 25280 4 bl1_55
port 223 nsew
rlabel metal1 s 33456 24240 33456 24240 4 vdd
port 513 nsew
rlabel metal1 s 33936 22369 33936 22369 4 vdd
port 513 nsew
rlabel metal1 s 34704 22660 34704 22660 4 vdd
port 513 nsew
rlabel metal1 s 33936 23949 33936 23949 4 vdd
port 513 nsew
rlabel metal1 s 32688 24739 32688 24739 4 vdd
port 513 nsew
rlabel metal1 s 33456 22660 33456 22660 4 vdd
port 513 nsew
rlabel metal1 s 33456 24739 33456 24739 4 vdd
port 513 nsew
rlabel metal1 s 34704 22369 34704 22369 4 vdd
port 513 nsew
rlabel metal1 s 32544 25280 32544 25280 4 bl0_52
port 209 nsew
rlabel metal1 s 32688 22660 32688 22660 4 vdd
port 513 nsew
rlabel metal1 s 33312 25280 33312 25280 4 br1_53
port 216 nsew
rlabel metal1 s 33456 23450 33456 23450 4 vdd
port 513 nsew
rlabel metal1 s 33792 25280 33792 25280 4 bl0_54
port 217 nsew
rlabel metal1 s 34080 25280 34080 25280 4 br1_54
port 220 nsew
rlabel metal1 s 32760 25280 32760 25280 4 bl1_52
port 211 nsew
rlabel metal1 s 33528 25280 33528 25280 4 br0_53
port 214 nsew
rlabel metal1 s 33936 22660 33936 22660 4 vdd
port 513 nsew
rlabel metal1 s 32616 25280 32616 25280 4 br0_52
port 210 nsew
rlabel metal1 s 33456 22369 33456 22369 4 vdd
port 513 nsew
rlabel metal1 s 34704 24739 34704 24739 4 vdd
port 513 nsew
rlabel metal1 s 33384 25280 33384 25280 4 bl1_53
port 215 nsew
rlabel metal1 s 33600 25280 33600 25280 4 bl0_53
port 213 nsew
rlabel metal1 s 34008 25280 34008 25280 4 bl1_54
port 219 nsew
rlabel metal1 s 30192 23949 30192 23949 4 vdd
port 513 nsew
rlabel metal1 s 30192 22369 30192 22369 4 vdd
port 513 nsew
rlabel metal1 s 30192 24240 30192 24240 4 vdd
port 513 nsew
rlabel metal1 s 30192 22660 30192 22660 4 vdd
port 513 nsew
rlabel metal1 s 31368 25280 31368 25280 4 br0_50
port 202 nsew
rlabel metal1 s 32208 23949 32208 23949 4 vdd
port 513 nsew
rlabel metal1 s 30192 24739 30192 24739 4 vdd
port 513 nsew
rlabel metal1 s 30960 25030 30960 25030 4 vdd
port 513 nsew
rlabel metal1 s 30192 25030 30192 25030 4 vdd
port 513 nsew
rlabel metal1 s 32208 22369 32208 22369 4 vdd
port 513 nsew
rlabel metal1 s 31032 25280 31032 25280 4 br0_49
port 198 nsew
rlabel metal1 s 30192 23159 30192 23159 4 vdd
port 513 nsew
rlabel metal1 s 31440 25030 31440 25030 4 vdd
port 513 nsew
rlabel metal1 s 30192 23450 30192 23450 4 vdd
port 513 nsew
rlabel metal1 s 31104 25280 31104 25280 4 bl0_49
port 197 nsew
rlabel metal1 s 31440 23450 31440 23450 4 vdd
port 513 nsew
rlabel metal1 s 31440 22660 31440 22660 4 vdd
port 513 nsew
rlabel metal1 s 30816 25280 30816 25280 4 br1_49
port 200 nsew
rlabel metal1 s 32208 24739 32208 24739 4 vdd
port 513 nsew
rlabel metal1 s 30960 24739 30960 24739 4 vdd
port 513 nsew
rlabel metal1 s 31440 24240 31440 24240 4 vdd
port 513 nsew
rlabel metal1 s 30048 25280 30048 25280 4 bl0_48
port 193 nsew
rlabel metal1 s 32136 25280 32136 25280 4 bl1_51
port 207 nsew
rlabel metal1 s 32208 23450 32208 23450 4 vdd
port 513 nsew
rlabel metal1 s 30960 22369 30960 22369 4 vdd
port 513 nsew
rlabel metal1 s 32208 22660 32208 22660 4 vdd
port 513 nsew
rlabel metal1 s 32208 23159 32208 23159 4 vdd
port 513 nsew
rlabel metal1 s 32280 25280 32280 25280 4 br0_51
port 206 nsew
rlabel metal1 s 31440 24739 31440 24739 4 vdd
port 513 nsew
rlabel metal1 s 31440 23949 31440 23949 4 vdd
port 513 nsew
rlabel metal1 s 30888 25280 30888 25280 4 bl1_49
port 199 nsew
rlabel metal1 s 30120 25280 30120 25280 4 br0_48
port 194 nsew
rlabel metal1 s 30960 24240 30960 24240 4 vdd
port 513 nsew
rlabel metal1 s 31584 25280 31584 25280 4 br1_50
port 204 nsew
rlabel metal1 s 31296 25280 31296 25280 4 bl0_50
port 201 nsew
rlabel metal1 s 30960 23949 30960 23949 4 vdd
port 513 nsew
rlabel metal1 s 31440 23159 31440 23159 4 vdd
port 513 nsew
rlabel metal1 s 31440 22369 31440 22369 4 vdd
port 513 nsew
rlabel metal1 s 30960 22660 30960 22660 4 vdd
port 513 nsew
rlabel metal1 s 30960 23159 30960 23159 4 vdd
port 513 nsew
rlabel metal1 s 32352 25280 32352 25280 4 bl0_51
port 205 nsew
rlabel metal1 s 31512 25280 31512 25280 4 bl1_50
port 203 nsew
rlabel metal1 s 32208 25030 32208 25030 4 vdd
port 513 nsew
rlabel metal1 s 30264 25280 30264 25280 4 bl1_48
port 195 nsew
rlabel metal1 s 30960 23450 30960 23450 4 vdd
port 513 nsew
rlabel metal1 s 32208 24240 32208 24240 4 vdd
port 513 nsew
rlabel metal1 s 30336 25280 30336 25280 4 br1_48
port 196 nsew
rlabel metal1 s 32064 25280 32064 25280 4 br1_51
port 208 nsew
rlabel metal1 s 30960 21870 30960 21870 4 vdd
port 513 nsew
rlabel metal1 s 32208 20789 32208 20789 4 vdd
port 513 nsew
rlabel metal1 s 30192 19209 30192 19209 4 vdd
port 513 nsew
rlabel metal1 s 30192 19500 30192 19500 4 vdd
port 513 nsew
rlabel metal1 s 30192 21870 30192 21870 4 vdd
port 513 nsew
rlabel metal1 s 30960 19209 30960 19209 4 vdd
port 513 nsew
rlabel metal1 s 30192 20789 30192 20789 4 vdd
port 513 nsew
rlabel metal1 s 32208 19500 32208 19500 4 vdd
port 513 nsew
rlabel metal1 s 30960 21080 30960 21080 4 vdd
port 513 nsew
rlabel metal1 s 32208 21080 32208 21080 4 vdd
port 513 nsew
rlabel metal1 s 30192 21080 30192 21080 4 vdd
port 513 nsew
rlabel metal1 s 32208 21870 32208 21870 4 vdd
port 513 nsew
rlabel metal1 s 32208 19209 32208 19209 4 vdd
port 513 nsew
rlabel metal1 s 30960 19999 30960 19999 4 vdd
port 513 nsew
rlabel metal1 s 31440 19500 31440 19500 4 vdd
port 513 nsew
rlabel metal1 s 31440 20789 31440 20789 4 vdd
port 513 nsew
rlabel metal1 s 30960 19500 30960 19500 4 vdd
port 513 nsew
rlabel metal1 s 31440 21080 31440 21080 4 vdd
port 513 nsew
rlabel metal1 s 31440 21870 31440 21870 4 vdd
port 513 nsew
rlabel metal1 s 30960 20290 30960 20290 4 vdd
port 513 nsew
rlabel metal1 s 30960 21579 30960 21579 4 vdd
port 513 nsew
rlabel metal1 s 30192 21579 30192 21579 4 vdd
port 513 nsew
rlabel metal1 s 32208 20290 32208 20290 4 vdd
port 513 nsew
rlabel metal1 s 30192 19999 30192 19999 4 vdd
port 513 nsew
rlabel metal1 s 31440 20290 31440 20290 4 vdd
port 513 nsew
rlabel metal1 s 30192 20290 30192 20290 4 vdd
port 513 nsew
rlabel metal1 s 30960 20789 30960 20789 4 vdd
port 513 nsew
rlabel metal1 s 32208 21579 32208 21579 4 vdd
port 513 nsew
rlabel metal1 s 32208 19999 32208 19999 4 vdd
port 513 nsew
rlabel metal1 s 31440 19999 31440 19999 4 vdd
port 513 nsew
rlabel metal1 s 31440 19209 31440 19209 4 vdd
port 513 nsew
rlabel metal1 s 31440 21579 31440 21579 4 vdd
port 513 nsew
rlabel metal1 s 34704 19500 34704 19500 4 vdd
port 513 nsew
rlabel metal1 s 34704 20789 34704 20789 4 vdd
port 513 nsew
rlabel metal1 s 32688 19999 32688 19999 4 vdd
port 513 nsew
rlabel metal1 s 33936 20290 33936 20290 4 vdd
port 513 nsew
rlabel metal1 s 34704 19209 34704 19209 4 vdd
port 513 nsew
rlabel metal1 s 33456 21080 33456 21080 4 vdd
port 513 nsew
rlabel metal1 s 34704 19999 34704 19999 4 vdd
port 513 nsew
rlabel metal1 s 32688 20789 32688 20789 4 vdd
port 513 nsew
rlabel metal1 s 34704 21080 34704 21080 4 vdd
port 513 nsew
rlabel metal1 s 33936 21579 33936 21579 4 vdd
port 513 nsew
rlabel metal1 s 32688 20290 32688 20290 4 vdd
port 513 nsew
rlabel metal1 s 32688 19500 32688 19500 4 vdd
port 513 nsew
rlabel metal1 s 33456 19500 33456 19500 4 vdd
port 513 nsew
rlabel metal1 s 33936 19209 33936 19209 4 vdd
port 513 nsew
rlabel metal1 s 33456 19999 33456 19999 4 vdd
port 513 nsew
rlabel metal1 s 33456 20290 33456 20290 4 vdd
port 513 nsew
rlabel metal1 s 33456 21579 33456 21579 4 vdd
port 513 nsew
rlabel metal1 s 33936 20789 33936 20789 4 vdd
port 513 nsew
rlabel metal1 s 33936 19500 33936 19500 4 vdd
port 513 nsew
rlabel metal1 s 33456 21870 33456 21870 4 vdd
port 513 nsew
rlabel metal1 s 34704 20290 34704 20290 4 vdd
port 513 nsew
rlabel metal1 s 34704 21579 34704 21579 4 vdd
port 513 nsew
rlabel metal1 s 33936 19999 33936 19999 4 vdd
port 513 nsew
rlabel metal1 s 33456 19209 33456 19209 4 vdd
port 513 nsew
rlabel metal1 s 32688 21870 32688 21870 4 vdd
port 513 nsew
rlabel metal1 s 32688 21080 32688 21080 4 vdd
port 513 nsew
rlabel metal1 s 33456 20789 33456 20789 4 vdd
port 513 nsew
rlabel metal1 s 33936 21080 33936 21080 4 vdd
port 513 nsew
rlabel metal1 s 32688 21579 32688 21579 4 vdd
port 513 nsew
rlabel metal1 s 34704 21870 34704 21870 4 vdd
port 513 nsew
rlabel metal1 s 33936 21870 33936 21870 4 vdd
port 513 nsew
rlabel metal1 s 32688 19209 32688 19209 4 vdd
port 513 nsew
rlabel metal1 s 33936 18710 33936 18710 4 vdd
port 513 nsew
rlabel metal1 s 32688 17130 32688 17130 4 vdd
port 513 nsew
rlabel metal1 s 33936 18419 33936 18419 4 vdd
port 513 nsew
rlabel metal1 s 33936 16340 33936 16340 4 vdd
port 513 nsew
rlabel metal1 s 33456 16049 33456 16049 4 vdd
port 513 nsew
rlabel metal1 s 33936 16839 33936 16839 4 vdd
port 513 nsew
rlabel metal1 s 33456 16839 33456 16839 4 vdd
port 513 nsew
rlabel metal1 s 32688 18419 32688 18419 4 vdd
port 513 nsew
rlabel metal1 s 34704 16839 34704 16839 4 vdd
port 513 nsew
rlabel metal1 s 33456 16340 33456 16340 4 vdd
port 513 nsew
rlabel metal1 s 33456 18419 33456 18419 4 vdd
port 513 nsew
rlabel metal1 s 33456 17130 33456 17130 4 vdd
port 513 nsew
rlabel metal1 s 32688 16049 32688 16049 4 vdd
port 513 nsew
rlabel metal1 s 32688 16839 32688 16839 4 vdd
port 513 nsew
rlabel metal1 s 32688 16340 32688 16340 4 vdd
port 513 nsew
rlabel metal1 s 34704 17920 34704 17920 4 vdd
port 513 nsew
rlabel metal1 s 33936 16049 33936 16049 4 vdd
port 513 nsew
rlabel metal1 s 32688 17629 32688 17629 4 vdd
port 513 nsew
rlabel metal1 s 33456 17629 33456 17629 4 vdd
port 513 nsew
rlabel metal1 s 34704 16340 34704 16340 4 vdd
port 513 nsew
rlabel metal1 s 33936 17920 33936 17920 4 vdd
port 513 nsew
rlabel metal1 s 33456 18710 33456 18710 4 vdd
port 513 nsew
rlabel metal1 s 34704 16049 34704 16049 4 vdd
port 513 nsew
rlabel metal1 s 34704 17629 34704 17629 4 vdd
port 513 nsew
rlabel metal1 s 33456 17920 33456 17920 4 vdd
port 513 nsew
rlabel metal1 s 34704 18419 34704 18419 4 vdd
port 513 nsew
rlabel metal1 s 34704 17130 34704 17130 4 vdd
port 513 nsew
rlabel metal1 s 33936 17629 33936 17629 4 vdd
port 513 nsew
rlabel metal1 s 32688 17920 32688 17920 4 vdd
port 513 nsew
rlabel metal1 s 33936 17130 33936 17130 4 vdd
port 513 nsew
rlabel metal1 s 34704 18710 34704 18710 4 vdd
port 513 nsew
rlabel metal1 s 32688 18710 32688 18710 4 vdd
port 513 nsew
rlabel metal1 s 30192 17920 30192 17920 4 vdd
port 513 nsew
rlabel metal1 s 31440 17920 31440 17920 4 vdd
port 513 nsew
rlabel metal1 s 32208 18419 32208 18419 4 vdd
port 513 nsew
rlabel metal1 s 32208 18710 32208 18710 4 vdd
port 513 nsew
rlabel metal1 s 31440 16049 31440 16049 4 vdd
port 513 nsew
rlabel metal1 s 32208 17130 32208 17130 4 vdd
port 513 nsew
rlabel metal1 s 31440 18710 31440 18710 4 vdd
port 513 nsew
rlabel metal1 s 31440 18419 31440 18419 4 vdd
port 513 nsew
rlabel metal1 s 30192 16340 30192 16340 4 vdd
port 513 nsew
rlabel metal1 s 30192 18710 30192 18710 4 vdd
port 513 nsew
rlabel metal1 s 32208 17920 32208 17920 4 vdd
port 513 nsew
rlabel metal1 s 32208 17629 32208 17629 4 vdd
port 513 nsew
rlabel metal1 s 30960 16839 30960 16839 4 vdd
port 513 nsew
rlabel metal1 s 30192 17629 30192 17629 4 vdd
port 513 nsew
rlabel metal1 s 30960 18710 30960 18710 4 vdd
port 513 nsew
rlabel metal1 s 30192 16839 30192 16839 4 vdd
port 513 nsew
rlabel metal1 s 30960 18419 30960 18419 4 vdd
port 513 nsew
rlabel metal1 s 30960 17130 30960 17130 4 vdd
port 513 nsew
rlabel metal1 s 31440 17130 31440 17130 4 vdd
port 513 nsew
rlabel metal1 s 32208 16049 32208 16049 4 vdd
port 513 nsew
rlabel metal1 s 31440 16340 31440 16340 4 vdd
port 513 nsew
rlabel metal1 s 30960 16049 30960 16049 4 vdd
port 513 nsew
rlabel metal1 s 30960 17920 30960 17920 4 vdd
port 513 nsew
rlabel metal1 s 32208 16839 32208 16839 4 vdd
port 513 nsew
rlabel metal1 s 32208 16340 32208 16340 4 vdd
port 513 nsew
rlabel metal1 s 31440 17629 31440 17629 4 vdd
port 513 nsew
rlabel metal1 s 30192 18419 30192 18419 4 vdd
port 513 nsew
rlabel metal1 s 30192 16049 30192 16049 4 vdd
port 513 nsew
rlabel metal1 s 30192 17130 30192 17130 4 vdd
port 513 nsew
rlabel metal1 s 30960 17629 30960 17629 4 vdd
port 513 nsew
rlabel metal1 s 31440 16839 31440 16839 4 vdd
port 513 nsew
rlabel metal1 s 30960 16340 30960 16340 4 vdd
port 513 nsew
rlabel metal1 s 30960 12889 30960 12889 4 vdd
port 513 nsew
rlabel metal1 s 30960 15259 30960 15259 4 vdd
port 513 nsew
rlabel metal1 s 32208 15550 32208 15550 4 vdd
port 513 nsew
rlabel metal1 s 30960 13679 30960 13679 4 vdd
port 513 nsew
rlabel metal1 s 31440 14469 31440 14469 4 vdd
port 513 nsew
rlabel metal1 s 32208 13180 32208 13180 4 vdd
port 513 nsew
rlabel metal1 s 30192 13679 30192 13679 4 vdd
port 513 nsew
rlabel metal1 s 30960 13180 30960 13180 4 vdd
port 513 nsew
rlabel metal1 s 32208 13970 32208 13970 4 vdd
port 513 nsew
rlabel metal1 s 30192 13180 30192 13180 4 vdd
port 513 nsew
rlabel metal1 s 30192 14760 30192 14760 4 vdd
port 513 nsew
rlabel metal1 s 30960 14760 30960 14760 4 vdd
port 513 nsew
rlabel metal1 s 31440 14760 31440 14760 4 vdd
port 513 nsew
rlabel metal1 s 30192 15259 30192 15259 4 vdd
port 513 nsew
rlabel metal1 s 30192 15550 30192 15550 4 vdd
port 513 nsew
rlabel metal1 s 30960 15550 30960 15550 4 vdd
port 513 nsew
rlabel metal1 s 32208 12889 32208 12889 4 vdd
port 513 nsew
rlabel metal1 s 32208 14469 32208 14469 4 vdd
port 513 nsew
rlabel metal1 s 31440 13180 31440 13180 4 vdd
port 513 nsew
rlabel metal1 s 31440 13970 31440 13970 4 vdd
port 513 nsew
rlabel metal1 s 31440 15550 31440 15550 4 vdd
port 513 nsew
rlabel metal1 s 30192 14469 30192 14469 4 vdd
port 513 nsew
rlabel metal1 s 31440 13679 31440 13679 4 vdd
port 513 nsew
rlabel metal1 s 32208 15259 32208 15259 4 vdd
port 513 nsew
rlabel metal1 s 31440 15259 31440 15259 4 vdd
port 513 nsew
rlabel metal1 s 32208 13679 32208 13679 4 vdd
port 513 nsew
rlabel metal1 s 30192 12889 30192 12889 4 vdd
port 513 nsew
rlabel metal1 s 32208 14760 32208 14760 4 vdd
port 513 nsew
rlabel metal1 s 30960 13970 30960 13970 4 vdd
port 513 nsew
rlabel metal1 s 31440 12889 31440 12889 4 vdd
port 513 nsew
rlabel metal1 s 30192 13970 30192 13970 4 vdd
port 513 nsew
rlabel metal1 s 30960 14469 30960 14469 4 vdd
port 513 nsew
rlabel metal1 s 33456 13180 33456 13180 4 vdd
port 513 nsew
rlabel metal1 s 33456 14760 33456 14760 4 vdd
port 513 nsew
rlabel metal1 s 32688 14760 32688 14760 4 vdd
port 513 nsew
rlabel metal1 s 32688 13679 32688 13679 4 vdd
port 513 nsew
rlabel metal1 s 33936 13180 33936 13180 4 vdd
port 513 nsew
rlabel metal1 s 34704 13970 34704 13970 4 vdd
port 513 nsew
rlabel metal1 s 32688 13180 32688 13180 4 vdd
port 513 nsew
rlabel metal1 s 33936 12889 33936 12889 4 vdd
port 513 nsew
rlabel metal1 s 34704 13180 34704 13180 4 vdd
port 513 nsew
rlabel metal1 s 33936 13679 33936 13679 4 vdd
port 513 nsew
rlabel metal1 s 33456 14469 33456 14469 4 vdd
port 513 nsew
rlabel metal1 s 34704 12889 34704 12889 4 vdd
port 513 nsew
rlabel metal1 s 34704 14760 34704 14760 4 vdd
port 513 nsew
rlabel metal1 s 33456 15259 33456 15259 4 vdd
port 513 nsew
rlabel metal1 s 33936 15550 33936 15550 4 vdd
port 513 nsew
rlabel metal1 s 33456 13679 33456 13679 4 vdd
port 513 nsew
rlabel metal1 s 33936 14760 33936 14760 4 vdd
port 513 nsew
rlabel metal1 s 32688 12889 32688 12889 4 vdd
port 513 nsew
rlabel metal1 s 33936 13970 33936 13970 4 vdd
port 513 nsew
rlabel metal1 s 33936 14469 33936 14469 4 vdd
port 513 nsew
rlabel metal1 s 34704 15550 34704 15550 4 vdd
port 513 nsew
rlabel metal1 s 32688 15259 32688 15259 4 vdd
port 513 nsew
rlabel metal1 s 33456 12889 33456 12889 4 vdd
port 513 nsew
rlabel metal1 s 34704 14469 34704 14469 4 vdd
port 513 nsew
rlabel metal1 s 34704 15259 34704 15259 4 vdd
port 513 nsew
rlabel metal1 s 33456 15550 33456 15550 4 vdd
port 513 nsew
rlabel metal1 s 33456 13970 33456 13970 4 vdd
port 513 nsew
rlabel metal1 s 32688 13970 32688 13970 4 vdd
port 513 nsew
rlabel metal1 s 33936 15259 33936 15259 4 vdd
port 513 nsew
rlabel metal1 s 32688 14469 32688 14469 4 vdd
port 513 nsew
rlabel metal1 s 32688 15550 32688 15550 4 vdd
port 513 nsew
rlabel metal1 s 34704 13679 34704 13679 4 vdd
port 513 nsew
rlabel metal1 s 39696 16340 39696 16340 4 vdd
port 513 nsew
rlabel metal1 s 39696 18419 39696 18419 4 vdd
port 513 nsew
rlabel metal1 s 38448 18710 38448 18710 4 vdd
port 513 nsew
rlabel metal1 s 38448 18419 38448 18419 4 vdd
port 513 nsew
rlabel metal1 s 39696 17130 39696 17130 4 vdd
port 513 nsew
rlabel metal1 s 38448 17629 38448 17629 4 vdd
port 513 nsew
rlabel metal1 s 39696 16839 39696 16839 4 vdd
port 513 nsew
rlabel metal1 s 38448 16049 38448 16049 4 vdd
port 513 nsew
rlabel metal1 s 39696 16049 39696 16049 4 vdd
port 513 nsew
rlabel metal1 s 39696 17629 39696 17629 4 vdd
port 513 nsew
rlabel metal1 s 37680 18419 37680 18419 4 vdd
port 513 nsew
rlabel metal1 s 37680 17920 37680 17920 4 vdd
port 513 nsew
rlabel metal1 s 37680 16340 37680 16340 4 vdd
port 513 nsew
rlabel metal1 s 38928 18710 38928 18710 4 vdd
port 513 nsew
rlabel metal1 s 39696 17920 39696 17920 4 vdd
port 513 nsew
rlabel metal1 s 38448 16839 38448 16839 4 vdd
port 513 nsew
rlabel metal1 s 37680 17130 37680 17130 4 vdd
port 513 nsew
rlabel metal1 s 38928 16049 38928 16049 4 vdd
port 513 nsew
rlabel metal1 s 38928 17130 38928 17130 4 vdd
port 513 nsew
rlabel metal1 s 38928 17629 38928 17629 4 vdd
port 513 nsew
rlabel metal1 s 38448 17920 38448 17920 4 vdd
port 513 nsew
rlabel metal1 s 37680 18710 37680 18710 4 vdd
port 513 nsew
rlabel metal1 s 38448 16340 38448 16340 4 vdd
port 513 nsew
rlabel metal1 s 37680 17629 37680 17629 4 vdd
port 513 nsew
rlabel metal1 s 37680 16839 37680 16839 4 vdd
port 513 nsew
rlabel metal1 s 38448 17130 38448 17130 4 vdd
port 513 nsew
rlabel metal1 s 39696 18710 39696 18710 4 vdd
port 513 nsew
rlabel metal1 s 38928 16340 38928 16340 4 vdd
port 513 nsew
rlabel metal1 s 38928 18419 38928 18419 4 vdd
port 513 nsew
rlabel metal1 s 37680 16049 37680 16049 4 vdd
port 513 nsew
rlabel metal1 s 38928 16839 38928 16839 4 vdd
port 513 nsew
rlabel metal1 s 38928 17920 38928 17920 4 vdd
port 513 nsew
rlabel metal1 s 36432 18419 36432 18419 4 vdd
port 513 nsew
rlabel metal1 s 35952 17920 35952 17920 4 vdd
port 513 nsew
rlabel metal1 s 35952 17130 35952 17130 4 vdd
port 513 nsew
rlabel metal1 s 35184 16049 35184 16049 4 vdd
port 513 nsew
rlabel metal1 s 36432 17920 36432 17920 4 vdd
port 513 nsew
rlabel metal1 s 36432 16839 36432 16839 4 vdd
port 513 nsew
rlabel metal1 s 35952 16839 35952 16839 4 vdd
port 513 nsew
rlabel metal1 s 35184 16839 35184 16839 4 vdd
port 513 nsew
rlabel metal1 s 35184 17629 35184 17629 4 vdd
port 513 nsew
rlabel metal1 s 35952 17629 35952 17629 4 vdd
port 513 nsew
rlabel metal1 s 35952 16049 35952 16049 4 vdd
port 513 nsew
rlabel metal1 s 35952 18710 35952 18710 4 vdd
port 513 nsew
rlabel metal1 s 35952 16340 35952 16340 4 vdd
port 513 nsew
rlabel metal1 s 37200 16049 37200 16049 4 vdd
port 513 nsew
rlabel metal1 s 36432 17629 36432 17629 4 vdd
port 513 nsew
rlabel metal1 s 36432 18710 36432 18710 4 vdd
port 513 nsew
rlabel metal1 s 35184 17920 35184 17920 4 vdd
port 513 nsew
rlabel metal1 s 37200 17920 37200 17920 4 vdd
port 513 nsew
rlabel metal1 s 35184 18710 35184 18710 4 vdd
port 513 nsew
rlabel metal1 s 37200 18419 37200 18419 4 vdd
port 513 nsew
rlabel metal1 s 35184 16340 35184 16340 4 vdd
port 513 nsew
rlabel metal1 s 36432 16049 36432 16049 4 vdd
port 513 nsew
rlabel metal1 s 37200 17130 37200 17130 4 vdd
port 513 nsew
rlabel metal1 s 36432 16340 36432 16340 4 vdd
port 513 nsew
rlabel metal1 s 37200 16340 37200 16340 4 vdd
port 513 nsew
rlabel metal1 s 35184 17130 35184 17130 4 vdd
port 513 nsew
rlabel metal1 s 37200 16839 37200 16839 4 vdd
port 513 nsew
rlabel metal1 s 35952 18419 35952 18419 4 vdd
port 513 nsew
rlabel metal1 s 37200 18710 37200 18710 4 vdd
port 513 nsew
rlabel metal1 s 35184 18419 35184 18419 4 vdd
port 513 nsew
rlabel metal1 s 37200 17629 37200 17629 4 vdd
port 513 nsew
rlabel metal1 s 36432 17130 36432 17130 4 vdd
port 513 nsew
rlabel metal1 s 35952 13180 35952 13180 4 vdd
port 513 nsew
rlabel metal1 s 35952 13679 35952 13679 4 vdd
port 513 nsew
rlabel metal1 s 35952 13970 35952 13970 4 vdd
port 513 nsew
rlabel metal1 s 37200 15259 37200 15259 4 vdd
port 513 nsew
rlabel metal1 s 35184 14760 35184 14760 4 vdd
port 513 nsew
rlabel metal1 s 35952 14469 35952 14469 4 vdd
port 513 nsew
rlabel metal1 s 35952 12889 35952 12889 4 vdd
port 513 nsew
rlabel metal1 s 35184 13970 35184 13970 4 vdd
port 513 nsew
rlabel metal1 s 37200 15550 37200 15550 4 vdd
port 513 nsew
rlabel metal1 s 35952 15550 35952 15550 4 vdd
port 513 nsew
rlabel metal1 s 36432 15550 36432 15550 4 vdd
port 513 nsew
rlabel metal1 s 37200 12889 37200 12889 4 vdd
port 513 nsew
rlabel metal1 s 36432 12889 36432 12889 4 vdd
port 513 nsew
rlabel metal1 s 36432 13970 36432 13970 4 vdd
port 513 nsew
rlabel metal1 s 35952 14760 35952 14760 4 vdd
port 513 nsew
rlabel metal1 s 35184 14469 35184 14469 4 vdd
port 513 nsew
rlabel metal1 s 37200 13679 37200 13679 4 vdd
port 513 nsew
rlabel metal1 s 36432 13679 36432 13679 4 vdd
port 513 nsew
rlabel metal1 s 35184 13679 35184 13679 4 vdd
port 513 nsew
rlabel metal1 s 37200 13180 37200 13180 4 vdd
port 513 nsew
rlabel metal1 s 36432 15259 36432 15259 4 vdd
port 513 nsew
rlabel metal1 s 37200 14469 37200 14469 4 vdd
port 513 nsew
rlabel metal1 s 35184 13180 35184 13180 4 vdd
port 513 nsew
rlabel metal1 s 35184 12889 35184 12889 4 vdd
port 513 nsew
rlabel metal1 s 35184 15550 35184 15550 4 vdd
port 513 nsew
rlabel metal1 s 37200 14760 37200 14760 4 vdd
port 513 nsew
rlabel metal1 s 36432 14760 36432 14760 4 vdd
port 513 nsew
rlabel metal1 s 37200 13970 37200 13970 4 vdd
port 513 nsew
rlabel metal1 s 36432 14469 36432 14469 4 vdd
port 513 nsew
rlabel metal1 s 35952 15259 35952 15259 4 vdd
port 513 nsew
rlabel metal1 s 36432 13180 36432 13180 4 vdd
port 513 nsew
rlabel metal1 s 35184 15259 35184 15259 4 vdd
port 513 nsew
rlabel metal1 s 38928 12889 38928 12889 4 vdd
port 513 nsew
rlabel metal1 s 38448 12889 38448 12889 4 vdd
port 513 nsew
rlabel metal1 s 38448 14469 38448 14469 4 vdd
port 513 nsew
rlabel metal1 s 38448 14760 38448 14760 4 vdd
port 513 nsew
rlabel metal1 s 37680 15259 37680 15259 4 vdd
port 513 nsew
rlabel metal1 s 38448 15259 38448 15259 4 vdd
port 513 nsew
rlabel metal1 s 37680 14469 37680 14469 4 vdd
port 513 nsew
rlabel metal1 s 37680 12889 37680 12889 4 vdd
port 513 nsew
rlabel metal1 s 38928 13970 38928 13970 4 vdd
port 513 nsew
rlabel metal1 s 38448 13180 38448 13180 4 vdd
port 513 nsew
rlabel metal1 s 39696 13970 39696 13970 4 vdd
port 513 nsew
rlabel metal1 s 39696 13180 39696 13180 4 vdd
port 513 nsew
rlabel metal1 s 38928 15550 38928 15550 4 vdd
port 513 nsew
rlabel metal1 s 38448 13679 38448 13679 4 vdd
port 513 nsew
rlabel metal1 s 38928 14760 38928 14760 4 vdd
port 513 nsew
rlabel metal1 s 37680 13679 37680 13679 4 vdd
port 513 nsew
rlabel metal1 s 39696 15550 39696 15550 4 vdd
port 513 nsew
rlabel metal1 s 38448 15550 38448 15550 4 vdd
port 513 nsew
rlabel metal1 s 37680 13970 37680 13970 4 vdd
port 513 nsew
rlabel metal1 s 38448 13970 38448 13970 4 vdd
port 513 nsew
rlabel metal1 s 38928 15259 38928 15259 4 vdd
port 513 nsew
rlabel metal1 s 39696 14760 39696 14760 4 vdd
port 513 nsew
rlabel metal1 s 37680 13180 37680 13180 4 vdd
port 513 nsew
rlabel metal1 s 37680 14760 37680 14760 4 vdd
port 513 nsew
rlabel metal1 s 39696 12889 39696 12889 4 vdd
port 513 nsew
rlabel metal1 s 39696 13679 39696 13679 4 vdd
port 513 nsew
rlabel metal1 s 38928 13679 38928 13679 4 vdd
port 513 nsew
rlabel metal1 s 37680 15550 37680 15550 4 vdd
port 513 nsew
rlabel metal1 s 38928 13180 38928 13180 4 vdd
port 513 nsew
rlabel metal1 s 39696 14469 39696 14469 4 vdd
port 513 nsew
rlabel metal1 s 38928 14469 38928 14469 4 vdd
port 513 nsew
rlabel metal1 s 39696 15259 39696 15259 4 vdd
port 513 nsew
rlabel metal1 s 27696 23159 27696 23159 4 vdd
port 513 nsew
rlabel metal1 s 29712 25030 29712 25030 4 vdd
port 513 nsew
rlabel metal1 s 27696 22660 27696 22660 4 vdd
port 513 nsew
rlabel metal1 s 27696 25030 27696 25030 4 vdd
port 513 nsew
rlabel metal1 s 29712 23450 29712 23450 4 vdd
port 513 nsew
rlabel metal1 s 28944 23159 28944 23159 4 vdd
port 513 nsew
rlabel metal1 s 29016 25280 29016 25280 4 bl1_46
port 187 nsew
rlabel metal1 s 28944 22660 28944 22660 4 vdd
port 513 nsew
rlabel metal1 s 28944 24240 28944 24240 4 vdd
port 513 nsew
rlabel metal1 s 29568 25280 29568 25280 4 br1_47
port 192 nsew
rlabel metal1 s 29712 23159 29712 23159 4 vdd
port 513 nsew
rlabel metal1 s 27840 25280 27840 25280 4 br1_44
port 180 nsew
rlabel metal1 s 27696 24240 27696 24240 4 vdd
port 513 nsew
rlabel metal1 s 28944 22369 28944 22369 4 vdd
port 513 nsew
rlabel metal1 s 27624 25280 27624 25280 4 br0_44
port 178 nsew
rlabel metal1 s 27552 25280 27552 25280 4 bl0_44
port 177 nsew
rlabel metal1 s 28944 23450 28944 23450 4 vdd
port 513 nsew
rlabel metal1 s 29712 24739 29712 24739 4 vdd
port 513 nsew
rlabel metal1 s 28464 24739 28464 24739 4 vdd
port 513 nsew
rlabel metal1 s 28464 25030 28464 25030 4 vdd
port 513 nsew
rlabel metal1 s 28608 25280 28608 25280 4 bl0_45
port 181 nsew
rlabel metal1 s 29712 23949 29712 23949 4 vdd
port 513 nsew
rlabel metal1 s 28464 23159 28464 23159 4 vdd
port 513 nsew
rlabel metal1 s 29640 25280 29640 25280 4 bl1_47
port 191 nsew
rlabel metal1 s 28944 23949 28944 23949 4 vdd
port 513 nsew
rlabel metal1 s 27696 24739 27696 24739 4 vdd
port 513 nsew
rlabel metal1 s 28464 23450 28464 23450 4 vdd
port 513 nsew
rlabel metal1 s 28320 25280 28320 25280 4 br1_45
port 184 nsew
rlabel metal1 s 28464 22369 28464 22369 4 vdd
port 513 nsew
rlabel metal1 s 28800 25280 28800 25280 4 bl0_46
port 185 nsew
rlabel metal1 s 27696 23949 27696 23949 4 vdd
port 513 nsew
rlabel metal1 s 28944 24739 28944 24739 4 vdd
port 513 nsew
rlabel metal1 s 27696 23450 27696 23450 4 vdd
port 513 nsew
rlabel metal1 s 28944 25030 28944 25030 4 vdd
port 513 nsew
rlabel metal1 s 29712 22369 29712 22369 4 vdd
port 513 nsew
rlabel metal1 s 29712 22660 29712 22660 4 vdd
port 513 nsew
rlabel metal1 s 29784 25280 29784 25280 4 br0_47
port 190 nsew
rlabel metal1 s 29856 25280 29856 25280 4 bl0_47
port 189 nsew
rlabel metal1 s 27696 22369 27696 22369 4 vdd
port 513 nsew
rlabel metal1 s 29088 25280 29088 25280 4 br1_46
port 188 nsew
rlabel metal1 s 28464 22660 28464 22660 4 vdd
port 513 nsew
rlabel metal1 s 28464 23949 28464 23949 4 vdd
port 513 nsew
rlabel metal1 s 28464 24240 28464 24240 4 vdd
port 513 nsew
rlabel metal1 s 27768 25280 27768 25280 4 bl1_44
port 179 nsew
rlabel metal1 s 28392 25280 28392 25280 4 bl1_45
port 183 nsew
rlabel metal1 s 29712 24240 29712 24240 4 vdd
port 513 nsew
rlabel metal1 s 28536 25280 28536 25280 4 br0_45
port 182 nsew
rlabel metal1 s 28872 25280 28872 25280 4 br0_46
port 186 nsew
rlabel metal1 s 26448 22369 26448 22369 4 vdd
port 513 nsew
rlabel metal1 s 26448 24240 26448 24240 4 vdd
port 513 nsew
rlabel metal1 s 25200 24739 25200 24739 4 vdd
port 513 nsew
rlabel metal1 s 27216 24240 27216 24240 4 vdd
port 513 nsew
rlabel metal1 s 25968 23949 25968 23949 4 vdd
port 513 nsew
rlabel metal1 s 27288 25280 27288 25280 4 br0_43
port 174 nsew
rlabel metal1 s 25200 24240 25200 24240 4 vdd
port 513 nsew
rlabel metal1 s 25200 23450 25200 23450 4 vdd
port 513 nsew
rlabel metal1 s 25968 23159 25968 23159 4 vdd
port 513 nsew
rlabel metal1 s 27216 23159 27216 23159 4 vdd
port 513 nsew
rlabel metal1 s 26448 25030 26448 25030 4 vdd
port 513 nsew
rlabel metal1 s 26376 25280 26376 25280 4 br0_42
port 170 nsew
rlabel metal1 s 26448 24739 26448 24739 4 vdd
port 513 nsew
rlabel metal1 s 26448 23159 26448 23159 4 vdd
port 513 nsew
rlabel metal1 s 26520 25280 26520 25280 4 bl1_42
port 171 nsew
rlabel metal1 s 27216 23450 27216 23450 4 vdd
port 513 nsew
rlabel metal1 s 27216 25030 27216 25030 4 vdd
port 513 nsew
rlabel metal1 s 26448 23450 26448 23450 4 vdd
port 513 nsew
rlabel metal1 s 27216 24739 27216 24739 4 vdd
port 513 nsew
rlabel metal1 s 25200 25030 25200 25030 4 vdd
port 513 nsew
rlabel metal1 s 25200 22660 25200 22660 4 vdd
port 513 nsew
rlabel metal1 s 25968 23450 25968 23450 4 vdd
port 513 nsew
rlabel metal1 s 25968 24240 25968 24240 4 vdd
port 513 nsew
rlabel metal1 s 25968 24739 25968 24739 4 vdd
port 513 nsew
rlabel metal1 s 27072 25280 27072 25280 4 br1_43
port 176 nsew
rlabel metal1 s 25200 23159 25200 23159 4 vdd
port 513 nsew
rlabel metal1 s 25128 25280 25128 25280 4 br0_40
port 162 nsew
rlabel metal1 s 25200 23949 25200 23949 4 vdd
port 513 nsew
rlabel metal1 s 25968 22660 25968 22660 4 vdd
port 513 nsew
rlabel metal1 s 25824 25280 25824 25280 4 br1_41
port 168 nsew
rlabel metal1 s 27360 25280 27360 25280 4 bl0_43
port 173 nsew
rlabel metal1 s 26040 25280 26040 25280 4 br0_41
port 166 nsew
rlabel metal1 s 25344 25280 25344 25280 4 br1_40
port 164 nsew
rlabel metal1 s 27216 23949 27216 23949 4 vdd
port 513 nsew
rlabel metal1 s 27216 22660 27216 22660 4 vdd
port 513 nsew
rlabel metal1 s 25968 22369 25968 22369 4 vdd
port 513 nsew
rlabel metal1 s 26448 23949 26448 23949 4 vdd
port 513 nsew
rlabel metal1 s 27216 22369 27216 22369 4 vdd
port 513 nsew
rlabel metal1 s 27144 25280 27144 25280 4 bl1_43
port 175 nsew
rlabel metal1 s 25200 22369 25200 22369 4 vdd
port 513 nsew
rlabel metal1 s 25272 25280 25272 25280 4 bl1_40
port 163 nsew
rlabel metal1 s 26112 25280 26112 25280 4 bl0_41
port 165 nsew
rlabel metal1 s 26592 25280 26592 25280 4 br1_42
port 172 nsew
rlabel metal1 s 26304 25280 26304 25280 4 bl0_42
port 169 nsew
rlabel metal1 s 26448 22660 26448 22660 4 vdd
port 513 nsew
rlabel metal1 s 25896 25280 25896 25280 4 bl1_41
port 167 nsew
rlabel metal1 s 25968 25030 25968 25030 4 vdd
port 513 nsew
rlabel metal1 s 25056 25280 25056 25280 4 bl0_40
port 161 nsew
rlabel metal1 s 25200 20789 25200 20789 4 vdd
port 513 nsew
rlabel metal1 s 26448 21579 26448 21579 4 vdd
port 513 nsew
rlabel metal1 s 27216 21080 27216 21080 4 vdd
port 513 nsew
rlabel metal1 s 25200 19209 25200 19209 4 vdd
port 513 nsew
rlabel metal1 s 25968 21579 25968 21579 4 vdd
port 513 nsew
rlabel metal1 s 26448 20290 26448 20290 4 vdd
port 513 nsew
rlabel metal1 s 27216 19500 27216 19500 4 vdd
port 513 nsew
rlabel metal1 s 25200 21870 25200 21870 4 vdd
port 513 nsew
rlabel metal1 s 27216 19209 27216 19209 4 vdd
port 513 nsew
rlabel metal1 s 26448 19999 26448 19999 4 vdd
port 513 nsew
rlabel metal1 s 26448 21080 26448 21080 4 vdd
port 513 nsew
rlabel metal1 s 25968 19999 25968 19999 4 vdd
port 513 nsew
rlabel metal1 s 25968 19209 25968 19209 4 vdd
port 513 nsew
rlabel metal1 s 25968 20290 25968 20290 4 vdd
port 513 nsew
rlabel metal1 s 27216 19999 27216 19999 4 vdd
port 513 nsew
rlabel metal1 s 27216 20789 27216 20789 4 vdd
port 513 nsew
rlabel metal1 s 25968 21080 25968 21080 4 vdd
port 513 nsew
rlabel metal1 s 25200 20290 25200 20290 4 vdd
port 513 nsew
rlabel metal1 s 26448 19209 26448 19209 4 vdd
port 513 nsew
rlabel metal1 s 26448 19500 26448 19500 4 vdd
port 513 nsew
rlabel metal1 s 25968 20789 25968 20789 4 vdd
port 513 nsew
rlabel metal1 s 25968 19500 25968 19500 4 vdd
port 513 nsew
rlabel metal1 s 26448 21870 26448 21870 4 vdd
port 513 nsew
rlabel metal1 s 25200 19500 25200 19500 4 vdd
port 513 nsew
rlabel metal1 s 25200 21080 25200 21080 4 vdd
port 513 nsew
rlabel metal1 s 25200 19999 25200 19999 4 vdd
port 513 nsew
rlabel metal1 s 26448 20789 26448 20789 4 vdd
port 513 nsew
rlabel metal1 s 27216 21579 27216 21579 4 vdd
port 513 nsew
rlabel metal1 s 27216 20290 27216 20290 4 vdd
port 513 nsew
rlabel metal1 s 27216 21870 27216 21870 4 vdd
port 513 nsew
rlabel metal1 s 25968 21870 25968 21870 4 vdd
port 513 nsew
rlabel metal1 s 25200 21579 25200 21579 4 vdd
port 513 nsew
rlabel metal1 s 28944 19999 28944 19999 4 vdd
port 513 nsew
rlabel metal1 s 29712 20290 29712 20290 4 vdd
port 513 nsew
rlabel metal1 s 27696 21579 27696 21579 4 vdd
port 513 nsew
rlabel metal1 s 28464 21870 28464 21870 4 vdd
port 513 nsew
rlabel metal1 s 29712 21870 29712 21870 4 vdd
port 513 nsew
rlabel metal1 s 28464 21579 28464 21579 4 vdd
port 513 nsew
rlabel metal1 s 28464 19999 28464 19999 4 vdd
port 513 nsew
rlabel metal1 s 29712 21579 29712 21579 4 vdd
port 513 nsew
rlabel metal1 s 28464 20290 28464 20290 4 vdd
port 513 nsew
rlabel metal1 s 29712 19999 29712 19999 4 vdd
port 513 nsew
rlabel metal1 s 27696 21080 27696 21080 4 vdd
port 513 nsew
rlabel metal1 s 28464 20789 28464 20789 4 vdd
port 513 nsew
rlabel metal1 s 29712 20789 29712 20789 4 vdd
port 513 nsew
rlabel metal1 s 27696 19500 27696 19500 4 vdd
port 513 nsew
rlabel metal1 s 27696 19209 27696 19209 4 vdd
port 513 nsew
rlabel metal1 s 27696 20290 27696 20290 4 vdd
port 513 nsew
rlabel metal1 s 29712 19500 29712 19500 4 vdd
port 513 nsew
rlabel metal1 s 27696 20789 27696 20789 4 vdd
port 513 nsew
rlabel metal1 s 29712 21080 29712 21080 4 vdd
port 513 nsew
rlabel metal1 s 28944 19500 28944 19500 4 vdd
port 513 nsew
rlabel metal1 s 28944 20290 28944 20290 4 vdd
port 513 nsew
rlabel metal1 s 28464 19209 28464 19209 4 vdd
port 513 nsew
rlabel metal1 s 28944 21870 28944 21870 4 vdd
port 513 nsew
rlabel metal1 s 27696 19999 27696 19999 4 vdd
port 513 nsew
rlabel metal1 s 28944 20789 28944 20789 4 vdd
port 513 nsew
rlabel metal1 s 27696 21870 27696 21870 4 vdd
port 513 nsew
rlabel metal1 s 28944 21579 28944 21579 4 vdd
port 513 nsew
rlabel metal1 s 28944 19209 28944 19209 4 vdd
port 513 nsew
rlabel metal1 s 28464 21080 28464 21080 4 vdd
port 513 nsew
rlabel metal1 s 28944 21080 28944 21080 4 vdd
port 513 nsew
rlabel metal1 s 29712 19209 29712 19209 4 vdd
port 513 nsew
rlabel metal1 s 28464 19500 28464 19500 4 vdd
port 513 nsew
rlabel metal1 s 24096 25280 24096 25280 4 br1_38
port 156 nsew
rlabel metal1 s 22776 25280 22776 25280 4 bl1_36
port 147 nsew
rlabel metal1 s 23472 25030 23472 25030 4 vdd
port 513 nsew
rlabel metal1 s 22704 23159 22704 23159 4 vdd
port 513 nsew
rlabel metal1 s 22704 24739 22704 24739 4 vdd
port 513 nsew
rlabel metal1 s 23472 23159 23472 23159 4 vdd
port 513 nsew
rlabel metal1 s 23544 25280 23544 25280 4 br0_37
port 150 nsew
rlabel metal1 s 23952 25030 23952 25030 4 vdd
port 513 nsew
rlabel metal1 s 22704 23450 22704 23450 4 vdd
port 513 nsew
rlabel metal1 s 22632 25280 22632 25280 4 br0_36
port 146 nsew
rlabel metal1 s 22704 22660 22704 22660 4 vdd
port 513 nsew
rlabel metal1 s 24648 25280 24648 25280 4 bl1_39
port 159 nsew
rlabel metal1 s 24720 24739 24720 24739 4 vdd
port 513 nsew
rlabel metal1 s 23472 22660 23472 22660 4 vdd
port 513 nsew
rlabel metal1 s 24792 25280 24792 25280 4 br0_39
port 158 nsew
rlabel metal1 s 22560 25280 22560 25280 4 bl0_36
port 145 nsew
rlabel metal1 s 23808 25280 23808 25280 4 bl0_38
port 153 nsew
rlabel metal1 s 23952 23450 23952 23450 4 vdd
port 513 nsew
rlabel metal1 s 24720 24240 24720 24240 4 vdd
port 513 nsew
rlabel metal1 s 23952 23949 23952 23949 4 vdd
port 513 nsew
rlabel metal1 s 24864 25280 24864 25280 4 bl0_39
port 157 nsew
rlabel metal1 s 24720 23949 24720 23949 4 vdd
port 513 nsew
rlabel metal1 s 23952 22660 23952 22660 4 vdd
port 513 nsew
rlabel metal1 s 23400 25280 23400 25280 4 bl1_37
port 151 nsew
rlabel metal1 s 23952 24739 23952 24739 4 vdd
port 513 nsew
rlabel metal1 s 23952 22369 23952 22369 4 vdd
port 513 nsew
rlabel metal1 s 24720 22660 24720 22660 4 vdd
port 513 nsew
rlabel metal1 s 23880 25280 23880 25280 4 br0_38
port 154 nsew
rlabel metal1 s 24720 23450 24720 23450 4 vdd
port 513 nsew
rlabel metal1 s 22704 23949 22704 23949 4 vdd
port 513 nsew
rlabel metal1 s 24024 25280 24024 25280 4 bl1_38
port 155 nsew
rlabel metal1 s 23616 25280 23616 25280 4 bl0_37
port 149 nsew
rlabel metal1 s 22704 22369 22704 22369 4 vdd
port 513 nsew
rlabel metal1 s 22848 25280 22848 25280 4 br1_36
port 148 nsew
rlabel metal1 s 23328 25280 23328 25280 4 br1_37
port 152 nsew
rlabel metal1 s 24576 25280 24576 25280 4 br1_39
port 160 nsew
rlabel metal1 s 23952 24240 23952 24240 4 vdd
port 513 nsew
rlabel metal1 s 23472 22369 23472 22369 4 vdd
port 513 nsew
rlabel metal1 s 23472 24240 23472 24240 4 vdd
port 513 nsew
rlabel metal1 s 24720 23159 24720 23159 4 vdd
port 513 nsew
rlabel metal1 s 24720 22369 24720 22369 4 vdd
port 513 nsew
rlabel metal1 s 23472 24739 23472 24739 4 vdd
port 513 nsew
rlabel metal1 s 22704 24240 22704 24240 4 vdd
port 513 nsew
rlabel metal1 s 23472 23450 23472 23450 4 vdd
port 513 nsew
rlabel metal1 s 23952 23159 23952 23159 4 vdd
port 513 nsew
rlabel metal1 s 24720 25030 24720 25030 4 vdd
port 513 nsew
rlabel metal1 s 23472 23949 23472 23949 4 vdd
port 513 nsew
rlabel metal1 s 22704 25030 22704 25030 4 vdd
port 513 nsew
rlabel metal1 s 21456 23450 21456 23450 4 vdd
port 513 nsew
rlabel metal1 s 22224 23949 22224 23949 4 vdd
port 513 nsew
rlabel metal1 s 22224 24240 22224 24240 4 vdd
port 513 nsew
rlabel metal1 s 22296 25280 22296 25280 4 br0_35
port 142 nsew
rlabel metal1 s 22224 25030 22224 25030 4 vdd
port 513 nsew
rlabel metal1 s 22224 23159 22224 23159 4 vdd
port 513 nsew
rlabel metal1 s 22224 22369 22224 22369 4 vdd
port 513 nsew
rlabel metal1 s 20976 24739 20976 24739 4 vdd
port 513 nsew
rlabel metal1 s 20280 25280 20280 25280 4 bl1_32
port 131 nsew
rlabel metal1 s 21456 23949 21456 23949 4 vdd
port 513 nsew
rlabel metal1 s 20208 23949 20208 23949 4 vdd
port 513 nsew
rlabel metal1 s 20208 23450 20208 23450 4 vdd
port 513 nsew
rlabel metal1 s 20976 25030 20976 25030 4 vdd
port 513 nsew
rlabel metal1 s 20208 23159 20208 23159 4 vdd
port 513 nsew
rlabel metal1 s 20976 23450 20976 23450 4 vdd
port 513 nsew
rlabel metal1 s 20136 25280 20136 25280 4 br0_32
port 130 nsew
rlabel metal1 s 20352 25280 20352 25280 4 br1_32
port 132 nsew
rlabel metal1 s 20976 23949 20976 23949 4 vdd
port 513 nsew
rlabel metal1 s 20976 22369 20976 22369 4 vdd
port 513 nsew
rlabel metal1 s 20976 23159 20976 23159 4 vdd
port 513 nsew
rlabel metal1 s 21600 25280 21600 25280 4 br1_34
port 140 nsew
rlabel metal1 s 21456 22660 21456 22660 4 vdd
port 513 nsew
rlabel metal1 s 21456 24240 21456 24240 4 vdd
port 513 nsew
rlabel metal1 s 20976 22660 20976 22660 4 vdd
port 513 nsew
rlabel metal1 s 21456 23159 21456 23159 4 vdd
port 513 nsew
rlabel metal1 s 21528 25280 21528 25280 4 bl1_34
port 139 nsew
rlabel metal1 s 20976 24240 20976 24240 4 vdd
port 513 nsew
rlabel metal1 s 21456 24739 21456 24739 4 vdd
port 513 nsew
rlabel metal1 s 21120 25280 21120 25280 4 bl0_33
port 133 nsew
rlabel metal1 s 20208 22369 20208 22369 4 vdd
port 513 nsew
rlabel metal1 s 21312 25280 21312 25280 4 bl0_34
port 137 nsew
rlabel metal1 s 22224 23450 22224 23450 4 vdd
port 513 nsew
rlabel metal1 s 20064 25280 20064 25280 4 bl0_32
port 129 nsew
rlabel metal1 s 21384 25280 21384 25280 4 br0_34
port 138 nsew
rlabel metal1 s 22152 25280 22152 25280 4 bl1_35
port 143 nsew
rlabel metal1 s 20208 22660 20208 22660 4 vdd
port 513 nsew
rlabel metal1 s 20208 24240 20208 24240 4 vdd
port 513 nsew
rlabel metal1 s 22368 25280 22368 25280 4 bl0_35
port 141 nsew
rlabel metal1 s 20208 24739 20208 24739 4 vdd
port 513 nsew
rlabel metal1 s 22224 24739 22224 24739 4 vdd
port 513 nsew
rlabel metal1 s 20208 25030 20208 25030 4 vdd
port 513 nsew
rlabel metal1 s 21456 22369 21456 22369 4 vdd
port 513 nsew
rlabel metal1 s 21048 25280 21048 25280 4 br0_33
port 134 nsew
rlabel metal1 s 22224 22660 22224 22660 4 vdd
port 513 nsew
rlabel metal1 s 22080 25280 22080 25280 4 br1_35
port 144 nsew
rlabel metal1 s 21456 25030 21456 25030 4 vdd
port 513 nsew
rlabel metal1 s 20832 25280 20832 25280 4 br1_33
port 136 nsew
rlabel metal1 s 20904 25280 20904 25280 4 bl1_33
port 135 nsew
rlabel metal1 s 20208 19209 20208 19209 4 vdd
port 513 nsew
rlabel metal1 s 20976 19999 20976 19999 4 vdd
port 513 nsew
rlabel metal1 s 21456 20789 21456 20789 4 vdd
port 513 nsew
rlabel metal1 s 22224 21579 22224 21579 4 vdd
port 513 nsew
rlabel metal1 s 20208 19999 20208 19999 4 vdd
port 513 nsew
rlabel metal1 s 22224 21870 22224 21870 4 vdd
port 513 nsew
rlabel metal1 s 20976 20789 20976 20789 4 vdd
port 513 nsew
rlabel metal1 s 20208 20290 20208 20290 4 vdd
port 513 nsew
rlabel metal1 s 20976 19209 20976 19209 4 vdd
port 513 nsew
rlabel metal1 s 21456 19999 21456 19999 4 vdd
port 513 nsew
rlabel metal1 s 22224 19999 22224 19999 4 vdd
port 513 nsew
rlabel metal1 s 21456 21080 21456 21080 4 vdd
port 513 nsew
rlabel metal1 s 20976 21579 20976 21579 4 vdd
port 513 nsew
rlabel metal1 s 20976 20290 20976 20290 4 vdd
port 513 nsew
rlabel metal1 s 21456 19209 21456 19209 4 vdd
port 513 nsew
rlabel metal1 s 21456 19500 21456 19500 4 vdd
port 513 nsew
rlabel metal1 s 22224 21080 22224 21080 4 vdd
port 513 nsew
rlabel metal1 s 22224 19500 22224 19500 4 vdd
port 513 nsew
rlabel metal1 s 20976 19500 20976 19500 4 vdd
port 513 nsew
rlabel metal1 s 21456 21579 21456 21579 4 vdd
port 513 nsew
rlabel metal1 s 21456 21870 21456 21870 4 vdd
port 513 nsew
rlabel metal1 s 20976 21080 20976 21080 4 vdd
port 513 nsew
rlabel metal1 s 20208 21579 20208 21579 4 vdd
port 513 nsew
rlabel metal1 s 22224 20290 22224 20290 4 vdd
port 513 nsew
rlabel metal1 s 20208 19500 20208 19500 4 vdd
port 513 nsew
rlabel metal1 s 20208 21870 20208 21870 4 vdd
port 513 nsew
rlabel metal1 s 20208 20789 20208 20789 4 vdd
port 513 nsew
rlabel metal1 s 22224 20789 22224 20789 4 vdd
port 513 nsew
rlabel metal1 s 20208 21080 20208 21080 4 vdd
port 513 nsew
rlabel metal1 s 21456 20290 21456 20290 4 vdd
port 513 nsew
rlabel metal1 s 20976 21870 20976 21870 4 vdd
port 513 nsew
rlabel metal1 s 22224 19209 22224 19209 4 vdd
port 513 nsew
rlabel metal1 s 23472 21579 23472 21579 4 vdd
port 513 nsew
rlabel metal1 s 23952 19209 23952 19209 4 vdd
port 513 nsew
rlabel metal1 s 23472 20789 23472 20789 4 vdd
port 513 nsew
rlabel metal1 s 23472 19209 23472 19209 4 vdd
port 513 nsew
rlabel metal1 s 22704 20290 22704 20290 4 vdd
port 513 nsew
rlabel metal1 s 23952 19999 23952 19999 4 vdd
port 513 nsew
rlabel metal1 s 22704 20789 22704 20789 4 vdd
port 513 nsew
rlabel metal1 s 23472 19500 23472 19500 4 vdd
port 513 nsew
rlabel metal1 s 23472 20290 23472 20290 4 vdd
port 513 nsew
rlabel metal1 s 24720 20290 24720 20290 4 vdd
port 513 nsew
rlabel metal1 s 23952 19500 23952 19500 4 vdd
port 513 nsew
rlabel metal1 s 23952 20290 23952 20290 4 vdd
port 513 nsew
rlabel metal1 s 22704 21870 22704 21870 4 vdd
port 513 nsew
rlabel metal1 s 22704 21080 22704 21080 4 vdd
port 513 nsew
rlabel metal1 s 22704 21579 22704 21579 4 vdd
port 513 nsew
rlabel metal1 s 24720 19500 24720 19500 4 vdd
port 513 nsew
rlabel metal1 s 23952 21870 23952 21870 4 vdd
port 513 nsew
rlabel metal1 s 22704 19209 22704 19209 4 vdd
port 513 nsew
rlabel metal1 s 23952 21080 23952 21080 4 vdd
port 513 nsew
rlabel metal1 s 24720 21579 24720 21579 4 vdd
port 513 nsew
rlabel metal1 s 22704 19999 22704 19999 4 vdd
port 513 nsew
rlabel metal1 s 24720 19999 24720 19999 4 vdd
port 513 nsew
rlabel metal1 s 22704 19500 22704 19500 4 vdd
port 513 nsew
rlabel metal1 s 23952 20789 23952 20789 4 vdd
port 513 nsew
rlabel metal1 s 24720 21870 24720 21870 4 vdd
port 513 nsew
rlabel metal1 s 24720 19209 24720 19209 4 vdd
port 513 nsew
rlabel metal1 s 23952 21579 23952 21579 4 vdd
port 513 nsew
rlabel metal1 s 23472 21870 23472 21870 4 vdd
port 513 nsew
rlabel metal1 s 24720 20789 24720 20789 4 vdd
port 513 nsew
rlabel metal1 s 23472 19999 23472 19999 4 vdd
port 513 nsew
rlabel metal1 s 23472 21080 23472 21080 4 vdd
port 513 nsew
rlabel metal1 s 24720 21080 24720 21080 4 vdd
port 513 nsew
rlabel metal1 s 23952 18710 23952 18710 4 vdd
port 513 nsew
rlabel metal1 s 23952 16340 23952 16340 4 vdd
port 513 nsew
rlabel metal1 s 23952 17130 23952 17130 4 vdd
port 513 nsew
rlabel metal1 s 24720 16839 24720 16839 4 vdd
port 513 nsew
rlabel metal1 s 22704 17920 22704 17920 4 vdd
port 513 nsew
rlabel metal1 s 24720 18419 24720 18419 4 vdd
port 513 nsew
rlabel metal1 s 23472 16340 23472 16340 4 vdd
port 513 nsew
rlabel metal1 s 24720 18710 24720 18710 4 vdd
port 513 nsew
rlabel metal1 s 24720 17130 24720 17130 4 vdd
port 513 nsew
rlabel metal1 s 22704 18419 22704 18419 4 vdd
port 513 nsew
rlabel metal1 s 22704 17130 22704 17130 4 vdd
port 513 nsew
rlabel metal1 s 24720 17629 24720 17629 4 vdd
port 513 nsew
rlabel metal1 s 24720 17920 24720 17920 4 vdd
port 513 nsew
rlabel metal1 s 23472 18710 23472 18710 4 vdd
port 513 nsew
rlabel metal1 s 22704 16049 22704 16049 4 vdd
port 513 nsew
rlabel metal1 s 23952 17920 23952 17920 4 vdd
port 513 nsew
rlabel metal1 s 23472 16049 23472 16049 4 vdd
port 513 nsew
rlabel metal1 s 23952 18419 23952 18419 4 vdd
port 513 nsew
rlabel metal1 s 23472 17629 23472 17629 4 vdd
port 513 nsew
rlabel metal1 s 23472 16839 23472 16839 4 vdd
port 513 nsew
rlabel metal1 s 24720 16049 24720 16049 4 vdd
port 513 nsew
rlabel metal1 s 22704 17629 22704 17629 4 vdd
port 513 nsew
rlabel metal1 s 23952 16839 23952 16839 4 vdd
port 513 nsew
rlabel metal1 s 22704 16340 22704 16340 4 vdd
port 513 nsew
rlabel metal1 s 23472 18419 23472 18419 4 vdd
port 513 nsew
rlabel metal1 s 24720 16340 24720 16340 4 vdd
port 513 nsew
rlabel metal1 s 22704 16839 22704 16839 4 vdd
port 513 nsew
rlabel metal1 s 23472 17130 23472 17130 4 vdd
port 513 nsew
rlabel metal1 s 23472 17920 23472 17920 4 vdd
port 513 nsew
rlabel metal1 s 23952 16049 23952 16049 4 vdd
port 513 nsew
rlabel metal1 s 22704 18710 22704 18710 4 vdd
port 513 nsew
rlabel metal1 s 23952 17629 23952 17629 4 vdd
port 513 nsew
rlabel metal1 s 22224 16340 22224 16340 4 vdd
port 513 nsew
rlabel metal1 s 20208 18419 20208 18419 4 vdd
port 513 nsew
rlabel metal1 s 20208 16839 20208 16839 4 vdd
port 513 nsew
rlabel metal1 s 22224 17920 22224 17920 4 vdd
port 513 nsew
rlabel metal1 s 21456 17130 21456 17130 4 vdd
port 513 nsew
rlabel metal1 s 20976 17130 20976 17130 4 vdd
port 513 nsew
rlabel metal1 s 20976 16340 20976 16340 4 vdd
port 513 nsew
rlabel metal1 s 20208 16340 20208 16340 4 vdd
port 513 nsew
rlabel metal1 s 20208 17629 20208 17629 4 vdd
port 513 nsew
rlabel metal1 s 20208 17130 20208 17130 4 vdd
port 513 nsew
rlabel metal1 s 22224 16839 22224 16839 4 vdd
port 513 nsew
rlabel metal1 s 22224 17130 22224 17130 4 vdd
port 513 nsew
rlabel metal1 s 22224 17629 22224 17629 4 vdd
port 513 nsew
rlabel metal1 s 21456 16049 21456 16049 4 vdd
port 513 nsew
rlabel metal1 s 21456 18710 21456 18710 4 vdd
port 513 nsew
rlabel metal1 s 20976 18419 20976 18419 4 vdd
port 513 nsew
rlabel metal1 s 21456 16340 21456 16340 4 vdd
port 513 nsew
rlabel metal1 s 20976 18710 20976 18710 4 vdd
port 513 nsew
rlabel metal1 s 21456 16839 21456 16839 4 vdd
port 513 nsew
rlabel metal1 s 21456 17629 21456 17629 4 vdd
port 513 nsew
rlabel metal1 s 21456 17920 21456 17920 4 vdd
port 513 nsew
rlabel metal1 s 20976 17629 20976 17629 4 vdd
port 513 nsew
rlabel metal1 s 20976 17920 20976 17920 4 vdd
port 513 nsew
rlabel metal1 s 22224 18710 22224 18710 4 vdd
port 513 nsew
rlabel metal1 s 21456 18419 21456 18419 4 vdd
port 513 nsew
rlabel metal1 s 20208 17920 20208 17920 4 vdd
port 513 nsew
rlabel metal1 s 20208 18710 20208 18710 4 vdd
port 513 nsew
rlabel metal1 s 20208 16049 20208 16049 4 vdd
port 513 nsew
rlabel metal1 s 22224 18419 22224 18419 4 vdd
port 513 nsew
rlabel metal1 s 22224 16049 22224 16049 4 vdd
port 513 nsew
rlabel metal1 s 20976 16839 20976 16839 4 vdd
port 513 nsew
rlabel metal1 s 20976 16049 20976 16049 4 vdd
port 513 nsew
rlabel metal1 s 21456 12889 21456 12889 4 vdd
port 513 nsew
rlabel metal1 s 20976 13970 20976 13970 4 vdd
port 513 nsew
rlabel metal1 s 22224 13679 22224 13679 4 vdd
port 513 nsew
rlabel metal1 s 20208 13970 20208 13970 4 vdd
port 513 nsew
rlabel metal1 s 21456 15259 21456 15259 4 vdd
port 513 nsew
rlabel metal1 s 20208 14469 20208 14469 4 vdd
port 513 nsew
rlabel metal1 s 20208 15550 20208 15550 4 vdd
port 513 nsew
rlabel metal1 s 20208 15259 20208 15259 4 vdd
port 513 nsew
rlabel metal1 s 22224 13970 22224 13970 4 vdd
port 513 nsew
rlabel metal1 s 22224 14469 22224 14469 4 vdd
port 513 nsew
rlabel metal1 s 21456 13180 21456 13180 4 vdd
port 513 nsew
rlabel metal1 s 20976 15550 20976 15550 4 vdd
port 513 nsew
rlabel metal1 s 20976 13180 20976 13180 4 vdd
port 513 nsew
rlabel metal1 s 21456 15550 21456 15550 4 vdd
port 513 nsew
rlabel metal1 s 20976 15259 20976 15259 4 vdd
port 513 nsew
rlabel metal1 s 20208 13679 20208 13679 4 vdd
port 513 nsew
rlabel metal1 s 20976 14469 20976 14469 4 vdd
port 513 nsew
rlabel metal1 s 22224 12889 22224 12889 4 vdd
port 513 nsew
rlabel metal1 s 22224 14760 22224 14760 4 vdd
port 513 nsew
rlabel metal1 s 22224 15550 22224 15550 4 vdd
port 513 nsew
rlabel metal1 s 21456 14760 21456 14760 4 vdd
port 513 nsew
rlabel metal1 s 20976 13679 20976 13679 4 vdd
port 513 nsew
rlabel metal1 s 22224 13180 22224 13180 4 vdd
port 513 nsew
rlabel metal1 s 20976 12889 20976 12889 4 vdd
port 513 nsew
rlabel metal1 s 21456 13970 21456 13970 4 vdd
port 513 nsew
rlabel metal1 s 20976 14760 20976 14760 4 vdd
port 513 nsew
rlabel metal1 s 21456 13679 21456 13679 4 vdd
port 513 nsew
rlabel metal1 s 22224 15259 22224 15259 4 vdd
port 513 nsew
rlabel metal1 s 20208 13180 20208 13180 4 vdd
port 513 nsew
rlabel metal1 s 20208 12889 20208 12889 4 vdd
port 513 nsew
rlabel metal1 s 21456 14469 21456 14469 4 vdd
port 513 nsew
rlabel metal1 s 20208 14760 20208 14760 4 vdd
port 513 nsew
rlabel metal1 s 23472 14760 23472 14760 4 vdd
port 513 nsew
rlabel metal1 s 23472 15550 23472 15550 4 vdd
port 513 nsew
rlabel metal1 s 23472 14469 23472 14469 4 vdd
port 513 nsew
rlabel metal1 s 23472 13679 23472 13679 4 vdd
port 513 nsew
rlabel metal1 s 24720 15259 24720 15259 4 vdd
port 513 nsew
rlabel metal1 s 23952 14760 23952 14760 4 vdd
port 513 nsew
rlabel metal1 s 22704 14469 22704 14469 4 vdd
port 513 nsew
rlabel metal1 s 22704 15550 22704 15550 4 vdd
port 513 nsew
rlabel metal1 s 22704 13970 22704 13970 4 vdd
port 513 nsew
rlabel metal1 s 22704 15259 22704 15259 4 vdd
port 513 nsew
rlabel metal1 s 23472 13970 23472 13970 4 vdd
port 513 nsew
rlabel metal1 s 23952 13180 23952 13180 4 vdd
port 513 nsew
rlabel metal1 s 22704 14760 22704 14760 4 vdd
port 513 nsew
rlabel metal1 s 23472 13180 23472 13180 4 vdd
port 513 nsew
rlabel metal1 s 24720 14760 24720 14760 4 vdd
port 513 nsew
rlabel metal1 s 24720 12889 24720 12889 4 vdd
port 513 nsew
rlabel metal1 s 22704 12889 22704 12889 4 vdd
port 513 nsew
rlabel metal1 s 24720 13679 24720 13679 4 vdd
port 513 nsew
rlabel metal1 s 24720 15550 24720 15550 4 vdd
port 513 nsew
rlabel metal1 s 24720 13180 24720 13180 4 vdd
port 513 nsew
rlabel metal1 s 23952 15550 23952 15550 4 vdd
port 513 nsew
rlabel metal1 s 24720 13970 24720 13970 4 vdd
port 513 nsew
rlabel metal1 s 22704 13679 22704 13679 4 vdd
port 513 nsew
rlabel metal1 s 23472 12889 23472 12889 4 vdd
port 513 nsew
rlabel metal1 s 23952 13679 23952 13679 4 vdd
port 513 nsew
rlabel metal1 s 24720 14469 24720 14469 4 vdd
port 513 nsew
rlabel metal1 s 23952 12889 23952 12889 4 vdd
port 513 nsew
rlabel metal1 s 23472 15259 23472 15259 4 vdd
port 513 nsew
rlabel metal1 s 23952 14469 23952 14469 4 vdd
port 513 nsew
rlabel metal1 s 23952 15259 23952 15259 4 vdd
port 513 nsew
rlabel metal1 s 23952 13970 23952 13970 4 vdd
port 513 nsew
rlabel metal1 s 22704 13180 22704 13180 4 vdd
port 513 nsew
rlabel metal1 s 29712 18710 29712 18710 4 vdd
port 513 nsew
rlabel metal1 s 27696 16340 27696 16340 4 vdd
port 513 nsew
rlabel metal1 s 28944 17130 28944 17130 4 vdd
port 513 nsew
rlabel metal1 s 29712 17130 29712 17130 4 vdd
port 513 nsew
rlabel metal1 s 27696 17629 27696 17629 4 vdd
port 513 nsew
rlabel metal1 s 28464 17130 28464 17130 4 vdd
port 513 nsew
rlabel metal1 s 29712 17920 29712 17920 4 vdd
port 513 nsew
rlabel metal1 s 28944 16839 28944 16839 4 vdd
port 513 nsew
rlabel metal1 s 29712 16839 29712 16839 4 vdd
port 513 nsew
rlabel metal1 s 27696 16839 27696 16839 4 vdd
port 513 nsew
rlabel metal1 s 28944 16049 28944 16049 4 vdd
port 513 nsew
rlabel metal1 s 28464 17920 28464 17920 4 vdd
port 513 nsew
rlabel metal1 s 27696 16049 27696 16049 4 vdd
port 513 nsew
rlabel metal1 s 28464 16839 28464 16839 4 vdd
port 513 nsew
rlabel metal1 s 28464 16340 28464 16340 4 vdd
port 513 nsew
rlabel metal1 s 28944 17920 28944 17920 4 vdd
port 513 nsew
rlabel metal1 s 28944 18419 28944 18419 4 vdd
port 513 nsew
rlabel metal1 s 29712 16340 29712 16340 4 vdd
port 513 nsew
rlabel metal1 s 27696 18710 27696 18710 4 vdd
port 513 nsew
rlabel metal1 s 28464 16049 28464 16049 4 vdd
port 513 nsew
rlabel metal1 s 28464 18710 28464 18710 4 vdd
port 513 nsew
rlabel metal1 s 27696 18419 27696 18419 4 vdd
port 513 nsew
rlabel metal1 s 27696 17130 27696 17130 4 vdd
port 513 nsew
rlabel metal1 s 29712 16049 29712 16049 4 vdd
port 513 nsew
rlabel metal1 s 28464 18419 28464 18419 4 vdd
port 513 nsew
rlabel metal1 s 28944 17629 28944 17629 4 vdd
port 513 nsew
rlabel metal1 s 28944 18710 28944 18710 4 vdd
port 513 nsew
rlabel metal1 s 29712 18419 29712 18419 4 vdd
port 513 nsew
rlabel metal1 s 28464 17629 28464 17629 4 vdd
port 513 nsew
rlabel metal1 s 28944 16340 28944 16340 4 vdd
port 513 nsew
rlabel metal1 s 27696 17920 27696 17920 4 vdd
port 513 nsew
rlabel metal1 s 29712 17629 29712 17629 4 vdd
port 513 nsew
rlabel metal1 s 25968 17629 25968 17629 4 vdd
port 513 nsew
rlabel metal1 s 26448 17920 26448 17920 4 vdd
port 513 nsew
rlabel metal1 s 25200 16340 25200 16340 4 vdd
port 513 nsew
rlabel metal1 s 27216 18419 27216 18419 4 vdd
port 513 nsew
rlabel metal1 s 27216 17130 27216 17130 4 vdd
port 513 nsew
rlabel metal1 s 25968 18710 25968 18710 4 vdd
port 513 nsew
rlabel metal1 s 27216 18710 27216 18710 4 vdd
port 513 nsew
rlabel metal1 s 25200 17130 25200 17130 4 vdd
port 513 nsew
rlabel metal1 s 26448 17130 26448 17130 4 vdd
port 513 nsew
rlabel metal1 s 25968 16340 25968 16340 4 vdd
port 513 nsew
rlabel metal1 s 27216 17920 27216 17920 4 vdd
port 513 nsew
rlabel metal1 s 26448 18710 26448 18710 4 vdd
port 513 nsew
rlabel metal1 s 25200 16049 25200 16049 4 vdd
port 513 nsew
rlabel metal1 s 25200 18419 25200 18419 4 vdd
port 513 nsew
rlabel metal1 s 26448 16340 26448 16340 4 vdd
port 513 nsew
rlabel metal1 s 27216 17629 27216 17629 4 vdd
port 513 nsew
rlabel metal1 s 25200 17920 25200 17920 4 vdd
port 513 nsew
rlabel metal1 s 25200 16839 25200 16839 4 vdd
port 513 nsew
rlabel metal1 s 25200 17629 25200 17629 4 vdd
port 513 nsew
rlabel metal1 s 26448 16839 26448 16839 4 vdd
port 513 nsew
rlabel metal1 s 27216 16340 27216 16340 4 vdd
port 513 nsew
rlabel metal1 s 25968 16839 25968 16839 4 vdd
port 513 nsew
rlabel metal1 s 26448 16049 26448 16049 4 vdd
port 513 nsew
rlabel metal1 s 26448 18419 26448 18419 4 vdd
port 513 nsew
rlabel metal1 s 26448 17629 26448 17629 4 vdd
port 513 nsew
rlabel metal1 s 25968 18419 25968 18419 4 vdd
port 513 nsew
rlabel metal1 s 27216 16049 27216 16049 4 vdd
port 513 nsew
rlabel metal1 s 25200 18710 25200 18710 4 vdd
port 513 nsew
rlabel metal1 s 25968 17920 25968 17920 4 vdd
port 513 nsew
rlabel metal1 s 25968 17130 25968 17130 4 vdd
port 513 nsew
rlabel metal1 s 25968 16049 25968 16049 4 vdd
port 513 nsew
rlabel metal1 s 27216 16839 27216 16839 4 vdd
port 513 nsew
rlabel metal1 s 26448 15259 26448 15259 4 vdd
port 513 nsew
rlabel metal1 s 26448 12889 26448 12889 4 vdd
port 513 nsew
rlabel metal1 s 25968 13679 25968 13679 4 vdd
port 513 nsew
rlabel metal1 s 27216 14469 27216 14469 4 vdd
port 513 nsew
rlabel metal1 s 27216 15259 27216 15259 4 vdd
port 513 nsew
rlabel metal1 s 25968 13180 25968 13180 4 vdd
port 513 nsew
rlabel metal1 s 25200 13180 25200 13180 4 vdd
port 513 nsew
rlabel metal1 s 25200 13679 25200 13679 4 vdd
port 513 nsew
rlabel metal1 s 27216 14760 27216 14760 4 vdd
port 513 nsew
rlabel metal1 s 26448 14760 26448 14760 4 vdd
port 513 nsew
rlabel metal1 s 27216 12889 27216 12889 4 vdd
port 513 nsew
rlabel metal1 s 27216 15550 27216 15550 4 vdd
port 513 nsew
rlabel metal1 s 27216 13970 27216 13970 4 vdd
port 513 nsew
rlabel metal1 s 25968 13970 25968 13970 4 vdd
port 513 nsew
rlabel metal1 s 26448 13180 26448 13180 4 vdd
port 513 nsew
rlabel metal1 s 25200 12889 25200 12889 4 vdd
port 513 nsew
rlabel metal1 s 25968 14469 25968 14469 4 vdd
port 513 nsew
rlabel metal1 s 27216 13679 27216 13679 4 vdd
port 513 nsew
rlabel metal1 s 26448 13970 26448 13970 4 vdd
port 513 nsew
rlabel metal1 s 25968 12889 25968 12889 4 vdd
port 513 nsew
rlabel metal1 s 25200 13970 25200 13970 4 vdd
port 513 nsew
rlabel metal1 s 26448 15550 26448 15550 4 vdd
port 513 nsew
rlabel metal1 s 25200 14760 25200 14760 4 vdd
port 513 nsew
rlabel metal1 s 25968 15259 25968 15259 4 vdd
port 513 nsew
rlabel metal1 s 26448 14469 26448 14469 4 vdd
port 513 nsew
rlabel metal1 s 26448 13679 26448 13679 4 vdd
port 513 nsew
rlabel metal1 s 25968 15550 25968 15550 4 vdd
port 513 nsew
rlabel metal1 s 25200 14469 25200 14469 4 vdd
port 513 nsew
rlabel metal1 s 25968 14760 25968 14760 4 vdd
port 513 nsew
rlabel metal1 s 25200 15259 25200 15259 4 vdd
port 513 nsew
rlabel metal1 s 27216 13180 27216 13180 4 vdd
port 513 nsew
rlabel metal1 s 25200 15550 25200 15550 4 vdd
port 513 nsew
rlabel metal1 s 28944 13970 28944 13970 4 vdd
port 513 nsew
rlabel metal1 s 29712 13180 29712 13180 4 vdd
port 513 nsew
rlabel metal1 s 27696 12889 27696 12889 4 vdd
port 513 nsew
rlabel metal1 s 28464 14760 28464 14760 4 vdd
port 513 nsew
rlabel metal1 s 28464 14469 28464 14469 4 vdd
port 513 nsew
rlabel metal1 s 28464 12889 28464 12889 4 vdd
port 513 nsew
rlabel metal1 s 28464 15259 28464 15259 4 vdd
port 513 nsew
rlabel metal1 s 29712 12889 29712 12889 4 vdd
port 513 nsew
rlabel metal1 s 28944 12889 28944 12889 4 vdd
port 513 nsew
rlabel metal1 s 27696 13180 27696 13180 4 vdd
port 513 nsew
rlabel metal1 s 28944 13679 28944 13679 4 vdd
port 513 nsew
rlabel metal1 s 29712 15550 29712 15550 4 vdd
port 513 nsew
rlabel metal1 s 29712 14469 29712 14469 4 vdd
port 513 nsew
rlabel metal1 s 27696 15259 27696 15259 4 vdd
port 513 nsew
rlabel metal1 s 28464 13180 28464 13180 4 vdd
port 513 nsew
rlabel metal1 s 28944 15550 28944 15550 4 vdd
port 513 nsew
rlabel metal1 s 28944 15259 28944 15259 4 vdd
port 513 nsew
rlabel metal1 s 27696 13679 27696 13679 4 vdd
port 513 nsew
rlabel metal1 s 28944 14469 28944 14469 4 vdd
port 513 nsew
rlabel metal1 s 29712 13970 29712 13970 4 vdd
port 513 nsew
rlabel metal1 s 27696 14760 27696 14760 4 vdd
port 513 nsew
rlabel metal1 s 28944 14760 28944 14760 4 vdd
port 513 nsew
rlabel metal1 s 27696 15550 27696 15550 4 vdd
port 513 nsew
rlabel metal1 s 29712 15259 29712 15259 4 vdd
port 513 nsew
rlabel metal1 s 28464 13970 28464 13970 4 vdd
port 513 nsew
rlabel metal1 s 28464 15550 28464 15550 4 vdd
port 513 nsew
rlabel metal1 s 27696 13970 27696 13970 4 vdd
port 513 nsew
rlabel metal1 s 27696 14469 27696 14469 4 vdd
port 513 nsew
rlabel metal1 s 29712 13679 29712 13679 4 vdd
port 513 nsew
rlabel metal1 s 28464 13679 28464 13679 4 vdd
port 513 nsew
rlabel metal1 s 29712 14760 29712 14760 4 vdd
port 513 nsew
rlabel metal1 s 28944 13180 28944 13180 4 vdd
port 513 nsew
rlabel metal1 s 28464 11600 28464 11600 4 vdd
port 513 nsew
rlabel metal1 s 29712 12099 29712 12099 4 vdd
port 513 nsew
rlabel metal1 s 28944 11309 28944 11309 4 vdd
port 513 nsew
rlabel metal1 s 29712 11309 29712 11309 4 vdd
port 513 nsew
rlabel metal1 s 28944 12390 28944 12390 4 vdd
port 513 nsew
rlabel metal1 s 29712 11600 29712 11600 4 vdd
port 513 nsew
rlabel metal1 s 28944 12099 28944 12099 4 vdd
port 513 nsew
rlabel metal1 s 27696 12099 27696 12099 4 vdd
port 513 nsew
rlabel metal1 s 28464 10519 28464 10519 4 vdd
port 513 nsew
rlabel metal1 s 27696 10519 27696 10519 4 vdd
port 513 nsew
rlabel metal1 s 29712 10810 29712 10810 4 vdd
port 513 nsew
rlabel metal1 s 28464 10020 28464 10020 4 vdd
port 513 nsew
rlabel metal1 s 29712 12390 29712 12390 4 vdd
port 513 nsew
rlabel metal1 s 27696 10020 27696 10020 4 vdd
port 513 nsew
rlabel metal1 s 28464 11309 28464 11309 4 vdd
port 513 nsew
rlabel metal1 s 27696 9729 27696 9729 4 vdd
port 513 nsew
rlabel metal1 s 28944 11600 28944 11600 4 vdd
port 513 nsew
rlabel metal1 s 29712 10020 29712 10020 4 vdd
port 513 nsew
rlabel metal1 s 28944 10519 28944 10519 4 vdd
port 513 nsew
rlabel metal1 s 28464 10810 28464 10810 4 vdd
port 513 nsew
rlabel metal1 s 27696 11309 27696 11309 4 vdd
port 513 nsew
rlabel metal1 s 28464 12390 28464 12390 4 vdd
port 513 nsew
rlabel metal1 s 29712 10519 29712 10519 4 vdd
port 513 nsew
rlabel metal1 s 27696 11600 27696 11600 4 vdd
port 513 nsew
rlabel metal1 s 27696 10810 27696 10810 4 vdd
port 513 nsew
rlabel metal1 s 29712 9729 29712 9729 4 vdd
port 513 nsew
rlabel metal1 s 27696 12390 27696 12390 4 vdd
port 513 nsew
rlabel metal1 s 28464 12099 28464 12099 4 vdd
port 513 nsew
rlabel metal1 s 28944 9729 28944 9729 4 vdd
port 513 nsew
rlabel metal1 s 28944 10810 28944 10810 4 vdd
port 513 nsew
rlabel metal1 s 28944 10020 28944 10020 4 vdd
port 513 nsew
rlabel metal1 s 28464 9729 28464 9729 4 vdd
port 513 nsew
rlabel metal1 s 25968 11600 25968 11600 4 vdd
port 513 nsew
rlabel metal1 s 25968 11309 25968 11309 4 vdd
port 513 nsew
rlabel metal1 s 27216 10810 27216 10810 4 vdd
port 513 nsew
rlabel metal1 s 25968 10519 25968 10519 4 vdd
port 513 nsew
rlabel metal1 s 25200 12099 25200 12099 4 vdd
port 513 nsew
rlabel metal1 s 25200 9729 25200 9729 4 vdd
port 513 nsew
rlabel metal1 s 26448 10519 26448 10519 4 vdd
port 513 nsew
rlabel metal1 s 25968 10020 25968 10020 4 vdd
port 513 nsew
rlabel metal1 s 25968 10810 25968 10810 4 vdd
port 513 nsew
rlabel metal1 s 26448 11309 26448 11309 4 vdd
port 513 nsew
rlabel metal1 s 25200 11600 25200 11600 4 vdd
port 513 nsew
rlabel metal1 s 25200 11309 25200 11309 4 vdd
port 513 nsew
rlabel metal1 s 27216 11309 27216 11309 4 vdd
port 513 nsew
rlabel metal1 s 26448 9729 26448 9729 4 vdd
port 513 nsew
rlabel metal1 s 27216 9729 27216 9729 4 vdd
port 513 nsew
rlabel metal1 s 27216 10020 27216 10020 4 vdd
port 513 nsew
rlabel metal1 s 25968 9729 25968 9729 4 vdd
port 513 nsew
rlabel metal1 s 27216 12390 27216 12390 4 vdd
port 513 nsew
rlabel metal1 s 25200 10020 25200 10020 4 vdd
port 513 nsew
rlabel metal1 s 25200 10810 25200 10810 4 vdd
port 513 nsew
rlabel metal1 s 27216 12099 27216 12099 4 vdd
port 513 nsew
rlabel metal1 s 26448 11600 26448 11600 4 vdd
port 513 nsew
rlabel metal1 s 25968 12099 25968 12099 4 vdd
port 513 nsew
rlabel metal1 s 25200 12390 25200 12390 4 vdd
port 513 nsew
rlabel metal1 s 26448 12390 26448 12390 4 vdd
port 513 nsew
rlabel metal1 s 26448 10020 26448 10020 4 vdd
port 513 nsew
rlabel metal1 s 27216 10519 27216 10519 4 vdd
port 513 nsew
rlabel metal1 s 27216 11600 27216 11600 4 vdd
port 513 nsew
rlabel metal1 s 25200 10519 25200 10519 4 vdd
port 513 nsew
rlabel metal1 s 26448 12099 26448 12099 4 vdd
port 513 nsew
rlabel metal1 s 25968 12390 25968 12390 4 vdd
port 513 nsew
rlabel metal1 s 26448 10810 26448 10810 4 vdd
port 513 nsew
rlabel metal1 s 26448 8939 26448 8939 4 vdd
port 513 nsew
rlabel metal1 s 27216 7359 27216 7359 4 vdd
port 513 nsew
rlabel metal1 s 25968 7359 25968 7359 4 vdd
port 513 nsew
rlabel metal1 s 27216 8939 27216 8939 4 vdd
port 513 nsew
rlabel metal1 s 25200 8149 25200 8149 4 vdd
port 513 nsew
rlabel metal1 s 27216 6860 27216 6860 4 vdd
port 513 nsew
rlabel metal1 s 25200 8939 25200 8939 4 vdd
port 513 nsew
rlabel metal1 s 25968 6569 25968 6569 4 vdd
port 513 nsew
rlabel metal1 s 26448 6860 26448 6860 4 vdd
port 513 nsew
rlabel metal1 s 25200 9230 25200 9230 4 vdd
port 513 nsew
rlabel metal1 s 25968 7650 25968 7650 4 vdd
port 513 nsew
rlabel metal1 s 26448 6569 26448 6569 4 vdd
port 513 nsew
rlabel metal1 s 25968 8440 25968 8440 4 vdd
port 513 nsew
rlabel metal1 s 27216 7650 27216 7650 4 vdd
port 513 nsew
rlabel metal1 s 26448 8149 26448 8149 4 vdd
port 513 nsew
rlabel metal1 s 25968 8149 25968 8149 4 vdd
port 513 nsew
rlabel metal1 s 26448 9230 26448 9230 4 vdd
port 513 nsew
rlabel metal1 s 25200 8440 25200 8440 4 vdd
port 513 nsew
rlabel metal1 s 25200 6569 25200 6569 4 vdd
port 513 nsew
rlabel metal1 s 26448 7359 26448 7359 4 vdd
port 513 nsew
rlabel metal1 s 27216 8149 27216 8149 4 vdd
port 513 nsew
rlabel metal1 s 25968 8939 25968 8939 4 vdd
port 513 nsew
rlabel metal1 s 27216 8440 27216 8440 4 vdd
port 513 nsew
rlabel metal1 s 25968 6860 25968 6860 4 vdd
port 513 nsew
rlabel metal1 s 25200 7650 25200 7650 4 vdd
port 513 nsew
rlabel metal1 s 27216 6569 27216 6569 4 vdd
port 513 nsew
rlabel metal1 s 25968 9230 25968 9230 4 vdd
port 513 nsew
rlabel metal1 s 26448 8440 26448 8440 4 vdd
port 513 nsew
rlabel metal1 s 27216 9230 27216 9230 4 vdd
port 513 nsew
rlabel metal1 s 26448 7650 26448 7650 4 vdd
port 513 nsew
rlabel metal1 s 25200 7359 25200 7359 4 vdd
port 513 nsew
rlabel metal1 s 25200 6860 25200 6860 4 vdd
port 513 nsew
rlabel metal1 s 29712 8149 29712 8149 4 vdd
port 513 nsew
rlabel metal1 s 28464 8440 28464 8440 4 vdd
port 513 nsew
rlabel metal1 s 28464 8149 28464 8149 4 vdd
port 513 nsew
rlabel metal1 s 29712 7359 29712 7359 4 vdd
port 513 nsew
rlabel metal1 s 28944 8939 28944 8939 4 vdd
port 513 nsew
rlabel metal1 s 29712 6860 29712 6860 4 vdd
port 513 nsew
rlabel metal1 s 29712 8440 29712 8440 4 vdd
port 513 nsew
rlabel metal1 s 27696 6569 27696 6569 4 vdd
port 513 nsew
rlabel metal1 s 27696 7650 27696 7650 4 vdd
port 513 nsew
rlabel metal1 s 27696 8440 27696 8440 4 vdd
port 513 nsew
rlabel metal1 s 27696 6860 27696 6860 4 vdd
port 513 nsew
rlabel metal1 s 29712 9230 29712 9230 4 vdd
port 513 nsew
rlabel metal1 s 28464 7359 28464 7359 4 vdd
port 513 nsew
rlabel metal1 s 27696 9230 27696 9230 4 vdd
port 513 nsew
rlabel metal1 s 27696 7359 27696 7359 4 vdd
port 513 nsew
rlabel metal1 s 29712 7650 29712 7650 4 vdd
port 513 nsew
rlabel metal1 s 27696 8149 27696 8149 4 vdd
port 513 nsew
rlabel metal1 s 27696 8939 27696 8939 4 vdd
port 513 nsew
rlabel metal1 s 28944 6569 28944 6569 4 vdd
port 513 nsew
rlabel metal1 s 28464 6860 28464 6860 4 vdd
port 513 nsew
rlabel metal1 s 29712 6569 29712 6569 4 vdd
port 513 nsew
rlabel metal1 s 28464 9230 28464 9230 4 vdd
port 513 nsew
rlabel metal1 s 28944 9230 28944 9230 4 vdd
port 513 nsew
rlabel metal1 s 28464 8939 28464 8939 4 vdd
port 513 nsew
rlabel metal1 s 28464 6569 28464 6569 4 vdd
port 513 nsew
rlabel metal1 s 29712 8939 29712 8939 4 vdd
port 513 nsew
rlabel metal1 s 28944 6860 28944 6860 4 vdd
port 513 nsew
rlabel metal1 s 28944 7650 28944 7650 4 vdd
port 513 nsew
rlabel metal1 s 28464 7650 28464 7650 4 vdd
port 513 nsew
rlabel metal1 s 28944 8440 28944 8440 4 vdd
port 513 nsew
rlabel metal1 s 28944 7359 28944 7359 4 vdd
port 513 nsew
rlabel metal1 s 28944 8149 28944 8149 4 vdd
port 513 nsew
rlabel metal1 s 24720 11600 24720 11600 4 vdd
port 513 nsew
rlabel metal1 s 24720 10519 24720 10519 4 vdd
port 513 nsew
rlabel metal1 s 24720 12099 24720 12099 4 vdd
port 513 nsew
rlabel metal1 s 23472 11600 23472 11600 4 vdd
port 513 nsew
rlabel metal1 s 23472 10810 23472 10810 4 vdd
port 513 nsew
rlabel metal1 s 22704 9729 22704 9729 4 vdd
port 513 nsew
rlabel metal1 s 23472 12390 23472 12390 4 vdd
port 513 nsew
rlabel metal1 s 24720 10020 24720 10020 4 vdd
port 513 nsew
rlabel metal1 s 23472 11309 23472 11309 4 vdd
port 513 nsew
rlabel metal1 s 23952 12099 23952 12099 4 vdd
port 513 nsew
rlabel metal1 s 23952 9729 23952 9729 4 vdd
port 513 nsew
rlabel metal1 s 24720 11309 24720 11309 4 vdd
port 513 nsew
rlabel metal1 s 24720 12390 24720 12390 4 vdd
port 513 nsew
rlabel metal1 s 22704 11600 22704 11600 4 vdd
port 513 nsew
rlabel metal1 s 22704 12390 22704 12390 4 vdd
port 513 nsew
rlabel metal1 s 23952 10020 23952 10020 4 vdd
port 513 nsew
rlabel metal1 s 23952 11309 23952 11309 4 vdd
port 513 nsew
rlabel metal1 s 24720 10810 24720 10810 4 vdd
port 513 nsew
rlabel metal1 s 23952 11600 23952 11600 4 vdd
port 513 nsew
rlabel metal1 s 23472 10519 23472 10519 4 vdd
port 513 nsew
rlabel metal1 s 23472 12099 23472 12099 4 vdd
port 513 nsew
rlabel metal1 s 23472 10020 23472 10020 4 vdd
port 513 nsew
rlabel metal1 s 22704 12099 22704 12099 4 vdd
port 513 nsew
rlabel metal1 s 24720 9729 24720 9729 4 vdd
port 513 nsew
rlabel metal1 s 23952 10519 23952 10519 4 vdd
port 513 nsew
rlabel metal1 s 22704 10519 22704 10519 4 vdd
port 513 nsew
rlabel metal1 s 22704 10020 22704 10020 4 vdd
port 513 nsew
rlabel metal1 s 23952 10810 23952 10810 4 vdd
port 513 nsew
rlabel metal1 s 23952 12390 23952 12390 4 vdd
port 513 nsew
rlabel metal1 s 23472 9729 23472 9729 4 vdd
port 513 nsew
rlabel metal1 s 22704 10810 22704 10810 4 vdd
port 513 nsew
rlabel metal1 s 22704 11309 22704 11309 4 vdd
port 513 nsew
rlabel metal1 s 20208 11309 20208 11309 4 vdd
port 513 nsew
rlabel metal1 s 22224 10810 22224 10810 4 vdd
port 513 nsew
rlabel metal1 s 20208 12099 20208 12099 4 vdd
port 513 nsew
rlabel metal1 s 21456 10020 21456 10020 4 vdd
port 513 nsew
rlabel metal1 s 20208 10810 20208 10810 4 vdd
port 513 nsew
rlabel metal1 s 20976 12099 20976 12099 4 vdd
port 513 nsew
rlabel metal1 s 20208 10519 20208 10519 4 vdd
port 513 nsew
rlabel metal1 s 22224 10519 22224 10519 4 vdd
port 513 nsew
rlabel metal1 s 20976 12390 20976 12390 4 vdd
port 513 nsew
rlabel metal1 s 20976 11309 20976 11309 4 vdd
port 513 nsew
rlabel metal1 s 21456 12099 21456 12099 4 vdd
port 513 nsew
rlabel metal1 s 21456 11309 21456 11309 4 vdd
port 513 nsew
rlabel metal1 s 20976 9729 20976 9729 4 vdd
port 513 nsew
rlabel metal1 s 20208 12390 20208 12390 4 vdd
port 513 nsew
rlabel metal1 s 22224 11309 22224 11309 4 vdd
port 513 nsew
rlabel metal1 s 21456 12390 21456 12390 4 vdd
port 513 nsew
rlabel metal1 s 22224 12390 22224 12390 4 vdd
port 513 nsew
rlabel metal1 s 20976 10810 20976 10810 4 vdd
port 513 nsew
rlabel metal1 s 21456 11600 21456 11600 4 vdd
port 513 nsew
rlabel metal1 s 20208 10020 20208 10020 4 vdd
port 513 nsew
rlabel metal1 s 20208 9729 20208 9729 4 vdd
port 513 nsew
rlabel metal1 s 20208 11600 20208 11600 4 vdd
port 513 nsew
rlabel metal1 s 21456 10810 21456 10810 4 vdd
port 513 nsew
rlabel metal1 s 22224 10020 22224 10020 4 vdd
port 513 nsew
rlabel metal1 s 22224 9729 22224 9729 4 vdd
port 513 nsew
rlabel metal1 s 22224 11600 22224 11600 4 vdd
port 513 nsew
rlabel metal1 s 20976 10519 20976 10519 4 vdd
port 513 nsew
rlabel metal1 s 22224 12099 22224 12099 4 vdd
port 513 nsew
rlabel metal1 s 21456 10519 21456 10519 4 vdd
port 513 nsew
rlabel metal1 s 20976 10020 20976 10020 4 vdd
port 513 nsew
rlabel metal1 s 21456 9729 21456 9729 4 vdd
port 513 nsew
rlabel metal1 s 20976 11600 20976 11600 4 vdd
port 513 nsew
rlabel metal1 s 21456 6569 21456 6569 4 vdd
port 513 nsew
rlabel metal1 s 20976 8149 20976 8149 4 vdd
port 513 nsew
rlabel metal1 s 20208 7359 20208 7359 4 vdd
port 513 nsew
rlabel metal1 s 21456 6860 21456 6860 4 vdd
port 513 nsew
rlabel metal1 s 22224 8149 22224 8149 4 vdd
port 513 nsew
rlabel metal1 s 21456 7650 21456 7650 4 vdd
port 513 nsew
rlabel metal1 s 20976 6860 20976 6860 4 vdd
port 513 nsew
rlabel metal1 s 20976 7359 20976 7359 4 vdd
port 513 nsew
rlabel metal1 s 21456 8440 21456 8440 4 vdd
port 513 nsew
rlabel metal1 s 20208 8149 20208 8149 4 vdd
port 513 nsew
rlabel metal1 s 22224 9230 22224 9230 4 vdd
port 513 nsew
rlabel metal1 s 20976 7650 20976 7650 4 vdd
port 513 nsew
rlabel metal1 s 22224 7650 22224 7650 4 vdd
port 513 nsew
rlabel metal1 s 20976 8939 20976 8939 4 vdd
port 513 nsew
rlabel metal1 s 21456 8939 21456 8939 4 vdd
port 513 nsew
rlabel metal1 s 21456 7359 21456 7359 4 vdd
port 513 nsew
rlabel metal1 s 20976 6569 20976 6569 4 vdd
port 513 nsew
rlabel metal1 s 20208 6569 20208 6569 4 vdd
port 513 nsew
rlabel metal1 s 20208 8939 20208 8939 4 vdd
port 513 nsew
rlabel metal1 s 22224 7359 22224 7359 4 vdd
port 513 nsew
rlabel metal1 s 20208 7650 20208 7650 4 vdd
port 513 nsew
rlabel metal1 s 20208 9230 20208 9230 4 vdd
port 513 nsew
rlabel metal1 s 22224 8939 22224 8939 4 vdd
port 513 nsew
rlabel metal1 s 22224 6569 22224 6569 4 vdd
port 513 nsew
rlabel metal1 s 22224 8440 22224 8440 4 vdd
port 513 nsew
rlabel metal1 s 20976 8440 20976 8440 4 vdd
port 513 nsew
rlabel metal1 s 20208 6860 20208 6860 4 vdd
port 513 nsew
rlabel metal1 s 21456 9230 21456 9230 4 vdd
port 513 nsew
rlabel metal1 s 20208 8440 20208 8440 4 vdd
port 513 nsew
rlabel metal1 s 22224 6860 22224 6860 4 vdd
port 513 nsew
rlabel metal1 s 20976 9230 20976 9230 4 vdd
port 513 nsew
rlabel metal1 s 21456 8149 21456 8149 4 vdd
port 513 nsew
rlabel metal1 s 24720 7650 24720 7650 4 vdd
port 513 nsew
rlabel metal1 s 23952 6569 23952 6569 4 vdd
port 513 nsew
rlabel metal1 s 23472 8149 23472 8149 4 vdd
port 513 nsew
rlabel metal1 s 23952 8939 23952 8939 4 vdd
port 513 nsew
rlabel metal1 s 24720 8440 24720 8440 4 vdd
port 513 nsew
rlabel metal1 s 22704 7650 22704 7650 4 vdd
port 513 nsew
rlabel metal1 s 22704 6860 22704 6860 4 vdd
port 513 nsew
rlabel metal1 s 24720 6569 24720 6569 4 vdd
port 513 nsew
rlabel metal1 s 23472 6860 23472 6860 4 vdd
port 513 nsew
rlabel metal1 s 24720 7359 24720 7359 4 vdd
port 513 nsew
rlabel metal1 s 22704 8149 22704 8149 4 vdd
port 513 nsew
rlabel metal1 s 22704 8939 22704 8939 4 vdd
port 513 nsew
rlabel metal1 s 22704 7359 22704 7359 4 vdd
port 513 nsew
rlabel metal1 s 23472 7650 23472 7650 4 vdd
port 513 nsew
rlabel metal1 s 22704 6569 22704 6569 4 vdd
port 513 nsew
rlabel metal1 s 23952 8149 23952 8149 4 vdd
port 513 nsew
rlabel metal1 s 24720 8149 24720 8149 4 vdd
port 513 nsew
rlabel metal1 s 23952 8440 23952 8440 4 vdd
port 513 nsew
rlabel metal1 s 23472 8939 23472 8939 4 vdd
port 513 nsew
rlabel metal1 s 23952 9230 23952 9230 4 vdd
port 513 nsew
rlabel metal1 s 23472 8440 23472 8440 4 vdd
port 513 nsew
rlabel metal1 s 24720 9230 24720 9230 4 vdd
port 513 nsew
rlabel metal1 s 23952 6860 23952 6860 4 vdd
port 513 nsew
rlabel metal1 s 23952 7359 23952 7359 4 vdd
port 513 nsew
rlabel metal1 s 22704 9230 22704 9230 4 vdd
port 513 nsew
rlabel metal1 s 23472 7359 23472 7359 4 vdd
port 513 nsew
rlabel metal1 s 24720 6860 24720 6860 4 vdd
port 513 nsew
rlabel metal1 s 23472 9230 23472 9230 4 vdd
port 513 nsew
rlabel metal1 s 22704 8440 22704 8440 4 vdd
port 513 nsew
rlabel metal1 s 23952 7650 23952 7650 4 vdd
port 513 nsew
rlabel metal1 s 23472 6569 23472 6569 4 vdd
port 513 nsew
rlabel metal1 s 24720 8939 24720 8939 4 vdd
port 513 nsew
rlabel metal1 s 22704 3409 22704 3409 4 vdd
port 513 nsew
rlabel metal1 s 23472 5280 23472 5280 4 vdd
port 513 nsew
rlabel metal1 s 23952 4490 23952 4490 4 vdd
port 513 nsew
rlabel metal1 s 23472 4989 23472 4989 4 vdd
port 513 nsew
rlabel metal1 s 24720 5779 24720 5779 4 vdd
port 513 nsew
rlabel metal1 s 23952 3700 23952 3700 4 vdd
port 513 nsew
rlabel metal1 s 22704 5280 22704 5280 4 vdd
port 513 nsew
rlabel metal1 s 24720 4490 24720 4490 4 vdd
port 513 nsew
rlabel metal1 s 23952 5280 23952 5280 4 vdd
port 513 nsew
rlabel metal1 s 23472 4490 23472 4490 4 vdd
port 513 nsew
rlabel metal1 s 22704 3700 22704 3700 4 vdd
port 513 nsew
rlabel metal1 s 23952 6070 23952 6070 4 vdd
port 513 nsew
rlabel metal1 s 23472 3700 23472 3700 4 vdd
port 513 nsew
rlabel metal1 s 23952 4989 23952 4989 4 vdd
port 513 nsew
rlabel metal1 s 22704 6070 22704 6070 4 vdd
port 513 nsew
rlabel metal1 s 23952 5779 23952 5779 4 vdd
port 513 nsew
rlabel metal1 s 22704 5779 22704 5779 4 vdd
port 513 nsew
rlabel metal1 s 24720 6070 24720 6070 4 vdd
port 513 nsew
rlabel metal1 s 23472 4199 23472 4199 4 vdd
port 513 nsew
rlabel metal1 s 24720 3700 24720 3700 4 vdd
port 513 nsew
rlabel metal1 s 23952 3409 23952 3409 4 vdd
port 513 nsew
rlabel metal1 s 24720 3409 24720 3409 4 vdd
port 513 nsew
rlabel metal1 s 24720 4199 24720 4199 4 vdd
port 513 nsew
rlabel metal1 s 23472 6070 23472 6070 4 vdd
port 513 nsew
rlabel metal1 s 24720 4989 24720 4989 4 vdd
port 513 nsew
rlabel metal1 s 23472 3409 23472 3409 4 vdd
port 513 nsew
rlabel metal1 s 23952 4199 23952 4199 4 vdd
port 513 nsew
rlabel metal1 s 22704 4490 22704 4490 4 vdd
port 513 nsew
rlabel metal1 s 22704 4199 22704 4199 4 vdd
port 513 nsew
rlabel metal1 s 24720 5280 24720 5280 4 vdd
port 513 nsew
rlabel metal1 s 23472 5779 23472 5779 4 vdd
port 513 nsew
rlabel metal1 s 22704 4989 22704 4989 4 vdd
port 513 nsew
rlabel metal1 s 21456 3409 21456 3409 4 vdd
port 513 nsew
rlabel metal1 s 20976 4199 20976 4199 4 vdd
port 513 nsew
rlabel metal1 s 21456 5280 21456 5280 4 vdd
port 513 nsew
rlabel metal1 s 20976 5779 20976 5779 4 vdd
port 513 nsew
rlabel metal1 s 20976 4490 20976 4490 4 vdd
port 513 nsew
rlabel metal1 s 20208 4490 20208 4490 4 vdd
port 513 nsew
rlabel metal1 s 20976 5280 20976 5280 4 vdd
port 513 nsew
rlabel metal1 s 21456 6070 21456 6070 4 vdd
port 513 nsew
rlabel metal1 s 20976 3700 20976 3700 4 vdd
port 513 nsew
rlabel metal1 s 20976 4989 20976 4989 4 vdd
port 513 nsew
rlabel metal1 s 22224 4490 22224 4490 4 vdd
port 513 nsew
rlabel metal1 s 22224 5779 22224 5779 4 vdd
port 513 nsew
rlabel metal1 s 20208 3409 20208 3409 4 vdd
port 513 nsew
rlabel metal1 s 20208 4199 20208 4199 4 vdd
port 513 nsew
rlabel metal1 s 20976 3409 20976 3409 4 vdd
port 513 nsew
rlabel metal1 s 21456 3700 21456 3700 4 vdd
port 513 nsew
rlabel metal1 s 21456 5779 21456 5779 4 vdd
port 513 nsew
rlabel metal1 s 21456 4989 21456 4989 4 vdd
port 513 nsew
rlabel metal1 s 20208 5779 20208 5779 4 vdd
port 513 nsew
rlabel metal1 s 20208 6070 20208 6070 4 vdd
port 513 nsew
rlabel metal1 s 21456 4199 21456 4199 4 vdd
port 513 nsew
rlabel metal1 s 22224 3409 22224 3409 4 vdd
port 513 nsew
rlabel metal1 s 22224 4199 22224 4199 4 vdd
port 513 nsew
rlabel metal1 s 22224 4989 22224 4989 4 vdd
port 513 nsew
rlabel metal1 s 20208 4989 20208 4989 4 vdd
port 513 nsew
rlabel metal1 s 20208 5280 20208 5280 4 vdd
port 513 nsew
rlabel metal1 s 22224 3700 22224 3700 4 vdd
port 513 nsew
rlabel metal1 s 22224 6070 22224 6070 4 vdd
port 513 nsew
rlabel metal1 s 21456 4490 21456 4490 4 vdd
port 513 nsew
rlabel metal1 s 20976 6070 20976 6070 4 vdd
port 513 nsew
rlabel metal1 s 22224 5280 22224 5280 4 vdd
port 513 nsew
rlabel metal1 s 20208 3700 20208 3700 4 vdd
port 513 nsew
rlabel metal1 s 20208 2619 20208 2619 4 vdd
port 513 nsew
rlabel metal1 s 21456 1330 21456 1330 4 vdd
port 513 nsew
rlabel metal1 s 21456 540 21456 540 4 vdd
port 513 nsew
rlabel metal1 s 20208 2910 20208 2910 4 vdd
port 513 nsew
rlabel metal1 s 22224 1039 22224 1039 4 vdd
port 513 nsew
rlabel metal1 s 22224 1330 22224 1330 4 vdd
port 513 nsew
rlabel metal1 s 21456 2619 21456 2619 4 vdd
port 513 nsew
rlabel metal1 s 20208 540 20208 540 4 vdd
port 513 nsew
rlabel metal1 s 20976 2120 20976 2120 4 vdd
port 513 nsew
rlabel metal1 s 22224 540 22224 540 4 vdd
port 513 nsew
rlabel metal1 s 20208 1829 20208 1829 4 vdd
port 513 nsew
rlabel metal1 s 22224 2619 22224 2619 4 vdd
port 513 nsew
rlabel metal1 s 20208 2120 20208 2120 4 vdd
port 513 nsew
rlabel metal1 s 20976 2910 20976 2910 4 vdd
port 513 nsew
rlabel metal1 s 21456 2120 21456 2120 4 vdd
port 513 nsew
rlabel metal1 s 20976 2619 20976 2619 4 vdd
port 513 nsew
rlabel metal1 s 22224 1829 22224 1829 4 vdd
port 513 nsew
rlabel metal1 s 22224 249 22224 249 4 vdd
port 513 nsew
rlabel metal1 s 21456 1829 21456 1829 4 vdd
port 513 nsew
rlabel metal1 s 20208 1330 20208 1330 4 vdd
port 513 nsew
rlabel metal1 s 20976 1039 20976 1039 4 vdd
port 513 nsew
rlabel metal1 s 21456 1039 21456 1039 4 vdd
port 513 nsew
rlabel metal1 s 21456 2910 21456 2910 4 vdd
port 513 nsew
rlabel metal1 s 21456 249 21456 249 4 vdd
port 513 nsew
rlabel metal1 s 20208 1039 20208 1039 4 vdd
port 513 nsew
rlabel metal1 s 22224 2910 22224 2910 4 vdd
port 513 nsew
rlabel metal1 s 20976 249 20976 249 4 vdd
port 513 nsew
rlabel metal1 s 20208 249 20208 249 4 vdd
port 513 nsew
rlabel metal1 s 20976 540 20976 540 4 vdd
port 513 nsew
rlabel metal1 s 22224 2120 22224 2120 4 vdd
port 513 nsew
rlabel metal1 s 20976 1330 20976 1330 4 vdd
port 513 nsew
rlabel metal1 s 20976 1829 20976 1829 4 vdd
port 513 nsew
rlabel metal1 s 23472 1829 23472 1829 4 vdd
port 513 nsew
rlabel metal1 s 23472 1039 23472 1039 4 vdd
port 513 nsew
rlabel metal1 s 22704 1330 22704 1330 4 vdd
port 513 nsew
rlabel metal1 s 23952 1039 23952 1039 4 vdd
port 513 nsew
rlabel metal1 s 24720 2619 24720 2619 4 vdd
port 513 nsew
rlabel metal1 s 24720 1829 24720 1829 4 vdd
port 513 nsew
rlabel metal1 s 23472 540 23472 540 4 vdd
port 513 nsew
rlabel metal1 s 22704 1039 22704 1039 4 vdd
port 513 nsew
rlabel metal1 s 22704 2910 22704 2910 4 vdd
port 513 nsew
rlabel metal1 s 22704 249 22704 249 4 vdd
port 513 nsew
rlabel metal1 s 24720 1330 24720 1330 4 vdd
port 513 nsew
rlabel metal1 s 23472 2120 23472 2120 4 vdd
port 513 nsew
rlabel metal1 s 24720 2120 24720 2120 4 vdd
port 513 nsew
rlabel metal1 s 22704 2120 22704 2120 4 vdd
port 513 nsew
rlabel metal1 s 22704 540 22704 540 4 vdd
port 513 nsew
rlabel metal1 s 23952 2120 23952 2120 4 vdd
port 513 nsew
rlabel metal1 s 22704 2619 22704 2619 4 vdd
port 513 nsew
rlabel metal1 s 23952 540 23952 540 4 vdd
port 513 nsew
rlabel metal1 s 23952 2910 23952 2910 4 vdd
port 513 nsew
rlabel metal1 s 23952 1330 23952 1330 4 vdd
port 513 nsew
rlabel metal1 s 24720 1039 24720 1039 4 vdd
port 513 nsew
rlabel metal1 s 23952 249 23952 249 4 vdd
port 513 nsew
rlabel metal1 s 23472 1330 23472 1330 4 vdd
port 513 nsew
rlabel metal1 s 23952 1829 23952 1829 4 vdd
port 513 nsew
rlabel metal1 s 22704 1829 22704 1829 4 vdd
port 513 nsew
rlabel metal1 s 24720 540 24720 540 4 vdd
port 513 nsew
rlabel metal1 s 23472 2619 23472 2619 4 vdd
port 513 nsew
rlabel metal1 s 24720 2910 24720 2910 4 vdd
port 513 nsew
rlabel metal1 s 23952 2619 23952 2619 4 vdd
port 513 nsew
rlabel metal1 s 23472 2910 23472 2910 4 vdd
port 513 nsew
rlabel metal1 s 23472 249 23472 249 4 vdd
port 513 nsew
rlabel metal1 s 24720 249 24720 249 4 vdd
port 513 nsew
rlabel metal1 s 28944 4490 28944 4490 4 vdd
port 513 nsew
rlabel metal1 s 27696 5280 27696 5280 4 vdd
port 513 nsew
rlabel metal1 s 27696 3409 27696 3409 4 vdd
port 513 nsew
rlabel metal1 s 28464 6070 28464 6070 4 vdd
port 513 nsew
rlabel metal1 s 27696 4989 27696 4989 4 vdd
port 513 nsew
rlabel metal1 s 28944 3409 28944 3409 4 vdd
port 513 nsew
rlabel metal1 s 28944 3700 28944 3700 4 vdd
port 513 nsew
rlabel metal1 s 28464 5779 28464 5779 4 vdd
port 513 nsew
rlabel metal1 s 29712 3409 29712 3409 4 vdd
port 513 nsew
rlabel metal1 s 29712 5280 29712 5280 4 vdd
port 513 nsew
rlabel metal1 s 28944 4199 28944 4199 4 vdd
port 513 nsew
rlabel metal1 s 28464 4199 28464 4199 4 vdd
port 513 nsew
rlabel metal1 s 29712 4490 29712 4490 4 vdd
port 513 nsew
rlabel metal1 s 29712 3700 29712 3700 4 vdd
port 513 nsew
rlabel metal1 s 29712 4989 29712 4989 4 vdd
port 513 nsew
rlabel metal1 s 27696 3700 27696 3700 4 vdd
port 513 nsew
rlabel metal1 s 28944 5779 28944 5779 4 vdd
port 513 nsew
rlabel metal1 s 29712 4199 29712 4199 4 vdd
port 513 nsew
rlabel metal1 s 28464 3409 28464 3409 4 vdd
port 513 nsew
rlabel metal1 s 27696 6070 27696 6070 4 vdd
port 513 nsew
rlabel metal1 s 29712 6070 29712 6070 4 vdd
port 513 nsew
rlabel metal1 s 28944 4989 28944 4989 4 vdd
port 513 nsew
rlabel metal1 s 29712 5779 29712 5779 4 vdd
port 513 nsew
rlabel metal1 s 27696 5779 27696 5779 4 vdd
port 513 nsew
rlabel metal1 s 27696 4199 27696 4199 4 vdd
port 513 nsew
rlabel metal1 s 28464 3700 28464 3700 4 vdd
port 513 nsew
rlabel metal1 s 28944 5280 28944 5280 4 vdd
port 513 nsew
rlabel metal1 s 28944 6070 28944 6070 4 vdd
port 513 nsew
rlabel metal1 s 28464 4989 28464 4989 4 vdd
port 513 nsew
rlabel metal1 s 27696 4490 27696 4490 4 vdd
port 513 nsew
rlabel metal1 s 28464 4490 28464 4490 4 vdd
port 513 nsew
rlabel metal1 s 28464 5280 28464 5280 4 vdd
port 513 nsew
rlabel metal1 s 25200 3409 25200 3409 4 vdd
port 513 nsew
rlabel metal1 s 25968 4989 25968 4989 4 vdd
port 513 nsew
rlabel metal1 s 26448 3409 26448 3409 4 vdd
port 513 nsew
rlabel metal1 s 26448 4199 26448 4199 4 vdd
port 513 nsew
rlabel metal1 s 26448 5280 26448 5280 4 vdd
port 513 nsew
rlabel metal1 s 26448 3700 26448 3700 4 vdd
port 513 nsew
rlabel metal1 s 27216 5779 27216 5779 4 vdd
port 513 nsew
rlabel metal1 s 27216 3409 27216 3409 4 vdd
port 513 nsew
rlabel metal1 s 25968 5779 25968 5779 4 vdd
port 513 nsew
rlabel metal1 s 26448 4490 26448 4490 4 vdd
port 513 nsew
rlabel metal1 s 27216 4989 27216 4989 4 vdd
port 513 nsew
rlabel metal1 s 25968 5280 25968 5280 4 vdd
port 513 nsew
rlabel metal1 s 26448 4989 26448 4989 4 vdd
port 513 nsew
rlabel metal1 s 25968 3409 25968 3409 4 vdd
port 513 nsew
rlabel metal1 s 25968 6070 25968 6070 4 vdd
port 513 nsew
rlabel metal1 s 25968 4199 25968 4199 4 vdd
port 513 nsew
rlabel metal1 s 27216 5280 27216 5280 4 vdd
port 513 nsew
rlabel metal1 s 25200 4989 25200 4989 4 vdd
port 513 nsew
rlabel metal1 s 25200 4199 25200 4199 4 vdd
port 513 nsew
rlabel metal1 s 25200 6070 25200 6070 4 vdd
port 513 nsew
rlabel metal1 s 27216 4490 27216 4490 4 vdd
port 513 nsew
rlabel metal1 s 26448 6070 26448 6070 4 vdd
port 513 nsew
rlabel metal1 s 25200 5280 25200 5280 4 vdd
port 513 nsew
rlabel metal1 s 27216 4199 27216 4199 4 vdd
port 513 nsew
rlabel metal1 s 25200 5779 25200 5779 4 vdd
port 513 nsew
rlabel metal1 s 25200 4490 25200 4490 4 vdd
port 513 nsew
rlabel metal1 s 25968 3700 25968 3700 4 vdd
port 513 nsew
rlabel metal1 s 25200 3700 25200 3700 4 vdd
port 513 nsew
rlabel metal1 s 26448 5779 26448 5779 4 vdd
port 513 nsew
rlabel metal1 s 25968 4490 25968 4490 4 vdd
port 513 nsew
rlabel metal1 s 27216 6070 27216 6070 4 vdd
port 513 nsew
rlabel metal1 s 27216 3700 27216 3700 4 vdd
port 513 nsew
rlabel metal1 s 27216 540 27216 540 4 vdd
port 513 nsew
rlabel metal1 s 26448 2910 26448 2910 4 vdd
port 513 nsew
rlabel metal1 s 27216 1039 27216 1039 4 vdd
port 513 nsew
rlabel metal1 s 25968 2619 25968 2619 4 vdd
port 513 nsew
rlabel metal1 s 27216 1829 27216 1829 4 vdd
port 513 nsew
rlabel metal1 s 25968 1330 25968 1330 4 vdd
port 513 nsew
rlabel metal1 s 26448 249 26448 249 4 vdd
port 513 nsew
rlabel metal1 s 27216 2120 27216 2120 4 vdd
port 513 nsew
rlabel metal1 s 25200 2619 25200 2619 4 vdd
port 513 nsew
rlabel metal1 s 26448 2120 26448 2120 4 vdd
port 513 nsew
rlabel metal1 s 27216 1330 27216 1330 4 vdd
port 513 nsew
rlabel metal1 s 26448 1330 26448 1330 4 vdd
port 513 nsew
rlabel metal1 s 27216 2619 27216 2619 4 vdd
port 513 nsew
rlabel metal1 s 25968 2120 25968 2120 4 vdd
port 513 nsew
rlabel metal1 s 25968 249 25968 249 4 vdd
port 513 nsew
rlabel metal1 s 27216 249 27216 249 4 vdd
port 513 nsew
rlabel metal1 s 26448 1829 26448 1829 4 vdd
port 513 nsew
rlabel metal1 s 25200 1330 25200 1330 4 vdd
port 513 nsew
rlabel metal1 s 25200 540 25200 540 4 vdd
port 513 nsew
rlabel metal1 s 26448 540 26448 540 4 vdd
port 513 nsew
rlabel metal1 s 25200 1829 25200 1829 4 vdd
port 513 nsew
rlabel metal1 s 25200 2120 25200 2120 4 vdd
port 513 nsew
rlabel metal1 s 25200 1039 25200 1039 4 vdd
port 513 nsew
rlabel metal1 s 27216 2910 27216 2910 4 vdd
port 513 nsew
rlabel metal1 s 25200 2910 25200 2910 4 vdd
port 513 nsew
rlabel metal1 s 25968 1039 25968 1039 4 vdd
port 513 nsew
rlabel metal1 s 25968 1829 25968 1829 4 vdd
port 513 nsew
rlabel metal1 s 26448 2619 26448 2619 4 vdd
port 513 nsew
rlabel metal1 s 25968 2910 25968 2910 4 vdd
port 513 nsew
rlabel metal1 s 25200 249 25200 249 4 vdd
port 513 nsew
rlabel metal1 s 26448 1039 26448 1039 4 vdd
port 513 nsew
rlabel metal1 s 25968 540 25968 540 4 vdd
port 513 nsew
rlabel metal1 s 27696 2120 27696 2120 4 vdd
port 513 nsew
rlabel metal1 s 29712 1039 29712 1039 4 vdd
port 513 nsew
rlabel metal1 s 28464 2120 28464 2120 4 vdd
port 513 nsew
rlabel metal1 s 28464 540 28464 540 4 vdd
port 513 nsew
rlabel metal1 s 28944 249 28944 249 4 vdd
port 513 nsew
rlabel metal1 s 28944 2910 28944 2910 4 vdd
port 513 nsew
rlabel metal1 s 28944 540 28944 540 4 vdd
port 513 nsew
rlabel metal1 s 27696 1330 27696 1330 4 vdd
port 513 nsew
rlabel metal1 s 29712 2910 29712 2910 4 vdd
port 513 nsew
rlabel metal1 s 28464 2619 28464 2619 4 vdd
port 513 nsew
rlabel metal1 s 28944 1330 28944 1330 4 vdd
port 513 nsew
rlabel metal1 s 27696 2910 27696 2910 4 vdd
port 513 nsew
rlabel metal1 s 29712 540 29712 540 4 vdd
port 513 nsew
rlabel metal1 s 28464 249 28464 249 4 vdd
port 513 nsew
rlabel metal1 s 27696 2619 27696 2619 4 vdd
port 513 nsew
rlabel metal1 s 27696 1039 27696 1039 4 vdd
port 513 nsew
rlabel metal1 s 29712 1829 29712 1829 4 vdd
port 513 nsew
rlabel metal1 s 28944 2619 28944 2619 4 vdd
port 513 nsew
rlabel metal1 s 28944 1829 28944 1829 4 vdd
port 513 nsew
rlabel metal1 s 27696 540 27696 540 4 vdd
port 513 nsew
rlabel metal1 s 29712 249 29712 249 4 vdd
port 513 nsew
rlabel metal1 s 28464 1039 28464 1039 4 vdd
port 513 nsew
rlabel metal1 s 27696 249 27696 249 4 vdd
port 513 nsew
rlabel metal1 s 29712 2619 29712 2619 4 vdd
port 513 nsew
rlabel metal1 s 29712 2120 29712 2120 4 vdd
port 513 nsew
rlabel metal1 s 28464 1330 28464 1330 4 vdd
port 513 nsew
rlabel metal1 s 28464 1829 28464 1829 4 vdd
port 513 nsew
rlabel metal1 s 28464 2910 28464 2910 4 vdd
port 513 nsew
rlabel metal1 s 27696 1829 27696 1829 4 vdd
port 513 nsew
rlabel metal1 s 28944 1039 28944 1039 4 vdd
port 513 nsew
rlabel metal1 s 29712 1330 29712 1330 4 vdd
port 513 nsew
rlabel metal1 s 28944 2120 28944 2120 4 vdd
port 513 nsew
rlabel metal1 s 38448 12390 38448 12390 4 vdd
port 513 nsew
rlabel metal1 s 39696 12390 39696 12390 4 vdd
port 513 nsew
rlabel metal1 s 38448 10810 38448 10810 4 vdd
port 513 nsew
rlabel metal1 s 38928 12099 38928 12099 4 vdd
port 513 nsew
rlabel metal1 s 38928 10519 38928 10519 4 vdd
port 513 nsew
rlabel metal1 s 37680 9729 37680 9729 4 vdd
port 513 nsew
rlabel metal1 s 39696 12099 39696 12099 4 vdd
port 513 nsew
rlabel metal1 s 38448 12099 38448 12099 4 vdd
port 513 nsew
rlabel metal1 s 38448 11309 38448 11309 4 vdd
port 513 nsew
rlabel metal1 s 37680 12390 37680 12390 4 vdd
port 513 nsew
rlabel metal1 s 39696 10810 39696 10810 4 vdd
port 513 nsew
rlabel metal1 s 39696 10020 39696 10020 4 vdd
port 513 nsew
rlabel metal1 s 38928 10810 38928 10810 4 vdd
port 513 nsew
rlabel metal1 s 38928 11600 38928 11600 4 vdd
port 513 nsew
rlabel metal1 s 39696 9729 39696 9729 4 vdd
port 513 nsew
rlabel metal1 s 39696 11600 39696 11600 4 vdd
port 513 nsew
rlabel metal1 s 38448 10020 38448 10020 4 vdd
port 513 nsew
rlabel metal1 s 37680 10810 37680 10810 4 vdd
port 513 nsew
rlabel metal1 s 37680 11600 37680 11600 4 vdd
port 513 nsew
rlabel metal1 s 39696 11309 39696 11309 4 vdd
port 513 nsew
rlabel metal1 s 37680 10020 37680 10020 4 vdd
port 513 nsew
rlabel metal1 s 38928 12390 38928 12390 4 vdd
port 513 nsew
rlabel metal1 s 37680 12099 37680 12099 4 vdd
port 513 nsew
rlabel metal1 s 37680 10519 37680 10519 4 vdd
port 513 nsew
rlabel metal1 s 38448 10519 38448 10519 4 vdd
port 513 nsew
rlabel metal1 s 39696 10519 39696 10519 4 vdd
port 513 nsew
rlabel metal1 s 38448 11600 38448 11600 4 vdd
port 513 nsew
rlabel metal1 s 38448 9729 38448 9729 4 vdd
port 513 nsew
rlabel metal1 s 38928 11309 38928 11309 4 vdd
port 513 nsew
rlabel metal1 s 38928 9729 38928 9729 4 vdd
port 513 nsew
rlabel metal1 s 38928 10020 38928 10020 4 vdd
port 513 nsew
rlabel metal1 s 37680 11309 37680 11309 4 vdd
port 513 nsew
rlabel metal1 s 35952 12390 35952 12390 4 vdd
port 513 nsew
rlabel metal1 s 36432 12390 36432 12390 4 vdd
port 513 nsew
rlabel metal1 s 35184 12390 35184 12390 4 vdd
port 513 nsew
rlabel metal1 s 37200 10020 37200 10020 4 vdd
port 513 nsew
rlabel metal1 s 35184 10810 35184 10810 4 vdd
port 513 nsew
rlabel metal1 s 37200 10810 37200 10810 4 vdd
port 513 nsew
rlabel metal1 s 35952 10810 35952 10810 4 vdd
port 513 nsew
rlabel metal1 s 35184 11309 35184 11309 4 vdd
port 513 nsew
rlabel metal1 s 37200 11309 37200 11309 4 vdd
port 513 nsew
rlabel metal1 s 37200 9729 37200 9729 4 vdd
port 513 nsew
rlabel metal1 s 35184 12099 35184 12099 4 vdd
port 513 nsew
rlabel metal1 s 35952 11600 35952 11600 4 vdd
port 513 nsew
rlabel metal1 s 36432 10020 36432 10020 4 vdd
port 513 nsew
rlabel metal1 s 35952 12099 35952 12099 4 vdd
port 513 nsew
rlabel metal1 s 36432 9729 36432 9729 4 vdd
port 513 nsew
rlabel metal1 s 35184 10519 35184 10519 4 vdd
port 513 nsew
rlabel metal1 s 37200 10519 37200 10519 4 vdd
port 513 nsew
rlabel metal1 s 35184 11600 35184 11600 4 vdd
port 513 nsew
rlabel metal1 s 36432 10810 36432 10810 4 vdd
port 513 nsew
rlabel metal1 s 35184 10020 35184 10020 4 vdd
port 513 nsew
rlabel metal1 s 36432 11309 36432 11309 4 vdd
port 513 nsew
rlabel metal1 s 35952 10020 35952 10020 4 vdd
port 513 nsew
rlabel metal1 s 37200 12099 37200 12099 4 vdd
port 513 nsew
rlabel metal1 s 37200 11600 37200 11600 4 vdd
port 513 nsew
rlabel metal1 s 35952 9729 35952 9729 4 vdd
port 513 nsew
rlabel metal1 s 37200 12390 37200 12390 4 vdd
port 513 nsew
rlabel metal1 s 36432 12099 36432 12099 4 vdd
port 513 nsew
rlabel metal1 s 35952 11309 35952 11309 4 vdd
port 513 nsew
rlabel metal1 s 36432 10519 36432 10519 4 vdd
port 513 nsew
rlabel metal1 s 35184 9729 35184 9729 4 vdd
port 513 nsew
rlabel metal1 s 36432 11600 36432 11600 4 vdd
port 513 nsew
rlabel metal1 s 35952 10519 35952 10519 4 vdd
port 513 nsew
rlabel metal1 s 37200 7359 37200 7359 4 vdd
port 513 nsew
rlabel metal1 s 35952 6569 35952 6569 4 vdd
port 513 nsew
rlabel metal1 s 35184 6569 35184 6569 4 vdd
port 513 nsew
rlabel metal1 s 35184 8440 35184 8440 4 vdd
port 513 nsew
rlabel metal1 s 37200 9230 37200 9230 4 vdd
port 513 nsew
rlabel metal1 s 35184 7650 35184 7650 4 vdd
port 513 nsew
rlabel metal1 s 35184 7359 35184 7359 4 vdd
port 513 nsew
rlabel metal1 s 35952 8939 35952 8939 4 vdd
port 513 nsew
rlabel metal1 s 37200 8440 37200 8440 4 vdd
port 513 nsew
rlabel metal1 s 36432 6860 36432 6860 4 vdd
port 513 nsew
rlabel metal1 s 35952 6860 35952 6860 4 vdd
port 513 nsew
rlabel metal1 s 35952 7359 35952 7359 4 vdd
port 513 nsew
rlabel metal1 s 35952 9230 35952 9230 4 vdd
port 513 nsew
rlabel metal1 s 36432 8149 36432 8149 4 vdd
port 513 nsew
rlabel metal1 s 36432 7650 36432 7650 4 vdd
port 513 nsew
rlabel metal1 s 35184 9230 35184 9230 4 vdd
port 513 nsew
rlabel metal1 s 36432 9230 36432 9230 4 vdd
port 513 nsew
rlabel metal1 s 35184 8939 35184 8939 4 vdd
port 513 nsew
rlabel metal1 s 35184 8149 35184 8149 4 vdd
port 513 nsew
rlabel metal1 s 35184 6860 35184 6860 4 vdd
port 513 nsew
rlabel metal1 s 37200 6569 37200 6569 4 vdd
port 513 nsew
rlabel metal1 s 36432 6569 36432 6569 4 vdd
port 513 nsew
rlabel metal1 s 35952 8440 35952 8440 4 vdd
port 513 nsew
rlabel metal1 s 37200 8939 37200 8939 4 vdd
port 513 nsew
rlabel metal1 s 37200 6860 37200 6860 4 vdd
port 513 nsew
rlabel metal1 s 36432 8440 36432 8440 4 vdd
port 513 nsew
rlabel metal1 s 35952 7650 35952 7650 4 vdd
port 513 nsew
rlabel metal1 s 37200 7650 37200 7650 4 vdd
port 513 nsew
rlabel metal1 s 35952 8149 35952 8149 4 vdd
port 513 nsew
rlabel metal1 s 37200 8149 37200 8149 4 vdd
port 513 nsew
rlabel metal1 s 36432 7359 36432 7359 4 vdd
port 513 nsew
rlabel metal1 s 36432 8939 36432 8939 4 vdd
port 513 nsew
rlabel metal1 s 37680 6569 37680 6569 4 vdd
port 513 nsew
rlabel metal1 s 38448 6860 38448 6860 4 vdd
port 513 nsew
rlabel metal1 s 38448 7359 38448 7359 4 vdd
port 513 nsew
rlabel metal1 s 38448 8149 38448 8149 4 vdd
port 513 nsew
rlabel metal1 s 38928 8939 38928 8939 4 vdd
port 513 nsew
rlabel metal1 s 38928 9230 38928 9230 4 vdd
port 513 nsew
rlabel metal1 s 38928 8440 38928 8440 4 vdd
port 513 nsew
rlabel metal1 s 38928 6569 38928 6569 4 vdd
port 513 nsew
rlabel metal1 s 39696 7650 39696 7650 4 vdd
port 513 nsew
rlabel metal1 s 37680 7359 37680 7359 4 vdd
port 513 nsew
rlabel metal1 s 37680 8440 37680 8440 4 vdd
port 513 nsew
rlabel metal1 s 39696 8939 39696 8939 4 vdd
port 513 nsew
rlabel metal1 s 37680 8939 37680 8939 4 vdd
port 513 nsew
rlabel metal1 s 38448 7650 38448 7650 4 vdd
port 513 nsew
rlabel metal1 s 37680 7650 37680 7650 4 vdd
port 513 nsew
rlabel metal1 s 38448 6569 38448 6569 4 vdd
port 513 nsew
rlabel metal1 s 38928 8149 38928 8149 4 vdd
port 513 nsew
rlabel metal1 s 39696 8149 39696 8149 4 vdd
port 513 nsew
rlabel metal1 s 38448 9230 38448 9230 4 vdd
port 513 nsew
rlabel metal1 s 37680 6860 37680 6860 4 vdd
port 513 nsew
rlabel metal1 s 38928 7359 38928 7359 4 vdd
port 513 nsew
rlabel metal1 s 39696 6569 39696 6569 4 vdd
port 513 nsew
rlabel metal1 s 39696 8440 39696 8440 4 vdd
port 513 nsew
rlabel metal1 s 39696 7359 39696 7359 4 vdd
port 513 nsew
rlabel metal1 s 38448 8939 38448 8939 4 vdd
port 513 nsew
rlabel metal1 s 39696 6860 39696 6860 4 vdd
port 513 nsew
rlabel metal1 s 38448 8440 38448 8440 4 vdd
port 513 nsew
rlabel metal1 s 37680 8149 37680 8149 4 vdd
port 513 nsew
rlabel metal1 s 38928 6860 38928 6860 4 vdd
port 513 nsew
rlabel metal1 s 37680 9230 37680 9230 4 vdd
port 513 nsew
rlabel metal1 s 38928 7650 38928 7650 4 vdd
port 513 nsew
rlabel metal1 s 39696 9230 39696 9230 4 vdd
port 513 nsew
rlabel metal1 s 33936 11600 33936 11600 4 vdd
port 513 nsew
rlabel metal1 s 33456 12390 33456 12390 4 vdd
port 513 nsew
rlabel metal1 s 33936 11309 33936 11309 4 vdd
port 513 nsew
rlabel metal1 s 34704 9729 34704 9729 4 vdd
port 513 nsew
rlabel metal1 s 34704 11600 34704 11600 4 vdd
port 513 nsew
rlabel metal1 s 33456 12099 33456 12099 4 vdd
port 513 nsew
rlabel metal1 s 32688 11600 32688 11600 4 vdd
port 513 nsew
rlabel metal1 s 33936 12099 33936 12099 4 vdd
port 513 nsew
rlabel metal1 s 33936 9729 33936 9729 4 vdd
port 513 nsew
rlabel metal1 s 34704 12099 34704 12099 4 vdd
port 513 nsew
rlabel metal1 s 33936 10519 33936 10519 4 vdd
port 513 nsew
rlabel metal1 s 33936 10810 33936 10810 4 vdd
port 513 nsew
rlabel metal1 s 32688 10519 32688 10519 4 vdd
port 513 nsew
rlabel metal1 s 32688 10020 32688 10020 4 vdd
port 513 nsew
rlabel metal1 s 33936 12390 33936 12390 4 vdd
port 513 nsew
rlabel metal1 s 32688 12390 32688 12390 4 vdd
port 513 nsew
rlabel metal1 s 34704 10020 34704 10020 4 vdd
port 513 nsew
rlabel metal1 s 34704 11309 34704 11309 4 vdd
port 513 nsew
rlabel metal1 s 32688 12099 32688 12099 4 vdd
port 513 nsew
rlabel metal1 s 32688 9729 32688 9729 4 vdd
port 513 nsew
rlabel metal1 s 33456 10519 33456 10519 4 vdd
port 513 nsew
rlabel metal1 s 33936 10020 33936 10020 4 vdd
port 513 nsew
rlabel metal1 s 33456 11309 33456 11309 4 vdd
port 513 nsew
rlabel metal1 s 34704 10519 34704 10519 4 vdd
port 513 nsew
rlabel metal1 s 33456 11600 33456 11600 4 vdd
port 513 nsew
rlabel metal1 s 34704 10810 34704 10810 4 vdd
port 513 nsew
rlabel metal1 s 32688 11309 32688 11309 4 vdd
port 513 nsew
rlabel metal1 s 32688 10810 32688 10810 4 vdd
port 513 nsew
rlabel metal1 s 33456 10810 33456 10810 4 vdd
port 513 nsew
rlabel metal1 s 33456 9729 33456 9729 4 vdd
port 513 nsew
rlabel metal1 s 33456 10020 33456 10020 4 vdd
port 513 nsew
rlabel metal1 s 34704 12390 34704 12390 4 vdd
port 513 nsew
rlabel metal1 s 31440 11600 31440 11600 4 vdd
port 513 nsew
rlabel metal1 s 30960 10020 30960 10020 4 vdd
port 513 nsew
rlabel metal1 s 30960 11600 30960 11600 4 vdd
port 513 nsew
rlabel metal1 s 31440 10020 31440 10020 4 vdd
port 513 nsew
rlabel metal1 s 32208 12099 32208 12099 4 vdd
port 513 nsew
rlabel metal1 s 32208 10020 32208 10020 4 vdd
port 513 nsew
rlabel metal1 s 31440 11309 31440 11309 4 vdd
port 513 nsew
rlabel metal1 s 32208 10519 32208 10519 4 vdd
port 513 nsew
rlabel metal1 s 32208 9729 32208 9729 4 vdd
port 513 nsew
rlabel metal1 s 30192 10519 30192 10519 4 vdd
port 513 nsew
rlabel metal1 s 31440 12390 31440 12390 4 vdd
port 513 nsew
rlabel metal1 s 32208 10810 32208 10810 4 vdd
port 513 nsew
rlabel metal1 s 31440 10810 31440 10810 4 vdd
port 513 nsew
rlabel metal1 s 30192 11309 30192 11309 4 vdd
port 513 nsew
rlabel metal1 s 30960 12099 30960 12099 4 vdd
port 513 nsew
rlabel metal1 s 30960 12390 30960 12390 4 vdd
port 513 nsew
rlabel metal1 s 30960 9729 30960 9729 4 vdd
port 513 nsew
rlabel metal1 s 30960 11309 30960 11309 4 vdd
port 513 nsew
rlabel metal1 s 32208 12390 32208 12390 4 vdd
port 513 nsew
rlabel metal1 s 32208 11309 32208 11309 4 vdd
port 513 nsew
rlabel metal1 s 30192 9729 30192 9729 4 vdd
port 513 nsew
rlabel metal1 s 30960 10519 30960 10519 4 vdd
port 513 nsew
rlabel metal1 s 30192 12390 30192 12390 4 vdd
port 513 nsew
rlabel metal1 s 30960 10810 30960 10810 4 vdd
port 513 nsew
rlabel metal1 s 30192 10020 30192 10020 4 vdd
port 513 nsew
rlabel metal1 s 30192 10810 30192 10810 4 vdd
port 513 nsew
rlabel metal1 s 32208 11600 32208 11600 4 vdd
port 513 nsew
rlabel metal1 s 30192 11600 30192 11600 4 vdd
port 513 nsew
rlabel metal1 s 31440 12099 31440 12099 4 vdd
port 513 nsew
rlabel metal1 s 30192 12099 30192 12099 4 vdd
port 513 nsew
rlabel metal1 s 31440 10519 31440 10519 4 vdd
port 513 nsew
rlabel metal1 s 31440 9729 31440 9729 4 vdd
port 513 nsew
rlabel metal1 s 31440 7359 31440 7359 4 vdd
port 513 nsew
rlabel metal1 s 30192 8149 30192 8149 4 vdd
port 513 nsew
rlabel metal1 s 30960 6569 30960 6569 4 vdd
port 513 nsew
rlabel metal1 s 31440 8440 31440 8440 4 vdd
port 513 nsew
rlabel metal1 s 32208 6860 32208 6860 4 vdd
port 513 nsew
rlabel metal1 s 31440 8149 31440 8149 4 vdd
port 513 nsew
rlabel metal1 s 30192 9230 30192 9230 4 vdd
port 513 nsew
rlabel metal1 s 32208 9230 32208 9230 4 vdd
port 513 nsew
rlabel metal1 s 30960 9230 30960 9230 4 vdd
port 513 nsew
rlabel metal1 s 30960 8440 30960 8440 4 vdd
port 513 nsew
rlabel metal1 s 30192 8440 30192 8440 4 vdd
port 513 nsew
rlabel metal1 s 31440 9230 31440 9230 4 vdd
port 513 nsew
rlabel metal1 s 32208 7650 32208 7650 4 vdd
port 513 nsew
rlabel metal1 s 30960 8149 30960 8149 4 vdd
port 513 nsew
rlabel metal1 s 31440 8939 31440 8939 4 vdd
port 513 nsew
rlabel metal1 s 30960 8939 30960 8939 4 vdd
port 513 nsew
rlabel metal1 s 32208 6569 32208 6569 4 vdd
port 513 nsew
rlabel metal1 s 30960 6860 30960 6860 4 vdd
port 513 nsew
rlabel metal1 s 32208 8149 32208 8149 4 vdd
port 513 nsew
rlabel metal1 s 30960 7650 30960 7650 4 vdd
port 513 nsew
rlabel metal1 s 32208 7359 32208 7359 4 vdd
port 513 nsew
rlabel metal1 s 32208 8440 32208 8440 4 vdd
port 513 nsew
rlabel metal1 s 30960 7359 30960 7359 4 vdd
port 513 nsew
rlabel metal1 s 32208 8939 32208 8939 4 vdd
port 513 nsew
rlabel metal1 s 30192 7359 30192 7359 4 vdd
port 513 nsew
rlabel metal1 s 31440 7650 31440 7650 4 vdd
port 513 nsew
rlabel metal1 s 30192 6860 30192 6860 4 vdd
port 513 nsew
rlabel metal1 s 30192 8939 30192 8939 4 vdd
port 513 nsew
rlabel metal1 s 31440 6860 31440 6860 4 vdd
port 513 nsew
rlabel metal1 s 30192 6569 30192 6569 4 vdd
port 513 nsew
rlabel metal1 s 30192 7650 30192 7650 4 vdd
port 513 nsew
rlabel metal1 s 31440 6569 31440 6569 4 vdd
port 513 nsew
rlabel metal1 s 34704 6569 34704 6569 4 vdd
port 513 nsew
rlabel metal1 s 34704 8939 34704 8939 4 vdd
port 513 nsew
rlabel metal1 s 34704 8149 34704 8149 4 vdd
port 513 nsew
rlabel metal1 s 33936 9230 33936 9230 4 vdd
port 513 nsew
rlabel metal1 s 34704 7650 34704 7650 4 vdd
port 513 nsew
rlabel metal1 s 33456 8939 33456 8939 4 vdd
port 513 nsew
rlabel metal1 s 33936 7650 33936 7650 4 vdd
port 513 nsew
rlabel metal1 s 33456 6860 33456 6860 4 vdd
port 513 nsew
rlabel metal1 s 33936 8149 33936 8149 4 vdd
port 513 nsew
rlabel metal1 s 33456 8149 33456 8149 4 vdd
port 513 nsew
rlabel metal1 s 33936 8440 33936 8440 4 vdd
port 513 nsew
rlabel metal1 s 33456 7359 33456 7359 4 vdd
port 513 nsew
rlabel metal1 s 33936 6860 33936 6860 4 vdd
port 513 nsew
rlabel metal1 s 32688 6569 32688 6569 4 vdd
port 513 nsew
rlabel metal1 s 34704 6860 34704 6860 4 vdd
port 513 nsew
rlabel metal1 s 33936 6569 33936 6569 4 vdd
port 513 nsew
rlabel metal1 s 32688 8149 32688 8149 4 vdd
port 513 nsew
rlabel metal1 s 34704 8440 34704 8440 4 vdd
port 513 nsew
rlabel metal1 s 33456 8440 33456 8440 4 vdd
port 513 nsew
rlabel metal1 s 33456 6569 33456 6569 4 vdd
port 513 nsew
rlabel metal1 s 32688 8939 32688 8939 4 vdd
port 513 nsew
rlabel metal1 s 33936 8939 33936 8939 4 vdd
port 513 nsew
rlabel metal1 s 32688 7359 32688 7359 4 vdd
port 513 nsew
rlabel metal1 s 32688 8440 32688 8440 4 vdd
port 513 nsew
rlabel metal1 s 34704 7359 34704 7359 4 vdd
port 513 nsew
rlabel metal1 s 34704 9230 34704 9230 4 vdd
port 513 nsew
rlabel metal1 s 32688 9230 32688 9230 4 vdd
port 513 nsew
rlabel metal1 s 32688 6860 32688 6860 4 vdd
port 513 nsew
rlabel metal1 s 32688 7650 32688 7650 4 vdd
port 513 nsew
rlabel metal1 s 33936 7359 33936 7359 4 vdd
port 513 nsew
rlabel metal1 s 33456 7650 33456 7650 4 vdd
port 513 nsew
rlabel metal1 s 33456 9230 33456 9230 4 vdd
port 513 nsew
rlabel metal1 s 32688 3409 32688 3409 4 vdd
port 513 nsew
rlabel metal1 s 32688 5280 32688 5280 4 vdd
port 513 nsew
rlabel metal1 s 33456 5779 33456 5779 4 vdd
port 513 nsew
rlabel metal1 s 32688 4490 32688 4490 4 vdd
port 513 nsew
rlabel metal1 s 32688 5779 32688 5779 4 vdd
port 513 nsew
rlabel metal1 s 33456 6070 33456 6070 4 vdd
port 513 nsew
rlabel metal1 s 33936 5779 33936 5779 4 vdd
port 513 nsew
rlabel metal1 s 34704 4199 34704 4199 4 vdd
port 513 nsew
rlabel metal1 s 33936 4199 33936 4199 4 vdd
port 513 nsew
rlabel metal1 s 33936 3409 33936 3409 4 vdd
port 513 nsew
rlabel metal1 s 34704 4490 34704 4490 4 vdd
port 513 nsew
rlabel metal1 s 33456 3409 33456 3409 4 vdd
port 513 nsew
rlabel metal1 s 34704 3700 34704 3700 4 vdd
port 513 nsew
rlabel metal1 s 34704 5779 34704 5779 4 vdd
port 513 nsew
rlabel metal1 s 33456 4490 33456 4490 4 vdd
port 513 nsew
rlabel metal1 s 32688 4199 32688 4199 4 vdd
port 513 nsew
rlabel metal1 s 33936 6070 33936 6070 4 vdd
port 513 nsew
rlabel metal1 s 34704 4989 34704 4989 4 vdd
port 513 nsew
rlabel metal1 s 33456 4199 33456 4199 4 vdd
port 513 nsew
rlabel metal1 s 32688 4989 32688 4989 4 vdd
port 513 nsew
rlabel metal1 s 34704 6070 34704 6070 4 vdd
port 513 nsew
rlabel metal1 s 34704 3409 34704 3409 4 vdd
port 513 nsew
rlabel metal1 s 33456 5280 33456 5280 4 vdd
port 513 nsew
rlabel metal1 s 33936 4989 33936 4989 4 vdd
port 513 nsew
rlabel metal1 s 33456 4989 33456 4989 4 vdd
port 513 nsew
rlabel metal1 s 32688 6070 32688 6070 4 vdd
port 513 nsew
rlabel metal1 s 33936 4490 33936 4490 4 vdd
port 513 nsew
rlabel metal1 s 33456 3700 33456 3700 4 vdd
port 513 nsew
rlabel metal1 s 33936 5280 33936 5280 4 vdd
port 513 nsew
rlabel metal1 s 34704 5280 34704 5280 4 vdd
port 513 nsew
rlabel metal1 s 33936 3700 33936 3700 4 vdd
port 513 nsew
rlabel metal1 s 32688 3700 32688 3700 4 vdd
port 513 nsew
rlabel metal1 s 32208 5280 32208 5280 4 vdd
port 513 nsew
rlabel metal1 s 31440 4989 31440 4989 4 vdd
port 513 nsew
rlabel metal1 s 32208 4490 32208 4490 4 vdd
port 513 nsew
rlabel metal1 s 30960 5280 30960 5280 4 vdd
port 513 nsew
rlabel metal1 s 32208 6070 32208 6070 4 vdd
port 513 nsew
rlabel metal1 s 30192 6070 30192 6070 4 vdd
port 513 nsew
rlabel metal1 s 32208 5779 32208 5779 4 vdd
port 513 nsew
rlabel metal1 s 32208 3700 32208 3700 4 vdd
port 513 nsew
rlabel metal1 s 31440 3700 31440 3700 4 vdd
port 513 nsew
rlabel metal1 s 31440 3409 31440 3409 4 vdd
port 513 nsew
rlabel metal1 s 30960 4989 30960 4989 4 vdd
port 513 nsew
rlabel metal1 s 31440 5779 31440 5779 4 vdd
port 513 nsew
rlabel metal1 s 31440 5280 31440 5280 4 vdd
port 513 nsew
rlabel metal1 s 30960 6070 30960 6070 4 vdd
port 513 nsew
rlabel metal1 s 30960 4490 30960 4490 4 vdd
port 513 nsew
rlabel metal1 s 31440 4490 31440 4490 4 vdd
port 513 nsew
rlabel metal1 s 30192 3700 30192 3700 4 vdd
port 513 nsew
rlabel metal1 s 30192 5280 30192 5280 4 vdd
port 513 nsew
rlabel metal1 s 30192 4490 30192 4490 4 vdd
port 513 nsew
rlabel metal1 s 30192 3409 30192 3409 4 vdd
port 513 nsew
rlabel metal1 s 30960 3700 30960 3700 4 vdd
port 513 nsew
rlabel metal1 s 30960 4199 30960 4199 4 vdd
port 513 nsew
rlabel metal1 s 32208 3409 32208 3409 4 vdd
port 513 nsew
rlabel metal1 s 32208 4989 32208 4989 4 vdd
port 513 nsew
rlabel metal1 s 30192 4989 30192 4989 4 vdd
port 513 nsew
rlabel metal1 s 32208 4199 32208 4199 4 vdd
port 513 nsew
rlabel metal1 s 30960 3409 30960 3409 4 vdd
port 513 nsew
rlabel metal1 s 30192 5779 30192 5779 4 vdd
port 513 nsew
rlabel metal1 s 31440 4199 31440 4199 4 vdd
port 513 nsew
rlabel metal1 s 30960 5779 30960 5779 4 vdd
port 513 nsew
rlabel metal1 s 31440 6070 31440 6070 4 vdd
port 513 nsew
rlabel metal1 s 30192 4199 30192 4199 4 vdd
port 513 nsew
rlabel metal1 s 30960 2120 30960 2120 4 vdd
port 513 nsew
rlabel metal1 s 30192 249 30192 249 4 vdd
port 513 nsew
rlabel metal1 s 31440 2120 31440 2120 4 vdd
port 513 nsew
rlabel metal1 s 30960 2619 30960 2619 4 vdd
port 513 nsew
rlabel metal1 s 32208 2619 32208 2619 4 vdd
port 513 nsew
rlabel metal1 s 31440 1039 31440 1039 4 vdd
port 513 nsew
rlabel metal1 s 30960 249 30960 249 4 vdd
port 513 nsew
rlabel metal1 s 32208 2120 32208 2120 4 vdd
port 513 nsew
rlabel metal1 s 31440 2910 31440 2910 4 vdd
port 513 nsew
rlabel metal1 s 32208 1039 32208 1039 4 vdd
port 513 nsew
rlabel metal1 s 31440 2619 31440 2619 4 vdd
port 513 nsew
rlabel metal1 s 30960 1039 30960 1039 4 vdd
port 513 nsew
rlabel metal1 s 30960 1330 30960 1330 4 vdd
port 513 nsew
rlabel metal1 s 30192 1829 30192 1829 4 vdd
port 513 nsew
rlabel metal1 s 32208 249 32208 249 4 vdd
port 513 nsew
rlabel metal1 s 31440 1829 31440 1829 4 vdd
port 513 nsew
rlabel metal1 s 31440 1330 31440 1330 4 vdd
port 513 nsew
rlabel metal1 s 31440 249 31440 249 4 vdd
port 513 nsew
rlabel metal1 s 32208 1330 32208 1330 4 vdd
port 513 nsew
rlabel metal1 s 30960 540 30960 540 4 vdd
port 513 nsew
rlabel metal1 s 32208 2910 32208 2910 4 vdd
port 513 nsew
rlabel metal1 s 32208 540 32208 540 4 vdd
port 513 nsew
rlabel metal1 s 30192 540 30192 540 4 vdd
port 513 nsew
rlabel metal1 s 30192 1039 30192 1039 4 vdd
port 513 nsew
rlabel metal1 s 30192 1330 30192 1330 4 vdd
port 513 nsew
rlabel metal1 s 32208 1829 32208 1829 4 vdd
port 513 nsew
rlabel metal1 s 30192 2619 30192 2619 4 vdd
port 513 nsew
rlabel metal1 s 31440 540 31440 540 4 vdd
port 513 nsew
rlabel metal1 s 30192 2120 30192 2120 4 vdd
port 513 nsew
rlabel metal1 s 30192 2910 30192 2910 4 vdd
port 513 nsew
rlabel metal1 s 30960 1829 30960 1829 4 vdd
port 513 nsew
rlabel metal1 s 30960 2910 30960 2910 4 vdd
port 513 nsew
rlabel metal1 s 34704 2120 34704 2120 4 vdd
port 513 nsew
rlabel metal1 s 32688 2910 32688 2910 4 vdd
port 513 nsew
rlabel metal1 s 33936 2910 33936 2910 4 vdd
port 513 nsew
rlabel metal1 s 33456 249 33456 249 4 vdd
port 513 nsew
rlabel metal1 s 34704 249 34704 249 4 vdd
port 513 nsew
rlabel metal1 s 32688 2619 32688 2619 4 vdd
port 513 nsew
rlabel metal1 s 33936 249 33936 249 4 vdd
port 513 nsew
rlabel metal1 s 33936 1330 33936 1330 4 vdd
port 513 nsew
rlabel metal1 s 34704 2910 34704 2910 4 vdd
port 513 nsew
rlabel metal1 s 32688 2120 32688 2120 4 vdd
port 513 nsew
rlabel metal1 s 33936 1829 33936 1829 4 vdd
port 513 nsew
rlabel metal1 s 33456 1829 33456 1829 4 vdd
port 513 nsew
rlabel metal1 s 32688 249 32688 249 4 vdd
port 513 nsew
rlabel metal1 s 33456 2910 33456 2910 4 vdd
port 513 nsew
rlabel metal1 s 33936 2120 33936 2120 4 vdd
port 513 nsew
rlabel metal1 s 33936 2619 33936 2619 4 vdd
port 513 nsew
rlabel metal1 s 34704 540 34704 540 4 vdd
port 513 nsew
rlabel metal1 s 34704 1829 34704 1829 4 vdd
port 513 nsew
rlabel metal1 s 33456 540 33456 540 4 vdd
port 513 nsew
rlabel metal1 s 34704 1330 34704 1330 4 vdd
port 513 nsew
rlabel metal1 s 33456 2619 33456 2619 4 vdd
port 513 nsew
rlabel metal1 s 33936 1039 33936 1039 4 vdd
port 513 nsew
rlabel metal1 s 33456 1039 33456 1039 4 vdd
port 513 nsew
rlabel metal1 s 32688 1039 32688 1039 4 vdd
port 513 nsew
rlabel metal1 s 34704 2619 34704 2619 4 vdd
port 513 nsew
rlabel metal1 s 33936 540 33936 540 4 vdd
port 513 nsew
rlabel metal1 s 33456 2120 33456 2120 4 vdd
port 513 nsew
rlabel metal1 s 33456 1330 33456 1330 4 vdd
port 513 nsew
rlabel metal1 s 32688 1330 32688 1330 4 vdd
port 513 nsew
rlabel metal1 s 34704 1039 34704 1039 4 vdd
port 513 nsew
rlabel metal1 s 32688 540 32688 540 4 vdd
port 513 nsew
rlabel metal1 s 32688 1829 32688 1829 4 vdd
port 513 nsew
rlabel metal1 s 38448 3409 38448 3409 4 vdd
port 513 nsew
rlabel metal1 s 38448 4199 38448 4199 4 vdd
port 513 nsew
rlabel metal1 s 39696 6070 39696 6070 4 vdd
port 513 nsew
rlabel metal1 s 37680 4199 37680 4199 4 vdd
port 513 nsew
rlabel metal1 s 39696 3700 39696 3700 4 vdd
port 513 nsew
rlabel metal1 s 38928 4199 38928 4199 4 vdd
port 513 nsew
rlabel metal1 s 38928 4989 38928 4989 4 vdd
port 513 nsew
rlabel metal1 s 37680 5280 37680 5280 4 vdd
port 513 nsew
rlabel metal1 s 38928 5280 38928 5280 4 vdd
port 513 nsew
rlabel metal1 s 38928 6070 38928 6070 4 vdd
port 513 nsew
rlabel metal1 s 38448 3700 38448 3700 4 vdd
port 513 nsew
rlabel metal1 s 38928 3409 38928 3409 4 vdd
port 513 nsew
rlabel metal1 s 37680 4989 37680 4989 4 vdd
port 513 nsew
rlabel metal1 s 37680 5779 37680 5779 4 vdd
port 513 nsew
rlabel metal1 s 39696 3409 39696 3409 4 vdd
port 513 nsew
rlabel metal1 s 37680 3409 37680 3409 4 vdd
port 513 nsew
rlabel metal1 s 39696 5280 39696 5280 4 vdd
port 513 nsew
rlabel metal1 s 37680 4490 37680 4490 4 vdd
port 513 nsew
rlabel metal1 s 38448 5779 38448 5779 4 vdd
port 513 nsew
rlabel metal1 s 38928 5779 38928 5779 4 vdd
port 513 nsew
rlabel metal1 s 39696 4199 39696 4199 4 vdd
port 513 nsew
rlabel metal1 s 38928 3700 38928 3700 4 vdd
port 513 nsew
rlabel metal1 s 38448 6070 38448 6070 4 vdd
port 513 nsew
rlabel metal1 s 38448 5280 38448 5280 4 vdd
port 513 nsew
rlabel metal1 s 38448 4989 38448 4989 4 vdd
port 513 nsew
rlabel metal1 s 37680 6070 37680 6070 4 vdd
port 513 nsew
rlabel metal1 s 39696 4989 39696 4989 4 vdd
port 513 nsew
rlabel metal1 s 38928 4490 38928 4490 4 vdd
port 513 nsew
rlabel metal1 s 39696 5779 39696 5779 4 vdd
port 513 nsew
rlabel metal1 s 39696 4490 39696 4490 4 vdd
port 513 nsew
rlabel metal1 s 37680 3700 37680 3700 4 vdd
port 513 nsew
rlabel metal1 s 38448 4490 38448 4490 4 vdd
port 513 nsew
rlabel metal1 s 36432 5779 36432 5779 4 vdd
port 513 nsew
rlabel metal1 s 36432 3700 36432 3700 4 vdd
port 513 nsew
rlabel metal1 s 35952 5280 35952 5280 4 vdd
port 513 nsew
rlabel metal1 s 35184 4199 35184 4199 4 vdd
port 513 nsew
rlabel metal1 s 35184 3409 35184 3409 4 vdd
port 513 nsew
rlabel metal1 s 35184 3700 35184 3700 4 vdd
port 513 nsew
rlabel metal1 s 35952 4989 35952 4989 4 vdd
port 513 nsew
rlabel metal1 s 36432 4490 36432 4490 4 vdd
port 513 nsew
rlabel metal1 s 35952 4199 35952 4199 4 vdd
port 513 nsew
rlabel metal1 s 35184 4490 35184 4490 4 vdd
port 513 nsew
rlabel metal1 s 37200 3409 37200 3409 4 vdd
port 513 nsew
rlabel metal1 s 35952 3409 35952 3409 4 vdd
port 513 nsew
rlabel metal1 s 35952 6070 35952 6070 4 vdd
port 513 nsew
rlabel metal1 s 37200 3700 37200 3700 4 vdd
port 513 nsew
rlabel metal1 s 36432 3409 36432 3409 4 vdd
port 513 nsew
rlabel metal1 s 36432 6070 36432 6070 4 vdd
port 513 nsew
rlabel metal1 s 36432 5280 36432 5280 4 vdd
port 513 nsew
rlabel metal1 s 35184 4989 35184 4989 4 vdd
port 513 nsew
rlabel metal1 s 35184 5779 35184 5779 4 vdd
port 513 nsew
rlabel metal1 s 35184 6070 35184 6070 4 vdd
port 513 nsew
rlabel metal1 s 35952 4490 35952 4490 4 vdd
port 513 nsew
rlabel metal1 s 37200 4490 37200 4490 4 vdd
port 513 nsew
rlabel metal1 s 35952 5779 35952 5779 4 vdd
port 513 nsew
rlabel metal1 s 36432 4989 36432 4989 4 vdd
port 513 nsew
rlabel metal1 s 37200 4199 37200 4199 4 vdd
port 513 nsew
rlabel metal1 s 35184 5280 35184 5280 4 vdd
port 513 nsew
rlabel metal1 s 35952 3700 35952 3700 4 vdd
port 513 nsew
rlabel metal1 s 37200 4989 37200 4989 4 vdd
port 513 nsew
rlabel metal1 s 37200 6070 37200 6070 4 vdd
port 513 nsew
rlabel metal1 s 36432 4199 36432 4199 4 vdd
port 513 nsew
rlabel metal1 s 37200 5779 37200 5779 4 vdd
port 513 nsew
rlabel metal1 s 37200 5280 37200 5280 4 vdd
port 513 nsew
rlabel metal1 s 36432 1829 36432 1829 4 vdd
port 513 nsew
rlabel metal1 s 35952 2619 35952 2619 4 vdd
port 513 nsew
rlabel metal1 s 35952 540 35952 540 4 vdd
port 513 nsew
rlabel metal1 s 37200 1829 37200 1829 4 vdd
port 513 nsew
rlabel metal1 s 35952 1330 35952 1330 4 vdd
port 513 nsew
rlabel metal1 s 35184 1330 35184 1330 4 vdd
port 513 nsew
rlabel metal1 s 37200 2619 37200 2619 4 vdd
port 513 nsew
rlabel metal1 s 35184 540 35184 540 4 vdd
port 513 nsew
rlabel metal1 s 35952 2120 35952 2120 4 vdd
port 513 nsew
rlabel metal1 s 35952 249 35952 249 4 vdd
port 513 nsew
rlabel metal1 s 35184 2619 35184 2619 4 vdd
port 513 nsew
rlabel metal1 s 36432 2120 36432 2120 4 vdd
port 513 nsew
rlabel metal1 s 36432 540 36432 540 4 vdd
port 513 nsew
rlabel metal1 s 35184 2910 35184 2910 4 vdd
port 513 nsew
rlabel metal1 s 37200 2910 37200 2910 4 vdd
port 513 nsew
rlabel metal1 s 36432 2619 36432 2619 4 vdd
port 513 nsew
rlabel metal1 s 35184 1039 35184 1039 4 vdd
port 513 nsew
rlabel metal1 s 35952 1829 35952 1829 4 vdd
port 513 nsew
rlabel metal1 s 37200 540 37200 540 4 vdd
port 513 nsew
rlabel metal1 s 35184 2120 35184 2120 4 vdd
port 513 nsew
rlabel metal1 s 36432 1039 36432 1039 4 vdd
port 513 nsew
rlabel metal1 s 37200 249 37200 249 4 vdd
port 513 nsew
rlabel metal1 s 35184 249 35184 249 4 vdd
port 513 nsew
rlabel metal1 s 36432 1330 36432 1330 4 vdd
port 513 nsew
rlabel metal1 s 36432 2910 36432 2910 4 vdd
port 513 nsew
rlabel metal1 s 35952 1039 35952 1039 4 vdd
port 513 nsew
rlabel metal1 s 37200 2120 37200 2120 4 vdd
port 513 nsew
rlabel metal1 s 37200 1330 37200 1330 4 vdd
port 513 nsew
rlabel metal1 s 36432 249 36432 249 4 vdd
port 513 nsew
rlabel metal1 s 35952 2910 35952 2910 4 vdd
port 513 nsew
rlabel metal1 s 37200 1039 37200 1039 4 vdd
port 513 nsew
rlabel metal1 s 35184 1829 35184 1829 4 vdd
port 513 nsew
rlabel metal1 s 37680 1829 37680 1829 4 vdd
port 513 nsew
rlabel metal1 s 39696 540 39696 540 4 vdd
port 513 nsew
rlabel metal1 s 39696 1829 39696 1829 4 vdd
port 513 nsew
rlabel metal1 s 38928 1829 38928 1829 4 vdd
port 513 nsew
rlabel metal1 s 37680 540 37680 540 4 vdd
port 513 nsew
rlabel metal1 s 37680 2910 37680 2910 4 vdd
port 513 nsew
rlabel metal1 s 38928 540 38928 540 4 vdd
port 513 nsew
rlabel metal1 s 39696 2619 39696 2619 4 vdd
port 513 nsew
rlabel metal1 s 38928 2120 38928 2120 4 vdd
port 513 nsew
rlabel metal1 s 39696 249 39696 249 4 vdd
port 513 nsew
rlabel metal1 s 38448 1330 38448 1330 4 vdd
port 513 nsew
rlabel metal1 s 37680 2120 37680 2120 4 vdd
port 513 nsew
rlabel metal1 s 38928 2910 38928 2910 4 vdd
port 513 nsew
rlabel metal1 s 38928 249 38928 249 4 vdd
port 513 nsew
rlabel metal1 s 38448 1829 38448 1829 4 vdd
port 513 nsew
rlabel metal1 s 38448 1039 38448 1039 4 vdd
port 513 nsew
rlabel metal1 s 38928 2619 38928 2619 4 vdd
port 513 nsew
rlabel metal1 s 38928 1039 38928 1039 4 vdd
port 513 nsew
rlabel metal1 s 37680 249 37680 249 4 vdd
port 513 nsew
rlabel metal1 s 39696 2120 39696 2120 4 vdd
port 513 nsew
rlabel metal1 s 38448 2910 38448 2910 4 vdd
port 513 nsew
rlabel metal1 s 37680 2619 37680 2619 4 vdd
port 513 nsew
rlabel metal1 s 37680 1330 37680 1330 4 vdd
port 513 nsew
rlabel metal1 s 37680 1039 37680 1039 4 vdd
port 513 nsew
rlabel metal1 s 39696 2910 39696 2910 4 vdd
port 513 nsew
rlabel metal1 s 38928 1330 38928 1330 4 vdd
port 513 nsew
rlabel metal1 s 38448 249 38448 249 4 vdd
port 513 nsew
rlabel metal1 s 39696 1039 39696 1039 4 vdd
port 513 nsew
rlabel metal1 s 38448 540 38448 540 4 vdd
port 513 nsew
rlabel metal1 s 38448 2619 38448 2619 4 vdd
port 513 nsew
rlabel metal1 s 38448 2120 38448 2120 4 vdd
port 513 nsew
rlabel metal1 s 39696 1330 39696 1330 4 vdd
port 513 nsew
rlabel metal2 s 38448 48190 38448 48190 4 gnd
port 514 nsew
rlabel metal2 s 37680 49533 37680 49533 4 gnd
port 514 nsew
rlabel metal2 s 38448 49217 38448 49217 4 gnd
port 514 nsew
rlabel metal2 s 38448 50323 38448 50323 4 gnd
port 514 nsew
rlabel metal2 s 37680 48743 37680 48743 4 gnd
port 514 nsew
rlabel metal2 s 38448 47953 38448 47953 4 gnd
port 514 nsew
rlabel metal2 s 37680 47953 37680 47953 4 gnd
port 514 nsew
rlabel metal2 s 39696 49770 39696 49770 4 gnd
port 514 nsew
rlabel metal2 s 38928 48980 38928 48980 4 gnd
port 514 nsew
rlabel metal2 s 38928 48427 38928 48427 4 gnd
port 514 nsew
rlabel metal2 s 39696 50323 39696 50323 4 gnd
port 514 nsew
rlabel metal2 s 39696 49533 39696 49533 4 gnd
port 514 nsew
rlabel metal2 s 37680 49217 37680 49217 4 gnd
port 514 nsew
rlabel metal2 s 38448 49770 38448 49770 4 gnd
port 514 nsew
rlabel metal2 s 38448 48980 38448 48980 4 gnd
port 514 nsew
rlabel metal2 s 39696 48743 39696 48743 4 gnd
port 514 nsew
rlabel metal2 s 38928 50007 38928 50007 4 gnd
port 514 nsew
rlabel metal2 s 38448 49533 38448 49533 4 gnd
port 514 nsew
rlabel metal2 s 38928 48743 38928 48743 4 gnd
port 514 nsew
rlabel metal2 s 39696 48980 39696 48980 4 gnd
port 514 nsew
rlabel metal2 s 38928 50323 38928 50323 4 gnd
port 514 nsew
rlabel metal2 s 38448 47637 38448 47637 4 gnd
port 514 nsew
rlabel metal2 s 39696 47637 39696 47637 4 gnd
port 514 nsew
rlabel metal2 s 38928 49217 38928 49217 4 gnd
port 514 nsew
rlabel metal2 s 37680 50007 37680 50007 4 gnd
port 514 nsew
rlabel metal2 s 37680 48190 37680 48190 4 gnd
port 514 nsew
rlabel metal2 s 38448 48427 38448 48427 4 gnd
port 514 nsew
rlabel metal2 s 38928 47953 38928 47953 4 gnd
port 514 nsew
rlabel metal2 s 39696 50007 39696 50007 4 gnd
port 514 nsew
rlabel metal2 s 39696 48190 39696 48190 4 gnd
port 514 nsew
rlabel metal2 s 37680 50560 37680 50560 4 gnd
port 514 nsew
rlabel metal2 s 38928 49533 38928 49533 4 gnd
port 514 nsew
rlabel metal2 s 38928 48190 38928 48190 4 gnd
port 514 nsew
rlabel metal2 s 39696 50560 39696 50560 4 gnd
port 514 nsew
rlabel metal2 s 38448 50007 38448 50007 4 gnd
port 514 nsew
rlabel metal2 s 38928 50560 38928 50560 4 gnd
port 514 nsew
rlabel metal2 s 39696 49217 39696 49217 4 gnd
port 514 nsew
rlabel metal2 s 37680 49770 37680 49770 4 gnd
port 514 nsew
rlabel metal2 s 39696 47953 39696 47953 4 gnd
port 514 nsew
rlabel metal2 s 37680 48980 37680 48980 4 gnd
port 514 nsew
rlabel metal2 s 37680 50323 37680 50323 4 gnd
port 514 nsew
rlabel metal2 s 38928 49770 38928 49770 4 gnd
port 514 nsew
rlabel metal2 s 37680 47637 37680 47637 4 gnd
port 514 nsew
rlabel metal2 s 38448 50560 38448 50560 4 gnd
port 514 nsew
rlabel metal2 s 39696 48427 39696 48427 4 gnd
port 514 nsew
rlabel metal2 s 37680 48427 37680 48427 4 gnd
port 514 nsew
rlabel metal2 s 38448 48743 38448 48743 4 gnd
port 514 nsew
rlabel metal2 s 38928 47637 38928 47637 4 gnd
port 514 nsew
rlabel metal2 s 36432 49770 36432 49770 4 gnd
port 514 nsew
rlabel metal2 s 35184 47953 35184 47953 4 gnd
port 514 nsew
rlabel metal2 s 35184 49533 35184 49533 4 gnd
port 514 nsew
rlabel metal2 s 37200 47637 37200 47637 4 gnd
port 514 nsew
rlabel metal2 s 35184 48743 35184 48743 4 gnd
port 514 nsew
rlabel metal2 s 37200 48190 37200 48190 4 gnd
port 514 nsew
rlabel metal2 s 35184 47637 35184 47637 4 gnd
port 514 nsew
rlabel metal2 s 36432 47953 36432 47953 4 gnd
port 514 nsew
rlabel metal2 s 35184 50323 35184 50323 4 gnd
port 514 nsew
rlabel metal2 s 37200 50560 37200 50560 4 gnd
port 514 nsew
rlabel metal2 s 35952 49217 35952 49217 4 gnd
port 514 nsew
rlabel metal2 s 37200 49533 37200 49533 4 gnd
port 514 nsew
rlabel metal2 s 35184 48190 35184 48190 4 gnd
port 514 nsew
rlabel metal2 s 35952 49533 35952 49533 4 gnd
port 514 nsew
rlabel metal2 s 35184 50560 35184 50560 4 gnd
port 514 nsew
rlabel metal2 s 35952 50007 35952 50007 4 gnd
port 514 nsew
rlabel metal2 s 35184 48980 35184 48980 4 gnd
port 514 nsew
rlabel metal2 s 35952 50560 35952 50560 4 gnd
port 514 nsew
rlabel metal2 s 36432 47637 36432 47637 4 gnd
port 514 nsew
rlabel metal2 s 36432 49217 36432 49217 4 gnd
port 514 nsew
rlabel metal2 s 36432 49533 36432 49533 4 gnd
port 514 nsew
rlabel metal2 s 37200 48427 37200 48427 4 gnd
port 514 nsew
rlabel metal2 s 37200 50007 37200 50007 4 gnd
port 514 nsew
rlabel metal2 s 37200 48743 37200 48743 4 gnd
port 514 nsew
rlabel metal2 s 36432 50323 36432 50323 4 gnd
port 514 nsew
rlabel metal2 s 36432 48980 36432 48980 4 gnd
port 514 nsew
rlabel metal2 s 35952 50323 35952 50323 4 gnd
port 514 nsew
rlabel metal2 s 37200 48980 37200 48980 4 gnd
port 514 nsew
rlabel metal2 s 35952 48190 35952 48190 4 gnd
port 514 nsew
rlabel metal2 s 36432 50007 36432 50007 4 gnd
port 514 nsew
rlabel metal2 s 37200 49217 37200 49217 4 gnd
port 514 nsew
rlabel metal2 s 36432 48427 36432 48427 4 gnd
port 514 nsew
rlabel metal2 s 35184 48427 35184 48427 4 gnd
port 514 nsew
rlabel metal2 s 35952 49770 35952 49770 4 gnd
port 514 nsew
rlabel metal2 s 35184 49217 35184 49217 4 gnd
port 514 nsew
rlabel metal2 s 36432 50560 36432 50560 4 gnd
port 514 nsew
rlabel metal2 s 35952 47953 35952 47953 4 gnd
port 514 nsew
rlabel metal2 s 35952 48980 35952 48980 4 gnd
port 514 nsew
rlabel metal2 s 36432 48190 36432 48190 4 gnd
port 514 nsew
rlabel metal2 s 37200 50323 37200 50323 4 gnd
port 514 nsew
rlabel metal2 s 35952 47637 35952 47637 4 gnd
port 514 nsew
rlabel metal2 s 37200 47953 37200 47953 4 gnd
port 514 nsew
rlabel metal2 s 35184 49770 35184 49770 4 gnd
port 514 nsew
rlabel metal2 s 35952 48743 35952 48743 4 gnd
port 514 nsew
rlabel metal2 s 36432 48743 36432 48743 4 gnd
port 514 nsew
rlabel metal2 s 35952 48427 35952 48427 4 gnd
port 514 nsew
rlabel metal2 s 37200 49770 37200 49770 4 gnd
port 514 nsew
rlabel metal2 s 35184 50007 35184 50007 4 gnd
port 514 nsew
rlabel metal2 s 36432 47163 36432 47163 4 gnd
port 514 nsew
rlabel metal2 s 37200 47400 37200 47400 4 gnd
port 514 nsew
rlabel metal2 s 35184 46847 35184 46847 4 gnd
port 514 nsew
rlabel metal2 s 37200 45030 37200 45030 4 gnd
port 514 nsew
rlabel metal2 s 35184 46057 35184 46057 4 gnd
port 514 nsew
rlabel metal2 s 36432 44793 36432 44793 4 gnd
port 514 nsew
rlabel metal2 s 35952 45583 35952 45583 4 gnd
port 514 nsew
rlabel metal2 s 35952 44793 35952 44793 4 gnd
port 514 nsew
rlabel metal2 s 37200 46610 37200 46610 4 gnd
port 514 nsew
rlabel metal2 s 36432 45030 36432 45030 4 gnd
port 514 nsew
rlabel metal2 s 35184 45030 35184 45030 4 gnd
port 514 nsew
rlabel metal2 s 37200 44477 37200 44477 4 gnd
port 514 nsew
rlabel metal2 s 35952 46373 35952 46373 4 gnd
port 514 nsew
rlabel metal2 s 37200 47163 37200 47163 4 gnd
port 514 nsew
rlabel metal2 s 36432 45267 36432 45267 4 gnd
port 514 nsew
rlabel metal2 s 35952 47163 35952 47163 4 gnd
port 514 nsew
rlabel metal2 s 37200 45267 37200 45267 4 gnd
port 514 nsew
rlabel metal2 s 35952 47400 35952 47400 4 gnd
port 514 nsew
rlabel metal2 s 35952 45030 35952 45030 4 gnd
port 514 nsew
rlabel metal2 s 36432 46847 36432 46847 4 gnd
port 514 nsew
rlabel metal2 s 37200 45820 37200 45820 4 gnd
port 514 nsew
rlabel metal2 s 36432 46373 36432 46373 4 gnd
port 514 nsew
rlabel metal2 s 36432 45583 36432 45583 4 gnd
port 514 nsew
rlabel metal2 s 35184 46610 35184 46610 4 gnd
port 514 nsew
rlabel metal2 s 35952 45820 35952 45820 4 gnd
port 514 nsew
rlabel metal2 s 35184 45583 35184 45583 4 gnd
port 514 nsew
rlabel metal2 s 36432 47400 36432 47400 4 gnd
port 514 nsew
rlabel metal2 s 35952 46610 35952 46610 4 gnd
port 514 nsew
rlabel metal2 s 35184 46373 35184 46373 4 gnd
port 514 nsew
rlabel metal2 s 37200 44793 37200 44793 4 gnd
port 514 nsew
rlabel metal2 s 36432 45820 36432 45820 4 gnd
port 514 nsew
rlabel metal2 s 37200 46847 37200 46847 4 gnd
port 514 nsew
rlabel metal2 s 35952 45267 35952 45267 4 gnd
port 514 nsew
rlabel metal2 s 35952 46057 35952 46057 4 gnd
port 514 nsew
rlabel metal2 s 36432 46610 36432 46610 4 gnd
port 514 nsew
rlabel metal2 s 35184 45820 35184 45820 4 gnd
port 514 nsew
rlabel metal2 s 35184 45267 35184 45267 4 gnd
port 514 nsew
rlabel metal2 s 35184 44477 35184 44477 4 gnd
port 514 nsew
rlabel metal2 s 35184 47400 35184 47400 4 gnd
port 514 nsew
rlabel metal2 s 36432 46057 36432 46057 4 gnd
port 514 nsew
rlabel metal2 s 35952 46847 35952 46847 4 gnd
port 514 nsew
rlabel metal2 s 35184 44793 35184 44793 4 gnd
port 514 nsew
rlabel metal2 s 37200 46057 37200 46057 4 gnd
port 514 nsew
rlabel metal2 s 35184 47163 35184 47163 4 gnd
port 514 nsew
rlabel metal2 s 35952 44477 35952 44477 4 gnd
port 514 nsew
rlabel metal2 s 37200 46373 37200 46373 4 gnd
port 514 nsew
rlabel metal2 s 36432 44477 36432 44477 4 gnd
port 514 nsew
rlabel metal2 s 37200 45583 37200 45583 4 gnd
port 514 nsew
rlabel metal2 s 38448 47163 38448 47163 4 gnd
port 514 nsew
rlabel metal2 s 37680 47163 37680 47163 4 gnd
port 514 nsew
rlabel metal2 s 39696 46610 39696 46610 4 gnd
port 514 nsew
rlabel metal2 s 38928 44793 38928 44793 4 gnd
port 514 nsew
rlabel metal2 s 38448 44477 38448 44477 4 gnd
port 514 nsew
rlabel metal2 s 38448 45267 38448 45267 4 gnd
port 514 nsew
rlabel metal2 s 38928 46610 38928 46610 4 gnd
port 514 nsew
rlabel metal2 s 38448 46373 38448 46373 4 gnd
port 514 nsew
rlabel metal2 s 38448 46610 38448 46610 4 gnd
port 514 nsew
rlabel metal2 s 38928 46373 38928 46373 4 gnd
port 514 nsew
rlabel metal2 s 37680 45267 37680 45267 4 gnd
port 514 nsew
rlabel metal2 s 39696 44477 39696 44477 4 gnd
port 514 nsew
rlabel metal2 s 38448 44793 38448 44793 4 gnd
port 514 nsew
rlabel metal2 s 37680 45030 37680 45030 4 gnd
port 514 nsew
rlabel metal2 s 39696 45267 39696 45267 4 gnd
port 514 nsew
rlabel metal2 s 38928 45267 38928 45267 4 gnd
port 514 nsew
rlabel metal2 s 39696 47163 39696 47163 4 gnd
port 514 nsew
rlabel metal2 s 37680 44793 37680 44793 4 gnd
port 514 nsew
rlabel metal2 s 38928 46847 38928 46847 4 gnd
port 514 nsew
rlabel metal2 s 37680 47400 37680 47400 4 gnd
port 514 nsew
rlabel metal2 s 38448 45820 38448 45820 4 gnd
port 514 nsew
rlabel metal2 s 39696 45030 39696 45030 4 gnd
port 514 nsew
rlabel metal2 s 38448 45030 38448 45030 4 gnd
port 514 nsew
rlabel metal2 s 39696 45583 39696 45583 4 gnd
port 514 nsew
rlabel metal2 s 38448 46847 38448 46847 4 gnd
port 514 nsew
rlabel metal2 s 38448 46057 38448 46057 4 gnd
port 514 nsew
rlabel metal2 s 37680 46610 37680 46610 4 gnd
port 514 nsew
rlabel metal2 s 38928 45820 38928 45820 4 gnd
port 514 nsew
rlabel metal2 s 39696 46373 39696 46373 4 gnd
port 514 nsew
rlabel metal2 s 38928 47400 38928 47400 4 gnd
port 514 nsew
rlabel metal2 s 39696 46847 39696 46847 4 gnd
port 514 nsew
rlabel metal2 s 39696 44793 39696 44793 4 gnd
port 514 nsew
rlabel metal2 s 37680 45820 37680 45820 4 gnd
port 514 nsew
rlabel metal2 s 39696 47400 39696 47400 4 gnd
port 514 nsew
rlabel metal2 s 38448 47400 38448 47400 4 gnd
port 514 nsew
rlabel metal2 s 38448 45583 38448 45583 4 gnd
port 514 nsew
rlabel metal2 s 38928 44477 38928 44477 4 gnd
port 514 nsew
rlabel metal2 s 38928 46057 38928 46057 4 gnd
port 514 nsew
rlabel metal2 s 38928 45030 38928 45030 4 gnd
port 514 nsew
rlabel metal2 s 37680 46847 37680 46847 4 gnd
port 514 nsew
rlabel metal2 s 39696 45820 39696 45820 4 gnd
port 514 nsew
rlabel metal2 s 38928 47163 38928 47163 4 gnd
port 514 nsew
rlabel metal2 s 38928 45583 38928 45583 4 gnd
port 514 nsew
rlabel metal2 s 39696 46057 39696 46057 4 gnd
port 514 nsew
rlabel metal2 s 37680 46057 37680 46057 4 gnd
port 514 nsew
rlabel metal2 s 37680 46373 37680 46373 4 gnd
port 514 nsew
rlabel metal2 s 37680 44477 37680 44477 4 gnd
port 514 nsew
rlabel metal2 s 37680 45583 37680 45583 4 gnd
port 514 nsew
rlabel metal2 s 34704 48743 34704 48743 4 gnd
port 514 nsew
rlabel metal2 s 33936 49770 33936 49770 4 gnd
port 514 nsew
rlabel metal2 s 32688 49533 32688 49533 4 gnd
port 514 nsew
rlabel metal2 s 33936 48427 33936 48427 4 gnd
port 514 nsew
rlabel metal2 s 34704 49217 34704 49217 4 gnd
port 514 nsew
rlabel metal2 s 34704 48980 34704 48980 4 gnd
port 514 nsew
rlabel metal2 s 34704 50007 34704 50007 4 gnd
port 514 nsew
rlabel metal2 s 34704 47637 34704 47637 4 gnd
port 514 nsew
rlabel metal2 s 34704 48190 34704 48190 4 gnd
port 514 nsew
rlabel metal2 s 33936 48980 33936 48980 4 gnd
port 514 nsew
rlabel metal2 s 33456 47637 33456 47637 4 gnd
port 514 nsew
rlabel metal2 s 33456 47953 33456 47953 4 gnd
port 514 nsew
rlabel metal2 s 32688 48190 32688 48190 4 gnd
port 514 nsew
rlabel metal2 s 32688 49770 32688 49770 4 gnd
port 514 nsew
rlabel metal2 s 32688 48743 32688 48743 4 gnd
port 514 nsew
rlabel metal2 s 33456 49533 33456 49533 4 gnd
port 514 nsew
rlabel metal2 s 33936 47637 33936 47637 4 gnd
port 514 nsew
rlabel metal2 s 33456 50560 33456 50560 4 gnd
port 514 nsew
rlabel metal2 s 34704 49770 34704 49770 4 gnd
port 514 nsew
rlabel metal2 s 34704 48427 34704 48427 4 gnd
port 514 nsew
rlabel metal2 s 34704 50560 34704 50560 4 gnd
port 514 nsew
rlabel metal2 s 33456 49217 33456 49217 4 gnd
port 514 nsew
rlabel metal2 s 34704 47953 34704 47953 4 gnd
port 514 nsew
rlabel metal2 s 33936 50323 33936 50323 4 gnd
port 514 nsew
rlabel metal2 s 32688 50007 32688 50007 4 gnd
port 514 nsew
rlabel metal2 s 34704 50323 34704 50323 4 gnd
port 514 nsew
rlabel metal2 s 32688 48980 32688 48980 4 gnd
port 514 nsew
rlabel metal2 s 34704 49533 34704 49533 4 gnd
port 514 nsew
rlabel metal2 s 33456 48427 33456 48427 4 gnd
port 514 nsew
rlabel metal2 s 32688 47637 32688 47637 4 gnd
port 514 nsew
rlabel metal2 s 33456 50323 33456 50323 4 gnd
port 514 nsew
rlabel metal2 s 33936 47953 33936 47953 4 gnd
port 514 nsew
rlabel metal2 s 33936 48743 33936 48743 4 gnd
port 514 nsew
rlabel metal2 s 33456 48980 33456 48980 4 gnd
port 514 nsew
rlabel metal2 s 33936 48190 33936 48190 4 gnd
port 514 nsew
rlabel metal2 s 32688 47953 32688 47953 4 gnd
port 514 nsew
rlabel metal2 s 33456 49770 33456 49770 4 gnd
port 514 nsew
rlabel metal2 s 32688 50323 32688 50323 4 gnd
port 514 nsew
rlabel metal2 s 33936 49217 33936 49217 4 gnd
port 514 nsew
rlabel metal2 s 32688 50560 32688 50560 4 gnd
port 514 nsew
rlabel metal2 s 32688 48427 32688 48427 4 gnd
port 514 nsew
rlabel metal2 s 33456 50007 33456 50007 4 gnd
port 514 nsew
rlabel metal2 s 33456 48190 33456 48190 4 gnd
port 514 nsew
rlabel metal2 s 33936 50007 33936 50007 4 gnd
port 514 nsew
rlabel metal2 s 33936 49533 33936 49533 4 gnd
port 514 nsew
rlabel metal2 s 33936 50560 33936 50560 4 gnd
port 514 nsew
rlabel metal2 s 32688 49217 32688 49217 4 gnd
port 514 nsew
rlabel metal2 s 33456 48743 33456 48743 4 gnd
port 514 nsew
rlabel metal2 s 30192 50323 30192 50323 4 gnd
port 514 nsew
rlabel metal2 s 30192 49770 30192 49770 4 gnd
port 514 nsew
rlabel metal2 s 30960 49217 30960 49217 4 gnd
port 514 nsew
rlabel metal2 s 32208 50560 32208 50560 4 gnd
port 514 nsew
rlabel metal2 s 31440 49533 31440 49533 4 gnd
port 514 nsew
rlabel metal2 s 30960 47637 30960 47637 4 gnd
port 514 nsew
rlabel metal2 s 32208 48427 32208 48427 4 gnd
port 514 nsew
rlabel metal2 s 30960 47953 30960 47953 4 gnd
port 514 nsew
rlabel metal2 s 30960 48743 30960 48743 4 gnd
port 514 nsew
rlabel metal2 s 30960 49533 30960 49533 4 gnd
port 514 nsew
rlabel metal2 s 31440 50007 31440 50007 4 gnd
port 514 nsew
rlabel metal2 s 30960 50007 30960 50007 4 gnd
port 514 nsew
rlabel metal2 s 31440 48743 31440 48743 4 gnd
port 514 nsew
rlabel metal2 s 32208 50007 32208 50007 4 gnd
port 514 nsew
rlabel metal2 s 30192 50560 30192 50560 4 gnd
port 514 nsew
rlabel metal2 s 31440 48427 31440 48427 4 gnd
port 514 nsew
rlabel metal2 s 30960 48980 30960 48980 4 gnd
port 514 nsew
rlabel metal2 s 31440 49770 31440 49770 4 gnd
port 514 nsew
rlabel metal2 s 32208 48743 32208 48743 4 gnd
port 514 nsew
rlabel metal2 s 31440 47953 31440 47953 4 gnd
port 514 nsew
rlabel metal2 s 32208 49770 32208 49770 4 gnd
port 514 nsew
rlabel metal2 s 31440 49217 31440 49217 4 gnd
port 514 nsew
rlabel metal2 s 31440 50323 31440 50323 4 gnd
port 514 nsew
rlabel metal2 s 32208 48190 32208 48190 4 gnd
port 514 nsew
rlabel metal2 s 30960 49770 30960 49770 4 gnd
port 514 nsew
rlabel metal2 s 30192 48743 30192 48743 4 gnd
port 514 nsew
rlabel metal2 s 30192 49533 30192 49533 4 gnd
port 514 nsew
rlabel metal2 s 30192 48427 30192 48427 4 gnd
port 514 nsew
rlabel metal2 s 32208 49533 32208 49533 4 gnd
port 514 nsew
rlabel metal2 s 31440 50560 31440 50560 4 gnd
port 514 nsew
rlabel metal2 s 30192 48980 30192 48980 4 gnd
port 514 nsew
rlabel metal2 s 30960 48427 30960 48427 4 gnd
port 514 nsew
rlabel metal2 s 30192 47953 30192 47953 4 gnd
port 514 nsew
rlabel metal2 s 31440 48980 31440 48980 4 gnd
port 514 nsew
rlabel metal2 s 30192 48190 30192 48190 4 gnd
port 514 nsew
rlabel metal2 s 32208 48980 32208 48980 4 gnd
port 514 nsew
rlabel metal2 s 30960 50560 30960 50560 4 gnd
port 514 nsew
rlabel metal2 s 32208 49217 32208 49217 4 gnd
port 514 nsew
rlabel metal2 s 30960 48190 30960 48190 4 gnd
port 514 nsew
rlabel metal2 s 32208 47637 32208 47637 4 gnd
port 514 nsew
rlabel metal2 s 31440 47637 31440 47637 4 gnd
port 514 nsew
rlabel metal2 s 30192 49217 30192 49217 4 gnd
port 514 nsew
rlabel metal2 s 31440 48190 31440 48190 4 gnd
port 514 nsew
rlabel metal2 s 30192 50007 30192 50007 4 gnd
port 514 nsew
rlabel metal2 s 32208 47953 32208 47953 4 gnd
port 514 nsew
rlabel metal2 s 32208 50323 32208 50323 4 gnd
port 514 nsew
rlabel metal2 s 30960 50323 30960 50323 4 gnd
port 514 nsew
rlabel metal2 s 30192 47637 30192 47637 4 gnd
port 514 nsew
rlabel metal2 s 31440 47163 31440 47163 4 gnd
port 514 nsew
rlabel metal2 s 30192 46847 30192 46847 4 gnd
port 514 nsew
rlabel metal2 s 32208 45820 32208 45820 4 gnd
port 514 nsew
rlabel metal2 s 31440 46373 31440 46373 4 gnd
port 514 nsew
rlabel metal2 s 31440 44477 31440 44477 4 gnd
port 514 nsew
rlabel metal2 s 30960 46847 30960 46847 4 gnd
port 514 nsew
rlabel metal2 s 30960 45583 30960 45583 4 gnd
port 514 nsew
rlabel metal2 s 32208 46057 32208 46057 4 gnd
port 514 nsew
rlabel metal2 s 30960 47400 30960 47400 4 gnd
port 514 nsew
rlabel metal2 s 31440 45030 31440 45030 4 gnd
port 514 nsew
rlabel metal2 s 30192 47163 30192 47163 4 gnd
port 514 nsew
rlabel metal2 s 31440 45820 31440 45820 4 gnd
port 514 nsew
rlabel metal2 s 31440 45267 31440 45267 4 gnd
port 514 nsew
rlabel metal2 s 30192 44793 30192 44793 4 gnd
port 514 nsew
rlabel metal2 s 30192 46610 30192 46610 4 gnd
port 514 nsew
rlabel metal2 s 32208 46847 32208 46847 4 gnd
port 514 nsew
rlabel metal2 s 31440 45583 31440 45583 4 gnd
port 514 nsew
rlabel metal2 s 30960 46057 30960 46057 4 gnd
port 514 nsew
rlabel metal2 s 31440 46610 31440 46610 4 gnd
port 514 nsew
rlabel metal2 s 31440 47400 31440 47400 4 gnd
port 514 nsew
rlabel metal2 s 32208 47163 32208 47163 4 gnd
port 514 nsew
rlabel metal2 s 30192 45267 30192 45267 4 gnd
port 514 nsew
rlabel metal2 s 30960 47163 30960 47163 4 gnd
port 514 nsew
rlabel metal2 s 31440 46057 31440 46057 4 gnd
port 514 nsew
rlabel metal2 s 30192 46373 30192 46373 4 gnd
port 514 nsew
rlabel metal2 s 31440 46847 31440 46847 4 gnd
port 514 nsew
rlabel metal2 s 30960 45820 30960 45820 4 gnd
port 514 nsew
rlabel metal2 s 30192 44477 30192 44477 4 gnd
port 514 nsew
rlabel metal2 s 32208 46610 32208 46610 4 gnd
port 514 nsew
rlabel metal2 s 30960 46373 30960 46373 4 gnd
port 514 nsew
rlabel metal2 s 32208 45030 32208 45030 4 gnd
port 514 nsew
rlabel metal2 s 30192 45030 30192 45030 4 gnd
port 514 nsew
rlabel metal2 s 32208 45267 32208 45267 4 gnd
port 514 nsew
rlabel metal2 s 32208 44477 32208 44477 4 gnd
port 514 nsew
rlabel metal2 s 30192 47400 30192 47400 4 gnd
port 514 nsew
rlabel metal2 s 32208 45583 32208 45583 4 gnd
port 514 nsew
rlabel metal2 s 30960 44477 30960 44477 4 gnd
port 514 nsew
rlabel metal2 s 32208 46373 32208 46373 4 gnd
port 514 nsew
rlabel metal2 s 30960 44793 30960 44793 4 gnd
port 514 nsew
rlabel metal2 s 30960 45030 30960 45030 4 gnd
port 514 nsew
rlabel metal2 s 32208 44793 32208 44793 4 gnd
port 514 nsew
rlabel metal2 s 32208 47400 32208 47400 4 gnd
port 514 nsew
rlabel metal2 s 31440 44793 31440 44793 4 gnd
port 514 nsew
rlabel metal2 s 30192 45583 30192 45583 4 gnd
port 514 nsew
rlabel metal2 s 30960 46610 30960 46610 4 gnd
port 514 nsew
rlabel metal2 s 30960 45267 30960 45267 4 gnd
port 514 nsew
rlabel metal2 s 30192 46057 30192 46057 4 gnd
port 514 nsew
rlabel metal2 s 30192 45820 30192 45820 4 gnd
port 514 nsew
rlabel metal2 s 33936 44477 33936 44477 4 gnd
port 514 nsew
rlabel metal2 s 32688 46610 32688 46610 4 gnd
port 514 nsew
rlabel metal2 s 32688 47163 32688 47163 4 gnd
port 514 nsew
rlabel metal2 s 34704 45267 34704 45267 4 gnd
port 514 nsew
rlabel metal2 s 32688 46847 32688 46847 4 gnd
port 514 nsew
rlabel metal2 s 32688 44793 32688 44793 4 gnd
port 514 nsew
rlabel metal2 s 33936 47163 33936 47163 4 gnd
port 514 nsew
rlabel metal2 s 33456 46373 33456 46373 4 gnd
port 514 nsew
rlabel metal2 s 34704 44477 34704 44477 4 gnd
port 514 nsew
rlabel metal2 s 33936 44793 33936 44793 4 gnd
port 514 nsew
rlabel metal2 s 34704 45820 34704 45820 4 gnd
port 514 nsew
rlabel metal2 s 33936 46847 33936 46847 4 gnd
port 514 nsew
rlabel metal2 s 33456 45267 33456 45267 4 gnd
port 514 nsew
rlabel metal2 s 33936 45820 33936 45820 4 gnd
port 514 nsew
rlabel metal2 s 33936 46610 33936 46610 4 gnd
port 514 nsew
rlabel metal2 s 33456 47163 33456 47163 4 gnd
port 514 nsew
rlabel metal2 s 33936 46373 33936 46373 4 gnd
port 514 nsew
rlabel metal2 s 33456 45583 33456 45583 4 gnd
port 514 nsew
rlabel metal2 s 32688 45583 32688 45583 4 gnd
port 514 nsew
rlabel metal2 s 33936 45030 33936 45030 4 gnd
port 514 nsew
rlabel metal2 s 33936 47400 33936 47400 4 gnd
port 514 nsew
rlabel metal2 s 34704 44793 34704 44793 4 gnd
port 514 nsew
rlabel metal2 s 33456 45820 33456 45820 4 gnd
port 514 nsew
rlabel metal2 s 33456 46847 33456 46847 4 gnd
port 514 nsew
rlabel metal2 s 33936 46057 33936 46057 4 gnd
port 514 nsew
rlabel metal2 s 33456 47400 33456 47400 4 gnd
port 514 nsew
rlabel metal2 s 33456 45030 33456 45030 4 gnd
port 514 nsew
rlabel metal2 s 32688 45030 32688 45030 4 gnd
port 514 nsew
rlabel metal2 s 33936 45267 33936 45267 4 gnd
port 514 nsew
rlabel metal2 s 32688 46373 32688 46373 4 gnd
port 514 nsew
rlabel metal2 s 33456 46057 33456 46057 4 gnd
port 514 nsew
rlabel metal2 s 34704 45583 34704 45583 4 gnd
port 514 nsew
rlabel metal2 s 33456 44477 33456 44477 4 gnd
port 514 nsew
rlabel metal2 s 32688 44477 32688 44477 4 gnd
port 514 nsew
rlabel metal2 s 33456 46610 33456 46610 4 gnd
port 514 nsew
rlabel metal2 s 32688 46057 32688 46057 4 gnd
port 514 nsew
rlabel metal2 s 32688 45820 32688 45820 4 gnd
port 514 nsew
rlabel metal2 s 34704 47163 34704 47163 4 gnd
port 514 nsew
rlabel metal2 s 34704 45030 34704 45030 4 gnd
port 514 nsew
rlabel metal2 s 33936 45583 33936 45583 4 gnd
port 514 nsew
rlabel metal2 s 32688 45267 32688 45267 4 gnd
port 514 nsew
rlabel metal2 s 34704 46373 34704 46373 4 gnd
port 514 nsew
rlabel metal2 s 34704 46057 34704 46057 4 gnd
port 514 nsew
rlabel metal2 s 33456 44793 33456 44793 4 gnd
port 514 nsew
rlabel metal2 s 32688 47400 32688 47400 4 gnd
port 514 nsew
rlabel metal2 s 34704 46847 34704 46847 4 gnd
port 514 nsew
rlabel metal2 s 34704 46610 34704 46610 4 gnd
port 514 nsew
rlabel metal2 s 34704 47400 34704 47400 4 gnd
port 514 nsew
rlabel metal2 s 33456 41317 33456 41317 4 gnd
port 514 nsew
rlabel metal2 s 33936 41870 33936 41870 4 gnd
port 514 nsew
rlabel metal2 s 34704 41870 34704 41870 4 gnd
port 514 nsew
rlabel metal2 s 33936 43213 33936 43213 4 gnd
port 514 nsew
rlabel metal2 s 32688 42107 32688 42107 4 gnd
port 514 nsew
rlabel metal2 s 33936 41317 33936 41317 4 gnd
port 514 nsew
rlabel metal2 s 32688 44003 32688 44003 4 gnd
port 514 nsew
rlabel metal2 s 32688 42897 32688 42897 4 gnd
port 514 nsew
rlabel metal2 s 34704 42660 34704 42660 4 gnd
port 514 nsew
rlabel metal2 s 33456 43213 33456 43213 4 gnd
port 514 nsew
rlabel metal2 s 34704 42107 34704 42107 4 gnd
port 514 nsew
rlabel metal2 s 33936 42423 33936 42423 4 gnd
port 514 nsew
rlabel metal2 s 32688 41317 32688 41317 4 gnd
port 514 nsew
rlabel metal2 s 34704 44003 34704 44003 4 gnd
port 514 nsew
rlabel metal2 s 32688 43450 32688 43450 4 gnd
port 514 nsew
rlabel metal2 s 32688 41870 32688 41870 4 gnd
port 514 nsew
rlabel metal2 s 33456 42897 33456 42897 4 gnd
port 514 nsew
rlabel metal2 s 33456 44240 33456 44240 4 gnd
port 514 nsew
rlabel metal2 s 34704 43687 34704 43687 4 gnd
port 514 nsew
rlabel metal2 s 33456 43450 33456 43450 4 gnd
port 514 nsew
rlabel metal2 s 33456 43687 33456 43687 4 gnd
port 514 nsew
rlabel metal2 s 34704 43450 34704 43450 4 gnd
port 514 nsew
rlabel metal2 s 32688 43213 32688 43213 4 gnd
port 514 nsew
rlabel metal2 s 32688 43687 32688 43687 4 gnd
port 514 nsew
rlabel metal2 s 34704 42897 34704 42897 4 gnd
port 514 nsew
rlabel metal2 s 32688 42660 32688 42660 4 gnd
port 514 nsew
rlabel metal2 s 34704 41317 34704 41317 4 gnd
port 514 nsew
rlabel metal2 s 33936 44003 33936 44003 4 gnd
port 514 nsew
rlabel metal2 s 34704 43213 34704 43213 4 gnd
port 514 nsew
rlabel metal2 s 33936 41633 33936 41633 4 gnd
port 514 nsew
rlabel metal2 s 32688 42423 32688 42423 4 gnd
port 514 nsew
rlabel metal2 s 33456 41633 33456 41633 4 gnd
port 514 nsew
rlabel metal2 s 33936 44240 33936 44240 4 gnd
port 514 nsew
rlabel metal2 s 33456 42660 33456 42660 4 gnd
port 514 nsew
rlabel metal2 s 34704 42423 34704 42423 4 gnd
port 514 nsew
rlabel metal2 s 33936 42660 33936 42660 4 gnd
port 514 nsew
rlabel metal2 s 33456 42423 33456 42423 4 gnd
port 514 nsew
rlabel metal2 s 33936 42897 33936 42897 4 gnd
port 514 nsew
rlabel metal2 s 32688 41633 32688 41633 4 gnd
port 514 nsew
rlabel metal2 s 33936 42107 33936 42107 4 gnd
port 514 nsew
rlabel metal2 s 33936 43450 33936 43450 4 gnd
port 514 nsew
rlabel metal2 s 32688 44240 32688 44240 4 gnd
port 514 nsew
rlabel metal2 s 33456 44003 33456 44003 4 gnd
port 514 nsew
rlabel metal2 s 33456 42107 33456 42107 4 gnd
port 514 nsew
rlabel metal2 s 33456 41870 33456 41870 4 gnd
port 514 nsew
rlabel metal2 s 33936 43687 33936 43687 4 gnd
port 514 nsew
rlabel metal2 s 34704 41633 34704 41633 4 gnd
port 514 nsew
rlabel metal2 s 34704 44240 34704 44240 4 gnd
port 514 nsew
rlabel metal2 s 30192 42660 30192 42660 4 gnd
port 514 nsew
rlabel metal2 s 31440 43687 31440 43687 4 gnd
port 514 nsew
rlabel metal2 s 32208 42107 32208 42107 4 gnd
port 514 nsew
rlabel metal2 s 30960 43213 30960 43213 4 gnd
port 514 nsew
rlabel metal2 s 31440 42423 31440 42423 4 gnd
port 514 nsew
rlabel metal2 s 30960 42107 30960 42107 4 gnd
port 514 nsew
rlabel metal2 s 32208 42423 32208 42423 4 gnd
port 514 nsew
rlabel metal2 s 31440 44240 31440 44240 4 gnd
port 514 nsew
rlabel metal2 s 30960 44240 30960 44240 4 gnd
port 514 nsew
rlabel metal2 s 30960 41317 30960 41317 4 gnd
port 514 nsew
rlabel metal2 s 30960 41870 30960 41870 4 gnd
port 514 nsew
rlabel metal2 s 30960 44003 30960 44003 4 gnd
port 514 nsew
rlabel metal2 s 32208 43687 32208 43687 4 gnd
port 514 nsew
rlabel metal2 s 30192 44240 30192 44240 4 gnd
port 514 nsew
rlabel metal2 s 32208 41633 32208 41633 4 gnd
port 514 nsew
rlabel metal2 s 31440 41633 31440 41633 4 gnd
port 514 nsew
rlabel metal2 s 32208 44003 32208 44003 4 gnd
port 514 nsew
rlabel metal2 s 30192 44003 30192 44003 4 gnd
port 514 nsew
rlabel metal2 s 30960 42897 30960 42897 4 gnd
port 514 nsew
rlabel metal2 s 30960 41633 30960 41633 4 gnd
port 514 nsew
rlabel metal2 s 30192 41633 30192 41633 4 gnd
port 514 nsew
rlabel metal2 s 30192 43213 30192 43213 4 gnd
port 514 nsew
rlabel metal2 s 30960 43687 30960 43687 4 gnd
port 514 nsew
rlabel metal2 s 32208 42660 32208 42660 4 gnd
port 514 nsew
rlabel metal2 s 30192 43687 30192 43687 4 gnd
port 514 nsew
rlabel metal2 s 31440 43450 31440 43450 4 gnd
port 514 nsew
rlabel metal2 s 30960 42660 30960 42660 4 gnd
port 514 nsew
rlabel metal2 s 32208 42897 32208 42897 4 gnd
port 514 nsew
rlabel metal2 s 31440 43213 31440 43213 4 gnd
port 514 nsew
rlabel metal2 s 30960 42423 30960 42423 4 gnd
port 514 nsew
rlabel metal2 s 31440 42897 31440 42897 4 gnd
port 514 nsew
rlabel metal2 s 30192 42107 30192 42107 4 gnd
port 514 nsew
rlabel metal2 s 31440 41317 31440 41317 4 gnd
port 514 nsew
rlabel metal2 s 31440 42107 31440 42107 4 gnd
port 514 nsew
rlabel metal2 s 30192 41870 30192 41870 4 gnd
port 514 nsew
rlabel metal2 s 31440 44003 31440 44003 4 gnd
port 514 nsew
rlabel metal2 s 30192 41317 30192 41317 4 gnd
port 514 nsew
rlabel metal2 s 32208 43450 32208 43450 4 gnd
port 514 nsew
rlabel metal2 s 31440 42660 31440 42660 4 gnd
port 514 nsew
rlabel metal2 s 32208 41317 32208 41317 4 gnd
port 514 nsew
rlabel metal2 s 30192 43450 30192 43450 4 gnd
port 514 nsew
rlabel metal2 s 31440 41870 31440 41870 4 gnd
port 514 nsew
rlabel metal2 s 30192 42897 30192 42897 4 gnd
port 514 nsew
rlabel metal2 s 30192 42423 30192 42423 4 gnd
port 514 nsew
rlabel metal2 s 30960 43450 30960 43450 4 gnd
port 514 nsew
rlabel metal2 s 32208 44240 32208 44240 4 gnd
port 514 nsew
rlabel metal2 s 32208 41870 32208 41870 4 gnd
port 514 nsew
rlabel metal2 s 32208 43213 32208 43213 4 gnd
port 514 nsew
rlabel metal2 s 32208 40527 32208 40527 4 gnd
port 514 nsew
rlabel metal2 s 30192 39737 30192 39737 4 gnd
port 514 nsew
rlabel metal2 s 30192 40527 30192 40527 4 gnd
port 514 nsew
rlabel metal2 s 32208 41080 32208 41080 4 gnd
port 514 nsew
rlabel metal2 s 30960 38473 30960 38473 4 gnd
port 514 nsew
rlabel metal2 s 32208 40053 32208 40053 4 gnd
port 514 nsew
rlabel metal2 s 31440 38947 31440 38947 4 gnd
port 514 nsew
rlabel metal2 s 31440 40527 31440 40527 4 gnd
port 514 nsew
rlabel metal2 s 30960 39500 30960 39500 4 gnd
port 514 nsew
rlabel metal2 s 30960 39737 30960 39737 4 gnd
port 514 nsew
rlabel metal2 s 32208 38473 32208 38473 4 gnd
port 514 nsew
rlabel metal2 s 30960 41080 30960 41080 4 gnd
port 514 nsew
rlabel metal2 s 32208 39263 32208 39263 4 gnd
port 514 nsew
rlabel metal2 s 32208 38710 32208 38710 4 gnd
port 514 nsew
rlabel metal2 s 31440 39500 31440 39500 4 gnd
port 514 nsew
rlabel metal2 s 32208 40290 32208 40290 4 gnd
port 514 nsew
rlabel metal2 s 30960 39263 30960 39263 4 gnd
port 514 nsew
rlabel metal2 s 30192 39263 30192 39263 4 gnd
port 514 nsew
rlabel metal2 s 30960 40527 30960 40527 4 gnd
port 514 nsew
rlabel metal2 s 30960 40053 30960 40053 4 gnd
port 514 nsew
rlabel metal2 s 31440 38157 31440 38157 4 gnd
port 514 nsew
rlabel metal2 s 31440 38473 31440 38473 4 gnd
port 514 nsew
rlabel metal2 s 30192 39500 30192 39500 4 gnd
port 514 nsew
rlabel metal2 s 31440 39737 31440 39737 4 gnd
port 514 nsew
rlabel metal2 s 31440 40843 31440 40843 4 gnd
port 514 nsew
rlabel metal2 s 31440 38710 31440 38710 4 gnd
port 514 nsew
rlabel metal2 s 30192 38157 30192 38157 4 gnd
port 514 nsew
rlabel metal2 s 30192 38710 30192 38710 4 gnd
port 514 nsew
rlabel metal2 s 32208 39500 32208 39500 4 gnd
port 514 nsew
rlabel metal2 s 30192 38473 30192 38473 4 gnd
port 514 nsew
rlabel metal2 s 30960 38947 30960 38947 4 gnd
port 514 nsew
rlabel metal2 s 32208 40843 32208 40843 4 gnd
port 514 nsew
rlabel metal2 s 30960 38157 30960 38157 4 gnd
port 514 nsew
rlabel metal2 s 30960 40843 30960 40843 4 gnd
port 514 nsew
rlabel metal2 s 30960 40290 30960 40290 4 gnd
port 514 nsew
rlabel metal2 s 31440 40053 31440 40053 4 gnd
port 514 nsew
rlabel metal2 s 30192 38947 30192 38947 4 gnd
port 514 nsew
rlabel metal2 s 30960 38710 30960 38710 4 gnd
port 514 nsew
rlabel metal2 s 32208 39737 32208 39737 4 gnd
port 514 nsew
rlabel metal2 s 31440 40290 31440 40290 4 gnd
port 514 nsew
rlabel metal2 s 30192 40053 30192 40053 4 gnd
port 514 nsew
rlabel metal2 s 30192 40290 30192 40290 4 gnd
port 514 nsew
rlabel metal2 s 31440 39263 31440 39263 4 gnd
port 514 nsew
rlabel metal2 s 32208 38947 32208 38947 4 gnd
port 514 nsew
rlabel metal2 s 31440 41080 31440 41080 4 gnd
port 514 nsew
rlabel metal2 s 30192 40843 30192 40843 4 gnd
port 514 nsew
rlabel metal2 s 32208 38157 32208 38157 4 gnd
port 514 nsew
rlabel metal2 s 30192 41080 30192 41080 4 gnd
port 514 nsew
rlabel metal2 s 33456 39500 33456 39500 4 gnd
port 514 nsew
rlabel metal2 s 33456 41080 33456 41080 4 gnd
port 514 nsew
rlabel metal2 s 33936 40843 33936 40843 4 gnd
port 514 nsew
rlabel metal2 s 33456 38947 33456 38947 4 gnd
port 514 nsew
rlabel metal2 s 33456 38473 33456 38473 4 gnd
port 514 nsew
rlabel metal2 s 34704 39737 34704 39737 4 gnd
port 514 nsew
rlabel metal2 s 34704 41080 34704 41080 4 gnd
port 514 nsew
rlabel metal2 s 33936 40053 33936 40053 4 gnd
port 514 nsew
rlabel metal2 s 32688 39263 32688 39263 4 gnd
port 514 nsew
rlabel metal2 s 33456 40843 33456 40843 4 gnd
port 514 nsew
rlabel metal2 s 33456 39737 33456 39737 4 gnd
port 514 nsew
rlabel metal2 s 32688 38157 32688 38157 4 gnd
port 514 nsew
rlabel metal2 s 34704 39500 34704 39500 4 gnd
port 514 nsew
rlabel metal2 s 32688 40053 32688 40053 4 gnd
port 514 nsew
rlabel metal2 s 33936 39500 33936 39500 4 gnd
port 514 nsew
rlabel metal2 s 32688 38473 32688 38473 4 gnd
port 514 nsew
rlabel metal2 s 32688 40527 32688 40527 4 gnd
port 514 nsew
rlabel metal2 s 33456 38157 33456 38157 4 gnd
port 514 nsew
rlabel metal2 s 34704 39263 34704 39263 4 gnd
port 514 nsew
rlabel metal2 s 34704 38473 34704 38473 4 gnd
port 514 nsew
rlabel metal2 s 33936 40527 33936 40527 4 gnd
port 514 nsew
rlabel metal2 s 33456 38710 33456 38710 4 gnd
port 514 nsew
rlabel metal2 s 33936 38710 33936 38710 4 gnd
port 514 nsew
rlabel metal2 s 33936 39737 33936 39737 4 gnd
port 514 nsew
rlabel metal2 s 34704 40290 34704 40290 4 gnd
port 514 nsew
rlabel metal2 s 32688 39737 32688 39737 4 gnd
port 514 nsew
rlabel metal2 s 32688 38947 32688 38947 4 gnd
port 514 nsew
rlabel metal2 s 34704 38157 34704 38157 4 gnd
port 514 nsew
rlabel metal2 s 33936 40290 33936 40290 4 gnd
port 514 nsew
rlabel metal2 s 33936 41080 33936 41080 4 gnd
port 514 nsew
rlabel metal2 s 33456 39263 33456 39263 4 gnd
port 514 nsew
rlabel metal2 s 33456 40053 33456 40053 4 gnd
port 514 nsew
rlabel metal2 s 32688 38710 32688 38710 4 gnd
port 514 nsew
rlabel metal2 s 33456 40290 33456 40290 4 gnd
port 514 nsew
rlabel metal2 s 33456 40527 33456 40527 4 gnd
port 514 nsew
rlabel metal2 s 32688 40843 32688 40843 4 gnd
port 514 nsew
rlabel metal2 s 34704 38710 34704 38710 4 gnd
port 514 nsew
rlabel metal2 s 32688 39500 32688 39500 4 gnd
port 514 nsew
rlabel metal2 s 33936 38947 33936 38947 4 gnd
port 514 nsew
rlabel metal2 s 33936 39263 33936 39263 4 gnd
port 514 nsew
rlabel metal2 s 32688 41080 32688 41080 4 gnd
port 514 nsew
rlabel metal2 s 34704 40053 34704 40053 4 gnd
port 514 nsew
rlabel metal2 s 33936 38473 33936 38473 4 gnd
port 514 nsew
rlabel metal2 s 33936 38157 33936 38157 4 gnd
port 514 nsew
rlabel metal2 s 34704 38947 34704 38947 4 gnd
port 514 nsew
rlabel metal2 s 34704 40527 34704 40527 4 gnd
port 514 nsew
rlabel metal2 s 34704 40843 34704 40843 4 gnd
port 514 nsew
rlabel metal2 s 32688 40290 32688 40290 4 gnd
port 514 nsew
rlabel metal2 s 37680 42423 37680 42423 4 gnd
port 514 nsew
rlabel metal2 s 38928 43687 38928 43687 4 gnd
port 514 nsew
rlabel metal2 s 38448 43450 38448 43450 4 gnd
port 514 nsew
rlabel metal2 s 38448 43687 38448 43687 4 gnd
port 514 nsew
rlabel metal2 s 38928 41870 38928 41870 4 gnd
port 514 nsew
rlabel metal2 s 38448 42107 38448 42107 4 gnd
port 514 nsew
rlabel metal2 s 38928 42107 38928 42107 4 gnd
port 514 nsew
rlabel metal2 s 38928 43450 38928 43450 4 gnd
port 514 nsew
rlabel metal2 s 37680 43687 37680 43687 4 gnd
port 514 nsew
rlabel metal2 s 38928 42897 38928 42897 4 gnd
port 514 nsew
rlabel metal2 s 38928 44240 38928 44240 4 gnd
port 514 nsew
rlabel metal2 s 38928 42660 38928 42660 4 gnd
port 514 nsew
rlabel metal2 s 38928 44003 38928 44003 4 gnd
port 514 nsew
rlabel metal2 s 38448 43213 38448 43213 4 gnd
port 514 nsew
rlabel metal2 s 39696 43213 39696 43213 4 gnd
port 514 nsew
rlabel metal2 s 37680 44003 37680 44003 4 gnd
port 514 nsew
rlabel metal2 s 37680 43450 37680 43450 4 gnd
port 514 nsew
rlabel metal2 s 37680 44240 37680 44240 4 gnd
port 514 nsew
rlabel metal2 s 37680 41317 37680 41317 4 gnd
port 514 nsew
rlabel metal2 s 37680 42107 37680 42107 4 gnd
port 514 nsew
rlabel metal2 s 38448 42897 38448 42897 4 gnd
port 514 nsew
rlabel metal2 s 39696 43450 39696 43450 4 gnd
port 514 nsew
rlabel metal2 s 38448 41870 38448 41870 4 gnd
port 514 nsew
rlabel metal2 s 38928 41317 38928 41317 4 gnd
port 514 nsew
rlabel metal2 s 39696 43687 39696 43687 4 gnd
port 514 nsew
rlabel metal2 s 38448 42423 38448 42423 4 gnd
port 514 nsew
rlabel metal2 s 38448 41633 38448 41633 4 gnd
port 514 nsew
rlabel metal2 s 39696 44240 39696 44240 4 gnd
port 514 nsew
rlabel metal2 s 37680 43213 37680 43213 4 gnd
port 514 nsew
rlabel metal2 s 38448 42660 38448 42660 4 gnd
port 514 nsew
rlabel metal2 s 39696 41633 39696 41633 4 gnd
port 514 nsew
rlabel metal2 s 39696 42660 39696 42660 4 gnd
port 514 nsew
rlabel metal2 s 37680 42660 37680 42660 4 gnd
port 514 nsew
rlabel metal2 s 39696 42423 39696 42423 4 gnd
port 514 nsew
rlabel metal2 s 38928 42423 38928 42423 4 gnd
port 514 nsew
rlabel metal2 s 39696 42897 39696 42897 4 gnd
port 514 nsew
rlabel metal2 s 39696 42107 39696 42107 4 gnd
port 514 nsew
rlabel metal2 s 38928 41633 38928 41633 4 gnd
port 514 nsew
rlabel metal2 s 38928 43213 38928 43213 4 gnd
port 514 nsew
rlabel metal2 s 39696 44003 39696 44003 4 gnd
port 514 nsew
rlabel metal2 s 37680 42897 37680 42897 4 gnd
port 514 nsew
rlabel metal2 s 37680 41870 37680 41870 4 gnd
port 514 nsew
rlabel metal2 s 38448 41317 38448 41317 4 gnd
port 514 nsew
rlabel metal2 s 39696 41317 39696 41317 4 gnd
port 514 nsew
rlabel metal2 s 38448 44003 38448 44003 4 gnd
port 514 nsew
rlabel metal2 s 38448 44240 38448 44240 4 gnd
port 514 nsew
rlabel metal2 s 39696 41870 39696 41870 4 gnd
port 514 nsew
rlabel metal2 s 37680 41633 37680 41633 4 gnd
port 514 nsew
rlabel metal2 s 37200 42660 37200 42660 4 gnd
port 514 nsew
rlabel metal2 s 35952 41633 35952 41633 4 gnd
port 514 nsew
rlabel metal2 s 36432 41317 36432 41317 4 gnd
port 514 nsew
rlabel metal2 s 35184 44003 35184 44003 4 gnd
port 514 nsew
rlabel metal2 s 35184 42107 35184 42107 4 gnd
port 514 nsew
rlabel metal2 s 35952 41317 35952 41317 4 gnd
port 514 nsew
rlabel metal2 s 35952 42423 35952 42423 4 gnd
port 514 nsew
rlabel metal2 s 35184 41317 35184 41317 4 gnd
port 514 nsew
rlabel metal2 s 35952 43687 35952 43687 4 gnd
port 514 nsew
rlabel metal2 s 36432 42107 36432 42107 4 gnd
port 514 nsew
rlabel metal2 s 35952 42897 35952 42897 4 gnd
port 514 nsew
rlabel metal2 s 36432 42660 36432 42660 4 gnd
port 514 nsew
rlabel metal2 s 36432 42423 36432 42423 4 gnd
port 514 nsew
rlabel metal2 s 35184 43687 35184 43687 4 gnd
port 514 nsew
rlabel metal2 s 35184 43450 35184 43450 4 gnd
port 514 nsew
rlabel metal2 s 35952 43213 35952 43213 4 gnd
port 514 nsew
rlabel metal2 s 35184 42660 35184 42660 4 gnd
port 514 nsew
rlabel metal2 s 37200 43687 37200 43687 4 gnd
port 514 nsew
rlabel metal2 s 35952 44240 35952 44240 4 gnd
port 514 nsew
rlabel metal2 s 37200 42107 37200 42107 4 gnd
port 514 nsew
rlabel metal2 s 36432 44240 36432 44240 4 gnd
port 514 nsew
rlabel metal2 s 37200 41633 37200 41633 4 gnd
port 514 nsew
rlabel metal2 s 35184 43213 35184 43213 4 gnd
port 514 nsew
rlabel metal2 s 35184 42897 35184 42897 4 gnd
port 514 nsew
rlabel metal2 s 35952 44003 35952 44003 4 gnd
port 514 nsew
rlabel metal2 s 36432 44003 36432 44003 4 gnd
port 514 nsew
rlabel metal2 s 36432 42897 36432 42897 4 gnd
port 514 nsew
rlabel metal2 s 35952 42107 35952 42107 4 gnd
port 514 nsew
rlabel metal2 s 36432 43687 36432 43687 4 gnd
port 514 nsew
rlabel metal2 s 37200 43450 37200 43450 4 gnd
port 514 nsew
rlabel metal2 s 35184 41633 35184 41633 4 gnd
port 514 nsew
rlabel metal2 s 35184 42423 35184 42423 4 gnd
port 514 nsew
rlabel metal2 s 36432 41633 36432 41633 4 gnd
port 514 nsew
rlabel metal2 s 36432 43450 36432 43450 4 gnd
port 514 nsew
rlabel metal2 s 35184 41870 35184 41870 4 gnd
port 514 nsew
rlabel metal2 s 36432 41870 36432 41870 4 gnd
port 514 nsew
rlabel metal2 s 37200 42897 37200 42897 4 gnd
port 514 nsew
rlabel metal2 s 37200 44003 37200 44003 4 gnd
port 514 nsew
rlabel metal2 s 37200 44240 37200 44240 4 gnd
port 514 nsew
rlabel metal2 s 36432 43213 36432 43213 4 gnd
port 514 nsew
rlabel metal2 s 37200 41870 37200 41870 4 gnd
port 514 nsew
rlabel metal2 s 35952 41870 35952 41870 4 gnd
port 514 nsew
rlabel metal2 s 35952 42660 35952 42660 4 gnd
port 514 nsew
rlabel metal2 s 37200 42423 37200 42423 4 gnd
port 514 nsew
rlabel metal2 s 35184 44240 35184 44240 4 gnd
port 514 nsew
rlabel metal2 s 37200 41317 37200 41317 4 gnd
port 514 nsew
rlabel metal2 s 37200 43213 37200 43213 4 gnd
port 514 nsew
rlabel metal2 s 35952 43450 35952 43450 4 gnd
port 514 nsew
rlabel metal2 s 36432 39500 36432 39500 4 gnd
port 514 nsew
rlabel metal2 s 37200 41080 37200 41080 4 gnd
port 514 nsew
rlabel metal2 s 35952 40290 35952 40290 4 gnd
port 514 nsew
rlabel metal2 s 35184 40843 35184 40843 4 gnd
port 514 nsew
rlabel metal2 s 37200 38157 37200 38157 4 gnd
port 514 nsew
rlabel metal2 s 35184 38473 35184 38473 4 gnd
port 514 nsew
rlabel metal2 s 35952 41080 35952 41080 4 gnd
port 514 nsew
rlabel metal2 s 35184 40053 35184 40053 4 gnd
port 514 nsew
rlabel metal2 s 35952 39263 35952 39263 4 gnd
port 514 nsew
rlabel metal2 s 35952 38157 35952 38157 4 gnd
port 514 nsew
rlabel metal2 s 36432 39737 36432 39737 4 gnd
port 514 nsew
rlabel metal2 s 36432 39263 36432 39263 4 gnd
port 514 nsew
rlabel metal2 s 37200 40053 37200 40053 4 gnd
port 514 nsew
rlabel metal2 s 37200 40843 37200 40843 4 gnd
port 514 nsew
rlabel metal2 s 35952 38473 35952 38473 4 gnd
port 514 nsew
rlabel metal2 s 37200 39263 37200 39263 4 gnd
port 514 nsew
rlabel metal2 s 35184 38947 35184 38947 4 gnd
port 514 nsew
rlabel metal2 s 35952 40053 35952 40053 4 gnd
port 514 nsew
rlabel metal2 s 35184 39500 35184 39500 4 gnd
port 514 nsew
rlabel metal2 s 35184 40527 35184 40527 4 gnd
port 514 nsew
rlabel metal2 s 35184 39263 35184 39263 4 gnd
port 514 nsew
rlabel metal2 s 35952 40843 35952 40843 4 gnd
port 514 nsew
rlabel metal2 s 36432 40290 36432 40290 4 gnd
port 514 nsew
rlabel metal2 s 35952 38947 35952 38947 4 gnd
port 514 nsew
rlabel metal2 s 35952 39500 35952 39500 4 gnd
port 514 nsew
rlabel metal2 s 36432 38947 36432 38947 4 gnd
port 514 nsew
rlabel metal2 s 36432 38157 36432 38157 4 gnd
port 514 nsew
rlabel metal2 s 35184 38157 35184 38157 4 gnd
port 514 nsew
rlabel metal2 s 35184 40290 35184 40290 4 gnd
port 514 nsew
rlabel metal2 s 37200 40290 37200 40290 4 gnd
port 514 nsew
rlabel metal2 s 36432 38473 36432 38473 4 gnd
port 514 nsew
rlabel metal2 s 35952 38710 35952 38710 4 gnd
port 514 nsew
rlabel metal2 s 37200 38710 37200 38710 4 gnd
port 514 nsew
rlabel metal2 s 35184 38710 35184 38710 4 gnd
port 514 nsew
rlabel metal2 s 37200 39500 37200 39500 4 gnd
port 514 nsew
rlabel metal2 s 37200 38947 37200 38947 4 gnd
port 514 nsew
rlabel metal2 s 36432 40053 36432 40053 4 gnd
port 514 nsew
rlabel metal2 s 35952 39737 35952 39737 4 gnd
port 514 nsew
rlabel metal2 s 35184 39737 35184 39737 4 gnd
port 514 nsew
rlabel metal2 s 36432 40843 36432 40843 4 gnd
port 514 nsew
rlabel metal2 s 35952 40527 35952 40527 4 gnd
port 514 nsew
rlabel metal2 s 35184 41080 35184 41080 4 gnd
port 514 nsew
rlabel metal2 s 36432 41080 36432 41080 4 gnd
port 514 nsew
rlabel metal2 s 36432 40527 36432 40527 4 gnd
port 514 nsew
rlabel metal2 s 37200 39737 37200 39737 4 gnd
port 514 nsew
rlabel metal2 s 37200 38473 37200 38473 4 gnd
port 514 nsew
rlabel metal2 s 36432 38710 36432 38710 4 gnd
port 514 nsew
rlabel metal2 s 37200 40527 37200 40527 4 gnd
port 514 nsew
rlabel metal2 s 38448 41080 38448 41080 4 gnd
port 514 nsew
rlabel metal2 s 39696 39500 39696 39500 4 gnd
port 514 nsew
rlabel metal2 s 39696 38710 39696 38710 4 gnd
port 514 nsew
rlabel metal2 s 39696 38473 39696 38473 4 gnd
port 514 nsew
rlabel metal2 s 38928 40843 38928 40843 4 gnd
port 514 nsew
rlabel metal2 s 38448 40527 38448 40527 4 gnd
port 514 nsew
rlabel metal2 s 37680 38947 37680 38947 4 gnd
port 514 nsew
rlabel metal2 s 38448 39263 38448 39263 4 gnd
port 514 nsew
rlabel metal2 s 38928 38710 38928 38710 4 gnd
port 514 nsew
rlabel metal2 s 38928 41080 38928 41080 4 gnd
port 514 nsew
rlabel metal2 s 38448 39500 38448 39500 4 gnd
port 514 nsew
rlabel metal2 s 38448 40290 38448 40290 4 gnd
port 514 nsew
rlabel metal2 s 37680 40527 37680 40527 4 gnd
port 514 nsew
rlabel metal2 s 38928 38947 38928 38947 4 gnd
port 514 nsew
rlabel metal2 s 37680 40053 37680 40053 4 gnd
port 514 nsew
rlabel metal2 s 38448 38157 38448 38157 4 gnd
port 514 nsew
rlabel metal2 s 37680 38473 37680 38473 4 gnd
port 514 nsew
rlabel metal2 s 37680 38157 37680 38157 4 gnd
port 514 nsew
rlabel metal2 s 37680 39500 37680 39500 4 gnd
port 514 nsew
rlabel metal2 s 38928 39737 38928 39737 4 gnd
port 514 nsew
rlabel metal2 s 38928 39500 38928 39500 4 gnd
port 514 nsew
rlabel metal2 s 39696 41080 39696 41080 4 gnd
port 514 nsew
rlabel metal2 s 38448 40053 38448 40053 4 gnd
port 514 nsew
rlabel metal2 s 39696 40290 39696 40290 4 gnd
port 514 nsew
rlabel metal2 s 38928 38157 38928 38157 4 gnd
port 514 nsew
rlabel metal2 s 38448 38947 38448 38947 4 gnd
port 514 nsew
rlabel metal2 s 38448 39737 38448 39737 4 gnd
port 514 nsew
rlabel metal2 s 37680 38710 37680 38710 4 gnd
port 514 nsew
rlabel metal2 s 38448 40843 38448 40843 4 gnd
port 514 nsew
rlabel metal2 s 39696 40527 39696 40527 4 gnd
port 514 nsew
rlabel metal2 s 37680 41080 37680 41080 4 gnd
port 514 nsew
rlabel metal2 s 39696 38947 39696 38947 4 gnd
port 514 nsew
rlabel metal2 s 38448 38710 38448 38710 4 gnd
port 514 nsew
rlabel metal2 s 38928 40527 38928 40527 4 gnd
port 514 nsew
rlabel metal2 s 38448 38473 38448 38473 4 gnd
port 514 nsew
rlabel metal2 s 39696 39263 39696 39263 4 gnd
port 514 nsew
rlabel metal2 s 39696 40843 39696 40843 4 gnd
port 514 nsew
rlabel metal2 s 37680 40290 37680 40290 4 gnd
port 514 nsew
rlabel metal2 s 37680 39737 37680 39737 4 gnd
port 514 nsew
rlabel metal2 s 39696 39737 39696 39737 4 gnd
port 514 nsew
rlabel metal2 s 39696 38157 39696 38157 4 gnd
port 514 nsew
rlabel metal2 s 37680 39263 37680 39263 4 gnd
port 514 nsew
rlabel metal2 s 38928 40290 38928 40290 4 gnd
port 514 nsew
rlabel metal2 s 38928 40053 38928 40053 4 gnd
port 514 nsew
rlabel metal2 s 37680 40843 37680 40843 4 gnd
port 514 nsew
rlabel metal2 s 39696 40053 39696 40053 4 gnd
port 514 nsew
rlabel metal2 s 38928 39263 38928 39263 4 gnd
port 514 nsew
rlabel metal2 s 38928 38473 38928 38473 4 gnd
port 514 nsew
rlabel metal2 s 27696 50007 27696 50007 4 gnd
port 514 nsew
rlabel metal2 s 29712 47637 29712 47637 4 gnd
port 514 nsew
rlabel metal2 s 27696 47953 27696 47953 4 gnd
port 514 nsew
rlabel metal2 s 28944 50007 28944 50007 4 gnd
port 514 nsew
rlabel metal2 s 29712 50323 29712 50323 4 gnd
port 514 nsew
rlabel metal2 s 28944 50323 28944 50323 4 gnd
port 514 nsew
rlabel metal2 s 29712 48743 29712 48743 4 gnd
port 514 nsew
rlabel metal2 s 28464 48427 28464 48427 4 gnd
port 514 nsew
rlabel metal2 s 27696 50560 27696 50560 4 gnd
port 514 nsew
rlabel metal2 s 28464 47637 28464 47637 4 gnd
port 514 nsew
rlabel metal2 s 27696 50323 27696 50323 4 gnd
port 514 nsew
rlabel metal2 s 28944 48190 28944 48190 4 gnd
port 514 nsew
rlabel metal2 s 27696 48980 27696 48980 4 gnd
port 514 nsew
rlabel metal2 s 29712 47953 29712 47953 4 gnd
port 514 nsew
rlabel metal2 s 27696 47637 27696 47637 4 gnd
port 514 nsew
rlabel metal2 s 28944 47637 28944 47637 4 gnd
port 514 nsew
rlabel metal2 s 29712 48190 29712 48190 4 gnd
port 514 nsew
rlabel metal2 s 29712 49217 29712 49217 4 gnd
port 514 nsew
rlabel metal2 s 29712 48980 29712 48980 4 gnd
port 514 nsew
rlabel metal2 s 28944 48980 28944 48980 4 gnd
port 514 nsew
rlabel metal2 s 28464 48190 28464 48190 4 gnd
port 514 nsew
rlabel metal2 s 28464 48743 28464 48743 4 gnd
port 514 nsew
rlabel metal2 s 29712 48427 29712 48427 4 gnd
port 514 nsew
rlabel metal2 s 28464 50323 28464 50323 4 gnd
port 514 nsew
rlabel metal2 s 28944 48743 28944 48743 4 gnd
port 514 nsew
rlabel metal2 s 28944 49533 28944 49533 4 gnd
port 514 nsew
rlabel metal2 s 28464 49533 28464 49533 4 gnd
port 514 nsew
rlabel metal2 s 28464 49770 28464 49770 4 gnd
port 514 nsew
rlabel metal2 s 28944 49770 28944 49770 4 gnd
port 514 nsew
rlabel metal2 s 28464 50560 28464 50560 4 gnd
port 514 nsew
rlabel metal2 s 29712 50007 29712 50007 4 gnd
port 514 nsew
rlabel metal2 s 28464 50007 28464 50007 4 gnd
port 514 nsew
rlabel metal2 s 28464 48980 28464 48980 4 gnd
port 514 nsew
rlabel metal2 s 27696 48743 27696 48743 4 gnd
port 514 nsew
rlabel metal2 s 27696 48190 27696 48190 4 gnd
port 514 nsew
rlabel metal2 s 28944 47953 28944 47953 4 gnd
port 514 nsew
rlabel metal2 s 28464 47953 28464 47953 4 gnd
port 514 nsew
rlabel metal2 s 29712 49770 29712 49770 4 gnd
port 514 nsew
rlabel metal2 s 29712 50560 29712 50560 4 gnd
port 514 nsew
rlabel metal2 s 29712 49533 29712 49533 4 gnd
port 514 nsew
rlabel metal2 s 27696 49770 27696 49770 4 gnd
port 514 nsew
rlabel metal2 s 28944 48427 28944 48427 4 gnd
port 514 nsew
rlabel metal2 s 27696 48427 27696 48427 4 gnd
port 514 nsew
rlabel metal2 s 28944 50560 28944 50560 4 gnd
port 514 nsew
rlabel metal2 s 27696 49217 27696 49217 4 gnd
port 514 nsew
rlabel metal2 s 28464 49217 28464 49217 4 gnd
port 514 nsew
rlabel metal2 s 28944 49217 28944 49217 4 gnd
port 514 nsew
rlabel metal2 s 27696 49533 27696 49533 4 gnd
port 514 nsew
rlabel metal2 s 25200 50007 25200 50007 4 gnd
port 514 nsew
rlabel metal2 s 26448 49217 26448 49217 4 gnd
port 514 nsew
rlabel metal2 s 25200 49770 25200 49770 4 gnd
port 514 nsew
rlabel metal2 s 25200 50323 25200 50323 4 gnd
port 514 nsew
rlabel metal2 s 27216 49217 27216 49217 4 gnd
port 514 nsew
rlabel metal2 s 27216 49770 27216 49770 4 gnd
port 514 nsew
rlabel metal2 s 25200 49217 25200 49217 4 gnd
port 514 nsew
rlabel metal2 s 27216 50560 27216 50560 4 gnd
port 514 nsew
rlabel metal2 s 25200 48980 25200 48980 4 gnd
port 514 nsew
rlabel metal2 s 25200 48427 25200 48427 4 gnd
port 514 nsew
rlabel metal2 s 25968 48743 25968 48743 4 gnd
port 514 nsew
rlabel metal2 s 25200 49533 25200 49533 4 gnd
port 514 nsew
rlabel metal2 s 25968 49217 25968 49217 4 gnd
port 514 nsew
rlabel metal2 s 25968 48980 25968 48980 4 gnd
port 514 nsew
rlabel metal2 s 25968 50007 25968 50007 4 gnd
port 514 nsew
rlabel metal2 s 27216 48743 27216 48743 4 gnd
port 514 nsew
rlabel metal2 s 26448 48743 26448 48743 4 gnd
port 514 nsew
rlabel metal2 s 27216 50323 27216 50323 4 gnd
port 514 nsew
rlabel metal2 s 25200 50560 25200 50560 4 gnd
port 514 nsew
rlabel metal2 s 26448 50323 26448 50323 4 gnd
port 514 nsew
rlabel metal2 s 26448 49533 26448 49533 4 gnd
port 514 nsew
rlabel metal2 s 26448 50007 26448 50007 4 gnd
port 514 nsew
rlabel metal2 s 25968 50560 25968 50560 4 gnd
port 514 nsew
rlabel metal2 s 27216 49533 27216 49533 4 gnd
port 514 nsew
rlabel metal2 s 25968 50323 25968 50323 4 gnd
port 514 nsew
rlabel metal2 s 26448 47953 26448 47953 4 gnd
port 514 nsew
rlabel metal2 s 26448 50560 26448 50560 4 gnd
port 514 nsew
rlabel metal2 s 25200 47637 25200 47637 4 gnd
port 514 nsew
rlabel metal2 s 27216 50007 27216 50007 4 gnd
port 514 nsew
rlabel metal2 s 27216 48190 27216 48190 4 gnd
port 514 nsew
rlabel metal2 s 27216 48980 27216 48980 4 gnd
port 514 nsew
rlabel metal2 s 26448 48190 26448 48190 4 gnd
port 514 nsew
rlabel metal2 s 25968 47637 25968 47637 4 gnd
port 514 nsew
rlabel metal2 s 26448 47637 26448 47637 4 gnd
port 514 nsew
rlabel metal2 s 27216 47637 27216 47637 4 gnd
port 514 nsew
rlabel metal2 s 25200 48743 25200 48743 4 gnd
port 514 nsew
rlabel metal2 s 27216 47953 27216 47953 4 gnd
port 514 nsew
rlabel metal2 s 25968 47953 25968 47953 4 gnd
port 514 nsew
rlabel metal2 s 27216 48427 27216 48427 4 gnd
port 514 nsew
rlabel metal2 s 25200 47953 25200 47953 4 gnd
port 514 nsew
rlabel metal2 s 26448 48427 26448 48427 4 gnd
port 514 nsew
rlabel metal2 s 25968 48190 25968 48190 4 gnd
port 514 nsew
rlabel metal2 s 26448 48980 26448 48980 4 gnd
port 514 nsew
rlabel metal2 s 25200 48190 25200 48190 4 gnd
port 514 nsew
rlabel metal2 s 25968 48427 25968 48427 4 gnd
port 514 nsew
rlabel metal2 s 26448 49770 26448 49770 4 gnd
port 514 nsew
rlabel metal2 s 25968 49533 25968 49533 4 gnd
port 514 nsew
rlabel metal2 s 25968 49770 25968 49770 4 gnd
port 514 nsew
rlabel metal2 s 26448 47163 26448 47163 4 gnd
port 514 nsew
rlabel metal2 s 27216 46610 27216 46610 4 gnd
port 514 nsew
rlabel metal2 s 26448 47400 26448 47400 4 gnd
port 514 nsew
rlabel metal2 s 25200 44793 25200 44793 4 gnd
port 514 nsew
rlabel metal2 s 25968 46373 25968 46373 4 gnd
port 514 nsew
rlabel metal2 s 25968 46610 25968 46610 4 gnd
port 514 nsew
rlabel metal2 s 25968 44793 25968 44793 4 gnd
port 514 nsew
rlabel metal2 s 27216 45820 27216 45820 4 gnd
port 514 nsew
rlabel metal2 s 26448 46847 26448 46847 4 gnd
port 514 nsew
rlabel metal2 s 26448 44477 26448 44477 4 gnd
port 514 nsew
rlabel metal2 s 25200 45820 25200 45820 4 gnd
port 514 nsew
rlabel metal2 s 27216 46373 27216 46373 4 gnd
port 514 nsew
rlabel metal2 s 26448 45583 26448 45583 4 gnd
port 514 nsew
rlabel metal2 s 26448 45267 26448 45267 4 gnd
port 514 nsew
rlabel metal2 s 26448 46057 26448 46057 4 gnd
port 514 nsew
rlabel metal2 s 25200 46373 25200 46373 4 gnd
port 514 nsew
rlabel metal2 s 25968 44477 25968 44477 4 gnd
port 514 nsew
rlabel metal2 s 27216 46847 27216 46847 4 gnd
port 514 nsew
rlabel metal2 s 25200 47163 25200 47163 4 gnd
port 514 nsew
rlabel metal2 s 27216 45583 27216 45583 4 gnd
port 514 nsew
rlabel metal2 s 27216 47400 27216 47400 4 gnd
port 514 nsew
rlabel metal2 s 25200 46057 25200 46057 4 gnd
port 514 nsew
rlabel metal2 s 25968 45583 25968 45583 4 gnd
port 514 nsew
rlabel metal2 s 25968 45820 25968 45820 4 gnd
port 514 nsew
rlabel metal2 s 25968 47400 25968 47400 4 gnd
port 514 nsew
rlabel metal2 s 26448 45030 26448 45030 4 gnd
port 514 nsew
rlabel metal2 s 25200 44477 25200 44477 4 gnd
port 514 nsew
rlabel metal2 s 27216 45267 27216 45267 4 gnd
port 514 nsew
rlabel metal2 s 26448 46610 26448 46610 4 gnd
port 514 nsew
rlabel metal2 s 27216 45030 27216 45030 4 gnd
port 514 nsew
rlabel metal2 s 26448 45820 26448 45820 4 gnd
port 514 nsew
rlabel metal2 s 27216 44477 27216 44477 4 gnd
port 514 nsew
rlabel metal2 s 25968 45030 25968 45030 4 gnd
port 514 nsew
rlabel metal2 s 25200 47400 25200 47400 4 gnd
port 514 nsew
rlabel metal2 s 25968 45267 25968 45267 4 gnd
port 514 nsew
rlabel metal2 s 25968 46057 25968 46057 4 gnd
port 514 nsew
rlabel metal2 s 27216 46057 27216 46057 4 gnd
port 514 nsew
rlabel metal2 s 27216 44793 27216 44793 4 gnd
port 514 nsew
rlabel metal2 s 26448 44793 26448 44793 4 gnd
port 514 nsew
rlabel metal2 s 25200 46847 25200 46847 4 gnd
port 514 nsew
rlabel metal2 s 25200 45030 25200 45030 4 gnd
port 514 nsew
rlabel metal2 s 25200 45267 25200 45267 4 gnd
port 514 nsew
rlabel metal2 s 27216 47163 27216 47163 4 gnd
port 514 nsew
rlabel metal2 s 25200 45583 25200 45583 4 gnd
port 514 nsew
rlabel metal2 s 25968 46847 25968 46847 4 gnd
port 514 nsew
rlabel metal2 s 25200 46610 25200 46610 4 gnd
port 514 nsew
rlabel metal2 s 25968 47163 25968 47163 4 gnd
port 514 nsew
rlabel metal2 s 26448 46373 26448 46373 4 gnd
port 514 nsew
rlabel metal2 s 28944 47163 28944 47163 4 gnd
port 514 nsew
rlabel metal2 s 28944 47400 28944 47400 4 gnd
port 514 nsew
rlabel metal2 s 28944 45267 28944 45267 4 gnd
port 514 nsew
rlabel metal2 s 28944 44477 28944 44477 4 gnd
port 514 nsew
rlabel metal2 s 29712 47400 29712 47400 4 gnd
port 514 nsew
rlabel metal2 s 27696 47400 27696 47400 4 gnd
port 514 nsew
rlabel metal2 s 28464 44793 28464 44793 4 gnd
port 514 nsew
rlabel metal2 s 29712 46610 29712 46610 4 gnd
port 514 nsew
rlabel metal2 s 28944 45030 28944 45030 4 gnd
port 514 nsew
rlabel metal2 s 28464 47400 28464 47400 4 gnd
port 514 nsew
rlabel metal2 s 28464 46057 28464 46057 4 gnd
port 514 nsew
rlabel metal2 s 29712 45030 29712 45030 4 gnd
port 514 nsew
rlabel metal2 s 28944 46847 28944 46847 4 gnd
port 514 nsew
rlabel metal2 s 29712 47163 29712 47163 4 gnd
port 514 nsew
rlabel metal2 s 27696 45583 27696 45583 4 gnd
port 514 nsew
rlabel metal2 s 28944 45583 28944 45583 4 gnd
port 514 nsew
rlabel metal2 s 28464 45583 28464 45583 4 gnd
port 514 nsew
rlabel metal2 s 28464 45030 28464 45030 4 gnd
port 514 nsew
rlabel metal2 s 29712 46847 29712 46847 4 gnd
port 514 nsew
rlabel metal2 s 28944 46610 28944 46610 4 gnd
port 514 nsew
rlabel metal2 s 28464 46847 28464 46847 4 gnd
port 514 nsew
rlabel metal2 s 29712 44793 29712 44793 4 gnd
port 514 nsew
rlabel metal2 s 27696 46373 27696 46373 4 gnd
port 514 nsew
rlabel metal2 s 29712 45583 29712 45583 4 gnd
port 514 nsew
rlabel metal2 s 29712 46057 29712 46057 4 gnd
port 514 nsew
rlabel metal2 s 27696 45030 27696 45030 4 gnd
port 514 nsew
rlabel metal2 s 28464 45267 28464 45267 4 gnd
port 514 nsew
rlabel metal2 s 27696 46610 27696 46610 4 gnd
port 514 nsew
rlabel metal2 s 27696 45820 27696 45820 4 gnd
port 514 nsew
rlabel metal2 s 27696 44793 27696 44793 4 gnd
port 514 nsew
rlabel metal2 s 28464 47163 28464 47163 4 gnd
port 514 nsew
rlabel metal2 s 29712 45820 29712 45820 4 gnd
port 514 nsew
rlabel metal2 s 29712 46373 29712 46373 4 gnd
port 514 nsew
rlabel metal2 s 27696 46057 27696 46057 4 gnd
port 514 nsew
rlabel metal2 s 28464 45820 28464 45820 4 gnd
port 514 nsew
rlabel metal2 s 28944 46057 28944 46057 4 gnd
port 514 nsew
rlabel metal2 s 28464 46373 28464 46373 4 gnd
port 514 nsew
rlabel metal2 s 28944 45820 28944 45820 4 gnd
port 514 nsew
rlabel metal2 s 27696 46847 27696 46847 4 gnd
port 514 nsew
rlabel metal2 s 27696 45267 27696 45267 4 gnd
port 514 nsew
rlabel metal2 s 29712 44477 29712 44477 4 gnd
port 514 nsew
rlabel metal2 s 29712 45267 29712 45267 4 gnd
port 514 nsew
rlabel metal2 s 27696 47163 27696 47163 4 gnd
port 514 nsew
rlabel metal2 s 28464 46610 28464 46610 4 gnd
port 514 nsew
rlabel metal2 s 28944 46373 28944 46373 4 gnd
port 514 nsew
rlabel metal2 s 28464 44477 28464 44477 4 gnd
port 514 nsew
rlabel metal2 s 28944 44793 28944 44793 4 gnd
port 514 nsew
rlabel metal2 s 27696 44477 27696 44477 4 gnd
port 514 nsew
rlabel metal2 s 23472 49770 23472 49770 4 gnd
port 514 nsew
rlabel metal2 s 23952 49770 23952 49770 4 gnd
port 514 nsew
rlabel metal2 s 22704 48190 22704 48190 4 gnd
port 514 nsew
rlabel metal2 s 22704 49533 22704 49533 4 gnd
port 514 nsew
rlabel metal2 s 23472 50560 23472 50560 4 gnd
port 514 nsew
rlabel metal2 s 24720 49770 24720 49770 4 gnd
port 514 nsew
rlabel metal2 s 23472 50323 23472 50323 4 gnd
port 514 nsew
rlabel metal2 s 24720 50323 24720 50323 4 gnd
port 514 nsew
rlabel metal2 s 23472 50007 23472 50007 4 gnd
port 514 nsew
rlabel metal2 s 22704 47953 22704 47953 4 gnd
port 514 nsew
rlabel metal2 s 24720 49217 24720 49217 4 gnd
port 514 nsew
rlabel metal2 s 23952 48190 23952 48190 4 gnd
port 514 nsew
rlabel metal2 s 24720 48427 24720 48427 4 gnd
port 514 nsew
rlabel metal2 s 22704 48743 22704 48743 4 gnd
port 514 nsew
rlabel metal2 s 24720 47953 24720 47953 4 gnd
port 514 nsew
rlabel metal2 s 22704 49217 22704 49217 4 gnd
port 514 nsew
rlabel metal2 s 23472 48743 23472 48743 4 gnd
port 514 nsew
rlabel metal2 s 22704 50560 22704 50560 4 gnd
port 514 nsew
rlabel metal2 s 24720 48980 24720 48980 4 gnd
port 514 nsew
rlabel metal2 s 23952 48743 23952 48743 4 gnd
port 514 nsew
rlabel metal2 s 23952 49217 23952 49217 4 gnd
port 514 nsew
rlabel metal2 s 22704 49770 22704 49770 4 gnd
port 514 nsew
rlabel metal2 s 24720 50007 24720 50007 4 gnd
port 514 nsew
rlabel metal2 s 23952 47953 23952 47953 4 gnd
port 514 nsew
rlabel metal2 s 22704 47637 22704 47637 4 gnd
port 514 nsew
rlabel metal2 s 24720 47637 24720 47637 4 gnd
port 514 nsew
rlabel metal2 s 23472 48980 23472 48980 4 gnd
port 514 nsew
rlabel metal2 s 24720 48743 24720 48743 4 gnd
port 514 nsew
rlabel metal2 s 23952 48980 23952 48980 4 gnd
port 514 nsew
rlabel metal2 s 24720 49533 24720 49533 4 gnd
port 514 nsew
rlabel metal2 s 23472 49217 23472 49217 4 gnd
port 514 nsew
rlabel metal2 s 23952 48427 23952 48427 4 gnd
port 514 nsew
rlabel metal2 s 22704 48427 22704 48427 4 gnd
port 514 nsew
rlabel metal2 s 22704 50007 22704 50007 4 gnd
port 514 nsew
rlabel metal2 s 23952 50007 23952 50007 4 gnd
port 514 nsew
rlabel metal2 s 23472 47953 23472 47953 4 gnd
port 514 nsew
rlabel metal2 s 23472 49533 23472 49533 4 gnd
port 514 nsew
rlabel metal2 s 22704 48980 22704 48980 4 gnd
port 514 nsew
rlabel metal2 s 24720 48190 24720 48190 4 gnd
port 514 nsew
rlabel metal2 s 23472 48190 23472 48190 4 gnd
port 514 nsew
rlabel metal2 s 23952 50560 23952 50560 4 gnd
port 514 nsew
rlabel metal2 s 23472 48427 23472 48427 4 gnd
port 514 nsew
rlabel metal2 s 24720 50560 24720 50560 4 gnd
port 514 nsew
rlabel metal2 s 23952 47637 23952 47637 4 gnd
port 514 nsew
rlabel metal2 s 23952 50323 23952 50323 4 gnd
port 514 nsew
rlabel metal2 s 23952 49533 23952 49533 4 gnd
port 514 nsew
rlabel metal2 s 23472 47637 23472 47637 4 gnd
port 514 nsew
rlabel metal2 s 22704 50323 22704 50323 4 gnd
port 514 nsew
rlabel metal2 s 20208 48427 20208 48427 4 gnd
port 514 nsew
rlabel metal2 s 20208 49770 20208 49770 4 gnd
port 514 nsew
rlabel metal2 s 20976 48743 20976 48743 4 gnd
port 514 nsew
rlabel metal2 s 21456 49217 21456 49217 4 gnd
port 514 nsew
rlabel metal2 s 21456 49533 21456 49533 4 gnd
port 514 nsew
rlabel metal2 s 21456 47637 21456 47637 4 gnd
port 514 nsew
rlabel metal2 s 21456 50323 21456 50323 4 gnd
port 514 nsew
rlabel metal2 s 22224 50323 22224 50323 4 gnd
port 514 nsew
rlabel metal2 s 20208 48980 20208 48980 4 gnd
port 514 nsew
rlabel metal2 s 20976 47953 20976 47953 4 gnd
port 514 nsew
rlabel metal2 s 21456 50007 21456 50007 4 gnd
port 514 nsew
rlabel metal2 s 21456 48190 21456 48190 4 gnd
port 514 nsew
rlabel metal2 s 20976 49770 20976 49770 4 gnd
port 514 nsew
rlabel metal2 s 22224 49770 22224 49770 4 gnd
port 514 nsew
rlabel metal2 s 20976 48427 20976 48427 4 gnd
port 514 nsew
rlabel metal2 s 20208 50007 20208 50007 4 gnd
port 514 nsew
rlabel metal2 s 22224 47953 22224 47953 4 gnd
port 514 nsew
rlabel metal2 s 21456 49770 21456 49770 4 gnd
port 514 nsew
rlabel metal2 s 20208 50560 20208 50560 4 gnd
port 514 nsew
rlabel metal2 s 21456 50560 21456 50560 4 gnd
port 514 nsew
rlabel metal2 s 20976 48980 20976 48980 4 gnd
port 514 nsew
rlabel metal2 s 22224 47637 22224 47637 4 gnd
port 514 nsew
rlabel metal2 s 21456 47953 21456 47953 4 gnd
port 514 nsew
rlabel metal2 s 22224 48980 22224 48980 4 gnd
port 514 nsew
rlabel metal2 s 21456 48743 21456 48743 4 gnd
port 514 nsew
rlabel metal2 s 22224 48427 22224 48427 4 gnd
port 514 nsew
rlabel metal2 s 21456 48980 21456 48980 4 gnd
port 514 nsew
rlabel metal2 s 20208 47637 20208 47637 4 gnd
port 514 nsew
rlabel metal2 s 20976 47637 20976 47637 4 gnd
port 514 nsew
rlabel metal2 s 22224 49533 22224 49533 4 gnd
port 514 nsew
rlabel metal2 s 20976 50007 20976 50007 4 gnd
port 514 nsew
rlabel metal2 s 20208 50323 20208 50323 4 gnd
port 514 nsew
rlabel metal2 s 20976 48190 20976 48190 4 gnd
port 514 nsew
rlabel metal2 s 20976 49217 20976 49217 4 gnd
port 514 nsew
rlabel metal2 s 22224 48743 22224 48743 4 gnd
port 514 nsew
rlabel metal2 s 22224 49217 22224 49217 4 gnd
port 514 nsew
rlabel metal2 s 20976 50323 20976 50323 4 gnd
port 514 nsew
rlabel metal2 s 20208 49217 20208 49217 4 gnd
port 514 nsew
rlabel metal2 s 20208 48190 20208 48190 4 gnd
port 514 nsew
rlabel metal2 s 20208 48743 20208 48743 4 gnd
port 514 nsew
rlabel metal2 s 20208 47953 20208 47953 4 gnd
port 514 nsew
rlabel metal2 s 21456 48427 21456 48427 4 gnd
port 514 nsew
rlabel metal2 s 20208 49533 20208 49533 4 gnd
port 514 nsew
rlabel metal2 s 22224 48190 22224 48190 4 gnd
port 514 nsew
rlabel metal2 s 20976 50560 20976 50560 4 gnd
port 514 nsew
rlabel metal2 s 22224 50560 22224 50560 4 gnd
port 514 nsew
rlabel metal2 s 22224 50007 22224 50007 4 gnd
port 514 nsew
rlabel metal2 s 20976 49533 20976 49533 4 gnd
port 514 nsew
rlabel metal2 s 21456 47400 21456 47400 4 gnd
port 514 nsew
rlabel metal2 s 22224 46373 22224 46373 4 gnd
port 514 nsew
rlabel metal2 s 20208 44477 20208 44477 4 gnd
port 514 nsew
rlabel metal2 s 22224 46847 22224 46847 4 gnd
port 514 nsew
rlabel metal2 s 20208 46610 20208 46610 4 gnd
port 514 nsew
rlabel metal2 s 20976 47163 20976 47163 4 gnd
port 514 nsew
rlabel metal2 s 21456 46847 21456 46847 4 gnd
port 514 nsew
rlabel metal2 s 20208 44793 20208 44793 4 gnd
port 514 nsew
rlabel metal2 s 20976 46610 20976 46610 4 gnd
port 514 nsew
rlabel metal2 s 21456 44793 21456 44793 4 gnd
port 514 nsew
rlabel metal2 s 22224 46057 22224 46057 4 gnd
port 514 nsew
rlabel metal2 s 20208 47163 20208 47163 4 gnd
port 514 nsew
rlabel metal2 s 21456 47163 21456 47163 4 gnd
port 514 nsew
rlabel metal2 s 21456 46373 21456 46373 4 gnd
port 514 nsew
rlabel metal2 s 22224 45583 22224 45583 4 gnd
port 514 nsew
rlabel metal2 s 20208 45583 20208 45583 4 gnd
port 514 nsew
rlabel metal2 s 20208 45820 20208 45820 4 gnd
port 514 nsew
rlabel metal2 s 21456 45583 21456 45583 4 gnd
port 514 nsew
rlabel metal2 s 21456 46610 21456 46610 4 gnd
port 514 nsew
rlabel metal2 s 20976 44793 20976 44793 4 gnd
port 514 nsew
rlabel metal2 s 20208 46373 20208 46373 4 gnd
port 514 nsew
rlabel metal2 s 22224 46610 22224 46610 4 gnd
port 514 nsew
rlabel metal2 s 20208 46057 20208 46057 4 gnd
port 514 nsew
rlabel metal2 s 20208 47400 20208 47400 4 gnd
port 514 nsew
rlabel metal2 s 20976 44477 20976 44477 4 gnd
port 514 nsew
rlabel metal2 s 21456 45030 21456 45030 4 gnd
port 514 nsew
rlabel metal2 s 20976 46847 20976 46847 4 gnd
port 514 nsew
rlabel metal2 s 20976 45820 20976 45820 4 gnd
port 514 nsew
rlabel metal2 s 20208 45030 20208 45030 4 gnd
port 514 nsew
rlabel metal2 s 20208 46847 20208 46847 4 gnd
port 514 nsew
rlabel metal2 s 21456 45267 21456 45267 4 gnd
port 514 nsew
rlabel metal2 s 22224 45267 22224 45267 4 gnd
port 514 nsew
rlabel metal2 s 20976 45583 20976 45583 4 gnd
port 514 nsew
rlabel metal2 s 22224 45820 22224 45820 4 gnd
port 514 nsew
rlabel metal2 s 22224 45030 22224 45030 4 gnd
port 514 nsew
rlabel metal2 s 20976 47400 20976 47400 4 gnd
port 514 nsew
rlabel metal2 s 22224 44477 22224 44477 4 gnd
port 514 nsew
rlabel metal2 s 22224 44793 22224 44793 4 gnd
port 514 nsew
rlabel metal2 s 20976 45267 20976 45267 4 gnd
port 514 nsew
rlabel metal2 s 20208 45267 20208 45267 4 gnd
port 514 nsew
rlabel metal2 s 21456 46057 21456 46057 4 gnd
port 514 nsew
rlabel metal2 s 21456 45820 21456 45820 4 gnd
port 514 nsew
rlabel metal2 s 22224 47163 22224 47163 4 gnd
port 514 nsew
rlabel metal2 s 21456 44477 21456 44477 4 gnd
port 514 nsew
rlabel metal2 s 20976 45030 20976 45030 4 gnd
port 514 nsew
rlabel metal2 s 20976 46373 20976 46373 4 gnd
port 514 nsew
rlabel metal2 s 20976 46057 20976 46057 4 gnd
port 514 nsew
rlabel metal2 s 22224 47400 22224 47400 4 gnd
port 514 nsew
rlabel metal2 s 24720 45267 24720 45267 4 gnd
port 514 nsew
rlabel metal2 s 23952 46847 23952 46847 4 gnd
port 514 nsew
rlabel metal2 s 23952 47400 23952 47400 4 gnd
port 514 nsew
rlabel metal2 s 24720 46057 24720 46057 4 gnd
port 514 nsew
rlabel metal2 s 24720 44793 24720 44793 4 gnd
port 514 nsew
rlabel metal2 s 24720 45030 24720 45030 4 gnd
port 514 nsew
rlabel metal2 s 22704 45267 22704 45267 4 gnd
port 514 nsew
rlabel metal2 s 23472 45267 23472 45267 4 gnd
port 514 nsew
rlabel metal2 s 23952 45583 23952 45583 4 gnd
port 514 nsew
rlabel metal2 s 23472 45583 23472 45583 4 gnd
port 514 nsew
rlabel metal2 s 24720 45820 24720 45820 4 gnd
port 514 nsew
rlabel metal2 s 22704 45030 22704 45030 4 gnd
port 514 nsew
rlabel metal2 s 23952 47163 23952 47163 4 gnd
port 514 nsew
rlabel metal2 s 23952 45030 23952 45030 4 gnd
port 514 nsew
rlabel metal2 s 23472 47400 23472 47400 4 gnd
port 514 nsew
rlabel metal2 s 22704 46057 22704 46057 4 gnd
port 514 nsew
rlabel metal2 s 23472 47163 23472 47163 4 gnd
port 514 nsew
rlabel metal2 s 23952 46610 23952 46610 4 gnd
port 514 nsew
rlabel metal2 s 23472 46610 23472 46610 4 gnd
port 514 nsew
rlabel metal2 s 22704 47400 22704 47400 4 gnd
port 514 nsew
rlabel metal2 s 23472 44477 23472 44477 4 gnd
port 514 nsew
rlabel metal2 s 22704 44477 22704 44477 4 gnd
port 514 nsew
rlabel metal2 s 24720 46847 24720 46847 4 gnd
port 514 nsew
rlabel metal2 s 22704 45820 22704 45820 4 gnd
port 514 nsew
rlabel metal2 s 24720 47400 24720 47400 4 gnd
port 514 nsew
rlabel metal2 s 23472 45030 23472 45030 4 gnd
port 514 nsew
rlabel metal2 s 22704 46373 22704 46373 4 gnd
port 514 nsew
rlabel metal2 s 24720 44477 24720 44477 4 gnd
port 514 nsew
rlabel metal2 s 22704 46610 22704 46610 4 gnd
port 514 nsew
rlabel metal2 s 24720 47163 24720 47163 4 gnd
port 514 nsew
rlabel metal2 s 23472 46373 23472 46373 4 gnd
port 514 nsew
rlabel metal2 s 22704 44793 22704 44793 4 gnd
port 514 nsew
rlabel metal2 s 23952 46373 23952 46373 4 gnd
port 514 nsew
rlabel metal2 s 23952 44793 23952 44793 4 gnd
port 514 nsew
rlabel metal2 s 23472 44793 23472 44793 4 gnd
port 514 nsew
rlabel metal2 s 24720 45583 24720 45583 4 gnd
port 514 nsew
rlabel metal2 s 23472 46057 23472 46057 4 gnd
port 514 nsew
rlabel metal2 s 23952 46057 23952 46057 4 gnd
port 514 nsew
rlabel metal2 s 22704 45583 22704 45583 4 gnd
port 514 nsew
rlabel metal2 s 22704 46847 22704 46847 4 gnd
port 514 nsew
rlabel metal2 s 23472 46847 23472 46847 4 gnd
port 514 nsew
rlabel metal2 s 22704 47163 22704 47163 4 gnd
port 514 nsew
rlabel metal2 s 23472 45820 23472 45820 4 gnd
port 514 nsew
rlabel metal2 s 23952 44477 23952 44477 4 gnd
port 514 nsew
rlabel metal2 s 24720 46610 24720 46610 4 gnd
port 514 nsew
rlabel metal2 s 23952 45267 23952 45267 4 gnd
port 514 nsew
rlabel metal2 s 23952 45820 23952 45820 4 gnd
port 514 nsew
rlabel metal2 s 24720 46373 24720 46373 4 gnd
port 514 nsew
rlabel metal2 s 22704 42897 22704 42897 4 gnd
port 514 nsew
rlabel metal2 s 23952 44240 23952 44240 4 gnd
port 514 nsew
rlabel metal2 s 23472 41870 23472 41870 4 gnd
port 514 nsew
rlabel metal2 s 22704 42423 22704 42423 4 gnd
port 514 nsew
rlabel metal2 s 24720 43450 24720 43450 4 gnd
port 514 nsew
rlabel metal2 s 23952 42660 23952 42660 4 gnd
port 514 nsew
rlabel metal2 s 23472 42660 23472 42660 4 gnd
port 514 nsew
rlabel metal2 s 22704 43450 22704 43450 4 gnd
port 514 nsew
rlabel metal2 s 23472 43450 23472 43450 4 gnd
port 514 nsew
rlabel metal2 s 22704 44240 22704 44240 4 gnd
port 514 nsew
rlabel metal2 s 24720 43213 24720 43213 4 gnd
port 514 nsew
rlabel metal2 s 23952 42897 23952 42897 4 gnd
port 514 nsew
rlabel metal2 s 23472 42107 23472 42107 4 gnd
port 514 nsew
rlabel metal2 s 23952 42107 23952 42107 4 gnd
port 514 nsew
rlabel metal2 s 24720 44003 24720 44003 4 gnd
port 514 nsew
rlabel metal2 s 23952 41317 23952 41317 4 gnd
port 514 nsew
rlabel metal2 s 24720 42423 24720 42423 4 gnd
port 514 nsew
rlabel metal2 s 23952 43450 23952 43450 4 gnd
port 514 nsew
rlabel metal2 s 22704 43687 22704 43687 4 gnd
port 514 nsew
rlabel metal2 s 23952 42423 23952 42423 4 gnd
port 514 nsew
rlabel metal2 s 23952 44003 23952 44003 4 gnd
port 514 nsew
rlabel metal2 s 22704 41317 22704 41317 4 gnd
port 514 nsew
rlabel metal2 s 23472 44003 23472 44003 4 gnd
port 514 nsew
rlabel metal2 s 23472 42897 23472 42897 4 gnd
port 514 nsew
rlabel metal2 s 22704 41633 22704 41633 4 gnd
port 514 nsew
rlabel metal2 s 24720 42897 24720 42897 4 gnd
port 514 nsew
rlabel metal2 s 24720 41633 24720 41633 4 gnd
port 514 nsew
rlabel metal2 s 24720 43687 24720 43687 4 gnd
port 514 nsew
rlabel metal2 s 24720 41317 24720 41317 4 gnd
port 514 nsew
rlabel metal2 s 22704 42660 22704 42660 4 gnd
port 514 nsew
rlabel metal2 s 22704 44003 22704 44003 4 gnd
port 514 nsew
rlabel metal2 s 23472 41317 23472 41317 4 gnd
port 514 nsew
rlabel metal2 s 23472 44240 23472 44240 4 gnd
port 514 nsew
rlabel metal2 s 22704 43213 22704 43213 4 gnd
port 514 nsew
rlabel metal2 s 22704 41870 22704 41870 4 gnd
port 514 nsew
rlabel metal2 s 24720 44240 24720 44240 4 gnd
port 514 nsew
rlabel metal2 s 24720 42660 24720 42660 4 gnd
port 514 nsew
rlabel metal2 s 22704 42107 22704 42107 4 gnd
port 514 nsew
rlabel metal2 s 24720 42107 24720 42107 4 gnd
port 514 nsew
rlabel metal2 s 23952 41870 23952 41870 4 gnd
port 514 nsew
rlabel metal2 s 23472 42423 23472 42423 4 gnd
port 514 nsew
rlabel metal2 s 23472 41633 23472 41633 4 gnd
port 514 nsew
rlabel metal2 s 23472 43213 23472 43213 4 gnd
port 514 nsew
rlabel metal2 s 23952 43687 23952 43687 4 gnd
port 514 nsew
rlabel metal2 s 23952 41633 23952 41633 4 gnd
port 514 nsew
rlabel metal2 s 24720 41870 24720 41870 4 gnd
port 514 nsew
rlabel metal2 s 23952 43213 23952 43213 4 gnd
port 514 nsew
rlabel metal2 s 23472 43687 23472 43687 4 gnd
port 514 nsew
rlabel metal2 s 22224 42660 22224 42660 4 gnd
port 514 nsew
rlabel metal2 s 20208 42660 20208 42660 4 gnd
port 514 nsew
rlabel metal2 s 22224 41633 22224 41633 4 gnd
port 514 nsew
rlabel metal2 s 20208 42107 20208 42107 4 gnd
port 514 nsew
rlabel metal2 s 20976 44003 20976 44003 4 gnd
port 514 nsew
rlabel metal2 s 22224 42897 22224 42897 4 gnd
port 514 nsew
rlabel metal2 s 21456 42423 21456 42423 4 gnd
port 514 nsew
rlabel metal2 s 20208 42897 20208 42897 4 gnd
port 514 nsew
rlabel metal2 s 21456 43213 21456 43213 4 gnd
port 514 nsew
rlabel metal2 s 22224 43450 22224 43450 4 gnd
port 514 nsew
rlabel metal2 s 20208 44003 20208 44003 4 gnd
port 514 nsew
rlabel metal2 s 22224 44240 22224 44240 4 gnd
port 514 nsew
rlabel metal2 s 21456 42897 21456 42897 4 gnd
port 514 nsew
rlabel metal2 s 20976 43213 20976 43213 4 gnd
port 514 nsew
rlabel metal2 s 20976 43687 20976 43687 4 gnd
port 514 nsew
rlabel metal2 s 21456 44003 21456 44003 4 gnd
port 514 nsew
rlabel metal2 s 22224 43687 22224 43687 4 gnd
port 514 nsew
rlabel metal2 s 20976 41317 20976 41317 4 gnd
port 514 nsew
rlabel metal2 s 22224 41870 22224 41870 4 gnd
port 514 nsew
rlabel metal2 s 20208 43450 20208 43450 4 gnd
port 514 nsew
rlabel metal2 s 20976 42897 20976 42897 4 gnd
port 514 nsew
rlabel metal2 s 21456 41870 21456 41870 4 gnd
port 514 nsew
rlabel metal2 s 20976 42423 20976 42423 4 gnd
port 514 nsew
rlabel metal2 s 22224 42423 22224 42423 4 gnd
port 514 nsew
rlabel metal2 s 20976 41633 20976 41633 4 gnd
port 514 nsew
rlabel metal2 s 22224 43213 22224 43213 4 gnd
port 514 nsew
rlabel metal2 s 20976 43450 20976 43450 4 gnd
port 514 nsew
rlabel metal2 s 21456 41317 21456 41317 4 gnd
port 514 nsew
rlabel metal2 s 20976 42660 20976 42660 4 gnd
port 514 nsew
rlabel metal2 s 22224 42107 22224 42107 4 gnd
port 514 nsew
rlabel metal2 s 20208 43687 20208 43687 4 gnd
port 514 nsew
rlabel metal2 s 20208 44240 20208 44240 4 gnd
port 514 nsew
rlabel metal2 s 20976 44240 20976 44240 4 gnd
port 514 nsew
rlabel metal2 s 20208 41317 20208 41317 4 gnd
port 514 nsew
rlabel metal2 s 21456 42107 21456 42107 4 gnd
port 514 nsew
rlabel metal2 s 21456 43687 21456 43687 4 gnd
port 514 nsew
rlabel metal2 s 22224 44003 22224 44003 4 gnd
port 514 nsew
rlabel metal2 s 21456 41633 21456 41633 4 gnd
port 514 nsew
rlabel metal2 s 21456 43450 21456 43450 4 gnd
port 514 nsew
rlabel metal2 s 21456 44240 21456 44240 4 gnd
port 514 nsew
rlabel metal2 s 20208 41870 20208 41870 4 gnd
port 514 nsew
rlabel metal2 s 22224 41317 22224 41317 4 gnd
port 514 nsew
rlabel metal2 s 21456 42660 21456 42660 4 gnd
port 514 nsew
rlabel metal2 s 20208 43213 20208 43213 4 gnd
port 514 nsew
rlabel metal2 s 20208 41633 20208 41633 4 gnd
port 514 nsew
rlabel metal2 s 20208 42423 20208 42423 4 gnd
port 514 nsew
rlabel metal2 s 20976 41870 20976 41870 4 gnd
port 514 nsew
rlabel metal2 s 20976 42107 20976 42107 4 gnd
port 514 nsew
rlabel metal2 s 20976 39737 20976 39737 4 gnd
port 514 nsew
rlabel metal2 s 22224 39737 22224 39737 4 gnd
port 514 nsew
rlabel metal2 s 20976 40843 20976 40843 4 gnd
port 514 nsew
rlabel metal2 s 20976 39263 20976 39263 4 gnd
port 514 nsew
rlabel metal2 s 20208 39263 20208 39263 4 gnd
port 514 nsew
rlabel metal2 s 22224 38473 22224 38473 4 gnd
port 514 nsew
rlabel metal2 s 20976 40053 20976 40053 4 gnd
port 514 nsew
rlabel metal2 s 22224 38947 22224 38947 4 gnd
port 514 nsew
rlabel metal2 s 22224 40527 22224 40527 4 gnd
port 514 nsew
rlabel metal2 s 21456 39263 21456 39263 4 gnd
port 514 nsew
rlabel metal2 s 21456 40290 21456 40290 4 gnd
port 514 nsew
rlabel metal2 s 20208 38947 20208 38947 4 gnd
port 514 nsew
rlabel metal2 s 20976 38157 20976 38157 4 gnd
port 514 nsew
rlabel metal2 s 21456 40527 21456 40527 4 gnd
port 514 nsew
rlabel metal2 s 22224 41080 22224 41080 4 gnd
port 514 nsew
rlabel metal2 s 21456 38157 21456 38157 4 gnd
port 514 nsew
rlabel metal2 s 20976 39500 20976 39500 4 gnd
port 514 nsew
rlabel metal2 s 20208 39500 20208 39500 4 gnd
port 514 nsew
rlabel metal2 s 22224 38710 22224 38710 4 gnd
port 514 nsew
rlabel metal2 s 20976 40527 20976 40527 4 gnd
port 514 nsew
rlabel metal2 s 21456 40843 21456 40843 4 gnd
port 514 nsew
rlabel metal2 s 20208 40290 20208 40290 4 gnd
port 514 nsew
rlabel metal2 s 20208 40843 20208 40843 4 gnd
port 514 nsew
rlabel metal2 s 22224 40843 22224 40843 4 gnd
port 514 nsew
rlabel metal2 s 20976 38710 20976 38710 4 gnd
port 514 nsew
rlabel metal2 s 20208 39737 20208 39737 4 gnd
port 514 nsew
rlabel metal2 s 20208 41080 20208 41080 4 gnd
port 514 nsew
rlabel metal2 s 20976 38473 20976 38473 4 gnd
port 514 nsew
rlabel metal2 s 22224 39263 22224 39263 4 gnd
port 514 nsew
rlabel metal2 s 20208 40053 20208 40053 4 gnd
port 514 nsew
rlabel metal2 s 21456 40053 21456 40053 4 gnd
port 514 nsew
rlabel metal2 s 21456 38473 21456 38473 4 gnd
port 514 nsew
rlabel metal2 s 21456 38947 21456 38947 4 gnd
port 514 nsew
rlabel metal2 s 21456 41080 21456 41080 4 gnd
port 514 nsew
rlabel metal2 s 20208 38157 20208 38157 4 gnd
port 514 nsew
rlabel metal2 s 22224 40053 22224 40053 4 gnd
port 514 nsew
rlabel metal2 s 22224 39500 22224 39500 4 gnd
port 514 nsew
rlabel metal2 s 21456 38710 21456 38710 4 gnd
port 514 nsew
rlabel metal2 s 20208 40527 20208 40527 4 gnd
port 514 nsew
rlabel metal2 s 22224 38157 22224 38157 4 gnd
port 514 nsew
rlabel metal2 s 20976 38947 20976 38947 4 gnd
port 514 nsew
rlabel metal2 s 20208 38473 20208 38473 4 gnd
port 514 nsew
rlabel metal2 s 20976 40290 20976 40290 4 gnd
port 514 nsew
rlabel metal2 s 20976 41080 20976 41080 4 gnd
port 514 nsew
rlabel metal2 s 21456 39737 21456 39737 4 gnd
port 514 nsew
rlabel metal2 s 20208 38710 20208 38710 4 gnd
port 514 nsew
rlabel metal2 s 21456 39500 21456 39500 4 gnd
port 514 nsew
rlabel metal2 s 22224 40290 22224 40290 4 gnd
port 514 nsew
rlabel metal2 s 23952 38947 23952 38947 4 gnd
port 514 nsew
rlabel metal2 s 24720 40053 24720 40053 4 gnd
port 514 nsew
rlabel metal2 s 23952 40843 23952 40843 4 gnd
port 514 nsew
rlabel metal2 s 24720 40290 24720 40290 4 gnd
port 514 nsew
rlabel metal2 s 23472 41080 23472 41080 4 gnd
port 514 nsew
rlabel metal2 s 22704 38157 22704 38157 4 gnd
port 514 nsew
rlabel metal2 s 24720 39737 24720 39737 4 gnd
port 514 nsew
rlabel metal2 s 23952 38710 23952 38710 4 gnd
port 514 nsew
rlabel metal2 s 24720 38947 24720 38947 4 gnd
port 514 nsew
rlabel metal2 s 23952 39500 23952 39500 4 gnd
port 514 nsew
rlabel metal2 s 22704 39737 22704 39737 4 gnd
port 514 nsew
rlabel metal2 s 23472 38157 23472 38157 4 gnd
port 514 nsew
rlabel metal2 s 24720 39500 24720 39500 4 gnd
port 514 nsew
rlabel metal2 s 23472 38947 23472 38947 4 gnd
port 514 nsew
rlabel metal2 s 22704 38473 22704 38473 4 gnd
port 514 nsew
rlabel metal2 s 22704 39500 22704 39500 4 gnd
port 514 nsew
rlabel metal2 s 24720 41080 24720 41080 4 gnd
port 514 nsew
rlabel metal2 s 23952 41080 23952 41080 4 gnd
port 514 nsew
rlabel metal2 s 22704 39263 22704 39263 4 gnd
port 514 nsew
rlabel metal2 s 24720 39263 24720 39263 4 gnd
port 514 nsew
rlabel metal2 s 23952 38473 23952 38473 4 gnd
port 514 nsew
rlabel metal2 s 23952 40527 23952 40527 4 gnd
port 514 nsew
rlabel metal2 s 23952 40053 23952 40053 4 gnd
port 514 nsew
rlabel metal2 s 23472 39737 23472 39737 4 gnd
port 514 nsew
rlabel metal2 s 22704 40843 22704 40843 4 gnd
port 514 nsew
rlabel metal2 s 24720 38157 24720 38157 4 gnd
port 514 nsew
rlabel metal2 s 23952 39263 23952 39263 4 gnd
port 514 nsew
rlabel metal2 s 22704 40053 22704 40053 4 gnd
port 514 nsew
rlabel metal2 s 24720 40843 24720 40843 4 gnd
port 514 nsew
rlabel metal2 s 24720 38473 24720 38473 4 gnd
port 514 nsew
rlabel metal2 s 22704 38710 22704 38710 4 gnd
port 514 nsew
rlabel metal2 s 23952 38157 23952 38157 4 gnd
port 514 nsew
rlabel metal2 s 23472 40527 23472 40527 4 gnd
port 514 nsew
rlabel metal2 s 23472 40053 23472 40053 4 gnd
port 514 nsew
rlabel metal2 s 23952 39737 23952 39737 4 gnd
port 514 nsew
rlabel metal2 s 23472 40843 23472 40843 4 gnd
port 514 nsew
rlabel metal2 s 22704 40527 22704 40527 4 gnd
port 514 nsew
rlabel metal2 s 23472 40290 23472 40290 4 gnd
port 514 nsew
rlabel metal2 s 23952 40290 23952 40290 4 gnd
port 514 nsew
rlabel metal2 s 23472 39263 23472 39263 4 gnd
port 514 nsew
rlabel metal2 s 22704 40290 22704 40290 4 gnd
port 514 nsew
rlabel metal2 s 23472 39500 23472 39500 4 gnd
port 514 nsew
rlabel metal2 s 23472 38473 23472 38473 4 gnd
port 514 nsew
rlabel metal2 s 23472 38710 23472 38710 4 gnd
port 514 nsew
rlabel metal2 s 24720 40527 24720 40527 4 gnd
port 514 nsew
rlabel metal2 s 22704 41080 22704 41080 4 gnd
port 514 nsew
rlabel metal2 s 22704 38947 22704 38947 4 gnd
port 514 nsew
rlabel metal2 s 24720 38710 24720 38710 4 gnd
port 514 nsew
rlabel metal2 s 28464 43213 28464 43213 4 gnd
port 514 nsew
rlabel metal2 s 27696 41633 27696 41633 4 gnd
port 514 nsew
rlabel metal2 s 27696 41870 27696 41870 4 gnd
port 514 nsew
rlabel metal2 s 27696 43687 27696 43687 4 gnd
port 514 nsew
rlabel metal2 s 28944 43687 28944 43687 4 gnd
port 514 nsew
rlabel metal2 s 28944 41633 28944 41633 4 gnd
port 514 nsew
rlabel metal2 s 27696 42897 27696 42897 4 gnd
port 514 nsew
rlabel metal2 s 29712 42423 29712 42423 4 gnd
port 514 nsew
rlabel metal2 s 27696 42423 27696 42423 4 gnd
port 514 nsew
rlabel metal2 s 28464 43687 28464 43687 4 gnd
port 514 nsew
rlabel metal2 s 29712 43213 29712 43213 4 gnd
port 514 nsew
rlabel metal2 s 28464 44003 28464 44003 4 gnd
port 514 nsew
rlabel metal2 s 29712 42897 29712 42897 4 gnd
port 514 nsew
rlabel metal2 s 27696 44240 27696 44240 4 gnd
port 514 nsew
rlabel metal2 s 28944 42660 28944 42660 4 gnd
port 514 nsew
rlabel metal2 s 27696 44003 27696 44003 4 gnd
port 514 nsew
rlabel metal2 s 28464 41870 28464 41870 4 gnd
port 514 nsew
rlabel metal2 s 27696 41317 27696 41317 4 gnd
port 514 nsew
rlabel metal2 s 28944 42897 28944 42897 4 gnd
port 514 nsew
rlabel metal2 s 28464 42660 28464 42660 4 gnd
port 514 nsew
rlabel metal2 s 28464 44240 28464 44240 4 gnd
port 514 nsew
rlabel metal2 s 28464 42897 28464 42897 4 gnd
port 514 nsew
rlabel metal2 s 28464 42423 28464 42423 4 gnd
port 514 nsew
rlabel metal2 s 29712 41870 29712 41870 4 gnd
port 514 nsew
rlabel metal2 s 28944 42423 28944 42423 4 gnd
port 514 nsew
rlabel metal2 s 29712 41317 29712 41317 4 gnd
port 514 nsew
rlabel metal2 s 28464 43450 28464 43450 4 gnd
port 514 nsew
rlabel metal2 s 28944 42107 28944 42107 4 gnd
port 514 nsew
rlabel metal2 s 29712 44003 29712 44003 4 gnd
port 514 nsew
rlabel metal2 s 28944 44003 28944 44003 4 gnd
port 514 nsew
rlabel metal2 s 28944 41870 28944 41870 4 gnd
port 514 nsew
rlabel metal2 s 28464 42107 28464 42107 4 gnd
port 514 nsew
rlabel metal2 s 29712 42107 29712 42107 4 gnd
port 514 nsew
rlabel metal2 s 29712 43687 29712 43687 4 gnd
port 514 nsew
rlabel metal2 s 28944 43213 28944 43213 4 gnd
port 514 nsew
rlabel metal2 s 29712 42660 29712 42660 4 gnd
port 514 nsew
rlabel metal2 s 28944 41317 28944 41317 4 gnd
port 514 nsew
rlabel metal2 s 27696 43213 27696 43213 4 gnd
port 514 nsew
rlabel metal2 s 29712 41633 29712 41633 4 gnd
port 514 nsew
rlabel metal2 s 27696 42107 27696 42107 4 gnd
port 514 nsew
rlabel metal2 s 28944 43450 28944 43450 4 gnd
port 514 nsew
rlabel metal2 s 28464 41633 28464 41633 4 gnd
port 514 nsew
rlabel metal2 s 27696 42660 27696 42660 4 gnd
port 514 nsew
rlabel metal2 s 29712 44240 29712 44240 4 gnd
port 514 nsew
rlabel metal2 s 27696 43450 27696 43450 4 gnd
port 514 nsew
rlabel metal2 s 28464 41317 28464 41317 4 gnd
port 514 nsew
rlabel metal2 s 29712 43450 29712 43450 4 gnd
port 514 nsew
rlabel metal2 s 28944 44240 28944 44240 4 gnd
port 514 nsew
rlabel metal2 s 25968 41317 25968 41317 4 gnd
port 514 nsew
rlabel metal2 s 27216 43687 27216 43687 4 gnd
port 514 nsew
rlabel metal2 s 25200 41633 25200 41633 4 gnd
port 514 nsew
rlabel metal2 s 25200 42660 25200 42660 4 gnd
port 514 nsew
rlabel metal2 s 25968 42897 25968 42897 4 gnd
port 514 nsew
rlabel metal2 s 27216 44003 27216 44003 4 gnd
port 514 nsew
rlabel metal2 s 25200 42897 25200 42897 4 gnd
port 514 nsew
rlabel metal2 s 26448 42423 26448 42423 4 gnd
port 514 nsew
rlabel metal2 s 26448 42897 26448 42897 4 gnd
port 514 nsew
rlabel metal2 s 25968 42107 25968 42107 4 gnd
port 514 nsew
rlabel metal2 s 26448 42660 26448 42660 4 gnd
port 514 nsew
rlabel metal2 s 25200 41317 25200 41317 4 gnd
port 514 nsew
rlabel metal2 s 26448 41870 26448 41870 4 gnd
port 514 nsew
rlabel metal2 s 25968 43450 25968 43450 4 gnd
port 514 nsew
rlabel metal2 s 26448 44003 26448 44003 4 gnd
port 514 nsew
rlabel metal2 s 25968 41870 25968 41870 4 gnd
port 514 nsew
rlabel metal2 s 26448 41317 26448 41317 4 gnd
port 514 nsew
rlabel metal2 s 25968 42423 25968 42423 4 gnd
port 514 nsew
rlabel metal2 s 27216 44240 27216 44240 4 gnd
port 514 nsew
rlabel metal2 s 25200 43687 25200 43687 4 gnd
port 514 nsew
rlabel metal2 s 25200 44240 25200 44240 4 gnd
port 514 nsew
rlabel metal2 s 26448 43213 26448 43213 4 gnd
port 514 nsew
rlabel metal2 s 25200 43450 25200 43450 4 gnd
port 514 nsew
rlabel metal2 s 27216 41633 27216 41633 4 gnd
port 514 nsew
rlabel metal2 s 27216 41870 27216 41870 4 gnd
port 514 nsew
rlabel metal2 s 25968 43213 25968 43213 4 gnd
port 514 nsew
rlabel metal2 s 27216 42107 27216 42107 4 gnd
port 514 nsew
rlabel metal2 s 25968 41633 25968 41633 4 gnd
port 514 nsew
rlabel metal2 s 27216 42897 27216 42897 4 gnd
port 514 nsew
rlabel metal2 s 27216 41317 27216 41317 4 gnd
port 514 nsew
rlabel metal2 s 25968 42660 25968 42660 4 gnd
port 514 nsew
rlabel metal2 s 26448 44240 26448 44240 4 gnd
port 514 nsew
rlabel metal2 s 25200 42107 25200 42107 4 gnd
port 514 nsew
rlabel metal2 s 25968 44003 25968 44003 4 gnd
port 514 nsew
rlabel metal2 s 25968 43687 25968 43687 4 gnd
port 514 nsew
rlabel metal2 s 25200 42423 25200 42423 4 gnd
port 514 nsew
rlabel metal2 s 25200 44003 25200 44003 4 gnd
port 514 nsew
rlabel metal2 s 26448 41633 26448 41633 4 gnd
port 514 nsew
rlabel metal2 s 25200 43213 25200 43213 4 gnd
port 514 nsew
rlabel metal2 s 25200 41870 25200 41870 4 gnd
port 514 nsew
rlabel metal2 s 27216 42660 27216 42660 4 gnd
port 514 nsew
rlabel metal2 s 25968 44240 25968 44240 4 gnd
port 514 nsew
rlabel metal2 s 27216 42423 27216 42423 4 gnd
port 514 nsew
rlabel metal2 s 26448 43450 26448 43450 4 gnd
port 514 nsew
rlabel metal2 s 27216 43213 27216 43213 4 gnd
port 514 nsew
rlabel metal2 s 26448 42107 26448 42107 4 gnd
port 514 nsew
rlabel metal2 s 27216 43450 27216 43450 4 gnd
port 514 nsew
rlabel metal2 s 26448 43687 26448 43687 4 gnd
port 514 nsew
rlabel metal2 s 26448 40290 26448 40290 4 gnd
port 514 nsew
rlabel metal2 s 27216 38157 27216 38157 4 gnd
port 514 nsew
rlabel metal2 s 25200 39737 25200 39737 4 gnd
port 514 nsew
rlabel metal2 s 25200 38710 25200 38710 4 gnd
port 514 nsew
rlabel metal2 s 26448 39737 26448 39737 4 gnd
port 514 nsew
rlabel metal2 s 25200 38157 25200 38157 4 gnd
port 514 nsew
rlabel metal2 s 26448 40053 26448 40053 4 gnd
port 514 nsew
rlabel metal2 s 26448 39500 26448 39500 4 gnd
port 514 nsew
rlabel metal2 s 26448 40527 26448 40527 4 gnd
port 514 nsew
rlabel metal2 s 25968 40527 25968 40527 4 gnd
port 514 nsew
rlabel metal2 s 25200 41080 25200 41080 4 gnd
port 514 nsew
rlabel metal2 s 26448 39263 26448 39263 4 gnd
port 514 nsew
rlabel metal2 s 27216 40290 27216 40290 4 gnd
port 514 nsew
rlabel metal2 s 27216 38947 27216 38947 4 gnd
port 514 nsew
rlabel metal2 s 25968 38947 25968 38947 4 gnd
port 514 nsew
rlabel metal2 s 25968 40290 25968 40290 4 gnd
port 514 nsew
rlabel metal2 s 27216 40053 27216 40053 4 gnd
port 514 nsew
rlabel metal2 s 25968 38710 25968 38710 4 gnd
port 514 nsew
rlabel metal2 s 26448 38473 26448 38473 4 gnd
port 514 nsew
rlabel metal2 s 27216 40843 27216 40843 4 gnd
port 514 nsew
rlabel metal2 s 27216 39263 27216 39263 4 gnd
port 514 nsew
rlabel metal2 s 25968 38473 25968 38473 4 gnd
port 514 nsew
rlabel metal2 s 25200 38473 25200 38473 4 gnd
port 514 nsew
rlabel metal2 s 26448 41080 26448 41080 4 gnd
port 514 nsew
rlabel metal2 s 25200 38947 25200 38947 4 gnd
port 514 nsew
rlabel metal2 s 25968 41080 25968 41080 4 gnd
port 514 nsew
rlabel metal2 s 26448 38157 26448 38157 4 gnd
port 514 nsew
rlabel metal2 s 27216 41080 27216 41080 4 gnd
port 514 nsew
rlabel metal2 s 25968 38157 25968 38157 4 gnd
port 514 nsew
rlabel metal2 s 26448 40843 26448 40843 4 gnd
port 514 nsew
rlabel metal2 s 25968 39263 25968 39263 4 gnd
port 514 nsew
rlabel metal2 s 25968 39737 25968 39737 4 gnd
port 514 nsew
rlabel metal2 s 27216 38710 27216 38710 4 gnd
port 514 nsew
rlabel metal2 s 25200 40527 25200 40527 4 gnd
port 514 nsew
rlabel metal2 s 25968 40843 25968 40843 4 gnd
port 514 nsew
rlabel metal2 s 26448 38710 26448 38710 4 gnd
port 514 nsew
rlabel metal2 s 25200 39500 25200 39500 4 gnd
port 514 nsew
rlabel metal2 s 27216 39500 27216 39500 4 gnd
port 514 nsew
rlabel metal2 s 26448 38947 26448 38947 4 gnd
port 514 nsew
rlabel metal2 s 27216 38473 27216 38473 4 gnd
port 514 nsew
rlabel metal2 s 25200 40053 25200 40053 4 gnd
port 514 nsew
rlabel metal2 s 25968 40053 25968 40053 4 gnd
port 514 nsew
rlabel metal2 s 27216 39737 27216 39737 4 gnd
port 514 nsew
rlabel metal2 s 25200 40290 25200 40290 4 gnd
port 514 nsew
rlabel metal2 s 25968 39500 25968 39500 4 gnd
port 514 nsew
rlabel metal2 s 25200 40843 25200 40843 4 gnd
port 514 nsew
rlabel metal2 s 25200 39263 25200 39263 4 gnd
port 514 nsew
rlabel metal2 s 27216 40527 27216 40527 4 gnd
port 514 nsew
rlabel metal2 s 28464 41080 28464 41080 4 gnd
port 514 nsew
rlabel metal2 s 27696 39500 27696 39500 4 gnd
port 514 nsew
rlabel metal2 s 28464 40290 28464 40290 4 gnd
port 514 nsew
rlabel metal2 s 27696 38157 27696 38157 4 gnd
port 514 nsew
rlabel metal2 s 29712 40053 29712 40053 4 gnd
port 514 nsew
rlabel metal2 s 28944 38473 28944 38473 4 gnd
port 514 nsew
rlabel metal2 s 27696 39263 27696 39263 4 gnd
port 514 nsew
rlabel metal2 s 29712 40290 29712 40290 4 gnd
port 514 nsew
rlabel metal2 s 28464 40843 28464 40843 4 gnd
port 514 nsew
rlabel metal2 s 27696 40290 27696 40290 4 gnd
port 514 nsew
rlabel metal2 s 29712 40527 29712 40527 4 gnd
port 514 nsew
rlabel metal2 s 28464 38157 28464 38157 4 gnd
port 514 nsew
rlabel metal2 s 28944 38157 28944 38157 4 gnd
port 514 nsew
rlabel metal2 s 27696 38710 27696 38710 4 gnd
port 514 nsew
rlabel metal2 s 28464 38947 28464 38947 4 gnd
port 514 nsew
rlabel metal2 s 28944 39737 28944 39737 4 gnd
port 514 nsew
rlabel metal2 s 28464 40527 28464 40527 4 gnd
port 514 nsew
rlabel metal2 s 29712 38473 29712 38473 4 gnd
port 514 nsew
rlabel metal2 s 28944 41080 28944 41080 4 gnd
port 514 nsew
rlabel metal2 s 29712 39263 29712 39263 4 gnd
port 514 nsew
rlabel metal2 s 27696 39737 27696 39737 4 gnd
port 514 nsew
rlabel metal2 s 27696 40843 27696 40843 4 gnd
port 514 nsew
rlabel metal2 s 27696 40053 27696 40053 4 gnd
port 514 nsew
rlabel metal2 s 28944 39500 28944 39500 4 gnd
port 514 nsew
rlabel metal2 s 27696 41080 27696 41080 4 gnd
port 514 nsew
rlabel metal2 s 29712 41080 29712 41080 4 gnd
port 514 nsew
rlabel metal2 s 28464 39263 28464 39263 4 gnd
port 514 nsew
rlabel metal2 s 28464 39737 28464 39737 4 gnd
port 514 nsew
rlabel metal2 s 29712 38157 29712 38157 4 gnd
port 514 nsew
rlabel metal2 s 28464 40053 28464 40053 4 gnd
port 514 nsew
rlabel metal2 s 28944 38947 28944 38947 4 gnd
port 514 nsew
rlabel metal2 s 28464 38473 28464 38473 4 gnd
port 514 nsew
rlabel metal2 s 28944 40527 28944 40527 4 gnd
port 514 nsew
rlabel metal2 s 28464 39500 28464 39500 4 gnd
port 514 nsew
rlabel metal2 s 28944 40843 28944 40843 4 gnd
port 514 nsew
rlabel metal2 s 27696 40527 27696 40527 4 gnd
port 514 nsew
rlabel metal2 s 29712 38710 29712 38710 4 gnd
port 514 nsew
rlabel metal2 s 28944 40053 28944 40053 4 gnd
port 514 nsew
rlabel metal2 s 28944 38710 28944 38710 4 gnd
port 514 nsew
rlabel metal2 s 28464 38710 28464 38710 4 gnd
port 514 nsew
rlabel metal2 s 29712 40843 29712 40843 4 gnd
port 514 nsew
rlabel metal2 s 29712 39500 29712 39500 4 gnd
port 514 nsew
rlabel metal2 s 28944 39263 28944 39263 4 gnd
port 514 nsew
rlabel metal2 s 29712 38947 29712 38947 4 gnd
port 514 nsew
rlabel metal2 s 27696 38473 27696 38473 4 gnd
port 514 nsew
rlabel metal2 s 28944 40290 28944 40290 4 gnd
port 514 nsew
rlabel metal2 s 29712 39737 29712 39737 4 gnd
port 514 nsew
rlabel metal2 s 27696 38947 27696 38947 4 gnd
port 514 nsew
rlabel metal2 s 28464 36893 28464 36893 4 gnd
port 514 nsew
rlabel metal2 s 27696 36577 27696 36577 4 gnd
port 514 nsew
rlabel metal2 s 28944 35787 28944 35787 4 gnd
port 514 nsew
rlabel metal2 s 27696 37367 27696 37367 4 gnd
port 514 nsew
rlabel metal2 s 28464 36577 28464 36577 4 gnd
port 514 nsew
rlabel metal2 s 29712 36103 29712 36103 4 gnd
port 514 nsew
rlabel metal2 s 28944 36577 28944 36577 4 gnd
port 514 nsew
rlabel metal2 s 28944 35313 28944 35313 4 gnd
port 514 nsew
rlabel metal2 s 28464 36340 28464 36340 4 gnd
port 514 nsew
rlabel metal2 s 29712 37130 29712 37130 4 gnd
port 514 nsew
rlabel metal2 s 27696 34997 27696 34997 4 gnd
port 514 nsew
rlabel metal2 s 28944 34997 28944 34997 4 gnd
port 514 nsew
rlabel metal2 s 29712 37683 29712 37683 4 gnd
port 514 nsew
rlabel metal2 s 28464 35550 28464 35550 4 gnd
port 514 nsew
rlabel metal2 s 27696 36340 27696 36340 4 gnd
port 514 nsew
rlabel metal2 s 29712 36340 29712 36340 4 gnd
port 514 nsew
rlabel metal2 s 28464 37920 28464 37920 4 gnd
port 514 nsew
rlabel metal2 s 28464 35787 28464 35787 4 gnd
port 514 nsew
rlabel metal2 s 29712 35550 29712 35550 4 gnd
port 514 nsew
rlabel metal2 s 28944 36103 28944 36103 4 gnd
port 514 nsew
rlabel metal2 s 28464 36103 28464 36103 4 gnd
port 514 nsew
rlabel metal2 s 28944 37683 28944 37683 4 gnd
port 514 nsew
rlabel metal2 s 27696 37920 27696 37920 4 gnd
port 514 nsew
rlabel metal2 s 29712 35313 29712 35313 4 gnd
port 514 nsew
rlabel metal2 s 27696 35550 27696 35550 4 gnd
port 514 nsew
rlabel metal2 s 28944 36893 28944 36893 4 gnd
port 514 nsew
rlabel metal2 s 29712 37367 29712 37367 4 gnd
port 514 nsew
rlabel metal2 s 27696 36103 27696 36103 4 gnd
port 514 nsew
rlabel metal2 s 28464 37130 28464 37130 4 gnd
port 514 nsew
rlabel metal2 s 28464 34997 28464 34997 4 gnd
port 514 nsew
rlabel metal2 s 28464 37683 28464 37683 4 gnd
port 514 nsew
rlabel metal2 s 28944 36340 28944 36340 4 gnd
port 514 nsew
rlabel metal2 s 28944 37367 28944 37367 4 gnd
port 514 nsew
rlabel metal2 s 29712 34997 29712 34997 4 gnd
port 514 nsew
rlabel metal2 s 28944 35550 28944 35550 4 gnd
port 514 nsew
rlabel metal2 s 28944 37920 28944 37920 4 gnd
port 514 nsew
rlabel metal2 s 27696 35787 27696 35787 4 gnd
port 514 nsew
rlabel metal2 s 27696 36893 27696 36893 4 gnd
port 514 nsew
rlabel metal2 s 28464 35313 28464 35313 4 gnd
port 514 nsew
rlabel metal2 s 29712 36893 29712 36893 4 gnd
port 514 nsew
rlabel metal2 s 27696 37130 27696 37130 4 gnd
port 514 nsew
rlabel metal2 s 27696 35313 27696 35313 4 gnd
port 514 nsew
rlabel metal2 s 28944 37130 28944 37130 4 gnd
port 514 nsew
rlabel metal2 s 28464 37367 28464 37367 4 gnd
port 514 nsew
rlabel metal2 s 27696 37683 27696 37683 4 gnd
port 514 nsew
rlabel metal2 s 29712 35787 29712 35787 4 gnd
port 514 nsew
rlabel metal2 s 29712 37920 29712 37920 4 gnd
port 514 nsew
rlabel metal2 s 29712 36577 29712 36577 4 gnd
port 514 nsew
rlabel metal2 s 27216 36893 27216 36893 4 gnd
port 514 nsew
rlabel metal2 s 26448 35550 26448 35550 4 gnd
port 514 nsew
rlabel metal2 s 25968 35313 25968 35313 4 gnd
port 514 nsew
rlabel metal2 s 27216 36340 27216 36340 4 gnd
port 514 nsew
rlabel metal2 s 26448 37920 26448 37920 4 gnd
port 514 nsew
rlabel metal2 s 26448 35787 26448 35787 4 gnd
port 514 nsew
rlabel metal2 s 26448 34997 26448 34997 4 gnd
port 514 nsew
rlabel metal2 s 25200 34997 25200 34997 4 gnd
port 514 nsew
rlabel metal2 s 27216 37683 27216 37683 4 gnd
port 514 nsew
rlabel metal2 s 27216 35550 27216 35550 4 gnd
port 514 nsew
rlabel metal2 s 27216 37367 27216 37367 4 gnd
port 514 nsew
rlabel metal2 s 25200 36340 25200 36340 4 gnd
port 514 nsew
rlabel metal2 s 27216 36103 27216 36103 4 gnd
port 514 nsew
rlabel metal2 s 27216 37130 27216 37130 4 gnd
port 514 nsew
rlabel metal2 s 26448 36893 26448 36893 4 gnd
port 514 nsew
rlabel metal2 s 25968 36893 25968 36893 4 gnd
port 514 nsew
rlabel metal2 s 25968 37920 25968 37920 4 gnd
port 514 nsew
rlabel metal2 s 26448 36340 26448 36340 4 gnd
port 514 nsew
rlabel metal2 s 26448 37130 26448 37130 4 gnd
port 514 nsew
rlabel metal2 s 25200 37920 25200 37920 4 gnd
port 514 nsew
rlabel metal2 s 25200 37367 25200 37367 4 gnd
port 514 nsew
rlabel metal2 s 25968 35787 25968 35787 4 gnd
port 514 nsew
rlabel metal2 s 25968 36340 25968 36340 4 gnd
port 514 nsew
rlabel metal2 s 25200 37683 25200 37683 4 gnd
port 514 nsew
rlabel metal2 s 25200 37130 25200 37130 4 gnd
port 514 nsew
rlabel metal2 s 25968 37367 25968 37367 4 gnd
port 514 nsew
rlabel metal2 s 25968 34997 25968 34997 4 gnd
port 514 nsew
rlabel metal2 s 25200 36577 25200 36577 4 gnd
port 514 nsew
rlabel metal2 s 26448 36103 26448 36103 4 gnd
port 514 nsew
rlabel metal2 s 25968 36577 25968 36577 4 gnd
port 514 nsew
rlabel metal2 s 26448 37367 26448 37367 4 gnd
port 514 nsew
rlabel metal2 s 26448 36577 26448 36577 4 gnd
port 514 nsew
rlabel metal2 s 27216 35313 27216 35313 4 gnd
port 514 nsew
rlabel metal2 s 27216 34997 27216 34997 4 gnd
port 514 nsew
rlabel metal2 s 26448 35313 26448 35313 4 gnd
port 514 nsew
rlabel metal2 s 25968 37683 25968 37683 4 gnd
port 514 nsew
rlabel metal2 s 25968 36103 25968 36103 4 gnd
port 514 nsew
rlabel metal2 s 25968 37130 25968 37130 4 gnd
port 514 nsew
rlabel metal2 s 25200 36893 25200 36893 4 gnd
port 514 nsew
rlabel metal2 s 27216 37920 27216 37920 4 gnd
port 514 nsew
rlabel metal2 s 27216 36577 27216 36577 4 gnd
port 514 nsew
rlabel metal2 s 25200 35550 25200 35550 4 gnd
port 514 nsew
rlabel metal2 s 25200 36103 25200 36103 4 gnd
port 514 nsew
rlabel metal2 s 27216 35787 27216 35787 4 gnd
port 514 nsew
rlabel metal2 s 26448 37683 26448 37683 4 gnd
port 514 nsew
rlabel metal2 s 25968 35550 25968 35550 4 gnd
port 514 nsew
rlabel metal2 s 25200 35313 25200 35313 4 gnd
port 514 nsew
rlabel metal2 s 25200 35787 25200 35787 4 gnd
port 514 nsew
rlabel metal2 s 25200 34523 25200 34523 4 gnd
port 514 nsew
rlabel metal2 s 27216 32627 27216 32627 4 gnd
port 514 nsew
rlabel metal2 s 26448 34207 26448 34207 4 gnd
port 514 nsew
rlabel metal2 s 27216 33417 27216 33417 4 gnd
port 514 nsew
rlabel metal2 s 25968 34760 25968 34760 4 gnd
port 514 nsew
rlabel metal2 s 26448 31837 26448 31837 4 gnd
port 514 nsew
rlabel metal2 s 25968 31837 25968 31837 4 gnd
port 514 nsew
rlabel metal2 s 26448 32153 26448 32153 4 gnd
port 514 nsew
rlabel metal2 s 26448 34523 26448 34523 4 gnd
port 514 nsew
rlabel metal2 s 26448 33970 26448 33970 4 gnd
port 514 nsew
rlabel metal2 s 25968 33417 25968 33417 4 gnd
port 514 nsew
rlabel metal2 s 27216 31837 27216 31837 4 gnd
port 514 nsew
rlabel metal2 s 25968 33970 25968 33970 4 gnd
port 514 nsew
rlabel metal2 s 26448 33733 26448 33733 4 gnd
port 514 nsew
rlabel metal2 s 25200 32943 25200 32943 4 gnd
port 514 nsew
rlabel metal2 s 25200 33417 25200 33417 4 gnd
port 514 nsew
rlabel metal2 s 25968 32943 25968 32943 4 gnd
port 514 nsew
rlabel metal2 s 26448 32390 26448 32390 4 gnd
port 514 nsew
rlabel metal2 s 25968 33180 25968 33180 4 gnd
port 514 nsew
rlabel metal2 s 25200 32153 25200 32153 4 gnd
port 514 nsew
rlabel metal2 s 27216 32153 27216 32153 4 gnd
port 514 nsew
rlabel metal2 s 25200 33970 25200 33970 4 gnd
port 514 nsew
rlabel metal2 s 27216 34760 27216 34760 4 gnd
port 514 nsew
rlabel metal2 s 25200 34760 25200 34760 4 gnd
port 514 nsew
rlabel metal2 s 27216 34207 27216 34207 4 gnd
port 514 nsew
rlabel metal2 s 27216 33970 27216 33970 4 gnd
port 514 nsew
rlabel metal2 s 25968 32153 25968 32153 4 gnd
port 514 nsew
rlabel metal2 s 25200 31837 25200 31837 4 gnd
port 514 nsew
rlabel metal2 s 26448 33417 26448 33417 4 gnd
port 514 nsew
rlabel metal2 s 25200 34207 25200 34207 4 gnd
port 514 nsew
rlabel metal2 s 25968 34207 25968 34207 4 gnd
port 514 nsew
rlabel metal2 s 25200 32627 25200 32627 4 gnd
port 514 nsew
rlabel metal2 s 26448 32943 26448 32943 4 gnd
port 514 nsew
rlabel metal2 s 25200 33733 25200 33733 4 gnd
port 514 nsew
rlabel metal2 s 25968 32627 25968 32627 4 gnd
port 514 nsew
rlabel metal2 s 25968 32390 25968 32390 4 gnd
port 514 nsew
rlabel metal2 s 25200 32390 25200 32390 4 gnd
port 514 nsew
rlabel metal2 s 26448 34760 26448 34760 4 gnd
port 514 nsew
rlabel metal2 s 25968 33733 25968 33733 4 gnd
port 514 nsew
rlabel metal2 s 27216 32943 27216 32943 4 gnd
port 514 nsew
rlabel metal2 s 27216 33733 27216 33733 4 gnd
port 514 nsew
rlabel metal2 s 27216 34523 27216 34523 4 gnd
port 514 nsew
rlabel metal2 s 26448 32627 26448 32627 4 gnd
port 514 nsew
rlabel metal2 s 27216 32390 27216 32390 4 gnd
port 514 nsew
rlabel metal2 s 25968 34523 25968 34523 4 gnd
port 514 nsew
rlabel metal2 s 26448 33180 26448 33180 4 gnd
port 514 nsew
rlabel metal2 s 25200 33180 25200 33180 4 gnd
port 514 nsew
rlabel metal2 s 27216 33180 27216 33180 4 gnd
port 514 nsew
rlabel metal2 s 28464 32390 28464 32390 4 gnd
port 514 nsew
rlabel metal2 s 28944 34523 28944 34523 4 gnd
port 514 nsew
rlabel metal2 s 28944 32390 28944 32390 4 gnd
port 514 nsew
rlabel metal2 s 28944 31837 28944 31837 4 gnd
port 514 nsew
rlabel metal2 s 28464 33970 28464 33970 4 gnd
port 514 nsew
rlabel metal2 s 29712 33417 29712 33417 4 gnd
port 514 nsew
rlabel metal2 s 27696 33970 27696 33970 4 gnd
port 514 nsew
rlabel metal2 s 27696 33180 27696 33180 4 gnd
port 514 nsew
rlabel metal2 s 29712 32627 29712 32627 4 gnd
port 514 nsew
rlabel metal2 s 27696 32390 27696 32390 4 gnd
port 514 nsew
rlabel metal2 s 28944 32627 28944 32627 4 gnd
port 514 nsew
rlabel metal2 s 29712 32390 29712 32390 4 gnd
port 514 nsew
rlabel metal2 s 27696 33417 27696 33417 4 gnd
port 514 nsew
rlabel metal2 s 29712 33970 29712 33970 4 gnd
port 514 nsew
rlabel metal2 s 28464 32153 28464 32153 4 gnd
port 514 nsew
rlabel metal2 s 28464 32943 28464 32943 4 gnd
port 514 nsew
rlabel metal2 s 27696 33733 27696 33733 4 gnd
port 514 nsew
rlabel metal2 s 28464 34207 28464 34207 4 gnd
port 514 nsew
rlabel metal2 s 29712 31837 29712 31837 4 gnd
port 514 nsew
rlabel metal2 s 28464 33733 28464 33733 4 gnd
port 514 nsew
rlabel metal2 s 29712 33733 29712 33733 4 gnd
port 514 nsew
rlabel metal2 s 28944 32153 28944 32153 4 gnd
port 514 nsew
rlabel metal2 s 28464 34760 28464 34760 4 gnd
port 514 nsew
rlabel metal2 s 28944 33733 28944 33733 4 gnd
port 514 nsew
rlabel metal2 s 28464 31837 28464 31837 4 gnd
port 514 nsew
rlabel metal2 s 28464 34523 28464 34523 4 gnd
port 514 nsew
rlabel metal2 s 27696 32153 27696 32153 4 gnd
port 514 nsew
rlabel metal2 s 29712 32153 29712 32153 4 gnd
port 514 nsew
rlabel metal2 s 29712 32943 29712 32943 4 gnd
port 514 nsew
rlabel metal2 s 27696 32627 27696 32627 4 gnd
port 514 nsew
rlabel metal2 s 28464 32627 28464 32627 4 gnd
port 514 nsew
rlabel metal2 s 29712 34760 29712 34760 4 gnd
port 514 nsew
rlabel metal2 s 28944 33180 28944 33180 4 gnd
port 514 nsew
rlabel metal2 s 27696 34207 27696 34207 4 gnd
port 514 nsew
rlabel metal2 s 29712 34523 29712 34523 4 gnd
port 514 nsew
rlabel metal2 s 28464 33180 28464 33180 4 gnd
port 514 nsew
rlabel metal2 s 27696 34760 27696 34760 4 gnd
port 514 nsew
rlabel metal2 s 28944 34760 28944 34760 4 gnd
port 514 nsew
rlabel metal2 s 29712 34207 29712 34207 4 gnd
port 514 nsew
rlabel metal2 s 28944 32943 28944 32943 4 gnd
port 514 nsew
rlabel metal2 s 27696 32943 27696 32943 4 gnd
port 514 nsew
rlabel metal2 s 29712 33180 29712 33180 4 gnd
port 514 nsew
rlabel metal2 s 27696 31837 27696 31837 4 gnd
port 514 nsew
rlabel metal2 s 28464 33417 28464 33417 4 gnd
port 514 nsew
rlabel metal2 s 28944 33417 28944 33417 4 gnd
port 514 nsew
rlabel metal2 s 28944 33970 28944 33970 4 gnd
port 514 nsew
rlabel metal2 s 28944 34207 28944 34207 4 gnd
port 514 nsew
rlabel metal2 s 27696 34523 27696 34523 4 gnd
port 514 nsew
rlabel metal2 s 23472 35313 23472 35313 4 gnd
port 514 nsew
rlabel metal2 s 24720 35313 24720 35313 4 gnd
port 514 nsew
rlabel metal2 s 23472 37367 23472 37367 4 gnd
port 514 nsew
rlabel metal2 s 22704 35550 22704 35550 4 gnd
port 514 nsew
rlabel metal2 s 23472 36893 23472 36893 4 gnd
port 514 nsew
rlabel metal2 s 23952 36103 23952 36103 4 gnd
port 514 nsew
rlabel metal2 s 22704 37920 22704 37920 4 gnd
port 514 nsew
rlabel metal2 s 24720 36577 24720 36577 4 gnd
port 514 nsew
rlabel metal2 s 23472 35550 23472 35550 4 gnd
port 514 nsew
rlabel metal2 s 24720 36893 24720 36893 4 gnd
port 514 nsew
rlabel metal2 s 23472 37920 23472 37920 4 gnd
port 514 nsew
rlabel metal2 s 24720 37683 24720 37683 4 gnd
port 514 nsew
rlabel metal2 s 22704 36893 22704 36893 4 gnd
port 514 nsew
rlabel metal2 s 23952 36893 23952 36893 4 gnd
port 514 nsew
rlabel metal2 s 24720 36103 24720 36103 4 gnd
port 514 nsew
rlabel metal2 s 22704 36103 22704 36103 4 gnd
port 514 nsew
rlabel metal2 s 22704 37130 22704 37130 4 gnd
port 514 nsew
rlabel metal2 s 24720 37130 24720 37130 4 gnd
port 514 nsew
rlabel metal2 s 23952 35313 23952 35313 4 gnd
port 514 nsew
rlabel metal2 s 23952 37130 23952 37130 4 gnd
port 514 nsew
rlabel metal2 s 23952 34997 23952 34997 4 gnd
port 514 nsew
rlabel metal2 s 24720 37920 24720 37920 4 gnd
port 514 nsew
rlabel metal2 s 23952 35550 23952 35550 4 gnd
port 514 nsew
rlabel metal2 s 23952 35787 23952 35787 4 gnd
port 514 nsew
rlabel metal2 s 24720 34997 24720 34997 4 gnd
port 514 nsew
rlabel metal2 s 24720 35787 24720 35787 4 gnd
port 514 nsew
rlabel metal2 s 23472 36103 23472 36103 4 gnd
port 514 nsew
rlabel metal2 s 23472 37130 23472 37130 4 gnd
port 514 nsew
rlabel metal2 s 23952 37367 23952 37367 4 gnd
port 514 nsew
rlabel metal2 s 23952 36340 23952 36340 4 gnd
port 514 nsew
rlabel metal2 s 23472 36577 23472 36577 4 gnd
port 514 nsew
rlabel metal2 s 22704 35787 22704 35787 4 gnd
port 514 nsew
rlabel metal2 s 22704 36340 22704 36340 4 gnd
port 514 nsew
rlabel metal2 s 22704 34997 22704 34997 4 gnd
port 514 nsew
rlabel metal2 s 24720 36340 24720 36340 4 gnd
port 514 nsew
rlabel metal2 s 23952 37920 23952 37920 4 gnd
port 514 nsew
rlabel metal2 s 24720 37367 24720 37367 4 gnd
port 514 nsew
rlabel metal2 s 22704 35313 22704 35313 4 gnd
port 514 nsew
rlabel metal2 s 23952 36577 23952 36577 4 gnd
port 514 nsew
rlabel metal2 s 22704 36577 22704 36577 4 gnd
port 514 nsew
rlabel metal2 s 23952 37683 23952 37683 4 gnd
port 514 nsew
rlabel metal2 s 22704 37683 22704 37683 4 gnd
port 514 nsew
rlabel metal2 s 23472 36340 23472 36340 4 gnd
port 514 nsew
rlabel metal2 s 23472 34997 23472 34997 4 gnd
port 514 nsew
rlabel metal2 s 23472 37683 23472 37683 4 gnd
port 514 nsew
rlabel metal2 s 24720 35550 24720 35550 4 gnd
port 514 nsew
rlabel metal2 s 22704 37367 22704 37367 4 gnd
port 514 nsew
rlabel metal2 s 23472 35787 23472 35787 4 gnd
port 514 nsew
rlabel metal2 s 22224 37683 22224 37683 4 gnd
port 514 nsew
rlabel metal2 s 20208 36340 20208 36340 4 gnd
port 514 nsew
rlabel metal2 s 20208 36893 20208 36893 4 gnd
port 514 nsew
rlabel metal2 s 21456 35787 21456 35787 4 gnd
port 514 nsew
rlabel metal2 s 20976 37920 20976 37920 4 gnd
port 514 nsew
rlabel metal2 s 20208 37920 20208 37920 4 gnd
port 514 nsew
rlabel metal2 s 21456 37920 21456 37920 4 gnd
port 514 nsew
rlabel metal2 s 22224 36340 22224 36340 4 gnd
port 514 nsew
rlabel metal2 s 20208 36577 20208 36577 4 gnd
port 514 nsew
rlabel metal2 s 20976 36103 20976 36103 4 gnd
port 514 nsew
rlabel metal2 s 20208 37130 20208 37130 4 gnd
port 514 nsew
rlabel metal2 s 22224 35787 22224 35787 4 gnd
port 514 nsew
rlabel metal2 s 20976 35787 20976 35787 4 gnd
port 514 nsew
rlabel metal2 s 20976 36577 20976 36577 4 gnd
port 514 nsew
rlabel metal2 s 20976 36340 20976 36340 4 gnd
port 514 nsew
rlabel metal2 s 21456 37683 21456 37683 4 gnd
port 514 nsew
rlabel metal2 s 20208 35313 20208 35313 4 gnd
port 514 nsew
rlabel metal2 s 20208 34997 20208 34997 4 gnd
port 514 nsew
rlabel metal2 s 20976 36893 20976 36893 4 gnd
port 514 nsew
rlabel metal2 s 20976 34997 20976 34997 4 gnd
port 514 nsew
rlabel metal2 s 22224 37130 22224 37130 4 gnd
port 514 nsew
rlabel metal2 s 21456 37367 21456 37367 4 gnd
port 514 nsew
rlabel metal2 s 20976 37683 20976 37683 4 gnd
port 514 nsew
rlabel metal2 s 20208 35550 20208 35550 4 gnd
port 514 nsew
rlabel metal2 s 21456 36340 21456 36340 4 gnd
port 514 nsew
rlabel metal2 s 22224 36893 22224 36893 4 gnd
port 514 nsew
rlabel metal2 s 20976 35550 20976 35550 4 gnd
port 514 nsew
rlabel metal2 s 20208 36103 20208 36103 4 gnd
port 514 nsew
rlabel metal2 s 22224 35550 22224 35550 4 gnd
port 514 nsew
rlabel metal2 s 22224 35313 22224 35313 4 gnd
port 514 nsew
rlabel metal2 s 20976 35313 20976 35313 4 gnd
port 514 nsew
rlabel metal2 s 21456 36103 21456 36103 4 gnd
port 514 nsew
rlabel metal2 s 21456 37130 21456 37130 4 gnd
port 514 nsew
rlabel metal2 s 22224 36577 22224 36577 4 gnd
port 514 nsew
rlabel metal2 s 20208 37683 20208 37683 4 gnd
port 514 nsew
rlabel metal2 s 22224 37920 22224 37920 4 gnd
port 514 nsew
rlabel metal2 s 20976 37130 20976 37130 4 gnd
port 514 nsew
rlabel metal2 s 21456 35550 21456 35550 4 gnd
port 514 nsew
rlabel metal2 s 22224 37367 22224 37367 4 gnd
port 514 nsew
rlabel metal2 s 21456 34997 21456 34997 4 gnd
port 514 nsew
rlabel metal2 s 20208 35787 20208 35787 4 gnd
port 514 nsew
rlabel metal2 s 21456 36577 21456 36577 4 gnd
port 514 nsew
rlabel metal2 s 22224 36103 22224 36103 4 gnd
port 514 nsew
rlabel metal2 s 21456 36893 21456 36893 4 gnd
port 514 nsew
rlabel metal2 s 21456 35313 21456 35313 4 gnd
port 514 nsew
rlabel metal2 s 20208 37367 20208 37367 4 gnd
port 514 nsew
rlabel metal2 s 22224 34997 22224 34997 4 gnd
port 514 nsew
rlabel metal2 s 20976 37367 20976 37367 4 gnd
port 514 nsew
rlabel metal2 s 20976 34760 20976 34760 4 gnd
port 514 nsew
rlabel metal2 s 21456 33180 21456 33180 4 gnd
port 514 nsew
rlabel metal2 s 20208 33417 20208 33417 4 gnd
port 514 nsew
rlabel metal2 s 20976 34207 20976 34207 4 gnd
port 514 nsew
rlabel metal2 s 21456 33733 21456 33733 4 gnd
port 514 nsew
rlabel metal2 s 20976 33180 20976 33180 4 gnd
port 514 nsew
rlabel metal2 s 20208 34523 20208 34523 4 gnd
port 514 nsew
rlabel metal2 s 21456 32627 21456 32627 4 gnd
port 514 nsew
rlabel metal2 s 20976 33733 20976 33733 4 gnd
port 514 nsew
rlabel metal2 s 20976 32153 20976 32153 4 gnd
port 514 nsew
rlabel metal2 s 20208 31837 20208 31837 4 gnd
port 514 nsew
rlabel metal2 s 20208 33970 20208 33970 4 gnd
port 514 nsew
rlabel metal2 s 22224 34760 22224 34760 4 gnd
port 514 nsew
rlabel metal2 s 21456 32153 21456 32153 4 gnd
port 514 nsew
rlabel metal2 s 20976 34523 20976 34523 4 gnd
port 514 nsew
rlabel metal2 s 20208 32390 20208 32390 4 gnd
port 514 nsew
rlabel metal2 s 20208 33733 20208 33733 4 gnd
port 514 nsew
rlabel metal2 s 21456 31837 21456 31837 4 gnd
port 514 nsew
rlabel metal2 s 22224 31837 22224 31837 4 gnd
port 514 nsew
rlabel metal2 s 20208 34760 20208 34760 4 gnd
port 514 nsew
rlabel metal2 s 21456 32943 21456 32943 4 gnd
port 514 nsew
rlabel metal2 s 22224 33970 22224 33970 4 gnd
port 514 nsew
rlabel metal2 s 21456 33970 21456 33970 4 gnd
port 514 nsew
rlabel metal2 s 22224 32390 22224 32390 4 gnd
port 514 nsew
rlabel metal2 s 22224 33417 22224 33417 4 gnd
port 514 nsew
rlabel metal2 s 20976 32627 20976 32627 4 gnd
port 514 nsew
rlabel metal2 s 20208 34207 20208 34207 4 gnd
port 514 nsew
rlabel metal2 s 22224 34207 22224 34207 4 gnd
port 514 nsew
rlabel metal2 s 22224 34523 22224 34523 4 gnd
port 514 nsew
rlabel metal2 s 20976 33417 20976 33417 4 gnd
port 514 nsew
rlabel metal2 s 20976 32943 20976 32943 4 gnd
port 514 nsew
rlabel metal2 s 21456 33417 21456 33417 4 gnd
port 514 nsew
rlabel metal2 s 20208 32153 20208 32153 4 gnd
port 514 nsew
rlabel metal2 s 21456 34523 21456 34523 4 gnd
port 514 nsew
rlabel metal2 s 20208 32943 20208 32943 4 gnd
port 514 nsew
rlabel metal2 s 21456 34207 21456 34207 4 gnd
port 514 nsew
rlabel metal2 s 20976 32390 20976 32390 4 gnd
port 514 nsew
rlabel metal2 s 21456 34760 21456 34760 4 gnd
port 514 nsew
rlabel metal2 s 20976 31837 20976 31837 4 gnd
port 514 nsew
rlabel metal2 s 20208 33180 20208 33180 4 gnd
port 514 nsew
rlabel metal2 s 22224 33733 22224 33733 4 gnd
port 514 nsew
rlabel metal2 s 22224 33180 22224 33180 4 gnd
port 514 nsew
rlabel metal2 s 22224 32943 22224 32943 4 gnd
port 514 nsew
rlabel metal2 s 20208 32627 20208 32627 4 gnd
port 514 nsew
rlabel metal2 s 22224 32153 22224 32153 4 gnd
port 514 nsew
rlabel metal2 s 21456 32390 21456 32390 4 gnd
port 514 nsew
rlabel metal2 s 20976 33970 20976 33970 4 gnd
port 514 nsew
rlabel metal2 s 22224 32627 22224 32627 4 gnd
port 514 nsew
rlabel metal2 s 22704 33970 22704 33970 4 gnd
port 514 nsew
rlabel metal2 s 24720 32627 24720 32627 4 gnd
port 514 nsew
rlabel metal2 s 24720 34760 24720 34760 4 gnd
port 514 nsew
rlabel metal2 s 22704 33733 22704 33733 4 gnd
port 514 nsew
rlabel metal2 s 23952 34523 23952 34523 4 gnd
port 514 nsew
rlabel metal2 s 22704 33180 22704 33180 4 gnd
port 514 nsew
rlabel metal2 s 23472 33180 23472 33180 4 gnd
port 514 nsew
rlabel metal2 s 23952 34760 23952 34760 4 gnd
port 514 nsew
rlabel metal2 s 22704 32943 22704 32943 4 gnd
port 514 nsew
rlabel metal2 s 23472 33970 23472 33970 4 gnd
port 514 nsew
rlabel metal2 s 23952 32390 23952 32390 4 gnd
port 514 nsew
rlabel metal2 s 22704 32153 22704 32153 4 gnd
port 514 nsew
rlabel metal2 s 24720 34207 24720 34207 4 gnd
port 514 nsew
rlabel metal2 s 22704 34207 22704 34207 4 gnd
port 514 nsew
rlabel metal2 s 24720 33417 24720 33417 4 gnd
port 514 nsew
rlabel metal2 s 23472 34760 23472 34760 4 gnd
port 514 nsew
rlabel metal2 s 23952 32153 23952 32153 4 gnd
port 514 nsew
rlabel metal2 s 24720 33970 24720 33970 4 gnd
port 514 nsew
rlabel metal2 s 22704 34760 22704 34760 4 gnd
port 514 nsew
rlabel metal2 s 24720 32943 24720 32943 4 gnd
port 514 nsew
rlabel metal2 s 22704 31837 22704 31837 4 gnd
port 514 nsew
rlabel metal2 s 22704 32627 22704 32627 4 gnd
port 514 nsew
rlabel metal2 s 23952 33417 23952 33417 4 gnd
port 514 nsew
rlabel metal2 s 24720 31837 24720 31837 4 gnd
port 514 nsew
rlabel metal2 s 23952 32943 23952 32943 4 gnd
port 514 nsew
rlabel metal2 s 23952 31837 23952 31837 4 gnd
port 514 nsew
rlabel metal2 s 23952 33970 23952 33970 4 gnd
port 514 nsew
rlabel metal2 s 23472 31837 23472 31837 4 gnd
port 514 nsew
rlabel metal2 s 23952 33180 23952 33180 4 gnd
port 514 nsew
rlabel metal2 s 23472 33733 23472 33733 4 gnd
port 514 nsew
rlabel metal2 s 23472 34207 23472 34207 4 gnd
port 514 nsew
rlabel metal2 s 23472 32153 23472 32153 4 gnd
port 514 nsew
rlabel metal2 s 23472 32943 23472 32943 4 gnd
port 514 nsew
rlabel metal2 s 24720 34523 24720 34523 4 gnd
port 514 nsew
rlabel metal2 s 23472 33417 23472 33417 4 gnd
port 514 nsew
rlabel metal2 s 24720 33733 24720 33733 4 gnd
port 514 nsew
rlabel metal2 s 23472 34523 23472 34523 4 gnd
port 514 nsew
rlabel metal2 s 23472 32390 23472 32390 4 gnd
port 514 nsew
rlabel metal2 s 22704 32390 22704 32390 4 gnd
port 514 nsew
rlabel metal2 s 23952 32627 23952 32627 4 gnd
port 514 nsew
rlabel metal2 s 23952 33733 23952 33733 4 gnd
port 514 nsew
rlabel metal2 s 24720 33180 24720 33180 4 gnd
port 514 nsew
rlabel metal2 s 24720 32390 24720 32390 4 gnd
port 514 nsew
rlabel metal2 s 22704 34523 22704 34523 4 gnd
port 514 nsew
rlabel metal2 s 24720 32153 24720 32153 4 gnd
port 514 nsew
rlabel metal2 s 23952 34207 23952 34207 4 gnd
port 514 nsew
rlabel metal2 s 22704 33417 22704 33417 4 gnd
port 514 nsew
rlabel metal2 s 23472 32627 23472 32627 4 gnd
port 514 nsew
rlabel metal2 s 23472 31363 23472 31363 4 gnd
port 514 nsew
rlabel metal2 s 23952 28677 23952 28677 4 gnd
port 514 nsew
rlabel metal2 s 23952 30257 23952 30257 4 gnd
port 514 nsew
rlabel metal2 s 23952 28993 23952 28993 4 gnd
port 514 nsew
rlabel metal2 s 24720 29783 24720 29783 4 gnd
port 514 nsew
rlabel metal2 s 23952 31047 23952 31047 4 gnd
port 514 nsew
rlabel metal2 s 22704 29783 22704 29783 4 gnd
port 514 nsew
rlabel metal2 s 24720 30257 24720 30257 4 gnd
port 514 nsew
rlabel metal2 s 22704 31047 22704 31047 4 gnd
port 514 nsew
rlabel metal2 s 22704 29230 22704 29230 4 gnd
port 514 nsew
rlabel metal2 s 23952 29783 23952 29783 4 gnd
port 514 nsew
rlabel metal2 s 24720 29467 24720 29467 4 gnd
port 514 nsew
rlabel metal2 s 23472 29783 23472 29783 4 gnd
port 514 nsew
rlabel metal2 s 23472 28677 23472 28677 4 gnd
port 514 nsew
rlabel metal2 s 22704 28993 22704 28993 4 gnd
port 514 nsew
rlabel metal2 s 24720 31600 24720 31600 4 gnd
port 514 nsew
rlabel metal2 s 24720 29230 24720 29230 4 gnd
port 514 nsew
rlabel metal2 s 23952 31363 23952 31363 4 gnd
port 514 nsew
rlabel metal2 s 24720 31363 24720 31363 4 gnd
port 514 nsew
rlabel metal2 s 23952 31600 23952 31600 4 gnd
port 514 nsew
rlabel metal2 s 23472 29467 23472 29467 4 gnd
port 514 nsew
rlabel metal2 s 23472 30020 23472 30020 4 gnd
port 514 nsew
rlabel metal2 s 22704 30257 22704 30257 4 gnd
port 514 nsew
rlabel metal2 s 23472 30257 23472 30257 4 gnd
port 514 nsew
rlabel metal2 s 24720 30810 24720 30810 4 gnd
port 514 nsew
rlabel metal2 s 23952 30810 23952 30810 4 gnd
port 514 nsew
rlabel metal2 s 22704 30573 22704 30573 4 gnd
port 514 nsew
rlabel metal2 s 22704 30810 22704 30810 4 gnd
port 514 nsew
rlabel metal2 s 23952 30020 23952 30020 4 gnd
port 514 nsew
rlabel metal2 s 24720 30573 24720 30573 4 gnd
port 514 nsew
rlabel metal2 s 24720 28677 24720 28677 4 gnd
port 514 nsew
rlabel metal2 s 23472 30573 23472 30573 4 gnd
port 514 nsew
rlabel metal2 s 23472 31047 23472 31047 4 gnd
port 514 nsew
rlabel metal2 s 23952 29467 23952 29467 4 gnd
port 514 nsew
rlabel metal2 s 23952 29230 23952 29230 4 gnd
port 514 nsew
rlabel metal2 s 23472 29230 23472 29230 4 gnd
port 514 nsew
rlabel metal2 s 22704 30020 22704 30020 4 gnd
port 514 nsew
rlabel metal2 s 23472 31600 23472 31600 4 gnd
port 514 nsew
rlabel metal2 s 22704 28677 22704 28677 4 gnd
port 514 nsew
rlabel metal2 s 22704 31363 22704 31363 4 gnd
port 514 nsew
rlabel metal2 s 24720 30020 24720 30020 4 gnd
port 514 nsew
rlabel metal2 s 23952 30573 23952 30573 4 gnd
port 514 nsew
rlabel metal2 s 24720 31047 24720 31047 4 gnd
port 514 nsew
rlabel metal2 s 24720 28993 24720 28993 4 gnd
port 514 nsew
rlabel metal2 s 22704 31600 22704 31600 4 gnd
port 514 nsew
rlabel metal2 s 23472 28993 23472 28993 4 gnd
port 514 nsew
rlabel metal2 s 22704 29467 22704 29467 4 gnd
port 514 nsew
rlabel metal2 s 23472 30810 23472 30810 4 gnd
port 514 nsew
rlabel metal2 s 20976 29467 20976 29467 4 gnd
port 514 nsew
rlabel metal2 s 22224 29467 22224 29467 4 gnd
port 514 nsew
rlabel metal2 s 20208 30257 20208 30257 4 gnd
port 514 nsew
rlabel metal2 s 22224 28677 22224 28677 4 gnd
port 514 nsew
rlabel metal2 s 20976 28677 20976 28677 4 gnd
port 514 nsew
rlabel metal2 s 20208 28993 20208 28993 4 gnd
port 514 nsew
rlabel metal2 s 20976 30810 20976 30810 4 gnd
port 514 nsew
rlabel metal2 s 21456 28993 21456 28993 4 gnd
port 514 nsew
rlabel metal2 s 20208 31047 20208 31047 4 gnd
port 514 nsew
rlabel metal2 s 21456 30573 21456 30573 4 gnd
port 514 nsew
rlabel metal2 s 21456 28677 21456 28677 4 gnd
port 514 nsew
rlabel metal2 s 20976 30257 20976 30257 4 gnd
port 514 nsew
rlabel metal2 s 22224 31600 22224 31600 4 gnd
port 514 nsew
rlabel metal2 s 22224 30257 22224 30257 4 gnd
port 514 nsew
rlabel metal2 s 20208 29783 20208 29783 4 gnd
port 514 nsew
rlabel metal2 s 20208 30020 20208 30020 4 gnd
port 514 nsew
rlabel metal2 s 20208 31363 20208 31363 4 gnd
port 514 nsew
rlabel metal2 s 21456 30020 21456 30020 4 gnd
port 514 nsew
rlabel metal2 s 20208 28677 20208 28677 4 gnd
port 514 nsew
rlabel metal2 s 22224 31047 22224 31047 4 gnd
port 514 nsew
rlabel metal2 s 21456 31047 21456 31047 4 gnd
port 514 nsew
rlabel metal2 s 20976 31363 20976 31363 4 gnd
port 514 nsew
rlabel metal2 s 20208 30573 20208 30573 4 gnd
port 514 nsew
rlabel metal2 s 22224 28993 22224 28993 4 gnd
port 514 nsew
rlabel metal2 s 21456 29783 21456 29783 4 gnd
port 514 nsew
rlabel metal2 s 20976 31600 20976 31600 4 gnd
port 514 nsew
rlabel metal2 s 20208 29230 20208 29230 4 gnd
port 514 nsew
rlabel metal2 s 20976 28993 20976 28993 4 gnd
port 514 nsew
rlabel metal2 s 21456 31363 21456 31363 4 gnd
port 514 nsew
rlabel metal2 s 21456 31600 21456 31600 4 gnd
port 514 nsew
rlabel metal2 s 22224 29230 22224 29230 4 gnd
port 514 nsew
rlabel metal2 s 22224 30810 22224 30810 4 gnd
port 514 nsew
rlabel metal2 s 20976 31047 20976 31047 4 gnd
port 514 nsew
rlabel metal2 s 20976 29783 20976 29783 4 gnd
port 514 nsew
rlabel metal2 s 22224 29783 22224 29783 4 gnd
port 514 nsew
rlabel metal2 s 21456 29467 21456 29467 4 gnd
port 514 nsew
rlabel metal2 s 22224 30573 22224 30573 4 gnd
port 514 nsew
rlabel metal2 s 20208 29467 20208 29467 4 gnd
port 514 nsew
rlabel metal2 s 21456 30257 21456 30257 4 gnd
port 514 nsew
rlabel metal2 s 20976 30573 20976 30573 4 gnd
port 514 nsew
rlabel metal2 s 20208 31600 20208 31600 4 gnd
port 514 nsew
rlabel metal2 s 20976 29230 20976 29230 4 gnd
port 514 nsew
rlabel metal2 s 20208 30810 20208 30810 4 gnd
port 514 nsew
rlabel metal2 s 22224 30020 22224 30020 4 gnd
port 514 nsew
rlabel metal2 s 21456 29230 21456 29230 4 gnd
port 514 nsew
rlabel metal2 s 21456 30810 21456 30810 4 gnd
port 514 nsew
rlabel metal2 s 22224 31363 22224 31363 4 gnd
port 514 nsew
rlabel metal2 s 20976 30020 20976 30020 4 gnd
port 514 nsew
rlabel metal2 s 21456 27413 21456 27413 4 gnd
port 514 nsew
rlabel metal2 s 21456 26623 21456 26623 4 gnd
port 514 nsew
rlabel metal2 s 21456 27097 21456 27097 4 gnd
port 514 nsew
rlabel metal2 s 22224 28203 22224 28203 4 gnd
port 514 nsew
rlabel metal2 s 20976 25833 20976 25833 4 gnd
port 514 nsew
rlabel metal2 s 20976 26860 20976 26860 4 gnd
port 514 nsew
rlabel metal2 s 22224 27097 22224 27097 4 gnd
port 514 nsew
rlabel metal2 s 21456 25517 21456 25517 4 gnd
port 514 nsew
rlabel metal2 s 22224 25833 22224 25833 4 gnd
port 514 nsew
rlabel metal2 s 20976 26623 20976 26623 4 gnd
port 514 nsew
rlabel metal2 s 20208 28440 20208 28440 4 gnd
port 514 nsew
rlabel metal2 s 22224 25517 22224 25517 4 gnd
port 514 nsew
rlabel metal2 s 20208 26623 20208 26623 4 gnd
port 514 nsew
rlabel metal2 s 20208 25517 20208 25517 4 gnd
port 514 nsew
rlabel metal2 s 20208 27650 20208 27650 4 gnd
port 514 nsew
rlabel metal2 s 20208 27413 20208 27413 4 gnd
port 514 nsew
rlabel metal2 s 20976 28203 20976 28203 4 gnd
port 514 nsew
rlabel metal2 s 22224 26307 22224 26307 4 gnd
port 514 nsew
rlabel metal2 s 20208 26070 20208 26070 4 gnd
port 514 nsew
rlabel metal2 s 20976 26307 20976 26307 4 gnd
port 514 nsew
rlabel metal2 s 22224 28440 22224 28440 4 gnd
port 514 nsew
rlabel metal2 s 20208 27097 20208 27097 4 gnd
port 514 nsew
rlabel metal2 s 21456 27650 21456 27650 4 gnd
port 514 nsew
rlabel metal2 s 20976 25517 20976 25517 4 gnd
port 514 nsew
rlabel metal2 s 20976 27650 20976 27650 4 gnd
port 514 nsew
rlabel metal2 s 21456 26860 21456 26860 4 gnd
port 514 nsew
rlabel metal2 s 22224 26623 22224 26623 4 gnd
port 514 nsew
rlabel metal2 s 22224 26070 22224 26070 4 gnd
port 514 nsew
rlabel metal2 s 20976 27887 20976 27887 4 gnd
port 514 nsew
rlabel metal2 s 20208 25833 20208 25833 4 gnd
port 514 nsew
rlabel metal2 s 20208 26860 20208 26860 4 gnd
port 514 nsew
rlabel metal2 s 20976 27097 20976 27097 4 gnd
port 514 nsew
rlabel metal2 s 21456 25833 21456 25833 4 gnd
port 514 nsew
rlabel metal2 s 20976 27413 20976 27413 4 gnd
port 514 nsew
rlabel metal2 s 21456 28203 21456 28203 4 gnd
port 514 nsew
rlabel metal2 s 21456 28440 21456 28440 4 gnd
port 514 nsew
rlabel metal2 s 22224 27887 22224 27887 4 gnd
port 514 nsew
rlabel metal2 s 21456 27887 21456 27887 4 gnd
port 514 nsew
rlabel metal2 s 20976 28440 20976 28440 4 gnd
port 514 nsew
rlabel metal2 s 21456 26307 21456 26307 4 gnd
port 514 nsew
rlabel metal2 s 22224 26860 22224 26860 4 gnd
port 514 nsew
rlabel metal2 s 22224 27413 22224 27413 4 gnd
port 514 nsew
rlabel metal2 s 20208 26307 20208 26307 4 gnd
port 514 nsew
rlabel metal2 s 20208 27887 20208 27887 4 gnd
port 514 nsew
rlabel metal2 s 21456 26070 21456 26070 4 gnd
port 514 nsew
rlabel metal2 s 20208 28203 20208 28203 4 gnd
port 514 nsew
rlabel metal2 s 22224 27650 22224 27650 4 gnd
port 514 nsew
rlabel metal2 s 20976 26070 20976 26070 4 gnd
port 514 nsew
rlabel metal2 s 23472 26070 23472 26070 4 gnd
port 514 nsew
rlabel metal2 s 24720 26307 24720 26307 4 gnd
port 514 nsew
rlabel metal2 s 22704 28203 22704 28203 4 gnd
port 514 nsew
rlabel metal2 s 22704 27887 22704 27887 4 gnd
port 514 nsew
rlabel metal2 s 23952 26623 23952 26623 4 gnd
port 514 nsew
rlabel metal2 s 23472 27413 23472 27413 4 gnd
port 514 nsew
rlabel metal2 s 23952 25833 23952 25833 4 gnd
port 514 nsew
rlabel metal2 s 23952 27097 23952 27097 4 gnd
port 514 nsew
rlabel metal2 s 24720 26623 24720 26623 4 gnd
port 514 nsew
rlabel metal2 s 23472 27097 23472 27097 4 gnd
port 514 nsew
rlabel metal2 s 23472 26623 23472 26623 4 gnd
port 514 nsew
rlabel metal2 s 24720 25517 24720 25517 4 gnd
port 514 nsew
rlabel metal2 s 23472 26307 23472 26307 4 gnd
port 514 nsew
rlabel metal2 s 22704 26307 22704 26307 4 gnd
port 514 nsew
rlabel metal2 s 24720 26860 24720 26860 4 gnd
port 514 nsew
rlabel metal2 s 23952 28440 23952 28440 4 gnd
port 514 nsew
rlabel metal2 s 22704 27650 22704 27650 4 gnd
port 514 nsew
rlabel metal2 s 23952 26307 23952 26307 4 gnd
port 514 nsew
rlabel metal2 s 22704 26623 22704 26623 4 gnd
port 514 nsew
rlabel metal2 s 23472 26860 23472 26860 4 gnd
port 514 nsew
rlabel metal2 s 24720 28440 24720 28440 4 gnd
port 514 nsew
rlabel metal2 s 23952 26070 23952 26070 4 gnd
port 514 nsew
rlabel metal2 s 24720 27650 24720 27650 4 gnd
port 514 nsew
rlabel metal2 s 24720 28203 24720 28203 4 gnd
port 514 nsew
rlabel metal2 s 23472 25517 23472 25517 4 gnd
port 514 nsew
rlabel metal2 s 24720 25833 24720 25833 4 gnd
port 514 nsew
rlabel metal2 s 23472 27650 23472 27650 4 gnd
port 514 nsew
rlabel metal2 s 24720 27887 24720 27887 4 gnd
port 514 nsew
rlabel metal2 s 23472 28440 23472 28440 4 gnd
port 514 nsew
rlabel metal2 s 22704 26860 22704 26860 4 gnd
port 514 nsew
rlabel metal2 s 23952 26860 23952 26860 4 gnd
port 514 nsew
rlabel metal2 s 22704 25833 22704 25833 4 gnd
port 514 nsew
rlabel metal2 s 23952 25517 23952 25517 4 gnd
port 514 nsew
rlabel metal2 s 24720 27413 24720 27413 4 gnd
port 514 nsew
rlabel metal2 s 23472 28203 23472 28203 4 gnd
port 514 nsew
rlabel metal2 s 22704 25517 22704 25517 4 gnd
port 514 nsew
rlabel metal2 s 23952 27650 23952 27650 4 gnd
port 514 nsew
rlabel metal2 s 24720 26070 24720 26070 4 gnd
port 514 nsew
rlabel metal2 s 22704 28440 22704 28440 4 gnd
port 514 nsew
rlabel metal2 s 22704 26070 22704 26070 4 gnd
port 514 nsew
rlabel metal2 s 23952 27887 23952 27887 4 gnd
port 514 nsew
rlabel metal2 s 23952 27413 23952 27413 4 gnd
port 514 nsew
rlabel metal2 s 22704 27097 22704 27097 4 gnd
port 514 nsew
rlabel metal2 s 23472 27887 23472 27887 4 gnd
port 514 nsew
rlabel metal2 s 24720 27097 24720 27097 4 gnd
port 514 nsew
rlabel metal2 s 22704 27413 22704 27413 4 gnd
port 514 nsew
rlabel metal2 s 23952 28203 23952 28203 4 gnd
port 514 nsew
rlabel metal2 s 23472 25833 23472 25833 4 gnd
port 514 nsew
rlabel metal2 s 27696 29783 27696 29783 4 gnd
port 514 nsew
rlabel metal2 s 28464 30020 28464 30020 4 gnd
port 514 nsew
rlabel metal2 s 28464 28993 28464 28993 4 gnd
port 514 nsew
rlabel metal2 s 28464 31600 28464 31600 4 gnd
port 514 nsew
rlabel metal2 s 28944 31047 28944 31047 4 gnd
port 514 nsew
rlabel metal2 s 28464 31047 28464 31047 4 gnd
port 514 nsew
rlabel metal2 s 28464 29467 28464 29467 4 gnd
port 514 nsew
rlabel metal2 s 27696 28993 27696 28993 4 gnd
port 514 nsew
rlabel metal2 s 28944 31363 28944 31363 4 gnd
port 514 nsew
rlabel metal2 s 27696 29230 27696 29230 4 gnd
port 514 nsew
rlabel metal2 s 28464 29783 28464 29783 4 gnd
port 514 nsew
rlabel metal2 s 27696 31363 27696 31363 4 gnd
port 514 nsew
rlabel metal2 s 28944 29230 28944 29230 4 gnd
port 514 nsew
rlabel metal2 s 28464 30573 28464 30573 4 gnd
port 514 nsew
rlabel metal2 s 28944 30020 28944 30020 4 gnd
port 514 nsew
rlabel metal2 s 28464 31363 28464 31363 4 gnd
port 514 nsew
rlabel metal2 s 27696 29467 27696 29467 4 gnd
port 514 nsew
rlabel metal2 s 29712 31600 29712 31600 4 gnd
port 514 nsew
rlabel metal2 s 28464 29230 28464 29230 4 gnd
port 514 nsew
rlabel metal2 s 27696 30810 27696 30810 4 gnd
port 514 nsew
rlabel metal2 s 29712 31047 29712 31047 4 gnd
port 514 nsew
rlabel metal2 s 29712 30810 29712 30810 4 gnd
port 514 nsew
rlabel metal2 s 29712 30257 29712 30257 4 gnd
port 514 nsew
rlabel metal2 s 29712 30573 29712 30573 4 gnd
port 514 nsew
rlabel metal2 s 27696 30573 27696 30573 4 gnd
port 514 nsew
rlabel metal2 s 29712 30020 29712 30020 4 gnd
port 514 nsew
rlabel metal2 s 27696 30020 27696 30020 4 gnd
port 514 nsew
rlabel metal2 s 28944 30257 28944 30257 4 gnd
port 514 nsew
rlabel metal2 s 28944 28993 28944 28993 4 gnd
port 514 nsew
rlabel metal2 s 28944 29467 28944 29467 4 gnd
port 514 nsew
rlabel metal2 s 27696 28677 27696 28677 4 gnd
port 514 nsew
rlabel metal2 s 27696 30257 27696 30257 4 gnd
port 514 nsew
rlabel metal2 s 28944 30573 28944 30573 4 gnd
port 514 nsew
rlabel metal2 s 27696 31600 27696 31600 4 gnd
port 514 nsew
rlabel metal2 s 28944 30810 28944 30810 4 gnd
port 514 nsew
rlabel metal2 s 27696 31047 27696 31047 4 gnd
port 514 nsew
rlabel metal2 s 29712 28677 29712 28677 4 gnd
port 514 nsew
rlabel metal2 s 28464 30810 28464 30810 4 gnd
port 514 nsew
rlabel metal2 s 29712 29230 29712 29230 4 gnd
port 514 nsew
rlabel metal2 s 28944 28677 28944 28677 4 gnd
port 514 nsew
rlabel metal2 s 29712 28993 29712 28993 4 gnd
port 514 nsew
rlabel metal2 s 29712 29467 29712 29467 4 gnd
port 514 nsew
rlabel metal2 s 28944 29783 28944 29783 4 gnd
port 514 nsew
rlabel metal2 s 29712 29783 29712 29783 4 gnd
port 514 nsew
rlabel metal2 s 29712 31363 29712 31363 4 gnd
port 514 nsew
rlabel metal2 s 28944 31600 28944 31600 4 gnd
port 514 nsew
rlabel metal2 s 28464 28677 28464 28677 4 gnd
port 514 nsew
rlabel metal2 s 28464 30257 28464 30257 4 gnd
port 514 nsew
rlabel metal2 s 25200 28677 25200 28677 4 gnd
port 514 nsew
rlabel metal2 s 25968 29230 25968 29230 4 gnd
port 514 nsew
rlabel metal2 s 27216 29783 27216 29783 4 gnd
port 514 nsew
rlabel metal2 s 27216 31363 27216 31363 4 gnd
port 514 nsew
rlabel metal2 s 26448 28993 26448 28993 4 gnd
port 514 nsew
rlabel metal2 s 25200 30020 25200 30020 4 gnd
port 514 nsew
rlabel metal2 s 27216 29467 27216 29467 4 gnd
port 514 nsew
rlabel metal2 s 26448 31047 26448 31047 4 gnd
port 514 nsew
rlabel metal2 s 25968 29467 25968 29467 4 gnd
port 514 nsew
rlabel metal2 s 26448 30020 26448 30020 4 gnd
port 514 nsew
rlabel metal2 s 26448 31363 26448 31363 4 gnd
port 514 nsew
rlabel metal2 s 27216 29230 27216 29230 4 gnd
port 514 nsew
rlabel metal2 s 26448 29467 26448 29467 4 gnd
port 514 nsew
rlabel metal2 s 26448 29783 26448 29783 4 gnd
port 514 nsew
rlabel metal2 s 26448 29230 26448 29230 4 gnd
port 514 nsew
rlabel metal2 s 25200 31600 25200 31600 4 gnd
port 514 nsew
rlabel metal2 s 25968 31600 25968 31600 4 gnd
port 514 nsew
rlabel metal2 s 25200 28993 25200 28993 4 gnd
port 514 nsew
rlabel metal2 s 25200 29783 25200 29783 4 gnd
port 514 nsew
rlabel metal2 s 27216 30810 27216 30810 4 gnd
port 514 nsew
rlabel metal2 s 27216 28677 27216 28677 4 gnd
port 514 nsew
rlabel metal2 s 27216 28993 27216 28993 4 gnd
port 514 nsew
rlabel metal2 s 25200 31363 25200 31363 4 gnd
port 514 nsew
rlabel metal2 s 25968 28993 25968 28993 4 gnd
port 514 nsew
rlabel metal2 s 26448 28677 26448 28677 4 gnd
port 514 nsew
rlabel metal2 s 25968 31363 25968 31363 4 gnd
port 514 nsew
rlabel metal2 s 25968 30810 25968 30810 4 gnd
port 514 nsew
rlabel metal2 s 26448 31600 26448 31600 4 gnd
port 514 nsew
rlabel metal2 s 25200 29230 25200 29230 4 gnd
port 514 nsew
rlabel metal2 s 25968 31047 25968 31047 4 gnd
port 514 nsew
rlabel metal2 s 26448 30810 26448 30810 4 gnd
port 514 nsew
rlabel metal2 s 25200 30573 25200 30573 4 gnd
port 514 nsew
rlabel metal2 s 27216 30573 27216 30573 4 gnd
port 514 nsew
rlabel metal2 s 27216 31047 27216 31047 4 gnd
port 514 nsew
rlabel metal2 s 25968 30020 25968 30020 4 gnd
port 514 nsew
rlabel metal2 s 26448 30573 26448 30573 4 gnd
port 514 nsew
rlabel metal2 s 25200 31047 25200 31047 4 gnd
port 514 nsew
rlabel metal2 s 26448 30257 26448 30257 4 gnd
port 514 nsew
rlabel metal2 s 25200 30810 25200 30810 4 gnd
port 514 nsew
rlabel metal2 s 25968 29783 25968 29783 4 gnd
port 514 nsew
rlabel metal2 s 27216 31600 27216 31600 4 gnd
port 514 nsew
rlabel metal2 s 27216 30020 27216 30020 4 gnd
port 514 nsew
rlabel metal2 s 25968 28677 25968 28677 4 gnd
port 514 nsew
rlabel metal2 s 25200 29467 25200 29467 4 gnd
port 514 nsew
rlabel metal2 s 25968 30573 25968 30573 4 gnd
port 514 nsew
rlabel metal2 s 25200 30257 25200 30257 4 gnd
port 514 nsew
rlabel metal2 s 27216 30257 27216 30257 4 gnd
port 514 nsew
rlabel metal2 s 25968 30257 25968 30257 4 gnd
port 514 nsew
rlabel metal2 s 25968 27887 25968 27887 4 gnd
port 514 nsew
rlabel metal2 s 27216 28203 27216 28203 4 gnd
port 514 nsew
rlabel metal2 s 25200 27887 25200 27887 4 gnd
port 514 nsew
rlabel metal2 s 26448 27650 26448 27650 4 gnd
port 514 nsew
rlabel metal2 s 27216 27650 27216 27650 4 gnd
port 514 nsew
rlabel metal2 s 27216 27097 27216 27097 4 gnd
port 514 nsew
rlabel metal2 s 26448 28440 26448 28440 4 gnd
port 514 nsew
rlabel metal2 s 25968 28440 25968 28440 4 gnd
port 514 nsew
rlabel metal2 s 25968 27097 25968 27097 4 gnd
port 514 nsew
rlabel metal2 s 26448 27413 26448 27413 4 gnd
port 514 nsew
rlabel metal2 s 25200 28440 25200 28440 4 gnd
port 514 nsew
rlabel metal2 s 26448 28203 26448 28203 4 gnd
port 514 nsew
rlabel metal2 s 27216 25517 27216 25517 4 gnd
port 514 nsew
rlabel metal2 s 27216 28440 27216 28440 4 gnd
port 514 nsew
rlabel metal2 s 25968 26860 25968 26860 4 gnd
port 514 nsew
rlabel metal2 s 25200 27650 25200 27650 4 gnd
port 514 nsew
rlabel metal2 s 26448 26860 26448 26860 4 gnd
port 514 nsew
rlabel metal2 s 26448 26623 26448 26623 4 gnd
port 514 nsew
rlabel metal2 s 25968 25517 25968 25517 4 gnd
port 514 nsew
rlabel metal2 s 25200 26623 25200 26623 4 gnd
port 514 nsew
rlabel metal2 s 25200 26307 25200 26307 4 gnd
port 514 nsew
rlabel metal2 s 25968 27650 25968 27650 4 gnd
port 514 nsew
rlabel metal2 s 25200 27413 25200 27413 4 gnd
port 514 nsew
rlabel metal2 s 27216 26307 27216 26307 4 gnd
port 514 nsew
rlabel metal2 s 25200 26070 25200 26070 4 gnd
port 514 nsew
rlabel metal2 s 25968 26623 25968 26623 4 gnd
port 514 nsew
rlabel metal2 s 25968 26070 25968 26070 4 gnd
port 514 nsew
rlabel metal2 s 25200 25517 25200 25517 4 gnd
port 514 nsew
rlabel metal2 s 27216 26623 27216 26623 4 gnd
port 514 nsew
rlabel metal2 s 26448 27887 26448 27887 4 gnd
port 514 nsew
rlabel metal2 s 26448 26070 26448 26070 4 gnd
port 514 nsew
rlabel metal2 s 25968 28203 25968 28203 4 gnd
port 514 nsew
rlabel metal2 s 27216 27887 27216 27887 4 gnd
port 514 nsew
rlabel metal2 s 26448 25517 26448 25517 4 gnd
port 514 nsew
rlabel metal2 s 25200 25833 25200 25833 4 gnd
port 514 nsew
rlabel metal2 s 27216 26070 27216 26070 4 gnd
port 514 nsew
rlabel metal2 s 27216 25833 27216 25833 4 gnd
port 514 nsew
rlabel metal2 s 26448 27097 26448 27097 4 gnd
port 514 nsew
rlabel metal2 s 25968 26307 25968 26307 4 gnd
port 514 nsew
rlabel metal2 s 26448 26307 26448 26307 4 gnd
port 514 nsew
rlabel metal2 s 27216 27413 27216 27413 4 gnd
port 514 nsew
rlabel metal2 s 26448 25833 26448 25833 4 gnd
port 514 nsew
rlabel metal2 s 25200 26860 25200 26860 4 gnd
port 514 nsew
rlabel metal2 s 25200 27097 25200 27097 4 gnd
port 514 nsew
rlabel metal2 s 25200 28203 25200 28203 4 gnd
port 514 nsew
rlabel metal2 s 25968 27413 25968 27413 4 gnd
port 514 nsew
rlabel metal2 s 27216 26860 27216 26860 4 gnd
port 514 nsew
rlabel metal2 s 25968 25833 25968 25833 4 gnd
port 514 nsew
rlabel metal2 s 27696 27097 27696 27097 4 gnd
port 514 nsew
rlabel metal2 s 28944 28440 28944 28440 4 gnd
port 514 nsew
rlabel metal2 s 28944 26623 28944 26623 4 gnd
port 514 nsew
rlabel metal2 s 27696 27413 27696 27413 4 gnd
port 514 nsew
rlabel metal2 s 28944 25833 28944 25833 4 gnd
port 514 nsew
rlabel metal2 s 29712 27097 29712 27097 4 gnd
port 514 nsew
rlabel metal2 s 28944 25517 28944 25517 4 gnd
port 514 nsew
rlabel metal2 s 28464 25517 28464 25517 4 gnd
port 514 nsew
rlabel metal2 s 29712 25833 29712 25833 4 gnd
port 514 nsew
rlabel metal2 s 27696 28440 27696 28440 4 gnd
port 514 nsew
rlabel metal2 s 28944 27887 28944 27887 4 gnd
port 514 nsew
rlabel metal2 s 27696 26860 27696 26860 4 gnd
port 514 nsew
rlabel metal2 s 28464 26070 28464 26070 4 gnd
port 514 nsew
rlabel metal2 s 27696 25517 27696 25517 4 gnd
port 514 nsew
rlabel metal2 s 29712 26623 29712 26623 4 gnd
port 514 nsew
rlabel metal2 s 29712 28440 29712 28440 4 gnd
port 514 nsew
rlabel metal2 s 28944 26860 28944 26860 4 gnd
port 514 nsew
rlabel metal2 s 29712 28203 29712 28203 4 gnd
port 514 nsew
rlabel metal2 s 28464 28440 28464 28440 4 gnd
port 514 nsew
rlabel metal2 s 28464 27413 28464 27413 4 gnd
port 514 nsew
rlabel metal2 s 29712 27887 29712 27887 4 gnd
port 514 nsew
rlabel metal2 s 29712 26860 29712 26860 4 gnd
port 514 nsew
rlabel metal2 s 27696 26623 27696 26623 4 gnd
port 514 nsew
rlabel metal2 s 27696 27887 27696 27887 4 gnd
port 514 nsew
rlabel metal2 s 28944 27413 28944 27413 4 gnd
port 514 nsew
rlabel metal2 s 29712 27413 29712 27413 4 gnd
port 514 nsew
rlabel metal2 s 28944 28203 28944 28203 4 gnd
port 514 nsew
rlabel metal2 s 28944 26307 28944 26307 4 gnd
port 514 nsew
rlabel metal2 s 29712 25517 29712 25517 4 gnd
port 514 nsew
rlabel metal2 s 27696 27650 27696 27650 4 gnd
port 514 nsew
rlabel metal2 s 28944 26070 28944 26070 4 gnd
port 514 nsew
rlabel metal2 s 28464 27097 28464 27097 4 gnd
port 514 nsew
rlabel metal2 s 28464 28203 28464 28203 4 gnd
port 514 nsew
rlabel metal2 s 28464 26623 28464 26623 4 gnd
port 514 nsew
rlabel metal2 s 28464 25833 28464 25833 4 gnd
port 514 nsew
rlabel metal2 s 28464 26307 28464 26307 4 gnd
port 514 nsew
rlabel metal2 s 27696 26307 27696 26307 4 gnd
port 514 nsew
rlabel metal2 s 29712 26070 29712 26070 4 gnd
port 514 nsew
rlabel metal2 s 29712 26307 29712 26307 4 gnd
port 514 nsew
rlabel metal2 s 28944 27650 28944 27650 4 gnd
port 514 nsew
rlabel metal2 s 28464 27650 28464 27650 4 gnd
port 514 nsew
rlabel metal2 s 28464 27887 28464 27887 4 gnd
port 514 nsew
rlabel metal2 s 29712 27650 29712 27650 4 gnd
port 514 nsew
rlabel metal2 s 28464 26860 28464 26860 4 gnd
port 514 nsew
rlabel metal2 s 27696 28203 27696 28203 4 gnd
port 514 nsew
rlabel metal2 s 27696 26070 27696 26070 4 gnd
port 514 nsew
rlabel metal2 s 28944 27097 28944 27097 4 gnd
port 514 nsew
rlabel metal2 s 27696 25833 27696 25833 4 gnd
port 514 nsew
rlabel metal2 s 38448 36893 38448 36893 4 gnd
port 514 nsew
rlabel metal2 s 38448 37920 38448 37920 4 gnd
port 514 nsew
rlabel metal2 s 39696 35550 39696 35550 4 gnd
port 514 nsew
rlabel metal2 s 38928 37130 38928 37130 4 gnd
port 514 nsew
rlabel metal2 s 38448 34997 38448 34997 4 gnd
port 514 nsew
rlabel metal2 s 37680 37130 37680 37130 4 gnd
port 514 nsew
rlabel metal2 s 39696 37367 39696 37367 4 gnd
port 514 nsew
rlabel metal2 s 39696 37920 39696 37920 4 gnd
port 514 nsew
rlabel metal2 s 38448 35787 38448 35787 4 gnd
port 514 nsew
rlabel metal2 s 37680 35313 37680 35313 4 gnd
port 514 nsew
rlabel metal2 s 38928 36577 38928 36577 4 gnd
port 514 nsew
rlabel metal2 s 37680 36103 37680 36103 4 gnd
port 514 nsew
rlabel metal2 s 38928 37683 38928 37683 4 gnd
port 514 nsew
rlabel metal2 s 39696 37130 39696 37130 4 gnd
port 514 nsew
rlabel metal2 s 38448 37683 38448 37683 4 gnd
port 514 nsew
rlabel metal2 s 39696 34997 39696 34997 4 gnd
port 514 nsew
rlabel metal2 s 38928 34997 38928 34997 4 gnd
port 514 nsew
rlabel metal2 s 39696 35313 39696 35313 4 gnd
port 514 nsew
rlabel metal2 s 39696 35787 39696 35787 4 gnd
port 514 nsew
rlabel metal2 s 37680 37367 37680 37367 4 gnd
port 514 nsew
rlabel metal2 s 38928 35313 38928 35313 4 gnd
port 514 nsew
rlabel metal2 s 38448 37367 38448 37367 4 gnd
port 514 nsew
rlabel metal2 s 38928 35787 38928 35787 4 gnd
port 514 nsew
rlabel metal2 s 38448 36103 38448 36103 4 gnd
port 514 nsew
rlabel metal2 s 37680 36340 37680 36340 4 gnd
port 514 nsew
rlabel metal2 s 38448 36577 38448 36577 4 gnd
port 514 nsew
rlabel metal2 s 37680 36577 37680 36577 4 gnd
port 514 nsew
rlabel metal2 s 39696 37683 39696 37683 4 gnd
port 514 nsew
rlabel metal2 s 39696 36340 39696 36340 4 gnd
port 514 nsew
rlabel metal2 s 38928 36103 38928 36103 4 gnd
port 514 nsew
rlabel metal2 s 39696 36103 39696 36103 4 gnd
port 514 nsew
rlabel metal2 s 37680 37920 37680 37920 4 gnd
port 514 nsew
rlabel metal2 s 38928 36340 38928 36340 4 gnd
port 514 nsew
rlabel metal2 s 38448 37130 38448 37130 4 gnd
port 514 nsew
rlabel metal2 s 39696 36893 39696 36893 4 gnd
port 514 nsew
rlabel metal2 s 37680 37683 37680 37683 4 gnd
port 514 nsew
rlabel metal2 s 37680 35550 37680 35550 4 gnd
port 514 nsew
rlabel metal2 s 39696 36577 39696 36577 4 gnd
port 514 nsew
rlabel metal2 s 37680 34997 37680 34997 4 gnd
port 514 nsew
rlabel metal2 s 38928 36893 38928 36893 4 gnd
port 514 nsew
rlabel metal2 s 38448 35550 38448 35550 4 gnd
port 514 nsew
rlabel metal2 s 37680 36893 37680 36893 4 gnd
port 514 nsew
rlabel metal2 s 38928 37920 38928 37920 4 gnd
port 514 nsew
rlabel metal2 s 37680 35787 37680 35787 4 gnd
port 514 nsew
rlabel metal2 s 38448 36340 38448 36340 4 gnd
port 514 nsew
rlabel metal2 s 38448 35313 38448 35313 4 gnd
port 514 nsew
rlabel metal2 s 38928 37367 38928 37367 4 gnd
port 514 nsew
rlabel metal2 s 38928 35550 38928 35550 4 gnd
port 514 nsew
rlabel metal2 s 36432 35550 36432 35550 4 gnd
port 514 nsew
rlabel metal2 s 36432 36893 36432 36893 4 gnd
port 514 nsew
rlabel metal2 s 35184 35550 35184 35550 4 gnd
port 514 nsew
rlabel metal2 s 35184 35313 35184 35313 4 gnd
port 514 nsew
rlabel metal2 s 37200 36340 37200 36340 4 gnd
port 514 nsew
rlabel metal2 s 35184 35787 35184 35787 4 gnd
port 514 nsew
rlabel metal2 s 37200 36893 37200 36893 4 gnd
port 514 nsew
rlabel metal2 s 36432 36103 36432 36103 4 gnd
port 514 nsew
rlabel metal2 s 35184 37130 35184 37130 4 gnd
port 514 nsew
rlabel metal2 s 36432 36577 36432 36577 4 gnd
port 514 nsew
rlabel metal2 s 37200 37130 37200 37130 4 gnd
port 514 nsew
rlabel metal2 s 35184 37920 35184 37920 4 gnd
port 514 nsew
rlabel metal2 s 35184 34997 35184 34997 4 gnd
port 514 nsew
rlabel metal2 s 36432 35313 36432 35313 4 gnd
port 514 nsew
rlabel metal2 s 35952 36577 35952 36577 4 gnd
port 514 nsew
rlabel metal2 s 35952 35550 35952 35550 4 gnd
port 514 nsew
rlabel metal2 s 37200 36103 37200 36103 4 gnd
port 514 nsew
rlabel metal2 s 35952 36340 35952 36340 4 gnd
port 514 nsew
rlabel metal2 s 37200 36577 37200 36577 4 gnd
port 514 nsew
rlabel metal2 s 35952 36893 35952 36893 4 gnd
port 514 nsew
rlabel metal2 s 35184 36340 35184 36340 4 gnd
port 514 nsew
rlabel metal2 s 37200 37920 37200 37920 4 gnd
port 514 nsew
rlabel metal2 s 36432 37920 36432 37920 4 gnd
port 514 nsew
rlabel metal2 s 35184 36893 35184 36893 4 gnd
port 514 nsew
rlabel metal2 s 36432 34997 36432 34997 4 gnd
port 514 nsew
rlabel metal2 s 35952 37920 35952 37920 4 gnd
port 514 nsew
rlabel metal2 s 35184 36103 35184 36103 4 gnd
port 514 nsew
rlabel metal2 s 35952 37683 35952 37683 4 gnd
port 514 nsew
rlabel metal2 s 37200 37683 37200 37683 4 gnd
port 514 nsew
rlabel metal2 s 37200 35313 37200 35313 4 gnd
port 514 nsew
rlabel metal2 s 36432 37683 36432 37683 4 gnd
port 514 nsew
rlabel metal2 s 36432 36340 36432 36340 4 gnd
port 514 nsew
rlabel metal2 s 35952 36103 35952 36103 4 gnd
port 514 nsew
rlabel metal2 s 35952 35787 35952 35787 4 gnd
port 514 nsew
rlabel metal2 s 37200 35787 37200 35787 4 gnd
port 514 nsew
rlabel metal2 s 37200 37367 37200 37367 4 gnd
port 514 nsew
rlabel metal2 s 35952 37367 35952 37367 4 gnd
port 514 nsew
rlabel metal2 s 35952 34997 35952 34997 4 gnd
port 514 nsew
rlabel metal2 s 37200 35550 37200 35550 4 gnd
port 514 nsew
rlabel metal2 s 37200 34997 37200 34997 4 gnd
port 514 nsew
rlabel metal2 s 36432 37367 36432 37367 4 gnd
port 514 nsew
rlabel metal2 s 35952 37130 35952 37130 4 gnd
port 514 nsew
rlabel metal2 s 35184 37683 35184 37683 4 gnd
port 514 nsew
rlabel metal2 s 35184 37367 35184 37367 4 gnd
port 514 nsew
rlabel metal2 s 36432 35787 36432 35787 4 gnd
port 514 nsew
rlabel metal2 s 35184 36577 35184 36577 4 gnd
port 514 nsew
rlabel metal2 s 36432 37130 36432 37130 4 gnd
port 514 nsew
rlabel metal2 s 35952 35313 35952 35313 4 gnd
port 514 nsew
rlabel metal2 s 35184 33733 35184 33733 4 gnd
port 514 nsew
rlabel metal2 s 36432 32627 36432 32627 4 gnd
port 514 nsew
rlabel metal2 s 37200 32627 37200 32627 4 gnd
port 514 nsew
rlabel metal2 s 37200 32943 37200 32943 4 gnd
port 514 nsew
rlabel metal2 s 35952 32627 35952 32627 4 gnd
port 514 nsew
rlabel metal2 s 36432 33180 36432 33180 4 gnd
port 514 nsew
rlabel metal2 s 35952 32943 35952 32943 4 gnd
port 514 nsew
rlabel metal2 s 35184 32390 35184 32390 4 gnd
port 514 nsew
rlabel metal2 s 35184 33180 35184 33180 4 gnd
port 514 nsew
rlabel metal2 s 36432 32153 36432 32153 4 gnd
port 514 nsew
rlabel metal2 s 35952 34207 35952 34207 4 gnd
port 514 nsew
rlabel metal2 s 37200 34760 37200 34760 4 gnd
port 514 nsew
rlabel metal2 s 36432 33417 36432 33417 4 gnd
port 514 nsew
rlabel metal2 s 37200 33970 37200 33970 4 gnd
port 514 nsew
rlabel metal2 s 36432 32943 36432 32943 4 gnd
port 514 nsew
rlabel metal2 s 37200 34523 37200 34523 4 gnd
port 514 nsew
rlabel metal2 s 35184 34207 35184 34207 4 gnd
port 514 nsew
rlabel metal2 s 35952 33970 35952 33970 4 gnd
port 514 nsew
rlabel metal2 s 36432 31837 36432 31837 4 gnd
port 514 nsew
rlabel metal2 s 36432 33733 36432 33733 4 gnd
port 514 nsew
rlabel metal2 s 36432 32390 36432 32390 4 gnd
port 514 nsew
rlabel metal2 s 37200 32390 37200 32390 4 gnd
port 514 nsew
rlabel metal2 s 35184 33417 35184 33417 4 gnd
port 514 nsew
rlabel metal2 s 37200 33417 37200 33417 4 gnd
port 514 nsew
rlabel metal2 s 37200 33180 37200 33180 4 gnd
port 514 nsew
rlabel metal2 s 37200 33733 37200 33733 4 gnd
port 514 nsew
rlabel metal2 s 35184 32153 35184 32153 4 gnd
port 514 nsew
rlabel metal2 s 35952 34760 35952 34760 4 gnd
port 514 nsew
rlabel metal2 s 37200 32153 37200 32153 4 gnd
port 514 nsew
rlabel metal2 s 35952 33180 35952 33180 4 gnd
port 514 nsew
rlabel metal2 s 37200 31837 37200 31837 4 gnd
port 514 nsew
rlabel metal2 s 35184 32943 35184 32943 4 gnd
port 514 nsew
rlabel metal2 s 35952 33417 35952 33417 4 gnd
port 514 nsew
rlabel metal2 s 36432 34760 36432 34760 4 gnd
port 514 nsew
rlabel metal2 s 35952 33733 35952 33733 4 gnd
port 514 nsew
rlabel metal2 s 35952 31837 35952 31837 4 gnd
port 514 nsew
rlabel metal2 s 36432 34207 36432 34207 4 gnd
port 514 nsew
rlabel metal2 s 35184 34760 35184 34760 4 gnd
port 514 nsew
rlabel metal2 s 37200 34207 37200 34207 4 gnd
port 514 nsew
rlabel metal2 s 35184 32627 35184 32627 4 gnd
port 514 nsew
rlabel metal2 s 35952 34523 35952 34523 4 gnd
port 514 nsew
rlabel metal2 s 35184 33970 35184 33970 4 gnd
port 514 nsew
rlabel metal2 s 36432 34523 36432 34523 4 gnd
port 514 nsew
rlabel metal2 s 35952 32390 35952 32390 4 gnd
port 514 nsew
rlabel metal2 s 35184 34523 35184 34523 4 gnd
port 514 nsew
rlabel metal2 s 36432 33970 36432 33970 4 gnd
port 514 nsew
rlabel metal2 s 35184 31837 35184 31837 4 gnd
port 514 nsew
rlabel metal2 s 35952 32153 35952 32153 4 gnd
port 514 nsew
rlabel metal2 s 38928 33733 38928 33733 4 gnd
port 514 nsew
rlabel metal2 s 38928 33970 38928 33970 4 gnd
port 514 nsew
rlabel metal2 s 37680 31837 37680 31837 4 gnd
port 514 nsew
rlabel metal2 s 38448 34760 38448 34760 4 gnd
port 514 nsew
rlabel metal2 s 38928 32153 38928 32153 4 gnd
port 514 nsew
rlabel metal2 s 38928 34523 38928 34523 4 gnd
port 514 nsew
rlabel metal2 s 37680 32390 37680 32390 4 gnd
port 514 nsew
rlabel metal2 s 37680 33970 37680 33970 4 gnd
port 514 nsew
rlabel metal2 s 39696 33180 39696 33180 4 gnd
port 514 nsew
rlabel metal2 s 38928 32943 38928 32943 4 gnd
port 514 nsew
rlabel metal2 s 38448 31837 38448 31837 4 gnd
port 514 nsew
rlabel metal2 s 39696 34207 39696 34207 4 gnd
port 514 nsew
rlabel metal2 s 39696 32627 39696 32627 4 gnd
port 514 nsew
rlabel metal2 s 38928 32390 38928 32390 4 gnd
port 514 nsew
rlabel metal2 s 37680 33180 37680 33180 4 gnd
port 514 nsew
rlabel metal2 s 39696 32153 39696 32153 4 gnd
port 514 nsew
rlabel metal2 s 37680 33733 37680 33733 4 gnd
port 514 nsew
rlabel metal2 s 38448 32390 38448 32390 4 gnd
port 514 nsew
rlabel metal2 s 37680 32627 37680 32627 4 gnd
port 514 nsew
rlabel metal2 s 39696 32390 39696 32390 4 gnd
port 514 nsew
rlabel metal2 s 38448 32153 38448 32153 4 gnd
port 514 nsew
rlabel metal2 s 38448 33970 38448 33970 4 gnd
port 514 nsew
rlabel metal2 s 37680 34207 37680 34207 4 gnd
port 514 nsew
rlabel metal2 s 39696 33733 39696 33733 4 gnd
port 514 nsew
rlabel metal2 s 37680 34523 37680 34523 4 gnd
port 514 nsew
rlabel metal2 s 38928 31837 38928 31837 4 gnd
port 514 nsew
rlabel metal2 s 37680 32943 37680 32943 4 gnd
port 514 nsew
rlabel metal2 s 38928 32627 38928 32627 4 gnd
port 514 nsew
rlabel metal2 s 38928 33417 38928 33417 4 gnd
port 514 nsew
rlabel metal2 s 37680 33417 37680 33417 4 gnd
port 514 nsew
rlabel metal2 s 38448 34207 38448 34207 4 gnd
port 514 nsew
rlabel metal2 s 39696 33417 39696 33417 4 gnd
port 514 nsew
rlabel metal2 s 38928 34760 38928 34760 4 gnd
port 514 nsew
rlabel metal2 s 39696 32943 39696 32943 4 gnd
port 514 nsew
rlabel metal2 s 38448 33180 38448 33180 4 gnd
port 514 nsew
rlabel metal2 s 38448 33733 38448 33733 4 gnd
port 514 nsew
rlabel metal2 s 39696 34760 39696 34760 4 gnd
port 514 nsew
rlabel metal2 s 38928 34207 38928 34207 4 gnd
port 514 nsew
rlabel metal2 s 38448 33417 38448 33417 4 gnd
port 514 nsew
rlabel metal2 s 39696 34523 39696 34523 4 gnd
port 514 nsew
rlabel metal2 s 37680 34760 37680 34760 4 gnd
port 514 nsew
rlabel metal2 s 38448 32627 38448 32627 4 gnd
port 514 nsew
rlabel metal2 s 38448 32943 38448 32943 4 gnd
port 514 nsew
rlabel metal2 s 39696 33970 39696 33970 4 gnd
port 514 nsew
rlabel metal2 s 38448 34523 38448 34523 4 gnd
port 514 nsew
rlabel metal2 s 39696 31837 39696 31837 4 gnd
port 514 nsew
rlabel metal2 s 38928 33180 38928 33180 4 gnd
port 514 nsew
rlabel metal2 s 37680 32153 37680 32153 4 gnd
port 514 nsew
rlabel metal2 s 32688 34997 32688 34997 4 gnd
port 514 nsew
rlabel metal2 s 33456 36103 33456 36103 4 gnd
port 514 nsew
rlabel metal2 s 34704 37920 34704 37920 4 gnd
port 514 nsew
rlabel metal2 s 32688 37367 32688 37367 4 gnd
port 514 nsew
rlabel metal2 s 33456 37683 33456 37683 4 gnd
port 514 nsew
rlabel metal2 s 33936 36340 33936 36340 4 gnd
port 514 nsew
rlabel metal2 s 33936 35313 33936 35313 4 gnd
port 514 nsew
rlabel metal2 s 34704 35550 34704 35550 4 gnd
port 514 nsew
rlabel metal2 s 33456 35313 33456 35313 4 gnd
port 514 nsew
rlabel metal2 s 32688 35313 32688 35313 4 gnd
port 514 nsew
rlabel metal2 s 32688 36103 32688 36103 4 gnd
port 514 nsew
rlabel metal2 s 33456 37920 33456 37920 4 gnd
port 514 nsew
rlabel metal2 s 33936 36893 33936 36893 4 gnd
port 514 nsew
rlabel metal2 s 33936 35550 33936 35550 4 gnd
port 514 nsew
rlabel metal2 s 33936 34997 33936 34997 4 gnd
port 514 nsew
rlabel metal2 s 33456 36577 33456 36577 4 gnd
port 514 nsew
rlabel metal2 s 33936 35787 33936 35787 4 gnd
port 514 nsew
rlabel metal2 s 33456 36340 33456 36340 4 gnd
port 514 nsew
rlabel metal2 s 34704 37683 34704 37683 4 gnd
port 514 nsew
rlabel metal2 s 33456 35550 33456 35550 4 gnd
port 514 nsew
rlabel metal2 s 32688 36340 32688 36340 4 gnd
port 514 nsew
rlabel metal2 s 32688 35550 32688 35550 4 gnd
port 514 nsew
rlabel metal2 s 34704 35313 34704 35313 4 gnd
port 514 nsew
rlabel metal2 s 32688 37920 32688 37920 4 gnd
port 514 nsew
rlabel metal2 s 33936 37683 33936 37683 4 gnd
port 514 nsew
rlabel metal2 s 33936 36577 33936 36577 4 gnd
port 514 nsew
rlabel metal2 s 32688 37130 32688 37130 4 gnd
port 514 nsew
rlabel metal2 s 32688 37683 32688 37683 4 gnd
port 514 nsew
rlabel metal2 s 34704 37130 34704 37130 4 gnd
port 514 nsew
rlabel metal2 s 34704 36893 34704 36893 4 gnd
port 514 nsew
rlabel metal2 s 34704 37367 34704 37367 4 gnd
port 514 nsew
rlabel metal2 s 33936 36103 33936 36103 4 gnd
port 514 nsew
rlabel metal2 s 34704 36577 34704 36577 4 gnd
port 514 nsew
rlabel metal2 s 32688 35787 32688 35787 4 gnd
port 514 nsew
rlabel metal2 s 34704 36340 34704 36340 4 gnd
port 514 nsew
rlabel metal2 s 34704 35787 34704 35787 4 gnd
port 514 nsew
rlabel metal2 s 33456 34997 33456 34997 4 gnd
port 514 nsew
rlabel metal2 s 33456 37130 33456 37130 4 gnd
port 514 nsew
rlabel metal2 s 32688 36577 32688 36577 4 gnd
port 514 nsew
rlabel metal2 s 34704 36103 34704 36103 4 gnd
port 514 nsew
rlabel metal2 s 34704 34997 34704 34997 4 gnd
port 514 nsew
rlabel metal2 s 33936 37130 33936 37130 4 gnd
port 514 nsew
rlabel metal2 s 33936 37367 33936 37367 4 gnd
port 514 nsew
rlabel metal2 s 33456 36893 33456 36893 4 gnd
port 514 nsew
rlabel metal2 s 33456 35787 33456 35787 4 gnd
port 514 nsew
rlabel metal2 s 33456 37367 33456 37367 4 gnd
port 514 nsew
rlabel metal2 s 33936 37920 33936 37920 4 gnd
port 514 nsew
rlabel metal2 s 32688 36893 32688 36893 4 gnd
port 514 nsew
rlabel metal2 s 32208 35313 32208 35313 4 gnd
port 514 nsew
rlabel metal2 s 32208 37920 32208 37920 4 gnd
port 514 nsew
rlabel metal2 s 31440 37130 31440 37130 4 gnd
port 514 nsew
rlabel metal2 s 30960 35550 30960 35550 4 gnd
port 514 nsew
rlabel metal2 s 30192 35550 30192 35550 4 gnd
port 514 nsew
rlabel metal2 s 30192 37920 30192 37920 4 gnd
port 514 nsew
rlabel metal2 s 30960 37130 30960 37130 4 gnd
port 514 nsew
rlabel metal2 s 30192 36340 30192 36340 4 gnd
port 514 nsew
rlabel metal2 s 31440 36103 31440 36103 4 gnd
port 514 nsew
rlabel metal2 s 30960 37920 30960 37920 4 gnd
port 514 nsew
rlabel metal2 s 32208 36103 32208 36103 4 gnd
port 514 nsew
rlabel metal2 s 32208 37130 32208 37130 4 gnd
port 514 nsew
rlabel metal2 s 30192 35313 30192 35313 4 gnd
port 514 nsew
rlabel metal2 s 31440 36893 31440 36893 4 gnd
port 514 nsew
rlabel metal2 s 30960 36103 30960 36103 4 gnd
port 514 nsew
rlabel metal2 s 31440 37683 31440 37683 4 gnd
port 514 nsew
rlabel metal2 s 32208 37683 32208 37683 4 gnd
port 514 nsew
rlabel metal2 s 30960 35313 30960 35313 4 gnd
port 514 nsew
rlabel metal2 s 32208 34997 32208 34997 4 gnd
port 514 nsew
rlabel metal2 s 30960 36577 30960 36577 4 gnd
port 514 nsew
rlabel metal2 s 30192 36577 30192 36577 4 gnd
port 514 nsew
rlabel metal2 s 30192 34997 30192 34997 4 gnd
port 514 nsew
rlabel metal2 s 30192 37683 30192 37683 4 gnd
port 514 nsew
rlabel metal2 s 32208 36340 32208 36340 4 gnd
port 514 nsew
rlabel metal2 s 30192 36893 30192 36893 4 gnd
port 514 nsew
rlabel metal2 s 32208 35787 32208 35787 4 gnd
port 514 nsew
rlabel metal2 s 30960 37367 30960 37367 4 gnd
port 514 nsew
rlabel metal2 s 30192 36103 30192 36103 4 gnd
port 514 nsew
rlabel metal2 s 31440 35313 31440 35313 4 gnd
port 514 nsew
rlabel metal2 s 30960 34997 30960 34997 4 gnd
port 514 nsew
rlabel metal2 s 32208 35550 32208 35550 4 gnd
port 514 nsew
rlabel metal2 s 30192 37367 30192 37367 4 gnd
port 514 nsew
rlabel metal2 s 32208 37367 32208 37367 4 gnd
port 514 nsew
rlabel metal2 s 30960 36893 30960 36893 4 gnd
port 514 nsew
rlabel metal2 s 31440 35787 31440 35787 4 gnd
port 514 nsew
rlabel metal2 s 30960 35787 30960 35787 4 gnd
port 514 nsew
rlabel metal2 s 31440 35550 31440 35550 4 gnd
port 514 nsew
rlabel metal2 s 31440 37367 31440 37367 4 gnd
port 514 nsew
rlabel metal2 s 30192 35787 30192 35787 4 gnd
port 514 nsew
rlabel metal2 s 31440 36340 31440 36340 4 gnd
port 514 nsew
rlabel metal2 s 32208 36893 32208 36893 4 gnd
port 514 nsew
rlabel metal2 s 30192 37130 30192 37130 4 gnd
port 514 nsew
rlabel metal2 s 31440 37920 31440 37920 4 gnd
port 514 nsew
rlabel metal2 s 30960 37683 30960 37683 4 gnd
port 514 nsew
rlabel metal2 s 31440 34997 31440 34997 4 gnd
port 514 nsew
rlabel metal2 s 31440 36577 31440 36577 4 gnd
port 514 nsew
rlabel metal2 s 30960 36340 30960 36340 4 gnd
port 514 nsew
rlabel metal2 s 32208 36577 32208 36577 4 gnd
port 514 nsew
rlabel metal2 s 32208 33733 32208 33733 4 gnd
port 514 nsew
rlabel metal2 s 30192 33417 30192 33417 4 gnd
port 514 nsew
rlabel metal2 s 30960 33970 30960 33970 4 gnd
port 514 nsew
rlabel metal2 s 31440 33970 31440 33970 4 gnd
port 514 nsew
rlabel metal2 s 30192 34760 30192 34760 4 gnd
port 514 nsew
rlabel metal2 s 30192 32390 30192 32390 4 gnd
port 514 nsew
rlabel metal2 s 30960 32153 30960 32153 4 gnd
port 514 nsew
rlabel metal2 s 31440 32627 31440 32627 4 gnd
port 514 nsew
rlabel metal2 s 30960 33417 30960 33417 4 gnd
port 514 nsew
rlabel metal2 s 30960 34760 30960 34760 4 gnd
port 514 nsew
rlabel metal2 s 32208 31837 32208 31837 4 gnd
port 514 nsew
rlabel metal2 s 30960 32943 30960 32943 4 gnd
port 514 nsew
rlabel metal2 s 30192 32627 30192 32627 4 gnd
port 514 nsew
rlabel metal2 s 32208 33417 32208 33417 4 gnd
port 514 nsew
rlabel metal2 s 31440 33417 31440 33417 4 gnd
port 514 nsew
rlabel metal2 s 32208 32627 32208 32627 4 gnd
port 514 nsew
rlabel metal2 s 31440 33180 31440 33180 4 gnd
port 514 nsew
rlabel metal2 s 32208 33970 32208 33970 4 gnd
port 514 nsew
rlabel metal2 s 31440 33733 31440 33733 4 gnd
port 514 nsew
rlabel metal2 s 30192 34207 30192 34207 4 gnd
port 514 nsew
rlabel metal2 s 30192 33733 30192 33733 4 gnd
port 514 nsew
rlabel metal2 s 30192 32943 30192 32943 4 gnd
port 514 nsew
rlabel metal2 s 32208 32943 32208 32943 4 gnd
port 514 nsew
rlabel metal2 s 32208 34523 32208 34523 4 gnd
port 514 nsew
rlabel metal2 s 32208 32390 32208 32390 4 gnd
port 514 nsew
rlabel metal2 s 32208 33180 32208 33180 4 gnd
port 514 nsew
rlabel metal2 s 31440 32153 31440 32153 4 gnd
port 514 nsew
rlabel metal2 s 32208 34207 32208 34207 4 gnd
port 514 nsew
rlabel metal2 s 30192 32153 30192 32153 4 gnd
port 514 nsew
rlabel metal2 s 30960 31837 30960 31837 4 gnd
port 514 nsew
rlabel metal2 s 31440 34207 31440 34207 4 gnd
port 514 nsew
rlabel metal2 s 30192 34523 30192 34523 4 gnd
port 514 nsew
rlabel metal2 s 30192 33970 30192 33970 4 gnd
port 514 nsew
rlabel metal2 s 30960 33180 30960 33180 4 gnd
port 514 nsew
rlabel metal2 s 31440 32390 31440 32390 4 gnd
port 514 nsew
rlabel metal2 s 30192 33180 30192 33180 4 gnd
port 514 nsew
rlabel metal2 s 30960 34523 30960 34523 4 gnd
port 514 nsew
rlabel metal2 s 30960 32390 30960 32390 4 gnd
port 514 nsew
rlabel metal2 s 31440 31837 31440 31837 4 gnd
port 514 nsew
rlabel metal2 s 31440 34760 31440 34760 4 gnd
port 514 nsew
rlabel metal2 s 32208 34760 32208 34760 4 gnd
port 514 nsew
rlabel metal2 s 30960 32627 30960 32627 4 gnd
port 514 nsew
rlabel metal2 s 30192 31837 30192 31837 4 gnd
port 514 nsew
rlabel metal2 s 30960 34207 30960 34207 4 gnd
port 514 nsew
rlabel metal2 s 32208 32153 32208 32153 4 gnd
port 514 nsew
rlabel metal2 s 30960 33733 30960 33733 4 gnd
port 514 nsew
rlabel metal2 s 31440 32943 31440 32943 4 gnd
port 514 nsew
rlabel metal2 s 31440 34523 31440 34523 4 gnd
port 514 nsew
rlabel metal2 s 33456 33417 33456 33417 4 gnd
port 514 nsew
rlabel metal2 s 33456 33970 33456 33970 4 gnd
port 514 nsew
rlabel metal2 s 33456 32943 33456 32943 4 gnd
port 514 nsew
rlabel metal2 s 33936 32627 33936 32627 4 gnd
port 514 nsew
rlabel metal2 s 32688 31837 32688 31837 4 gnd
port 514 nsew
rlabel metal2 s 34704 32943 34704 32943 4 gnd
port 514 nsew
rlabel metal2 s 32688 33970 32688 33970 4 gnd
port 514 nsew
rlabel metal2 s 34704 34523 34704 34523 4 gnd
port 514 nsew
rlabel metal2 s 33456 34523 33456 34523 4 gnd
port 514 nsew
rlabel metal2 s 32688 33180 32688 33180 4 gnd
port 514 nsew
rlabel metal2 s 33456 34760 33456 34760 4 gnd
port 514 nsew
rlabel metal2 s 32688 33417 32688 33417 4 gnd
port 514 nsew
rlabel metal2 s 33936 32390 33936 32390 4 gnd
port 514 nsew
rlabel metal2 s 34704 34207 34704 34207 4 gnd
port 514 nsew
rlabel metal2 s 33456 33180 33456 33180 4 gnd
port 514 nsew
rlabel metal2 s 34704 33180 34704 33180 4 gnd
port 514 nsew
rlabel metal2 s 33936 33180 33936 33180 4 gnd
port 514 nsew
rlabel metal2 s 34704 32153 34704 32153 4 gnd
port 514 nsew
rlabel metal2 s 33456 34207 33456 34207 4 gnd
port 514 nsew
rlabel metal2 s 33936 33733 33936 33733 4 gnd
port 514 nsew
rlabel metal2 s 34704 34760 34704 34760 4 gnd
port 514 nsew
rlabel metal2 s 33936 31837 33936 31837 4 gnd
port 514 nsew
rlabel metal2 s 34704 32390 34704 32390 4 gnd
port 514 nsew
rlabel metal2 s 33456 32390 33456 32390 4 gnd
port 514 nsew
rlabel metal2 s 32688 32627 32688 32627 4 gnd
port 514 nsew
rlabel metal2 s 34704 33417 34704 33417 4 gnd
port 514 nsew
rlabel metal2 s 33936 34207 33936 34207 4 gnd
port 514 nsew
rlabel metal2 s 33456 32153 33456 32153 4 gnd
port 514 nsew
rlabel metal2 s 32688 32943 32688 32943 4 gnd
port 514 nsew
rlabel metal2 s 33936 33417 33936 33417 4 gnd
port 514 nsew
rlabel metal2 s 32688 32390 32688 32390 4 gnd
port 514 nsew
rlabel metal2 s 33456 31837 33456 31837 4 gnd
port 514 nsew
rlabel metal2 s 32688 34760 32688 34760 4 gnd
port 514 nsew
rlabel metal2 s 32688 32153 32688 32153 4 gnd
port 514 nsew
rlabel metal2 s 33456 33733 33456 33733 4 gnd
port 514 nsew
rlabel metal2 s 33936 32943 33936 32943 4 gnd
port 514 nsew
rlabel metal2 s 34704 33970 34704 33970 4 gnd
port 514 nsew
rlabel metal2 s 33936 34760 33936 34760 4 gnd
port 514 nsew
rlabel metal2 s 33936 32153 33936 32153 4 gnd
port 514 nsew
rlabel metal2 s 32688 34523 32688 34523 4 gnd
port 514 nsew
rlabel metal2 s 34704 32627 34704 32627 4 gnd
port 514 nsew
rlabel metal2 s 34704 31837 34704 31837 4 gnd
port 514 nsew
rlabel metal2 s 32688 34207 32688 34207 4 gnd
port 514 nsew
rlabel metal2 s 32688 33733 32688 33733 4 gnd
port 514 nsew
rlabel metal2 s 33936 34523 33936 34523 4 gnd
port 514 nsew
rlabel metal2 s 34704 33733 34704 33733 4 gnd
port 514 nsew
rlabel metal2 s 33456 32627 33456 32627 4 gnd
port 514 nsew
rlabel metal2 s 33936 33970 33936 33970 4 gnd
port 514 nsew
rlabel metal2 s 34704 31047 34704 31047 4 gnd
port 514 nsew
rlabel metal2 s 32688 28993 32688 28993 4 gnd
port 514 nsew
rlabel metal2 s 33936 28993 33936 28993 4 gnd
port 514 nsew
rlabel metal2 s 33456 29467 33456 29467 4 gnd
port 514 nsew
rlabel metal2 s 33936 30257 33936 30257 4 gnd
port 514 nsew
rlabel metal2 s 33456 31363 33456 31363 4 gnd
port 514 nsew
rlabel metal2 s 33456 28993 33456 28993 4 gnd
port 514 nsew
rlabel metal2 s 33456 28677 33456 28677 4 gnd
port 514 nsew
rlabel metal2 s 32688 31047 32688 31047 4 gnd
port 514 nsew
rlabel metal2 s 33936 30810 33936 30810 4 gnd
port 514 nsew
rlabel metal2 s 33456 29783 33456 29783 4 gnd
port 514 nsew
rlabel metal2 s 33936 28677 33936 28677 4 gnd
port 514 nsew
rlabel metal2 s 34704 30020 34704 30020 4 gnd
port 514 nsew
rlabel metal2 s 32688 29467 32688 29467 4 gnd
port 514 nsew
rlabel metal2 s 33456 30020 33456 30020 4 gnd
port 514 nsew
rlabel metal2 s 34704 29230 34704 29230 4 gnd
port 514 nsew
rlabel metal2 s 33936 30573 33936 30573 4 gnd
port 514 nsew
rlabel metal2 s 33456 31600 33456 31600 4 gnd
port 514 nsew
rlabel metal2 s 32688 30573 32688 30573 4 gnd
port 514 nsew
rlabel metal2 s 32688 30020 32688 30020 4 gnd
port 514 nsew
rlabel metal2 s 34704 28993 34704 28993 4 gnd
port 514 nsew
rlabel metal2 s 34704 30810 34704 30810 4 gnd
port 514 nsew
rlabel metal2 s 32688 28677 32688 28677 4 gnd
port 514 nsew
rlabel metal2 s 33936 31047 33936 31047 4 gnd
port 514 nsew
rlabel metal2 s 33456 29230 33456 29230 4 gnd
port 514 nsew
rlabel metal2 s 33936 30020 33936 30020 4 gnd
port 514 nsew
rlabel metal2 s 33936 29783 33936 29783 4 gnd
port 514 nsew
rlabel metal2 s 34704 31363 34704 31363 4 gnd
port 514 nsew
rlabel metal2 s 33456 30573 33456 30573 4 gnd
port 514 nsew
rlabel metal2 s 32688 30810 32688 30810 4 gnd
port 514 nsew
rlabel metal2 s 33936 29467 33936 29467 4 gnd
port 514 nsew
rlabel metal2 s 33936 31600 33936 31600 4 gnd
port 514 nsew
rlabel metal2 s 34704 28677 34704 28677 4 gnd
port 514 nsew
rlabel metal2 s 33456 30810 33456 30810 4 gnd
port 514 nsew
rlabel metal2 s 33936 31363 33936 31363 4 gnd
port 514 nsew
rlabel metal2 s 32688 30257 32688 30257 4 gnd
port 514 nsew
rlabel metal2 s 34704 31600 34704 31600 4 gnd
port 514 nsew
rlabel metal2 s 33456 31047 33456 31047 4 gnd
port 514 nsew
rlabel metal2 s 34704 30257 34704 30257 4 gnd
port 514 nsew
rlabel metal2 s 33936 29230 33936 29230 4 gnd
port 514 nsew
rlabel metal2 s 34704 30573 34704 30573 4 gnd
port 514 nsew
rlabel metal2 s 32688 29230 32688 29230 4 gnd
port 514 nsew
rlabel metal2 s 32688 31363 32688 31363 4 gnd
port 514 nsew
rlabel metal2 s 34704 29467 34704 29467 4 gnd
port 514 nsew
rlabel metal2 s 32688 31600 32688 31600 4 gnd
port 514 nsew
rlabel metal2 s 34704 29783 34704 29783 4 gnd
port 514 nsew
rlabel metal2 s 32688 29783 32688 29783 4 gnd
port 514 nsew
rlabel metal2 s 33456 30257 33456 30257 4 gnd
port 514 nsew
rlabel metal2 s 32208 29783 32208 29783 4 gnd
port 514 nsew
rlabel metal2 s 32208 29230 32208 29230 4 gnd
port 514 nsew
rlabel metal2 s 31440 30810 31440 30810 4 gnd
port 514 nsew
rlabel metal2 s 30192 31047 30192 31047 4 gnd
port 514 nsew
rlabel metal2 s 30960 29230 30960 29230 4 gnd
port 514 nsew
rlabel metal2 s 30960 30810 30960 30810 4 gnd
port 514 nsew
rlabel metal2 s 32208 30020 32208 30020 4 gnd
port 514 nsew
rlabel metal2 s 31440 30257 31440 30257 4 gnd
port 514 nsew
rlabel metal2 s 30192 31363 30192 31363 4 gnd
port 514 nsew
rlabel metal2 s 30960 30573 30960 30573 4 gnd
port 514 nsew
rlabel metal2 s 31440 30020 31440 30020 4 gnd
port 514 nsew
rlabel metal2 s 30960 28993 30960 28993 4 gnd
port 514 nsew
rlabel metal2 s 32208 30810 32208 30810 4 gnd
port 514 nsew
rlabel metal2 s 30960 30257 30960 30257 4 gnd
port 514 nsew
rlabel metal2 s 31440 30573 31440 30573 4 gnd
port 514 nsew
rlabel metal2 s 32208 30257 32208 30257 4 gnd
port 514 nsew
rlabel metal2 s 32208 30573 32208 30573 4 gnd
port 514 nsew
rlabel metal2 s 30192 30810 30192 30810 4 gnd
port 514 nsew
rlabel metal2 s 30960 29467 30960 29467 4 gnd
port 514 nsew
rlabel metal2 s 31440 31600 31440 31600 4 gnd
port 514 nsew
rlabel metal2 s 31440 29783 31440 29783 4 gnd
port 514 nsew
rlabel metal2 s 31440 29467 31440 29467 4 gnd
port 514 nsew
rlabel metal2 s 31440 28677 31440 28677 4 gnd
port 514 nsew
rlabel metal2 s 31440 29230 31440 29230 4 gnd
port 514 nsew
rlabel metal2 s 31440 31047 31440 31047 4 gnd
port 514 nsew
rlabel metal2 s 30960 31047 30960 31047 4 gnd
port 514 nsew
rlabel metal2 s 32208 31047 32208 31047 4 gnd
port 514 nsew
rlabel metal2 s 30192 31600 30192 31600 4 gnd
port 514 nsew
rlabel metal2 s 30192 30257 30192 30257 4 gnd
port 514 nsew
rlabel metal2 s 32208 28677 32208 28677 4 gnd
port 514 nsew
rlabel metal2 s 30960 31600 30960 31600 4 gnd
port 514 nsew
rlabel metal2 s 30192 30573 30192 30573 4 gnd
port 514 nsew
rlabel metal2 s 30960 31363 30960 31363 4 gnd
port 514 nsew
rlabel metal2 s 30192 29783 30192 29783 4 gnd
port 514 nsew
rlabel metal2 s 32208 29467 32208 29467 4 gnd
port 514 nsew
rlabel metal2 s 32208 28993 32208 28993 4 gnd
port 514 nsew
rlabel metal2 s 32208 31600 32208 31600 4 gnd
port 514 nsew
rlabel metal2 s 31440 28993 31440 28993 4 gnd
port 514 nsew
rlabel metal2 s 30192 28993 30192 28993 4 gnd
port 514 nsew
rlabel metal2 s 30192 29230 30192 29230 4 gnd
port 514 nsew
rlabel metal2 s 30192 29467 30192 29467 4 gnd
port 514 nsew
rlabel metal2 s 30192 30020 30192 30020 4 gnd
port 514 nsew
rlabel metal2 s 30960 29783 30960 29783 4 gnd
port 514 nsew
rlabel metal2 s 31440 31363 31440 31363 4 gnd
port 514 nsew
rlabel metal2 s 30960 30020 30960 30020 4 gnd
port 514 nsew
rlabel metal2 s 30192 28677 30192 28677 4 gnd
port 514 nsew
rlabel metal2 s 32208 31363 32208 31363 4 gnd
port 514 nsew
rlabel metal2 s 30960 28677 30960 28677 4 gnd
port 514 nsew
rlabel metal2 s 30960 26623 30960 26623 4 gnd
port 514 nsew
rlabel metal2 s 31440 27887 31440 27887 4 gnd
port 514 nsew
rlabel metal2 s 31440 26623 31440 26623 4 gnd
port 514 nsew
rlabel metal2 s 30960 25833 30960 25833 4 gnd
port 514 nsew
rlabel metal2 s 30192 27887 30192 27887 4 gnd
port 514 nsew
rlabel metal2 s 30192 26860 30192 26860 4 gnd
port 514 nsew
rlabel metal2 s 31440 27650 31440 27650 4 gnd
port 514 nsew
rlabel metal2 s 30960 28203 30960 28203 4 gnd
port 514 nsew
rlabel metal2 s 30960 27413 30960 27413 4 gnd
port 514 nsew
rlabel metal2 s 31440 25517 31440 25517 4 gnd
port 514 nsew
rlabel metal2 s 30192 27650 30192 27650 4 gnd
port 514 nsew
rlabel metal2 s 32208 26860 32208 26860 4 gnd
port 514 nsew
rlabel metal2 s 31440 26070 31440 26070 4 gnd
port 514 nsew
rlabel metal2 s 30192 28203 30192 28203 4 gnd
port 514 nsew
rlabel metal2 s 32208 26307 32208 26307 4 gnd
port 514 nsew
rlabel metal2 s 30960 26860 30960 26860 4 gnd
port 514 nsew
rlabel metal2 s 31440 28440 31440 28440 4 gnd
port 514 nsew
rlabel metal2 s 31440 26307 31440 26307 4 gnd
port 514 nsew
rlabel metal2 s 32208 28203 32208 28203 4 gnd
port 514 nsew
rlabel metal2 s 30192 27097 30192 27097 4 gnd
port 514 nsew
rlabel metal2 s 30960 26070 30960 26070 4 gnd
port 514 nsew
rlabel metal2 s 30192 26070 30192 26070 4 gnd
port 514 nsew
rlabel metal2 s 31440 28203 31440 28203 4 gnd
port 514 nsew
rlabel metal2 s 30960 28440 30960 28440 4 gnd
port 514 nsew
rlabel metal2 s 31440 27413 31440 27413 4 gnd
port 514 nsew
rlabel metal2 s 30960 25517 30960 25517 4 gnd
port 514 nsew
rlabel metal2 s 30192 26623 30192 26623 4 gnd
port 514 nsew
rlabel metal2 s 30192 26307 30192 26307 4 gnd
port 514 nsew
rlabel metal2 s 31440 25833 31440 25833 4 gnd
port 514 nsew
rlabel metal2 s 32208 26623 32208 26623 4 gnd
port 514 nsew
rlabel metal2 s 32208 25833 32208 25833 4 gnd
port 514 nsew
rlabel metal2 s 30192 25833 30192 25833 4 gnd
port 514 nsew
rlabel metal2 s 32208 26070 32208 26070 4 gnd
port 514 nsew
rlabel metal2 s 30192 28440 30192 28440 4 gnd
port 514 nsew
rlabel metal2 s 30192 27413 30192 27413 4 gnd
port 514 nsew
rlabel metal2 s 32208 27097 32208 27097 4 gnd
port 514 nsew
rlabel metal2 s 30960 26307 30960 26307 4 gnd
port 514 nsew
rlabel metal2 s 32208 25517 32208 25517 4 gnd
port 514 nsew
rlabel metal2 s 30960 27887 30960 27887 4 gnd
port 514 nsew
rlabel metal2 s 30960 27650 30960 27650 4 gnd
port 514 nsew
rlabel metal2 s 30192 25517 30192 25517 4 gnd
port 514 nsew
rlabel metal2 s 32208 28440 32208 28440 4 gnd
port 514 nsew
rlabel metal2 s 32208 27887 32208 27887 4 gnd
port 514 nsew
rlabel metal2 s 31440 26860 31440 26860 4 gnd
port 514 nsew
rlabel metal2 s 31440 27097 31440 27097 4 gnd
port 514 nsew
rlabel metal2 s 32208 27413 32208 27413 4 gnd
port 514 nsew
rlabel metal2 s 30960 27097 30960 27097 4 gnd
port 514 nsew
rlabel metal2 s 32208 27650 32208 27650 4 gnd
port 514 nsew
rlabel metal2 s 34704 25517 34704 25517 4 gnd
port 514 nsew
rlabel metal2 s 34704 27887 34704 27887 4 gnd
port 514 nsew
rlabel metal2 s 32688 28203 32688 28203 4 gnd
port 514 nsew
rlabel metal2 s 32688 26623 32688 26623 4 gnd
port 514 nsew
rlabel metal2 s 34704 27650 34704 27650 4 gnd
port 514 nsew
rlabel metal2 s 34704 27413 34704 27413 4 gnd
port 514 nsew
rlabel metal2 s 32688 25833 32688 25833 4 gnd
port 514 nsew
rlabel metal2 s 32688 28440 32688 28440 4 gnd
port 514 nsew
rlabel metal2 s 33936 26623 33936 26623 4 gnd
port 514 nsew
rlabel metal2 s 32688 27097 32688 27097 4 gnd
port 514 nsew
rlabel metal2 s 33936 25833 33936 25833 4 gnd
port 514 nsew
rlabel metal2 s 33456 26070 33456 26070 4 gnd
port 514 nsew
rlabel metal2 s 33456 26307 33456 26307 4 gnd
port 514 nsew
rlabel metal2 s 33456 26623 33456 26623 4 gnd
port 514 nsew
rlabel metal2 s 34704 26307 34704 26307 4 gnd
port 514 nsew
rlabel metal2 s 34704 26070 34704 26070 4 gnd
port 514 nsew
rlabel metal2 s 33456 27097 33456 27097 4 gnd
port 514 nsew
rlabel metal2 s 34704 28440 34704 28440 4 gnd
port 514 nsew
rlabel metal2 s 33936 26070 33936 26070 4 gnd
port 514 nsew
rlabel metal2 s 33456 27887 33456 27887 4 gnd
port 514 nsew
rlabel metal2 s 32688 27413 32688 27413 4 gnd
port 514 nsew
rlabel metal2 s 34704 25833 34704 25833 4 gnd
port 514 nsew
rlabel metal2 s 33456 26860 33456 26860 4 gnd
port 514 nsew
rlabel metal2 s 33936 28440 33936 28440 4 gnd
port 514 nsew
rlabel metal2 s 33456 25517 33456 25517 4 gnd
port 514 nsew
rlabel metal2 s 32688 27650 32688 27650 4 gnd
port 514 nsew
rlabel metal2 s 34704 26623 34704 26623 4 gnd
port 514 nsew
rlabel metal2 s 33936 27650 33936 27650 4 gnd
port 514 nsew
rlabel metal2 s 33936 27887 33936 27887 4 gnd
port 514 nsew
rlabel metal2 s 32688 27887 32688 27887 4 gnd
port 514 nsew
rlabel metal2 s 32688 26070 32688 26070 4 gnd
port 514 nsew
rlabel metal2 s 34704 26860 34704 26860 4 gnd
port 514 nsew
rlabel metal2 s 33936 27413 33936 27413 4 gnd
port 514 nsew
rlabel metal2 s 33936 25517 33936 25517 4 gnd
port 514 nsew
rlabel metal2 s 33456 27650 33456 27650 4 gnd
port 514 nsew
rlabel metal2 s 34704 27097 34704 27097 4 gnd
port 514 nsew
rlabel metal2 s 32688 26307 32688 26307 4 gnd
port 514 nsew
rlabel metal2 s 33456 28440 33456 28440 4 gnd
port 514 nsew
rlabel metal2 s 33936 28203 33936 28203 4 gnd
port 514 nsew
rlabel metal2 s 33936 26307 33936 26307 4 gnd
port 514 nsew
rlabel metal2 s 33936 26860 33936 26860 4 gnd
port 514 nsew
rlabel metal2 s 34704 28203 34704 28203 4 gnd
port 514 nsew
rlabel metal2 s 32688 25517 32688 25517 4 gnd
port 514 nsew
rlabel metal2 s 33456 28203 33456 28203 4 gnd
port 514 nsew
rlabel metal2 s 33456 27413 33456 27413 4 gnd
port 514 nsew
rlabel metal2 s 33456 25833 33456 25833 4 gnd
port 514 nsew
rlabel metal2 s 32688 26860 32688 26860 4 gnd
port 514 nsew
rlabel metal2 s 33936 27097 33936 27097 4 gnd
port 514 nsew
rlabel metal2 s 37680 31600 37680 31600 4 gnd
port 514 nsew
rlabel metal2 s 38928 30020 38928 30020 4 gnd
port 514 nsew
rlabel metal2 s 38928 31047 38928 31047 4 gnd
port 514 nsew
rlabel metal2 s 38448 29783 38448 29783 4 gnd
port 514 nsew
rlabel metal2 s 38928 28993 38928 28993 4 gnd
port 514 nsew
rlabel metal2 s 37680 29230 37680 29230 4 gnd
port 514 nsew
rlabel metal2 s 39696 30020 39696 30020 4 gnd
port 514 nsew
rlabel metal2 s 38448 29230 38448 29230 4 gnd
port 514 nsew
rlabel metal2 s 38928 29467 38928 29467 4 gnd
port 514 nsew
rlabel metal2 s 38448 31363 38448 31363 4 gnd
port 514 nsew
rlabel metal2 s 38928 30573 38928 30573 4 gnd
port 514 nsew
rlabel metal2 s 39696 29230 39696 29230 4 gnd
port 514 nsew
rlabel metal2 s 38448 28993 38448 28993 4 gnd
port 514 nsew
rlabel metal2 s 37680 29783 37680 29783 4 gnd
port 514 nsew
rlabel metal2 s 39696 29467 39696 29467 4 gnd
port 514 nsew
rlabel metal2 s 37680 31363 37680 31363 4 gnd
port 514 nsew
rlabel metal2 s 38928 30257 38928 30257 4 gnd
port 514 nsew
rlabel metal2 s 37680 30573 37680 30573 4 gnd
port 514 nsew
rlabel metal2 s 37680 30020 37680 30020 4 gnd
port 514 nsew
rlabel metal2 s 38928 31363 38928 31363 4 gnd
port 514 nsew
rlabel metal2 s 38448 28677 38448 28677 4 gnd
port 514 nsew
rlabel metal2 s 38448 30020 38448 30020 4 gnd
port 514 nsew
rlabel metal2 s 38448 29467 38448 29467 4 gnd
port 514 nsew
rlabel metal2 s 37680 28993 37680 28993 4 gnd
port 514 nsew
rlabel metal2 s 38448 30573 38448 30573 4 gnd
port 514 nsew
rlabel metal2 s 39696 30573 39696 30573 4 gnd
port 514 nsew
rlabel metal2 s 38448 30810 38448 30810 4 gnd
port 514 nsew
rlabel metal2 s 38448 30257 38448 30257 4 gnd
port 514 nsew
rlabel metal2 s 38928 29783 38928 29783 4 gnd
port 514 nsew
rlabel metal2 s 39696 28677 39696 28677 4 gnd
port 514 nsew
rlabel metal2 s 37680 30810 37680 30810 4 gnd
port 514 nsew
rlabel metal2 s 37680 29467 37680 29467 4 gnd
port 514 nsew
rlabel metal2 s 38928 31600 38928 31600 4 gnd
port 514 nsew
rlabel metal2 s 37680 28677 37680 28677 4 gnd
port 514 nsew
rlabel metal2 s 38928 28677 38928 28677 4 gnd
port 514 nsew
rlabel metal2 s 38448 31047 38448 31047 4 gnd
port 514 nsew
rlabel metal2 s 37680 30257 37680 30257 4 gnd
port 514 nsew
rlabel metal2 s 37680 31047 37680 31047 4 gnd
port 514 nsew
rlabel metal2 s 39696 30257 39696 30257 4 gnd
port 514 nsew
rlabel metal2 s 39696 30810 39696 30810 4 gnd
port 514 nsew
rlabel metal2 s 39696 31363 39696 31363 4 gnd
port 514 nsew
rlabel metal2 s 38448 31600 38448 31600 4 gnd
port 514 nsew
rlabel metal2 s 39696 29783 39696 29783 4 gnd
port 514 nsew
rlabel metal2 s 38928 29230 38928 29230 4 gnd
port 514 nsew
rlabel metal2 s 38928 30810 38928 30810 4 gnd
port 514 nsew
rlabel metal2 s 39696 28993 39696 28993 4 gnd
port 514 nsew
rlabel metal2 s 39696 31047 39696 31047 4 gnd
port 514 nsew
rlabel metal2 s 39696 31600 39696 31600 4 gnd
port 514 nsew
rlabel metal2 s 36432 30810 36432 30810 4 gnd
port 514 nsew
rlabel metal2 s 35952 28993 35952 28993 4 gnd
port 514 nsew
rlabel metal2 s 37200 30573 37200 30573 4 gnd
port 514 nsew
rlabel metal2 s 35184 28993 35184 28993 4 gnd
port 514 nsew
rlabel metal2 s 35184 28677 35184 28677 4 gnd
port 514 nsew
rlabel metal2 s 36432 31363 36432 31363 4 gnd
port 514 nsew
rlabel metal2 s 36432 28677 36432 28677 4 gnd
port 514 nsew
rlabel metal2 s 37200 30257 37200 30257 4 gnd
port 514 nsew
rlabel metal2 s 35952 30020 35952 30020 4 gnd
port 514 nsew
rlabel metal2 s 37200 30020 37200 30020 4 gnd
port 514 nsew
rlabel metal2 s 36432 30257 36432 30257 4 gnd
port 514 nsew
rlabel metal2 s 36432 29467 36432 29467 4 gnd
port 514 nsew
rlabel metal2 s 35184 30573 35184 30573 4 gnd
port 514 nsew
rlabel metal2 s 35184 31363 35184 31363 4 gnd
port 514 nsew
rlabel metal2 s 36432 30573 36432 30573 4 gnd
port 514 nsew
rlabel metal2 s 35184 30020 35184 30020 4 gnd
port 514 nsew
rlabel metal2 s 37200 31047 37200 31047 4 gnd
port 514 nsew
rlabel metal2 s 35184 31600 35184 31600 4 gnd
port 514 nsew
rlabel metal2 s 35952 30810 35952 30810 4 gnd
port 514 nsew
rlabel metal2 s 36432 31600 36432 31600 4 gnd
port 514 nsew
rlabel metal2 s 35184 31047 35184 31047 4 gnd
port 514 nsew
rlabel metal2 s 35952 29783 35952 29783 4 gnd
port 514 nsew
rlabel metal2 s 36432 30020 36432 30020 4 gnd
port 514 nsew
rlabel metal2 s 35184 29230 35184 29230 4 gnd
port 514 nsew
rlabel metal2 s 35952 30257 35952 30257 4 gnd
port 514 nsew
rlabel metal2 s 36432 31047 36432 31047 4 gnd
port 514 nsew
rlabel metal2 s 35184 30810 35184 30810 4 gnd
port 514 nsew
rlabel metal2 s 35952 30573 35952 30573 4 gnd
port 514 nsew
rlabel metal2 s 35952 31600 35952 31600 4 gnd
port 514 nsew
rlabel metal2 s 35184 30257 35184 30257 4 gnd
port 514 nsew
rlabel metal2 s 35952 29230 35952 29230 4 gnd
port 514 nsew
rlabel metal2 s 37200 28677 37200 28677 4 gnd
port 514 nsew
rlabel metal2 s 37200 29230 37200 29230 4 gnd
port 514 nsew
rlabel metal2 s 37200 28993 37200 28993 4 gnd
port 514 nsew
rlabel metal2 s 37200 31600 37200 31600 4 gnd
port 514 nsew
rlabel metal2 s 35952 31363 35952 31363 4 gnd
port 514 nsew
rlabel metal2 s 35952 31047 35952 31047 4 gnd
port 514 nsew
rlabel metal2 s 37200 29783 37200 29783 4 gnd
port 514 nsew
rlabel metal2 s 35952 29467 35952 29467 4 gnd
port 514 nsew
rlabel metal2 s 35952 28677 35952 28677 4 gnd
port 514 nsew
rlabel metal2 s 37200 29467 37200 29467 4 gnd
port 514 nsew
rlabel metal2 s 35184 29467 35184 29467 4 gnd
port 514 nsew
rlabel metal2 s 36432 29230 36432 29230 4 gnd
port 514 nsew
rlabel metal2 s 36432 28993 36432 28993 4 gnd
port 514 nsew
rlabel metal2 s 37200 31363 37200 31363 4 gnd
port 514 nsew
rlabel metal2 s 37200 30810 37200 30810 4 gnd
port 514 nsew
rlabel metal2 s 36432 29783 36432 29783 4 gnd
port 514 nsew
rlabel metal2 s 35184 29783 35184 29783 4 gnd
port 514 nsew
rlabel metal2 s 37200 27413 37200 27413 4 gnd
port 514 nsew
rlabel metal2 s 36432 25517 36432 25517 4 gnd
port 514 nsew
rlabel metal2 s 35952 25517 35952 25517 4 gnd
port 514 nsew
rlabel metal2 s 35952 28440 35952 28440 4 gnd
port 514 nsew
rlabel metal2 s 35184 27650 35184 27650 4 gnd
port 514 nsew
rlabel metal2 s 36432 26860 36432 26860 4 gnd
port 514 nsew
rlabel metal2 s 36432 26307 36432 26307 4 gnd
port 514 nsew
rlabel metal2 s 35184 26307 35184 26307 4 gnd
port 514 nsew
rlabel metal2 s 35952 27887 35952 27887 4 gnd
port 514 nsew
rlabel metal2 s 35952 26860 35952 26860 4 gnd
port 514 nsew
rlabel metal2 s 36432 27097 36432 27097 4 gnd
port 514 nsew
rlabel metal2 s 35952 26623 35952 26623 4 gnd
port 514 nsew
rlabel metal2 s 35952 25833 35952 25833 4 gnd
port 514 nsew
rlabel metal2 s 35184 28440 35184 28440 4 gnd
port 514 nsew
rlabel metal2 s 35184 26070 35184 26070 4 gnd
port 514 nsew
rlabel metal2 s 35184 25833 35184 25833 4 gnd
port 514 nsew
rlabel metal2 s 36432 27413 36432 27413 4 gnd
port 514 nsew
rlabel metal2 s 37200 26860 37200 26860 4 gnd
port 514 nsew
rlabel metal2 s 35952 27650 35952 27650 4 gnd
port 514 nsew
rlabel metal2 s 35184 26860 35184 26860 4 gnd
port 514 nsew
rlabel metal2 s 36432 28203 36432 28203 4 gnd
port 514 nsew
rlabel metal2 s 35184 27413 35184 27413 4 gnd
port 514 nsew
rlabel metal2 s 35952 27097 35952 27097 4 gnd
port 514 nsew
rlabel metal2 s 35184 28203 35184 28203 4 gnd
port 514 nsew
rlabel metal2 s 35184 26623 35184 26623 4 gnd
port 514 nsew
rlabel metal2 s 36432 26623 36432 26623 4 gnd
port 514 nsew
rlabel metal2 s 37200 27097 37200 27097 4 gnd
port 514 nsew
rlabel metal2 s 36432 27650 36432 27650 4 gnd
port 514 nsew
rlabel metal2 s 37200 28440 37200 28440 4 gnd
port 514 nsew
rlabel metal2 s 37200 26307 37200 26307 4 gnd
port 514 nsew
rlabel metal2 s 35952 27413 35952 27413 4 gnd
port 514 nsew
rlabel metal2 s 35184 27887 35184 27887 4 gnd
port 514 nsew
rlabel metal2 s 35952 28203 35952 28203 4 gnd
port 514 nsew
rlabel metal2 s 35952 26070 35952 26070 4 gnd
port 514 nsew
rlabel metal2 s 36432 28440 36432 28440 4 gnd
port 514 nsew
rlabel metal2 s 36432 27887 36432 27887 4 gnd
port 514 nsew
rlabel metal2 s 36432 26070 36432 26070 4 gnd
port 514 nsew
rlabel metal2 s 36432 25833 36432 25833 4 gnd
port 514 nsew
rlabel metal2 s 35184 27097 35184 27097 4 gnd
port 514 nsew
rlabel metal2 s 37200 25833 37200 25833 4 gnd
port 514 nsew
rlabel metal2 s 37200 27650 37200 27650 4 gnd
port 514 nsew
rlabel metal2 s 37200 26623 37200 26623 4 gnd
port 514 nsew
rlabel metal2 s 35184 25517 35184 25517 4 gnd
port 514 nsew
rlabel metal2 s 37200 26070 37200 26070 4 gnd
port 514 nsew
rlabel metal2 s 37200 28203 37200 28203 4 gnd
port 514 nsew
rlabel metal2 s 35952 26307 35952 26307 4 gnd
port 514 nsew
rlabel metal2 s 37200 25517 37200 25517 4 gnd
port 514 nsew
rlabel metal2 s 37200 27887 37200 27887 4 gnd
port 514 nsew
rlabel metal2 s 38928 28203 38928 28203 4 gnd
port 514 nsew
rlabel metal2 s 39696 25833 39696 25833 4 gnd
port 514 nsew
rlabel metal2 s 37680 26070 37680 26070 4 gnd
port 514 nsew
rlabel metal2 s 38928 26860 38928 26860 4 gnd
port 514 nsew
rlabel metal2 s 39696 26860 39696 26860 4 gnd
port 514 nsew
rlabel metal2 s 38928 26070 38928 26070 4 gnd
port 514 nsew
rlabel metal2 s 38928 26623 38928 26623 4 gnd
port 514 nsew
rlabel metal2 s 38448 26307 38448 26307 4 gnd
port 514 nsew
rlabel metal2 s 39696 28203 39696 28203 4 gnd
port 514 nsew
rlabel metal2 s 38928 25833 38928 25833 4 gnd
port 514 nsew
rlabel metal2 s 37680 26307 37680 26307 4 gnd
port 514 nsew
rlabel metal2 s 37680 25833 37680 25833 4 gnd
port 514 nsew
rlabel metal2 s 39696 27413 39696 27413 4 gnd
port 514 nsew
rlabel metal2 s 37680 27887 37680 27887 4 gnd
port 514 nsew
rlabel metal2 s 38448 28203 38448 28203 4 gnd
port 514 nsew
rlabel metal2 s 38448 25833 38448 25833 4 gnd
port 514 nsew
rlabel metal2 s 39696 27650 39696 27650 4 gnd
port 514 nsew
rlabel metal2 s 37680 25517 37680 25517 4 gnd
port 514 nsew
rlabel metal2 s 37680 26623 37680 26623 4 gnd
port 514 nsew
rlabel metal2 s 37680 26860 37680 26860 4 gnd
port 514 nsew
rlabel metal2 s 38928 28440 38928 28440 4 gnd
port 514 nsew
rlabel metal2 s 38448 28440 38448 28440 4 gnd
port 514 nsew
rlabel metal2 s 37680 28203 37680 28203 4 gnd
port 514 nsew
rlabel metal2 s 38928 27650 38928 27650 4 gnd
port 514 nsew
rlabel metal2 s 38448 26070 38448 26070 4 gnd
port 514 nsew
rlabel metal2 s 38448 26623 38448 26623 4 gnd
port 514 nsew
rlabel metal2 s 37680 27097 37680 27097 4 gnd
port 514 nsew
rlabel metal2 s 38448 26860 38448 26860 4 gnd
port 514 nsew
rlabel metal2 s 39696 26307 39696 26307 4 gnd
port 514 nsew
rlabel metal2 s 38928 25517 38928 25517 4 gnd
port 514 nsew
rlabel metal2 s 39696 27097 39696 27097 4 gnd
port 514 nsew
rlabel metal2 s 38448 27887 38448 27887 4 gnd
port 514 nsew
rlabel metal2 s 38928 27097 38928 27097 4 gnd
port 514 nsew
rlabel metal2 s 38448 27650 38448 27650 4 gnd
port 514 nsew
rlabel metal2 s 37680 27650 37680 27650 4 gnd
port 514 nsew
rlabel metal2 s 37680 28440 37680 28440 4 gnd
port 514 nsew
rlabel metal2 s 39696 26070 39696 26070 4 gnd
port 514 nsew
rlabel metal2 s 39696 28440 39696 28440 4 gnd
port 514 nsew
rlabel metal2 s 38448 27413 38448 27413 4 gnd
port 514 nsew
rlabel metal2 s 39696 27887 39696 27887 4 gnd
port 514 nsew
rlabel metal2 s 38928 27413 38928 27413 4 gnd
port 514 nsew
rlabel metal2 s 39696 26623 39696 26623 4 gnd
port 514 nsew
rlabel metal2 s 39696 25517 39696 25517 4 gnd
port 514 nsew
rlabel metal2 s 38928 26307 38928 26307 4 gnd
port 514 nsew
rlabel metal2 s 38928 27887 38928 27887 4 gnd
port 514 nsew
rlabel metal2 s 38448 25517 38448 25517 4 gnd
port 514 nsew
rlabel metal2 s 37680 27413 37680 27413 4 gnd
port 514 nsew
rlabel metal2 s 38448 27097 38448 27097 4 gnd
port 514 nsew
rlabel metal2 s 18480 49533 18480 49533 4 gnd
port 514 nsew
rlabel metal2 s 18480 50007 18480 50007 4 gnd
port 514 nsew
rlabel metal2 s 18480 49770 18480 49770 4 gnd
port 514 nsew
rlabel metal2 s 19728 50007 19728 50007 4 gnd
port 514 nsew
rlabel metal2 s 17712 50560 17712 50560 4 gnd
port 514 nsew
rlabel metal2 s 18480 47637 18480 47637 4 gnd
port 514 nsew
rlabel metal2 s 19968 49643 19968 49643 4 wl1_125
port 508 nsew
rlabel metal2 s 17712 48980 17712 48980 4 gnd
port 514 nsew
rlabel metal2 s 19728 50323 19728 50323 4 gnd
port 514 nsew
rlabel metal2 s 17712 47637 17712 47637 4 gnd
port 514 nsew
rlabel metal2 s 18960 48980 18960 48980 4 gnd
port 514 nsew
rlabel metal2 s 17712 49770 17712 49770 4 gnd
port 514 nsew
rlabel metal2 s 19968 50433 19968 50433 4 wl1_127
port 512 nsew
rlabel metal2 s 19968 49423 19968 49423 4 wl0_125
port 507 nsew
rlabel metal2 s 19728 49533 19728 49533 4 gnd
port 514 nsew
rlabel metal2 s 18960 48743 18960 48743 4 gnd
port 514 nsew
rlabel metal2 s 19728 47637 19728 47637 4 gnd
port 514 nsew
rlabel metal2 s 17712 48743 17712 48743 4 gnd
port 514 nsew
rlabel metal2 s 18480 48743 18480 48743 4 gnd
port 514 nsew
rlabel metal2 s 19728 48427 19728 48427 4 gnd
port 514 nsew
rlabel metal2 s 17712 48190 17712 48190 4 gnd
port 514 nsew
rlabel metal2 s 19728 48743 19728 48743 4 gnd
port 514 nsew
rlabel metal2 s 18480 48427 18480 48427 4 gnd
port 514 nsew
rlabel metal2 s 18960 49217 18960 49217 4 gnd
port 514 nsew
rlabel metal2 s 19728 48190 19728 48190 4 gnd
port 514 nsew
rlabel metal2 s 17712 50007 17712 50007 4 gnd
port 514 nsew
rlabel metal2 s 19728 49217 19728 49217 4 gnd
port 514 nsew
rlabel metal2 s 18480 49217 18480 49217 4 gnd
port 514 nsew
rlabel metal2 s 18960 47953 18960 47953 4 gnd
port 514 nsew
rlabel metal2 s 18960 48190 18960 48190 4 gnd
port 514 nsew
rlabel metal2 s 19968 47747 19968 47747 4 wl0_120
port 497 nsew
rlabel metal2 s 18480 48980 18480 48980 4 gnd
port 514 nsew
rlabel metal2 s 17712 50323 17712 50323 4 gnd
port 514 nsew
rlabel metal2 s 18960 50007 18960 50007 4 gnd
port 514 nsew
rlabel metal2 s 18960 49533 18960 49533 4 gnd
port 514 nsew
rlabel metal2 s 19728 50560 19728 50560 4 gnd
port 514 nsew
rlabel metal2 s 18480 48190 18480 48190 4 gnd
port 514 nsew
rlabel metal2 s 19728 49770 19728 49770 4 gnd
port 514 nsew
rlabel metal2 s 17712 48427 17712 48427 4 gnd
port 514 nsew
rlabel metal2 s 18960 50560 18960 50560 4 gnd
port 514 nsew
rlabel metal2 s 18960 48427 18960 48427 4 gnd
port 514 nsew
rlabel metal2 s 18960 49770 18960 49770 4 gnd
port 514 nsew
rlabel metal2 s 18480 47953 18480 47953 4 gnd
port 514 nsew
rlabel metal2 s 19728 48980 19728 48980 4 gnd
port 514 nsew
rlabel metal2 s 19968 50117 19968 50117 4 wl0_126
port 509 nsew
rlabel metal2 s 18960 47637 18960 47637 4 gnd
port 514 nsew
rlabel metal2 s 18960 50323 18960 50323 4 gnd
port 514 nsew
rlabel metal2 s 17712 47953 17712 47953 4 gnd
port 514 nsew
rlabel metal2 s 17712 49217 17712 49217 4 gnd
port 514 nsew
rlabel metal2 s 19728 47953 19728 47953 4 gnd
port 514 nsew
rlabel metal2 s 18480 50323 18480 50323 4 gnd
port 514 nsew
rlabel metal2 s 17712 49533 17712 49533 4 gnd
port 514 nsew
rlabel metal2 s 18480 50560 18480 50560 4 gnd
port 514 nsew
rlabel metal2 s 19968 50213 19968 50213 4 wl0_127
port 511 nsew
rlabel metal2 s 19968 49897 19968 49897 4 wl1_126
port 510 nsew
rlabel metal2 s 19968 48633 19968 48633 4 wl0_123
port 503 nsew
rlabel metal2 s 19968 48537 19968 48537 4 wl0_122
port 501 nsew
rlabel metal2 s 19968 48853 19968 48853 4 wl1_123
port 504 nsew
rlabel metal2 s 19968 49107 19968 49107 4 wl1_124
port 506 nsew
rlabel metal2 s 19968 47843 19968 47843 4 wl0_121
port 499 nsew
rlabel metal2 s 19968 49327 19968 49327 4 wl0_124
port 505 nsew
rlabel metal2 s 19968 48063 19968 48063 4 wl1_121
port 500 nsew
rlabel metal2 s 19968 48317 19968 48317 4 wl1_122
port 502 nsew
rlabel metal2 s 19968 47527 19968 47527 4 wl1_120
port 498 nsew
rlabel metal2 s 17232 48190 17232 48190 4 gnd
port 514 nsew
rlabel metal2 s 17232 50323 17232 50323 4 gnd
port 514 nsew
rlabel metal2 s 15216 50323 15216 50323 4 gnd
port 514 nsew
rlabel metal2 s 17232 49217 17232 49217 4 gnd
port 514 nsew
rlabel metal2 s 15216 49217 15216 49217 4 gnd
port 514 nsew
rlabel metal2 s 15984 50560 15984 50560 4 gnd
port 514 nsew
rlabel metal2 s 17232 50007 17232 50007 4 gnd
port 514 nsew
rlabel metal2 s 15984 49217 15984 49217 4 gnd
port 514 nsew
rlabel metal2 s 15216 47953 15216 47953 4 gnd
port 514 nsew
rlabel metal2 s 15216 48190 15216 48190 4 gnd
port 514 nsew
rlabel metal2 s 15984 48743 15984 48743 4 gnd
port 514 nsew
rlabel metal2 s 15984 48427 15984 48427 4 gnd
port 514 nsew
rlabel metal2 s 15984 50007 15984 50007 4 gnd
port 514 nsew
rlabel metal2 s 16464 48743 16464 48743 4 gnd
port 514 nsew
rlabel metal2 s 17232 48980 17232 48980 4 gnd
port 514 nsew
rlabel metal2 s 15984 49533 15984 49533 4 gnd
port 514 nsew
rlabel metal2 s 16464 48980 16464 48980 4 gnd
port 514 nsew
rlabel metal2 s 17232 48427 17232 48427 4 gnd
port 514 nsew
rlabel metal2 s 16464 50560 16464 50560 4 gnd
port 514 nsew
rlabel metal2 s 17232 49770 17232 49770 4 gnd
port 514 nsew
rlabel metal2 s 17232 49533 17232 49533 4 gnd
port 514 nsew
rlabel metal2 s 17232 47637 17232 47637 4 gnd
port 514 nsew
rlabel metal2 s 16464 48427 16464 48427 4 gnd
port 514 nsew
rlabel metal2 s 15216 48980 15216 48980 4 gnd
port 514 nsew
rlabel metal2 s 16464 47637 16464 47637 4 gnd
port 514 nsew
rlabel metal2 s 15216 50007 15216 50007 4 gnd
port 514 nsew
rlabel metal2 s 15984 49770 15984 49770 4 gnd
port 514 nsew
rlabel metal2 s 15216 50560 15216 50560 4 gnd
port 514 nsew
rlabel metal2 s 16464 50007 16464 50007 4 gnd
port 514 nsew
rlabel metal2 s 15216 48427 15216 48427 4 gnd
port 514 nsew
rlabel metal2 s 15984 50323 15984 50323 4 gnd
port 514 nsew
rlabel metal2 s 15984 47953 15984 47953 4 gnd
port 514 nsew
rlabel metal2 s 15984 48190 15984 48190 4 gnd
port 514 nsew
rlabel metal2 s 17232 50560 17232 50560 4 gnd
port 514 nsew
rlabel metal2 s 17232 48743 17232 48743 4 gnd
port 514 nsew
rlabel metal2 s 15984 48980 15984 48980 4 gnd
port 514 nsew
rlabel metal2 s 15216 49533 15216 49533 4 gnd
port 514 nsew
rlabel metal2 s 15216 49770 15216 49770 4 gnd
port 514 nsew
rlabel metal2 s 16464 50323 16464 50323 4 gnd
port 514 nsew
rlabel metal2 s 15984 47637 15984 47637 4 gnd
port 514 nsew
rlabel metal2 s 17232 47953 17232 47953 4 gnd
port 514 nsew
rlabel metal2 s 16464 47953 16464 47953 4 gnd
port 514 nsew
rlabel metal2 s 16464 49217 16464 49217 4 gnd
port 514 nsew
rlabel metal2 s 16464 49770 16464 49770 4 gnd
port 514 nsew
rlabel metal2 s 16464 48190 16464 48190 4 gnd
port 514 nsew
rlabel metal2 s 15216 48743 15216 48743 4 gnd
port 514 nsew
rlabel metal2 s 16464 49533 16464 49533 4 gnd
port 514 nsew
rlabel metal2 s 15216 47637 15216 47637 4 gnd
port 514 nsew
rlabel metal2 s 15216 45030 15216 45030 4 gnd
port 514 nsew
rlabel metal2 s 16464 46847 16464 46847 4 gnd
port 514 nsew
rlabel metal2 s 15216 45267 15216 45267 4 gnd
port 514 nsew
rlabel metal2 s 17232 46057 17232 46057 4 gnd
port 514 nsew
rlabel metal2 s 17232 47163 17232 47163 4 gnd
port 514 nsew
rlabel metal2 s 15216 46847 15216 46847 4 gnd
port 514 nsew
rlabel metal2 s 16464 46373 16464 46373 4 gnd
port 514 nsew
rlabel metal2 s 15984 47163 15984 47163 4 gnd
port 514 nsew
rlabel metal2 s 15216 46373 15216 46373 4 gnd
port 514 nsew
rlabel metal2 s 17232 47400 17232 47400 4 gnd
port 514 nsew
rlabel metal2 s 15984 46373 15984 46373 4 gnd
port 514 nsew
rlabel metal2 s 16464 45583 16464 45583 4 gnd
port 514 nsew
rlabel metal2 s 16464 44793 16464 44793 4 gnd
port 514 nsew
rlabel metal2 s 15216 45583 15216 45583 4 gnd
port 514 nsew
rlabel metal2 s 15216 44793 15216 44793 4 gnd
port 514 nsew
rlabel metal2 s 15216 47163 15216 47163 4 gnd
port 514 nsew
rlabel metal2 s 17232 44793 17232 44793 4 gnd
port 514 nsew
rlabel metal2 s 15984 46057 15984 46057 4 gnd
port 514 nsew
rlabel metal2 s 16464 47400 16464 47400 4 gnd
port 514 nsew
rlabel metal2 s 15984 46847 15984 46847 4 gnd
port 514 nsew
rlabel metal2 s 15216 47400 15216 47400 4 gnd
port 514 nsew
rlabel metal2 s 17232 46373 17232 46373 4 gnd
port 514 nsew
rlabel metal2 s 16464 44477 16464 44477 4 gnd
port 514 nsew
rlabel metal2 s 17232 45583 17232 45583 4 gnd
port 514 nsew
rlabel metal2 s 17232 45030 17232 45030 4 gnd
port 514 nsew
rlabel metal2 s 15216 46610 15216 46610 4 gnd
port 514 nsew
rlabel metal2 s 16464 45030 16464 45030 4 gnd
port 514 nsew
rlabel metal2 s 15216 45820 15216 45820 4 gnd
port 514 nsew
rlabel metal2 s 15216 46057 15216 46057 4 gnd
port 514 nsew
rlabel metal2 s 15984 44477 15984 44477 4 gnd
port 514 nsew
rlabel metal2 s 15216 44477 15216 44477 4 gnd
port 514 nsew
rlabel metal2 s 17232 46610 17232 46610 4 gnd
port 514 nsew
rlabel metal2 s 17232 44477 17232 44477 4 gnd
port 514 nsew
rlabel metal2 s 15984 45030 15984 45030 4 gnd
port 514 nsew
rlabel metal2 s 16464 47163 16464 47163 4 gnd
port 514 nsew
rlabel metal2 s 16464 45820 16464 45820 4 gnd
port 514 nsew
rlabel metal2 s 15984 44793 15984 44793 4 gnd
port 514 nsew
rlabel metal2 s 16464 46610 16464 46610 4 gnd
port 514 nsew
rlabel metal2 s 17232 45267 17232 45267 4 gnd
port 514 nsew
rlabel metal2 s 15984 46610 15984 46610 4 gnd
port 514 nsew
rlabel metal2 s 15984 45820 15984 45820 4 gnd
port 514 nsew
rlabel metal2 s 17232 46847 17232 46847 4 gnd
port 514 nsew
rlabel metal2 s 16464 46057 16464 46057 4 gnd
port 514 nsew
rlabel metal2 s 15984 45267 15984 45267 4 gnd
port 514 nsew
rlabel metal2 s 16464 45267 16464 45267 4 gnd
port 514 nsew
rlabel metal2 s 15984 47400 15984 47400 4 gnd
port 514 nsew
rlabel metal2 s 15984 45583 15984 45583 4 gnd
port 514 nsew
rlabel metal2 s 17232 45820 17232 45820 4 gnd
port 514 nsew
rlabel metal2 s 18960 45267 18960 45267 4 gnd
port 514 nsew
rlabel metal2 s 17712 47400 17712 47400 4 gnd
port 514 nsew
rlabel metal2 s 19728 44477 19728 44477 4 gnd
port 514 nsew
rlabel metal2 s 18960 44477 18960 44477 4 gnd
port 514 nsew
rlabel metal2 s 18480 45583 18480 45583 4 gnd
port 514 nsew
rlabel metal2 s 17712 47163 17712 47163 4 gnd
port 514 nsew
rlabel metal2 s 17712 45820 17712 45820 4 gnd
port 514 nsew
rlabel metal2 s 18480 47163 18480 47163 4 gnd
port 514 nsew
rlabel metal2 s 18480 45820 18480 45820 4 gnd
port 514 nsew
rlabel metal2 s 19728 46057 19728 46057 4 gnd
port 514 nsew
rlabel metal2 s 18480 45267 18480 45267 4 gnd
port 514 nsew
rlabel metal2 s 17712 45030 17712 45030 4 gnd
port 514 nsew
rlabel metal2 s 19728 46373 19728 46373 4 gnd
port 514 nsew
rlabel metal2 s 18960 46373 18960 46373 4 gnd
port 514 nsew
rlabel metal2 s 18480 44477 18480 44477 4 gnd
port 514 nsew
rlabel metal2 s 18480 46847 18480 46847 4 gnd
port 514 nsew
rlabel metal2 s 18960 44793 18960 44793 4 gnd
port 514 nsew
rlabel metal2 s 17712 46057 17712 46057 4 gnd
port 514 nsew
rlabel metal2 s 19728 45820 19728 45820 4 gnd
port 514 nsew
rlabel metal2 s 17712 45267 17712 45267 4 gnd
port 514 nsew
rlabel metal2 s 19968 44903 19968 44903 4 wl1_113
port 484 nsew
rlabel metal2 s 19968 46263 19968 46263 4 wl0_117
port 491 nsew
rlabel metal2 s 18960 47400 18960 47400 4 gnd
port 514 nsew
rlabel metal2 s 18960 46610 18960 46610 4 gnd
port 514 nsew
rlabel metal2 s 18480 46057 18480 46057 4 gnd
port 514 nsew
rlabel metal2 s 18480 46373 18480 46373 4 gnd
port 514 nsew
rlabel metal2 s 17712 46610 17712 46610 4 gnd
port 514 nsew
rlabel metal2 s 18960 46847 18960 46847 4 gnd
port 514 nsew
rlabel metal2 s 18960 47163 18960 47163 4 gnd
port 514 nsew
rlabel metal2 s 18480 47400 18480 47400 4 gnd
port 514 nsew
rlabel metal2 s 17712 45583 17712 45583 4 gnd
port 514 nsew
rlabel metal2 s 17712 44477 17712 44477 4 gnd
port 514 nsew
rlabel metal2 s 18960 45583 18960 45583 4 gnd
port 514 nsew
rlabel metal2 s 19728 45030 19728 45030 4 gnd
port 514 nsew
rlabel metal2 s 18960 45030 18960 45030 4 gnd
port 514 nsew
rlabel metal2 s 18480 45030 18480 45030 4 gnd
port 514 nsew
rlabel metal2 s 19728 46610 19728 46610 4 gnd
port 514 nsew
rlabel metal2 s 18960 46057 18960 46057 4 gnd
port 514 nsew
rlabel metal2 s 19728 47400 19728 47400 4 gnd
port 514 nsew
rlabel metal2 s 19728 47163 19728 47163 4 gnd
port 514 nsew
rlabel metal2 s 19728 45583 19728 45583 4 gnd
port 514 nsew
rlabel metal2 s 19968 46957 19968 46957 4 wl0_118
port 493 nsew
rlabel metal2 s 19968 46167 19968 46167 4 wl0_116
port 489 nsew
rlabel metal2 s 19968 44367 19968 44367 4 wl1_112
port 482 nsew
rlabel metal2 s 18480 44793 18480 44793 4 gnd
port 514 nsew
rlabel metal2 s 19728 46847 19728 46847 4 gnd
port 514 nsew
rlabel metal2 s 19728 45267 19728 45267 4 gnd
port 514 nsew
rlabel metal2 s 19968 47053 19968 47053 4 wl0_119
port 495 nsew
rlabel metal2 s 19968 47273 19968 47273 4 wl1_119
port 496 nsew
rlabel metal2 s 19968 44683 19968 44683 4 wl0_113
port 483 nsew
rlabel metal2 s 17712 46847 17712 46847 4 gnd
port 514 nsew
rlabel metal2 s 19968 45947 19968 45947 4 wl1_116
port 490 nsew
rlabel metal2 s 17712 46373 17712 46373 4 gnd
port 514 nsew
rlabel metal2 s 17712 44793 17712 44793 4 gnd
port 514 nsew
rlabel metal2 s 19728 44793 19728 44793 4 gnd
port 514 nsew
rlabel metal2 s 19968 45473 19968 45473 4 wl0_115
port 487 nsew
rlabel metal2 s 19968 45157 19968 45157 4 wl1_114
port 486 nsew
rlabel metal2 s 19968 45377 19968 45377 4 wl0_114
port 485 nsew
rlabel metal2 s 18960 45820 18960 45820 4 gnd
port 514 nsew
rlabel metal2 s 19968 45693 19968 45693 4 wl1_115
port 488 nsew
rlabel metal2 s 19968 46737 19968 46737 4 wl1_118
port 494 nsew
rlabel metal2 s 19968 46483 19968 46483 4 wl1_117
port 492 nsew
rlabel metal2 s 19968 44587 19968 44587 4 wl0_112
port 481 nsew
rlabel metal2 s 18480 46610 18480 46610 4 gnd
port 514 nsew
rlabel metal2 s 14736 49217 14736 49217 4 gnd
port 514 nsew
rlabel metal2 s 12720 48427 12720 48427 4 gnd
port 514 nsew
rlabel metal2 s 12720 50007 12720 50007 4 gnd
port 514 nsew
rlabel metal2 s 13488 48980 13488 48980 4 gnd
port 514 nsew
rlabel metal2 s 13968 50007 13968 50007 4 gnd
port 514 nsew
rlabel metal2 s 13968 49217 13968 49217 4 gnd
port 514 nsew
rlabel metal2 s 13488 49533 13488 49533 4 gnd
port 514 nsew
rlabel metal2 s 12720 49533 12720 49533 4 gnd
port 514 nsew
rlabel metal2 s 14736 49770 14736 49770 4 gnd
port 514 nsew
rlabel metal2 s 13488 49770 13488 49770 4 gnd
port 514 nsew
rlabel metal2 s 12720 47637 12720 47637 4 gnd
port 514 nsew
rlabel metal2 s 13488 47953 13488 47953 4 gnd
port 514 nsew
rlabel metal2 s 14736 50323 14736 50323 4 gnd
port 514 nsew
rlabel metal2 s 13968 50323 13968 50323 4 gnd
port 514 nsew
rlabel metal2 s 14736 47637 14736 47637 4 gnd
port 514 nsew
rlabel metal2 s 13488 50007 13488 50007 4 gnd
port 514 nsew
rlabel metal2 s 14736 50560 14736 50560 4 gnd
port 514 nsew
rlabel metal2 s 14736 48427 14736 48427 4 gnd
port 514 nsew
rlabel metal2 s 12720 50323 12720 50323 4 gnd
port 514 nsew
rlabel metal2 s 13488 50323 13488 50323 4 gnd
port 514 nsew
rlabel metal2 s 14736 49533 14736 49533 4 gnd
port 514 nsew
rlabel metal2 s 12720 49770 12720 49770 4 gnd
port 514 nsew
rlabel metal2 s 14736 47953 14736 47953 4 gnd
port 514 nsew
rlabel metal2 s 12720 48190 12720 48190 4 gnd
port 514 nsew
rlabel metal2 s 13488 48427 13488 48427 4 gnd
port 514 nsew
rlabel metal2 s 13968 48190 13968 48190 4 gnd
port 514 nsew
rlabel metal2 s 13488 49217 13488 49217 4 gnd
port 514 nsew
rlabel metal2 s 12720 48980 12720 48980 4 gnd
port 514 nsew
rlabel metal2 s 13968 48743 13968 48743 4 gnd
port 514 nsew
rlabel metal2 s 12720 50560 12720 50560 4 gnd
port 514 nsew
rlabel metal2 s 13488 48743 13488 48743 4 gnd
port 514 nsew
rlabel metal2 s 12720 49217 12720 49217 4 gnd
port 514 nsew
rlabel metal2 s 13488 48190 13488 48190 4 gnd
port 514 nsew
rlabel metal2 s 12720 48743 12720 48743 4 gnd
port 514 nsew
rlabel metal2 s 14736 48743 14736 48743 4 gnd
port 514 nsew
rlabel metal2 s 14736 48190 14736 48190 4 gnd
port 514 nsew
rlabel metal2 s 14736 48980 14736 48980 4 gnd
port 514 nsew
rlabel metal2 s 13968 50560 13968 50560 4 gnd
port 514 nsew
rlabel metal2 s 13968 48980 13968 48980 4 gnd
port 514 nsew
rlabel metal2 s 13968 49533 13968 49533 4 gnd
port 514 nsew
rlabel metal2 s 13968 47637 13968 47637 4 gnd
port 514 nsew
rlabel metal2 s 12720 47953 12720 47953 4 gnd
port 514 nsew
rlabel metal2 s 13968 47953 13968 47953 4 gnd
port 514 nsew
rlabel metal2 s 13488 50560 13488 50560 4 gnd
port 514 nsew
rlabel metal2 s 13488 47637 13488 47637 4 gnd
port 514 nsew
rlabel metal2 s 13968 49770 13968 49770 4 gnd
port 514 nsew
rlabel metal2 s 13968 48427 13968 48427 4 gnd
port 514 nsew
rlabel metal2 s 14736 50007 14736 50007 4 gnd
port 514 nsew
rlabel metal2 s 11472 50007 11472 50007 4 gnd
port 514 nsew
rlabel metal2 s 12240 49217 12240 49217 4 gnd
port 514 nsew
rlabel metal2 s 11472 50560 11472 50560 4 gnd
port 514 nsew
rlabel metal2 s 11472 48190 11472 48190 4 gnd
port 514 nsew
rlabel metal2 s 12240 47953 12240 47953 4 gnd
port 514 nsew
rlabel metal2 s 10992 49217 10992 49217 4 gnd
port 514 nsew
rlabel metal2 s 10992 50007 10992 50007 4 gnd
port 514 nsew
rlabel metal2 s 10992 47637 10992 47637 4 gnd
port 514 nsew
rlabel metal2 s 10992 49533 10992 49533 4 gnd
port 514 nsew
rlabel metal2 s 10224 49533 10224 49533 4 gnd
port 514 nsew
rlabel metal2 s 10224 47637 10224 47637 4 gnd
port 514 nsew
rlabel metal2 s 10224 48980 10224 48980 4 gnd
port 514 nsew
rlabel metal2 s 12240 48980 12240 48980 4 gnd
port 514 nsew
rlabel metal2 s 10224 47953 10224 47953 4 gnd
port 514 nsew
rlabel metal2 s 10224 50560 10224 50560 4 gnd
port 514 nsew
rlabel metal2 s 11472 50323 11472 50323 4 gnd
port 514 nsew
rlabel metal2 s 12240 48743 12240 48743 4 gnd
port 514 nsew
rlabel metal2 s 11472 48980 11472 48980 4 gnd
port 514 nsew
rlabel metal2 s 10992 50560 10992 50560 4 gnd
port 514 nsew
rlabel metal2 s 10224 49770 10224 49770 4 gnd
port 514 nsew
rlabel metal2 s 12240 50323 12240 50323 4 gnd
port 514 nsew
rlabel metal2 s 12240 47637 12240 47637 4 gnd
port 514 nsew
rlabel metal2 s 10992 50323 10992 50323 4 gnd
port 514 nsew
rlabel metal2 s 12240 49533 12240 49533 4 gnd
port 514 nsew
rlabel metal2 s 11472 49770 11472 49770 4 gnd
port 514 nsew
rlabel metal2 s 12240 50560 12240 50560 4 gnd
port 514 nsew
rlabel metal2 s 11472 47637 11472 47637 4 gnd
port 514 nsew
rlabel metal2 s 12240 48427 12240 48427 4 gnd
port 514 nsew
rlabel metal2 s 10224 50323 10224 50323 4 gnd
port 514 nsew
rlabel metal2 s 11472 49217 11472 49217 4 gnd
port 514 nsew
rlabel metal2 s 10992 48190 10992 48190 4 gnd
port 514 nsew
rlabel metal2 s 11472 48427 11472 48427 4 gnd
port 514 nsew
rlabel metal2 s 10992 48980 10992 48980 4 gnd
port 514 nsew
rlabel metal2 s 10992 47953 10992 47953 4 gnd
port 514 nsew
rlabel metal2 s 10224 48427 10224 48427 4 gnd
port 514 nsew
rlabel metal2 s 12240 48190 12240 48190 4 gnd
port 514 nsew
rlabel metal2 s 10224 48743 10224 48743 4 gnd
port 514 nsew
rlabel metal2 s 10992 48743 10992 48743 4 gnd
port 514 nsew
rlabel metal2 s 10992 48427 10992 48427 4 gnd
port 514 nsew
rlabel metal2 s 10224 48190 10224 48190 4 gnd
port 514 nsew
rlabel metal2 s 10992 49770 10992 49770 4 gnd
port 514 nsew
rlabel metal2 s 11472 48743 11472 48743 4 gnd
port 514 nsew
rlabel metal2 s 12240 50007 12240 50007 4 gnd
port 514 nsew
rlabel metal2 s 11472 47953 11472 47953 4 gnd
port 514 nsew
rlabel metal2 s 12240 49770 12240 49770 4 gnd
port 514 nsew
rlabel metal2 s 10224 49217 10224 49217 4 gnd
port 514 nsew
rlabel metal2 s 11472 49533 11472 49533 4 gnd
port 514 nsew
rlabel metal2 s 10224 50007 10224 50007 4 gnd
port 514 nsew
rlabel metal2 s 10224 46057 10224 46057 4 gnd
port 514 nsew
rlabel metal2 s 11472 45267 11472 45267 4 gnd
port 514 nsew
rlabel metal2 s 12240 44477 12240 44477 4 gnd
port 514 nsew
rlabel metal2 s 10992 45583 10992 45583 4 gnd
port 514 nsew
rlabel metal2 s 10224 47163 10224 47163 4 gnd
port 514 nsew
rlabel metal2 s 10992 46057 10992 46057 4 gnd
port 514 nsew
rlabel metal2 s 11472 45820 11472 45820 4 gnd
port 514 nsew
rlabel metal2 s 11472 46610 11472 46610 4 gnd
port 514 nsew
rlabel metal2 s 10992 45820 10992 45820 4 gnd
port 514 nsew
rlabel metal2 s 10224 44477 10224 44477 4 gnd
port 514 nsew
rlabel metal2 s 10224 46847 10224 46847 4 gnd
port 514 nsew
rlabel metal2 s 10224 45583 10224 45583 4 gnd
port 514 nsew
rlabel metal2 s 10224 45030 10224 45030 4 gnd
port 514 nsew
rlabel metal2 s 10224 44793 10224 44793 4 gnd
port 514 nsew
rlabel metal2 s 12240 46057 12240 46057 4 gnd
port 514 nsew
rlabel metal2 s 10224 45820 10224 45820 4 gnd
port 514 nsew
rlabel metal2 s 12240 46610 12240 46610 4 gnd
port 514 nsew
rlabel metal2 s 10224 45267 10224 45267 4 gnd
port 514 nsew
rlabel metal2 s 11472 47163 11472 47163 4 gnd
port 514 nsew
rlabel metal2 s 12240 47400 12240 47400 4 gnd
port 514 nsew
rlabel metal2 s 12240 45820 12240 45820 4 gnd
port 514 nsew
rlabel metal2 s 11472 46847 11472 46847 4 gnd
port 514 nsew
rlabel metal2 s 10224 46610 10224 46610 4 gnd
port 514 nsew
rlabel metal2 s 12240 46847 12240 46847 4 gnd
port 514 nsew
rlabel metal2 s 11472 45030 11472 45030 4 gnd
port 514 nsew
rlabel metal2 s 12240 45267 12240 45267 4 gnd
port 514 nsew
rlabel metal2 s 11472 45583 11472 45583 4 gnd
port 514 nsew
rlabel metal2 s 10992 44477 10992 44477 4 gnd
port 514 nsew
rlabel metal2 s 11472 46057 11472 46057 4 gnd
port 514 nsew
rlabel metal2 s 10992 45267 10992 45267 4 gnd
port 514 nsew
rlabel metal2 s 12240 44793 12240 44793 4 gnd
port 514 nsew
rlabel metal2 s 10224 47400 10224 47400 4 gnd
port 514 nsew
rlabel metal2 s 12240 47163 12240 47163 4 gnd
port 514 nsew
rlabel metal2 s 10992 45030 10992 45030 4 gnd
port 514 nsew
rlabel metal2 s 11472 44477 11472 44477 4 gnd
port 514 nsew
rlabel metal2 s 12240 45030 12240 45030 4 gnd
port 514 nsew
rlabel metal2 s 12240 46373 12240 46373 4 gnd
port 514 nsew
rlabel metal2 s 11472 44793 11472 44793 4 gnd
port 514 nsew
rlabel metal2 s 12240 45583 12240 45583 4 gnd
port 514 nsew
rlabel metal2 s 11472 46373 11472 46373 4 gnd
port 514 nsew
rlabel metal2 s 10992 46847 10992 46847 4 gnd
port 514 nsew
rlabel metal2 s 11472 47400 11472 47400 4 gnd
port 514 nsew
rlabel metal2 s 10992 47400 10992 47400 4 gnd
port 514 nsew
rlabel metal2 s 10992 44793 10992 44793 4 gnd
port 514 nsew
rlabel metal2 s 10992 46373 10992 46373 4 gnd
port 514 nsew
rlabel metal2 s 10992 46610 10992 46610 4 gnd
port 514 nsew
rlabel metal2 s 10992 47163 10992 47163 4 gnd
port 514 nsew
rlabel metal2 s 10224 46373 10224 46373 4 gnd
port 514 nsew
rlabel metal2 s 12720 45820 12720 45820 4 gnd
port 514 nsew
rlabel metal2 s 14736 47163 14736 47163 4 gnd
port 514 nsew
rlabel metal2 s 14736 46373 14736 46373 4 gnd
port 514 nsew
rlabel metal2 s 12720 44477 12720 44477 4 gnd
port 514 nsew
rlabel metal2 s 14736 44793 14736 44793 4 gnd
port 514 nsew
rlabel metal2 s 13968 47400 13968 47400 4 gnd
port 514 nsew
rlabel metal2 s 14736 45267 14736 45267 4 gnd
port 514 nsew
rlabel metal2 s 13968 46057 13968 46057 4 gnd
port 514 nsew
rlabel metal2 s 12720 47163 12720 47163 4 gnd
port 514 nsew
rlabel metal2 s 14736 47400 14736 47400 4 gnd
port 514 nsew
rlabel metal2 s 13488 46373 13488 46373 4 gnd
port 514 nsew
rlabel metal2 s 12720 46373 12720 46373 4 gnd
port 514 nsew
rlabel metal2 s 13968 45267 13968 45267 4 gnd
port 514 nsew
rlabel metal2 s 14736 44477 14736 44477 4 gnd
port 514 nsew
rlabel metal2 s 12720 44793 12720 44793 4 gnd
port 514 nsew
rlabel metal2 s 12720 45583 12720 45583 4 gnd
port 514 nsew
rlabel metal2 s 14736 46847 14736 46847 4 gnd
port 514 nsew
rlabel metal2 s 13488 46057 13488 46057 4 gnd
port 514 nsew
rlabel metal2 s 13488 47163 13488 47163 4 gnd
port 514 nsew
rlabel metal2 s 13968 46373 13968 46373 4 gnd
port 514 nsew
rlabel metal2 s 14736 45583 14736 45583 4 gnd
port 514 nsew
rlabel metal2 s 12720 46847 12720 46847 4 gnd
port 514 nsew
rlabel metal2 s 13968 45820 13968 45820 4 gnd
port 514 nsew
rlabel metal2 s 13488 45267 13488 45267 4 gnd
port 514 nsew
rlabel metal2 s 13968 45030 13968 45030 4 gnd
port 514 nsew
rlabel metal2 s 14736 45030 14736 45030 4 gnd
port 514 nsew
rlabel metal2 s 14736 45820 14736 45820 4 gnd
port 514 nsew
rlabel metal2 s 13968 44477 13968 44477 4 gnd
port 514 nsew
rlabel metal2 s 13968 46610 13968 46610 4 gnd
port 514 nsew
rlabel metal2 s 12720 45267 12720 45267 4 gnd
port 514 nsew
rlabel metal2 s 14736 46610 14736 46610 4 gnd
port 514 nsew
rlabel metal2 s 13488 47400 13488 47400 4 gnd
port 514 nsew
rlabel metal2 s 12720 46057 12720 46057 4 gnd
port 514 nsew
rlabel metal2 s 13488 45820 13488 45820 4 gnd
port 514 nsew
rlabel metal2 s 12720 45030 12720 45030 4 gnd
port 514 nsew
rlabel metal2 s 13968 45583 13968 45583 4 gnd
port 514 nsew
rlabel metal2 s 13488 44477 13488 44477 4 gnd
port 514 nsew
rlabel metal2 s 13488 45030 13488 45030 4 gnd
port 514 nsew
rlabel metal2 s 12720 47400 12720 47400 4 gnd
port 514 nsew
rlabel metal2 s 13968 46847 13968 46847 4 gnd
port 514 nsew
rlabel metal2 s 13488 46610 13488 46610 4 gnd
port 514 nsew
rlabel metal2 s 13488 45583 13488 45583 4 gnd
port 514 nsew
rlabel metal2 s 13968 44793 13968 44793 4 gnd
port 514 nsew
rlabel metal2 s 13968 47163 13968 47163 4 gnd
port 514 nsew
rlabel metal2 s 14736 46057 14736 46057 4 gnd
port 514 nsew
rlabel metal2 s 12720 46610 12720 46610 4 gnd
port 514 nsew
rlabel metal2 s 13488 44793 13488 44793 4 gnd
port 514 nsew
rlabel metal2 s 13488 46847 13488 46847 4 gnd
port 514 nsew
rlabel metal2 s 12720 43687 12720 43687 4 gnd
port 514 nsew
rlabel metal2 s 14736 41870 14736 41870 4 gnd
port 514 nsew
rlabel metal2 s 13968 41870 13968 41870 4 gnd
port 514 nsew
rlabel metal2 s 13968 41633 13968 41633 4 gnd
port 514 nsew
rlabel metal2 s 14736 42897 14736 42897 4 gnd
port 514 nsew
rlabel metal2 s 13968 44003 13968 44003 4 gnd
port 514 nsew
rlabel metal2 s 12720 41633 12720 41633 4 gnd
port 514 nsew
rlabel metal2 s 13968 42423 13968 42423 4 gnd
port 514 nsew
rlabel metal2 s 12720 42107 12720 42107 4 gnd
port 514 nsew
rlabel metal2 s 14736 43687 14736 43687 4 gnd
port 514 nsew
rlabel metal2 s 12720 42660 12720 42660 4 gnd
port 514 nsew
rlabel metal2 s 13488 44003 13488 44003 4 gnd
port 514 nsew
rlabel metal2 s 13968 43450 13968 43450 4 gnd
port 514 nsew
rlabel metal2 s 13488 42423 13488 42423 4 gnd
port 514 nsew
rlabel metal2 s 13968 44240 13968 44240 4 gnd
port 514 nsew
rlabel metal2 s 12720 41317 12720 41317 4 gnd
port 514 nsew
rlabel metal2 s 14736 42107 14736 42107 4 gnd
port 514 nsew
rlabel metal2 s 12720 43450 12720 43450 4 gnd
port 514 nsew
rlabel metal2 s 13488 44240 13488 44240 4 gnd
port 514 nsew
rlabel metal2 s 13488 42660 13488 42660 4 gnd
port 514 nsew
rlabel metal2 s 14736 43450 14736 43450 4 gnd
port 514 nsew
rlabel metal2 s 13488 42107 13488 42107 4 gnd
port 514 nsew
rlabel metal2 s 12720 44240 12720 44240 4 gnd
port 514 nsew
rlabel metal2 s 12720 43213 12720 43213 4 gnd
port 514 nsew
rlabel metal2 s 12720 42897 12720 42897 4 gnd
port 514 nsew
rlabel metal2 s 14736 42660 14736 42660 4 gnd
port 514 nsew
rlabel metal2 s 14736 41633 14736 41633 4 gnd
port 514 nsew
rlabel metal2 s 13968 41317 13968 41317 4 gnd
port 514 nsew
rlabel metal2 s 13968 43213 13968 43213 4 gnd
port 514 nsew
rlabel metal2 s 13968 42107 13968 42107 4 gnd
port 514 nsew
rlabel metal2 s 13488 43213 13488 43213 4 gnd
port 514 nsew
rlabel metal2 s 13488 43450 13488 43450 4 gnd
port 514 nsew
rlabel metal2 s 13968 42897 13968 42897 4 gnd
port 514 nsew
rlabel metal2 s 14736 42423 14736 42423 4 gnd
port 514 nsew
rlabel metal2 s 13488 41633 13488 41633 4 gnd
port 514 nsew
rlabel metal2 s 14736 44240 14736 44240 4 gnd
port 514 nsew
rlabel metal2 s 12720 44003 12720 44003 4 gnd
port 514 nsew
rlabel metal2 s 14736 41317 14736 41317 4 gnd
port 514 nsew
rlabel metal2 s 13968 42660 13968 42660 4 gnd
port 514 nsew
rlabel metal2 s 13488 42897 13488 42897 4 gnd
port 514 nsew
rlabel metal2 s 13488 43687 13488 43687 4 gnd
port 514 nsew
rlabel metal2 s 14736 43213 14736 43213 4 gnd
port 514 nsew
rlabel metal2 s 13488 41870 13488 41870 4 gnd
port 514 nsew
rlabel metal2 s 13488 41317 13488 41317 4 gnd
port 514 nsew
rlabel metal2 s 13968 43687 13968 43687 4 gnd
port 514 nsew
rlabel metal2 s 14736 44003 14736 44003 4 gnd
port 514 nsew
rlabel metal2 s 12720 41870 12720 41870 4 gnd
port 514 nsew
rlabel metal2 s 12720 42423 12720 42423 4 gnd
port 514 nsew
rlabel metal2 s 10224 41870 10224 41870 4 gnd
port 514 nsew
rlabel metal2 s 12240 44240 12240 44240 4 gnd
port 514 nsew
rlabel metal2 s 11472 42107 11472 42107 4 gnd
port 514 nsew
rlabel metal2 s 10224 43213 10224 43213 4 gnd
port 514 nsew
rlabel metal2 s 12240 41870 12240 41870 4 gnd
port 514 nsew
rlabel metal2 s 12240 41317 12240 41317 4 gnd
port 514 nsew
rlabel metal2 s 11472 42897 11472 42897 4 gnd
port 514 nsew
rlabel metal2 s 11472 44240 11472 44240 4 gnd
port 514 nsew
rlabel metal2 s 10224 42897 10224 42897 4 gnd
port 514 nsew
rlabel metal2 s 10992 41870 10992 41870 4 gnd
port 514 nsew
rlabel metal2 s 11472 43450 11472 43450 4 gnd
port 514 nsew
rlabel metal2 s 11472 43213 11472 43213 4 gnd
port 514 nsew
rlabel metal2 s 10224 41633 10224 41633 4 gnd
port 514 nsew
rlabel metal2 s 10992 41633 10992 41633 4 gnd
port 514 nsew
rlabel metal2 s 10992 43687 10992 43687 4 gnd
port 514 nsew
rlabel metal2 s 12240 43450 12240 43450 4 gnd
port 514 nsew
rlabel metal2 s 10224 44240 10224 44240 4 gnd
port 514 nsew
rlabel metal2 s 12240 42897 12240 42897 4 gnd
port 514 nsew
rlabel metal2 s 10992 44240 10992 44240 4 gnd
port 514 nsew
rlabel metal2 s 10224 42107 10224 42107 4 gnd
port 514 nsew
rlabel metal2 s 10224 42423 10224 42423 4 gnd
port 514 nsew
rlabel metal2 s 11472 42660 11472 42660 4 gnd
port 514 nsew
rlabel metal2 s 10992 42107 10992 42107 4 gnd
port 514 nsew
rlabel metal2 s 12240 44003 12240 44003 4 gnd
port 514 nsew
rlabel metal2 s 11472 44003 11472 44003 4 gnd
port 514 nsew
rlabel metal2 s 10224 43450 10224 43450 4 gnd
port 514 nsew
rlabel metal2 s 10224 44003 10224 44003 4 gnd
port 514 nsew
rlabel metal2 s 10992 43450 10992 43450 4 gnd
port 514 nsew
rlabel metal2 s 12240 43687 12240 43687 4 gnd
port 514 nsew
rlabel metal2 s 11472 43687 11472 43687 4 gnd
port 514 nsew
rlabel metal2 s 10992 42897 10992 42897 4 gnd
port 514 nsew
rlabel metal2 s 10992 42423 10992 42423 4 gnd
port 514 nsew
rlabel metal2 s 11472 41317 11472 41317 4 gnd
port 514 nsew
rlabel metal2 s 12240 42107 12240 42107 4 gnd
port 514 nsew
rlabel metal2 s 11472 41633 11472 41633 4 gnd
port 514 nsew
rlabel metal2 s 11472 41870 11472 41870 4 gnd
port 514 nsew
rlabel metal2 s 10224 43687 10224 43687 4 gnd
port 514 nsew
rlabel metal2 s 12240 42660 12240 42660 4 gnd
port 514 nsew
rlabel metal2 s 12240 41633 12240 41633 4 gnd
port 514 nsew
rlabel metal2 s 12240 42423 12240 42423 4 gnd
port 514 nsew
rlabel metal2 s 10992 43213 10992 43213 4 gnd
port 514 nsew
rlabel metal2 s 10992 42660 10992 42660 4 gnd
port 514 nsew
rlabel metal2 s 10224 41317 10224 41317 4 gnd
port 514 nsew
rlabel metal2 s 10992 41317 10992 41317 4 gnd
port 514 nsew
rlabel metal2 s 12240 43213 12240 43213 4 gnd
port 514 nsew
rlabel metal2 s 10224 42660 10224 42660 4 gnd
port 514 nsew
rlabel metal2 s 11472 42423 11472 42423 4 gnd
port 514 nsew
rlabel metal2 s 10992 44003 10992 44003 4 gnd
port 514 nsew
rlabel metal2 s 10992 41080 10992 41080 4 gnd
port 514 nsew
rlabel metal2 s 10224 39500 10224 39500 4 gnd
port 514 nsew
rlabel metal2 s 11472 40527 11472 40527 4 gnd
port 514 nsew
rlabel metal2 s 10224 40053 10224 40053 4 gnd
port 514 nsew
rlabel metal2 s 10224 38473 10224 38473 4 gnd
port 514 nsew
rlabel metal2 s 10992 39263 10992 39263 4 gnd
port 514 nsew
rlabel metal2 s 10992 39500 10992 39500 4 gnd
port 514 nsew
rlabel metal2 s 10224 38947 10224 38947 4 gnd
port 514 nsew
rlabel metal2 s 10992 40053 10992 40053 4 gnd
port 514 nsew
rlabel metal2 s 10992 38947 10992 38947 4 gnd
port 514 nsew
rlabel metal2 s 12240 38710 12240 38710 4 gnd
port 514 nsew
rlabel metal2 s 10992 38710 10992 38710 4 gnd
port 514 nsew
rlabel metal2 s 12240 41080 12240 41080 4 gnd
port 514 nsew
rlabel metal2 s 11472 40053 11472 40053 4 gnd
port 514 nsew
rlabel metal2 s 11472 38157 11472 38157 4 gnd
port 514 nsew
rlabel metal2 s 10992 40290 10992 40290 4 gnd
port 514 nsew
rlabel metal2 s 12240 40843 12240 40843 4 gnd
port 514 nsew
rlabel metal2 s 12240 38157 12240 38157 4 gnd
port 514 nsew
rlabel metal2 s 10224 39737 10224 39737 4 gnd
port 514 nsew
rlabel metal2 s 12240 40053 12240 40053 4 gnd
port 514 nsew
rlabel metal2 s 10224 38710 10224 38710 4 gnd
port 514 nsew
rlabel metal2 s 10992 40843 10992 40843 4 gnd
port 514 nsew
rlabel metal2 s 11472 39737 11472 39737 4 gnd
port 514 nsew
rlabel metal2 s 11472 39263 11472 39263 4 gnd
port 514 nsew
rlabel metal2 s 11472 40843 11472 40843 4 gnd
port 514 nsew
rlabel metal2 s 11472 38710 11472 38710 4 gnd
port 514 nsew
rlabel metal2 s 11472 40290 11472 40290 4 gnd
port 514 nsew
rlabel metal2 s 12240 39500 12240 39500 4 gnd
port 514 nsew
rlabel metal2 s 10224 40843 10224 40843 4 gnd
port 514 nsew
rlabel metal2 s 11472 38473 11472 38473 4 gnd
port 514 nsew
rlabel metal2 s 12240 39263 12240 39263 4 gnd
port 514 nsew
rlabel metal2 s 10224 39263 10224 39263 4 gnd
port 514 nsew
rlabel metal2 s 10224 38157 10224 38157 4 gnd
port 514 nsew
rlabel metal2 s 12240 39737 12240 39737 4 gnd
port 514 nsew
rlabel metal2 s 11472 38947 11472 38947 4 gnd
port 514 nsew
rlabel metal2 s 10224 40527 10224 40527 4 gnd
port 514 nsew
rlabel metal2 s 10992 39737 10992 39737 4 gnd
port 514 nsew
rlabel metal2 s 10224 40290 10224 40290 4 gnd
port 514 nsew
rlabel metal2 s 12240 38473 12240 38473 4 gnd
port 514 nsew
rlabel metal2 s 10992 38157 10992 38157 4 gnd
port 514 nsew
rlabel metal2 s 12240 38947 12240 38947 4 gnd
port 514 nsew
rlabel metal2 s 10992 38473 10992 38473 4 gnd
port 514 nsew
rlabel metal2 s 11472 41080 11472 41080 4 gnd
port 514 nsew
rlabel metal2 s 10224 41080 10224 41080 4 gnd
port 514 nsew
rlabel metal2 s 11472 39500 11472 39500 4 gnd
port 514 nsew
rlabel metal2 s 12240 40290 12240 40290 4 gnd
port 514 nsew
rlabel metal2 s 12240 40527 12240 40527 4 gnd
port 514 nsew
rlabel metal2 s 10992 40527 10992 40527 4 gnd
port 514 nsew
rlabel metal2 s 13488 40290 13488 40290 4 gnd
port 514 nsew
rlabel metal2 s 13488 38473 13488 38473 4 gnd
port 514 nsew
rlabel metal2 s 14736 39263 14736 39263 4 gnd
port 514 nsew
rlabel metal2 s 12720 40053 12720 40053 4 gnd
port 514 nsew
rlabel metal2 s 13488 39500 13488 39500 4 gnd
port 514 nsew
rlabel metal2 s 13968 40527 13968 40527 4 gnd
port 514 nsew
rlabel metal2 s 12720 38473 12720 38473 4 gnd
port 514 nsew
rlabel metal2 s 12720 38710 12720 38710 4 gnd
port 514 nsew
rlabel metal2 s 13488 40527 13488 40527 4 gnd
port 514 nsew
rlabel metal2 s 13968 38947 13968 38947 4 gnd
port 514 nsew
rlabel metal2 s 12720 39737 12720 39737 4 gnd
port 514 nsew
rlabel metal2 s 12720 40843 12720 40843 4 gnd
port 514 nsew
rlabel metal2 s 13968 39263 13968 39263 4 gnd
port 514 nsew
rlabel metal2 s 13968 38473 13968 38473 4 gnd
port 514 nsew
rlabel metal2 s 12720 39263 12720 39263 4 gnd
port 514 nsew
rlabel metal2 s 12720 39500 12720 39500 4 gnd
port 514 nsew
rlabel metal2 s 13968 38710 13968 38710 4 gnd
port 514 nsew
rlabel metal2 s 13488 39737 13488 39737 4 gnd
port 514 nsew
rlabel metal2 s 13488 38157 13488 38157 4 gnd
port 514 nsew
rlabel metal2 s 12720 38947 12720 38947 4 gnd
port 514 nsew
rlabel metal2 s 12720 38157 12720 38157 4 gnd
port 514 nsew
rlabel metal2 s 12720 41080 12720 41080 4 gnd
port 514 nsew
rlabel metal2 s 13968 39737 13968 39737 4 gnd
port 514 nsew
rlabel metal2 s 14736 38710 14736 38710 4 gnd
port 514 nsew
rlabel metal2 s 13488 38947 13488 38947 4 gnd
port 514 nsew
rlabel metal2 s 14736 38473 14736 38473 4 gnd
port 514 nsew
rlabel metal2 s 13968 40053 13968 40053 4 gnd
port 514 nsew
rlabel metal2 s 14736 39737 14736 39737 4 gnd
port 514 nsew
rlabel metal2 s 13968 41080 13968 41080 4 gnd
port 514 nsew
rlabel metal2 s 14736 40843 14736 40843 4 gnd
port 514 nsew
rlabel metal2 s 14736 40527 14736 40527 4 gnd
port 514 nsew
rlabel metal2 s 12720 40290 12720 40290 4 gnd
port 514 nsew
rlabel metal2 s 14736 40290 14736 40290 4 gnd
port 514 nsew
rlabel metal2 s 13488 40843 13488 40843 4 gnd
port 514 nsew
rlabel metal2 s 14736 38947 14736 38947 4 gnd
port 514 nsew
rlabel metal2 s 14736 41080 14736 41080 4 gnd
port 514 nsew
rlabel metal2 s 13488 39263 13488 39263 4 gnd
port 514 nsew
rlabel metal2 s 12720 40527 12720 40527 4 gnd
port 514 nsew
rlabel metal2 s 14736 39500 14736 39500 4 gnd
port 514 nsew
rlabel metal2 s 14736 40053 14736 40053 4 gnd
port 514 nsew
rlabel metal2 s 13968 40843 13968 40843 4 gnd
port 514 nsew
rlabel metal2 s 13488 40053 13488 40053 4 gnd
port 514 nsew
rlabel metal2 s 13968 38157 13968 38157 4 gnd
port 514 nsew
rlabel metal2 s 13488 38710 13488 38710 4 gnd
port 514 nsew
rlabel metal2 s 13968 40290 13968 40290 4 gnd
port 514 nsew
rlabel metal2 s 13968 39500 13968 39500 4 gnd
port 514 nsew
rlabel metal2 s 13488 41080 13488 41080 4 gnd
port 514 nsew
rlabel metal2 s 14736 38157 14736 38157 4 gnd
port 514 nsew
rlabel metal2 s 18960 44240 18960 44240 4 gnd
port 514 nsew
rlabel metal2 s 17712 42897 17712 42897 4 gnd
port 514 nsew
rlabel metal2 s 18960 41633 18960 41633 4 gnd
port 514 nsew
rlabel metal2 s 17712 41870 17712 41870 4 gnd
port 514 nsew
rlabel metal2 s 17712 42423 17712 42423 4 gnd
port 514 nsew
rlabel metal2 s 19728 42897 19728 42897 4 gnd
port 514 nsew
rlabel metal2 s 19728 42107 19728 42107 4 gnd
port 514 nsew
rlabel metal2 s 19728 43450 19728 43450 4 gnd
port 514 nsew
rlabel metal2 s 18960 42423 18960 42423 4 gnd
port 514 nsew
rlabel metal2 s 19728 41870 19728 41870 4 gnd
port 514 nsew
rlabel metal2 s 17712 42660 17712 42660 4 gnd
port 514 nsew
rlabel metal2 s 18480 42660 18480 42660 4 gnd
port 514 nsew
rlabel metal2 s 18480 42897 18480 42897 4 gnd
port 514 nsew
rlabel metal2 s 18480 43687 18480 43687 4 gnd
port 514 nsew
rlabel metal2 s 18960 42107 18960 42107 4 gnd
port 514 nsew
rlabel metal2 s 19728 41633 19728 41633 4 gnd
port 514 nsew
rlabel metal2 s 18960 44003 18960 44003 4 gnd
port 514 nsew
rlabel metal2 s 19728 41317 19728 41317 4 gnd
port 514 nsew
rlabel metal2 s 17712 42107 17712 42107 4 gnd
port 514 nsew
rlabel metal2 s 18480 44240 18480 44240 4 gnd
port 514 nsew
rlabel metal2 s 18480 42423 18480 42423 4 gnd
port 514 nsew
rlabel metal2 s 18480 42107 18480 42107 4 gnd
port 514 nsew
rlabel metal2 s 19728 42423 19728 42423 4 gnd
port 514 nsew
rlabel metal2 s 17712 41633 17712 41633 4 gnd
port 514 nsew
rlabel metal2 s 17712 41317 17712 41317 4 gnd
port 514 nsew
rlabel metal2 s 19728 42660 19728 42660 4 gnd
port 514 nsew
rlabel metal2 s 18960 43213 18960 43213 4 gnd
port 514 nsew
rlabel metal2 s 19728 44240 19728 44240 4 gnd
port 514 nsew
rlabel metal2 s 17712 43213 17712 43213 4 gnd
port 514 nsew
rlabel metal2 s 18960 43450 18960 43450 4 gnd
port 514 nsew
rlabel metal2 s 19728 43213 19728 43213 4 gnd
port 514 nsew
rlabel metal2 s 18480 41870 18480 41870 4 gnd
port 514 nsew
rlabel metal2 s 19728 44003 19728 44003 4 gnd
port 514 nsew
rlabel metal2 s 18960 42660 18960 42660 4 gnd
port 514 nsew
rlabel metal2 s 19728 43687 19728 43687 4 gnd
port 514 nsew
rlabel metal2 s 18480 41633 18480 41633 4 gnd
port 514 nsew
rlabel metal2 s 18480 44003 18480 44003 4 gnd
port 514 nsew
rlabel metal2 s 18960 41870 18960 41870 4 gnd
port 514 nsew
rlabel metal2 s 18960 43687 18960 43687 4 gnd
port 514 nsew
rlabel metal2 s 18960 41317 18960 41317 4 gnd
port 514 nsew
rlabel metal2 s 17712 43450 17712 43450 4 gnd
port 514 nsew
rlabel metal2 s 17712 44003 17712 44003 4 gnd
port 514 nsew
rlabel metal2 s 17712 44240 17712 44240 4 gnd
port 514 nsew
rlabel metal2 s 18960 42897 18960 42897 4 gnd
port 514 nsew
rlabel metal2 s 18480 43213 18480 43213 4 gnd
port 514 nsew
rlabel metal2 s 19968 43797 19968 43797 4 wl0_110
port 477 nsew
rlabel metal2 s 19968 43103 19968 43103 4 wl0_109
port 475 nsew
rlabel metal2 s 19968 43323 19968 43323 4 wl1_109
port 476 nsew
rlabel metal2 s 19968 41427 19968 41427 4 wl0_104
port 465 nsew
rlabel metal2 s 19968 43893 19968 43893 4 wl0_111
port 479 nsew
rlabel metal2 s 19968 42313 19968 42313 4 wl0_107
port 471 nsew
rlabel metal2 s 19968 42217 19968 42217 4 wl0_106
port 469 nsew
rlabel metal2 s 19968 42787 19968 42787 4 wl1_108
port 474 nsew
rlabel metal2 s 19968 41743 19968 41743 4 wl1_105
port 468 nsew
rlabel metal2 s 19968 43007 19968 43007 4 wl0_108
port 473 nsew
rlabel metal2 s 19968 44113 19968 44113 4 wl1_111
port 480 nsew
rlabel metal2 s 19968 42533 19968 42533 4 wl1_107
port 472 nsew
rlabel metal2 s 19968 41523 19968 41523 4 wl0_105
port 467 nsew
rlabel metal2 s 18480 43450 18480 43450 4 gnd
port 514 nsew
rlabel metal2 s 19968 43577 19968 43577 4 wl1_110
port 478 nsew
rlabel metal2 s 17712 43687 17712 43687 4 gnd
port 514 nsew
rlabel metal2 s 19968 41997 19968 41997 4 wl1_106
port 470 nsew
rlabel metal2 s 18480 41317 18480 41317 4 gnd
port 514 nsew
rlabel metal2 s 19968 41207 19968 41207 4 wl1_104
port 466 nsew
rlabel metal2 s 17232 41870 17232 41870 4 gnd
port 514 nsew
rlabel metal2 s 16464 42660 16464 42660 4 gnd
port 514 nsew
rlabel metal2 s 15216 41633 15216 41633 4 gnd
port 514 nsew
rlabel metal2 s 15984 43687 15984 43687 4 gnd
port 514 nsew
rlabel metal2 s 15216 44003 15216 44003 4 gnd
port 514 nsew
rlabel metal2 s 16464 43450 16464 43450 4 gnd
port 514 nsew
rlabel metal2 s 16464 41870 16464 41870 4 gnd
port 514 nsew
rlabel metal2 s 17232 44240 17232 44240 4 gnd
port 514 nsew
rlabel metal2 s 15216 42660 15216 42660 4 gnd
port 514 nsew
rlabel metal2 s 15984 41633 15984 41633 4 gnd
port 514 nsew
rlabel metal2 s 15984 42107 15984 42107 4 gnd
port 514 nsew
rlabel metal2 s 16464 42423 16464 42423 4 gnd
port 514 nsew
rlabel metal2 s 16464 42897 16464 42897 4 gnd
port 514 nsew
rlabel metal2 s 15984 41870 15984 41870 4 gnd
port 514 nsew
rlabel metal2 s 15984 43450 15984 43450 4 gnd
port 514 nsew
rlabel metal2 s 17232 41317 17232 41317 4 gnd
port 514 nsew
rlabel metal2 s 15984 44240 15984 44240 4 gnd
port 514 nsew
rlabel metal2 s 17232 44003 17232 44003 4 gnd
port 514 nsew
rlabel metal2 s 16464 43213 16464 43213 4 gnd
port 514 nsew
rlabel metal2 s 17232 41633 17232 41633 4 gnd
port 514 nsew
rlabel metal2 s 17232 42423 17232 42423 4 gnd
port 514 nsew
rlabel metal2 s 15984 42897 15984 42897 4 gnd
port 514 nsew
rlabel metal2 s 15216 41870 15216 41870 4 gnd
port 514 nsew
rlabel metal2 s 15984 41317 15984 41317 4 gnd
port 514 nsew
rlabel metal2 s 15216 42107 15216 42107 4 gnd
port 514 nsew
rlabel metal2 s 16464 44003 16464 44003 4 gnd
port 514 nsew
rlabel metal2 s 15216 42897 15216 42897 4 gnd
port 514 nsew
rlabel metal2 s 15216 43450 15216 43450 4 gnd
port 514 nsew
rlabel metal2 s 15984 44003 15984 44003 4 gnd
port 514 nsew
rlabel metal2 s 16464 41633 16464 41633 4 gnd
port 514 nsew
rlabel metal2 s 15984 42660 15984 42660 4 gnd
port 514 nsew
rlabel metal2 s 15216 42423 15216 42423 4 gnd
port 514 nsew
rlabel metal2 s 15984 42423 15984 42423 4 gnd
port 514 nsew
rlabel metal2 s 17232 42660 17232 42660 4 gnd
port 514 nsew
rlabel metal2 s 15216 44240 15216 44240 4 gnd
port 514 nsew
rlabel metal2 s 17232 42107 17232 42107 4 gnd
port 514 nsew
rlabel metal2 s 15216 43687 15216 43687 4 gnd
port 514 nsew
rlabel metal2 s 15216 41317 15216 41317 4 gnd
port 514 nsew
rlabel metal2 s 16464 41317 16464 41317 4 gnd
port 514 nsew
rlabel metal2 s 15216 43213 15216 43213 4 gnd
port 514 nsew
rlabel metal2 s 17232 43687 17232 43687 4 gnd
port 514 nsew
rlabel metal2 s 16464 44240 16464 44240 4 gnd
port 514 nsew
rlabel metal2 s 17232 43213 17232 43213 4 gnd
port 514 nsew
rlabel metal2 s 17232 43450 17232 43450 4 gnd
port 514 nsew
rlabel metal2 s 16464 43687 16464 43687 4 gnd
port 514 nsew
rlabel metal2 s 15984 43213 15984 43213 4 gnd
port 514 nsew
rlabel metal2 s 17232 42897 17232 42897 4 gnd
port 514 nsew
rlabel metal2 s 16464 42107 16464 42107 4 gnd
port 514 nsew
rlabel metal2 s 16464 39737 16464 39737 4 gnd
port 514 nsew
rlabel metal2 s 17232 40053 17232 40053 4 gnd
port 514 nsew
rlabel metal2 s 15216 38710 15216 38710 4 gnd
port 514 nsew
rlabel metal2 s 15216 38157 15216 38157 4 gnd
port 514 nsew
rlabel metal2 s 16464 40290 16464 40290 4 gnd
port 514 nsew
rlabel metal2 s 15216 39263 15216 39263 4 gnd
port 514 nsew
rlabel metal2 s 17232 40527 17232 40527 4 gnd
port 514 nsew
rlabel metal2 s 15216 39500 15216 39500 4 gnd
port 514 nsew
rlabel metal2 s 15216 39737 15216 39737 4 gnd
port 514 nsew
rlabel metal2 s 16464 39263 16464 39263 4 gnd
port 514 nsew
rlabel metal2 s 16464 39500 16464 39500 4 gnd
port 514 nsew
rlabel metal2 s 16464 38710 16464 38710 4 gnd
port 514 nsew
rlabel metal2 s 16464 38157 16464 38157 4 gnd
port 514 nsew
rlabel metal2 s 15984 40053 15984 40053 4 gnd
port 514 nsew
rlabel metal2 s 15984 41080 15984 41080 4 gnd
port 514 nsew
rlabel metal2 s 17232 38473 17232 38473 4 gnd
port 514 nsew
rlabel metal2 s 17232 39500 17232 39500 4 gnd
port 514 nsew
rlabel metal2 s 17232 38947 17232 38947 4 gnd
port 514 nsew
rlabel metal2 s 17232 40290 17232 40290 4 gnd
port 514 nsew
rlabel metal2 s 15984 40290 15984 40290 4 gnd
port 514 nsew
rlabel metal2 s 15984 39263 15984 39263 4 gnd
port 514 nsew
rlabel metal2 s 15984 40527 15984 40527 4 gnd
port 514 nsew
rlabel metal2 s 17232 41080 17232 41080 4 gnd
port 514 nsew
rlabel metal2 s 15216 40527 15216 40527 4 gnd
port 514 nsew
rlabel metal2 s 15984 38710 15984 38710 4 gnd
port 514 nsew
rlabel metal2 s 17232 39737 17232 39737 4 gnd
port 514 nsew
rlabel metal2 s 15984 38947 15984 38947 4 gnd
port 514 nsew
rlabel metal2 s 17232 38710 17232 38710 4 gnd
port 514 nsew
rlabel metal2 s 16464 40843 16464 40843 4 gnd
port 514 nsew
rlabel metal2 s 15984 40843 15984 40843 4 gnd
port 514 nsew
rlabel metal2 s 17232 40843 17232 40843 4 gnd
port 514 nsew
rlabel metal2 s 17232 38157 17232 38157 4 gnd
port 514 nsew
rlabel metal2 s 15216 40843 15216 40843 4 gnd
port 514 nsew
rlabel metal2 s 16464 38947 16464 38947 4 gnd
port 514 nsew
rlabel metal2 s 15216 41080 15216 41080 4 gnd
port 514 nsew
rlabel metal2 s 15216 38473 15216 38473 4 gnd
port 514 nsew
rlabel metal2 s 15216 40290 15216 40290 4 gnd
port 514 nsew
rlabel metal2 s 15984 39500 15984 39500 4 gnd
port 514 nsew
rlabel metal2 s 16464 41080 16464 41080 4 gnd
port 514 nsew
rlabel metal2 s 15984 38157 15984 38157 4 gnd
port 514 nsew
rlabel metal2 s 15216 38947 15216 38947 4 gnd
port 514 nsew
rlabel metal2 s 15216 40053 15216 40053 4 gnd
port 514 nsew
rlabel metal2 s 16464 40527 16464 40527 4 gnd
port 514 nsew
rlabel metal2 s 15984 39737 15984 39737 4 gnd
port 514 nsew
rlabel metal2 s 15984 38473 15984 38473 4 gnd
port 514 nsew
rlabel metal2 s 16464 38473 16464 38473 4 gnd
port 514 nsew
rlabel metal2 s 17232 39263 17232 39263 4 gnd
port 514 nsew
rlabel metal2 s 16464 40053 16464 40053 4 gnd
port 514 nsew
rlabel metal2 s 18480 39500 18480 39500 4 gnd
port 514 nsew
rlabel metal2 s 19728 41080 19728 41080 4 gnd
port 514 nsew
rlabel metal2 s 18480 38473 18480 38473 4 gnd
port 514 nsew
rlabel metal2 s 18480 39737 18480 39737 4 gnd
port 514 nsew
rlabel metal2 s 17712 39737 17712 39737 4 gnd
port 514 nsew
rlabel metal2 s 19728 39737 19728 39737 4 gnd
port 514 nsew
rlabel metal2 s 18960 40053 18960 40053 4 gnd
port 514 nsew
rlabel metal2 s 18480 40843 18480 40843 4 gnd
port 514 nsew
rlabel metal2 s 18960 40290 18960 40290 4 gnd
port 514 nsew
rlabel metal2 s 19728 38473 19728 38473 4 gnd
port 514 nsew
rlabel metal2 s 18960 38710 18960 38710 4 gnd
port 514 nsew
rlabel metal2 s 18480 39263 18480 39263 4 gnd
port 514 nsew
rlabel metal2 s 18480 38710 18480 38710 4 gnd
port 514 nsew
rlabel metal2 s 18960 39263 18960 39263 4 gnd
port 514 nsew
rlabel metal2 s 19728 40527 19728 40527 4 gnd
port 514 nsew
rlabel metal2 s 18960 41080 18960 41080 4 gnd
port 514 nsew
rlabel metal2 s 19968 40733 19968 40733 4 wl0_103
port 463 nsew
rlabel metal2 s 19728 40053 19728 40053 4 gnd
port 514 nsew
rlabel metal2 s 19728 40290 19728 40290 4 gnd
port 514 nsew
rlabel metal2 s 18480 40053 18480 40053 4 gnd
port 514 nsew
rlabel metal2 s 19968 39373 19968 39373 4 wl1_99
port 456 nsew
rlabel metal2 s 18480 38947 18480 38947 4 gnd
port 514 nsew
rlabel metal2 s 17712 39263 17712 39263 4 gnd
port 514 nsew
rlabel metal2 s 18480 38157 18480 38157 4 gnd
port 514 nsew
rlabel metal2 s 18960 40527 18960 40527 4 gnd
port 514 nsew
rlabel metal2 s 17712 41080 17712 41080 4 gnd
port 514 nsew
rlabel metal2 s 17712 38710 17712 38710 4 gnd
port 514 nsew
rlabel metal2 s 17712 38157 17712 38157 4 gnd
port 514 nsew
rlabel metal2 s 17712 40527 17712 40527 4 gnd
port 514 nsew
rlabel metal2 s 19968 39847 19968 39847 4 wl0_100
port 457 nsew
rlabel metal2 s 19968 40637 19968 40637 4 wl0_102
port 461 nsew
rlabel metal2 s 18480 41080 18480 41080 4 gnd
port 514 nsew
rlabel metal2 s 18480 40527 18480 40527 4 gnd
port 514 nsew
rlabel metal2 s 17712 39500 17712 39500 4 gnd
port 514 nsew
rlabel metal2 s 19968 40417 19968 40417 4 wl1_102
port 462 nsew
rlabel metal2 s 19968 38267 19968 38267 4 wl0_96
port 449 nsew
rlabel metal2 s 19968 39627 19968 39627 4 wl1_100
port 458 nsew
rlabel metal2 s 19968 39057 19968 39057 4 wl0_98
port 453 nsew
rlabel metal2 s 18960 38157 18960 38157 4 gnd
port 514 nsew
rlabel metal2 s 17712 40290 17712 40290 4 gnd
port 514 nsew
rlabel metal2 s 19968 39943 19968 39943 4 wl0_101
port 459 nsew
rlabel metal2 s 19728 38947 19728 38947 4 gnd
port 514 nsew
rlabel metal2 s 19728 38710 19728 38710 4 gnd
port 514 nsew
rlabel metal2 s 19728 40843 19728 40843 4 gnd
port 514 nsew
rlabel metal2 s 18960 38473 18960 38473 4 gnd
port 514 nsew
rlabel metal2 s 17712 38947 17712 38947 4 gnd
port 514 nsew
rlabel metal2 s 19968 38837 19968 38837 4 wl1_98
port 454 nsew
rlabel metal2 s 19968 38047 19968 38047 4 wl1_96
port 450 nsew
rlabel metal2 s 19728 39263 19728 39263 4 gnd
port 514 nsew
rlabel metal2 s 18480 40290 18480 40290 4 gnd
port 514 nsew
rlabel metal2 s 19728 38157 19728 38157 4 gnd
port 514 nsew
rlabel metal2 s 18960 40843 18960 40843 4 gnd
port 514 nsew
rlabel metal2 s 19728 39500 19728 39500 4 gnd
port 514 nsew
rlabel metal2 s 19968 38583 19968 38583 4 wl1_97
port 452 nsew
rlabel metal2 s 19968 40163 19968 40163 4 wl1_101
port 460 nsew
rlabel metal2 s 19968 40953 19968 40953 4 wl1_103
port 464 nsew
rlabel metal2 s 19968 39153 19968 39153 4 wl0_99
port 455 nsew
rlabel metal2 s 19968 38363 19968 38363 4 wl0_97
port 451 nsew
rlabel metal2 s 17712 40053 17712 40053 4 gnd
port 514 nsew
rlabel metal2 s 18960 39737 18960 39737 4 gnd
port 514 nsew
rlabel metal2 s 17712 40843 17712 40843 4 gnd
port 514 nsew
rlabel metal2 s 18960 39500 18960 39500 4 gnd
port 514 nsew
rlabel metal2 s 17712 38473 17712 38473 4 gnd
port 514 nsew
rlabel metal2 s 18960 38947 18960 38947 4 gnd
port 514 nsew
rlabel metal2 s 9744 47637 9744 47637 4 gnd
port 514 nsew
rlabel metal2 s 8976 50007 8976 50007 4 gnd
port 514 nsew
rlabel metal2 s 7728 49217 7728 49217 4 gnd
port 514 nsew
rlabel metal2 s 8976 47953 8976 47953 4 gnd
port 514 nsew
rlabel metal2 s 9744 48190 9744 48190 4 gnd
port 514 nsew
rlabel metal2 s 8976 49770 8976 49770 4 gnd
port 514 nsew
rlabel metal2 s 8496 50323 8496 50323 4 gnd
port 514 nsew
rlabel metal2 s 9744 50007 9744 50007 4 gnd
port 514 nsew
rlabel metal2 s 9744 48980 9744 48980 4 gnd
port 514 nsew
rlabel metal2 s 8496 48190 8496 48190 4 gnd
port 514 nsew
rlabel metal2 s 7728 48427 7728 48427 4 gnd
port 514 nsew
rlabel metal2 s 8976 47637 8976 47637 4 gnd
port 514 nsew
rlabel metal2 s 7728 49533 7728 49533 4 gnd
port 514 nsew
rlabel metal2 s 7728 48980 7728 48980 4 gnd
port 514 nsew
rlabel metal2 s 8496 50007 8496 50007 4 gnd
port 514 nsew
rlabel metal2 s 9744 47953 9744 47953 4 gnd
port 514 nsew
rlabel metal2 s 7728 48190 7728 48190 4 gnd
port 514 nsew
rlabel metal2 s 8976 49533 8976 49533 4 gnd
port 514 nsew
rlabel metal2 s 8976 50323 8976 50323 4 gnd
port 514 nsew
rlabel metal2 s 7728 50007 7728 50007 4 gnd
port 514 nsew
rlabel metal2 s 8496 47953 8496 47953 4 gnd
port 514 nsew
rlabel metal2 s 8496 48427 8496 48427 4 gnd
port 514 nsew
rlabel metal2 s 8496 47637 8496 47637 4 gnd
port 514 nsew
rlabel metal2 s 9744 48743 9744 48743 4 gnd
port 514 nsew
rlabel metal2 s 7728 49770 7728 49770 4 gnd
port 514 nsew
rlabel metal2 s 7728 50560 7728 50560 4 gnd
port 514 nsew
rlabel metal2 s 8976 48427 8976 48427 4 gnd
port 514 nsew
rlabel metal2 s 8496 49770 8496 49770 4 gnd
port 514 nsew
rlabel metal2 s 9744 49533 9744 49533 4 gnd
port 514 nsew
rlabel metal2 s 8976 48980 8976 48980 4 gnd
port 514 nsew
rlabel metal2 s 9744 50560 9744 50560 4 gnd
port 514 nsew
rlabel metal2 s 8496 49533 8496 49533 4 gnd
port 514 nsew
rlabel metal2 s 8496 48743 8496 48743 4 gnd
port 514 nsew
rlabel metal2 s 8976 48190 8976 48190 4 gnd
port 514 nsew
rlabel metal2 s 9744 48427 9744 48427 4 gnd
port 514 nsew
rlabel metal2 s 7728 48743 7728 48743 4 gnd
port 514 nsew
rlabel metal2 s 9744 49770 9744 49770 4 gnd
port 514 nsew
rlabel metal2 s 8496 48980 8496 48980 4 gnd
port 514 nsew
rlabel metal2 s 7728 50323 7728 50323 4 gnd
port 514 nsew
rlabel metal2 s 7728 47637 7728 47637 4 gnd
port 514 nsew
rlabel metal2 s 8496 49217 8496 49217 4 gnd
port 514 nsew
rlabel metal2 s 9744 50323 9744 50323 4 gnd
port 514 nsew
rlabel metal2 s 8496 50560 8496 50560 4 gnd
port 514 nsew
rlabel metal2 s 8976 50560 8976 50560 4 gnd
port 514 nsew
rlabel metal2 s 7728 47953 7728 47953 4 gnd
port 514 nsew
rlabel metal2 s 8976 48743 8976 48743 4 gnd
port 514 nsew
rlabel metal2 s 9744 49217 9744 49217 4 gnd
port 514 nsew
rlabel metal2 s 8976 49217 8976 49217 4 gnd
port 514 nsew
rlabel metal2 s 6480 50560 6480 50560 4 gnd
port 514 nsew
rlabel metal2 s 6480 47953 6480 47953 4 gnd
port 514 nsew
rlabel metal2 s 6000 47953 6000 47953 4 gnd
port 514 nsew
rlabel metal2 s 7248 50560 7248 50560 4 gnd
port 514 nsew
rlabel metal2 s 6000 50323 6000 50323 4 gnd
port 514 nsew
rlabel metal2 s 7248 48980 7248 48980 4 gnd
port 514 nsew
rlabel metal2 s 5232 47953 5232 47953 4 gnd
port 514 nsew
rlabel metal2 s 5232 49217 5232 49217 4 gnd
port 514 nsew
rlabel metal2 s 6480 49770 6480 49770 4 gnd
port 514 nsew
rlabel metal2 s 7248 49770 7248 49770 4 gnd
port 514 nsew
rlabel metal2 s 6000 48743 6000 48743 4 gnd
port 514 nsew
rlabel metal2 s 5232 48190 5232 48190 4 gnd
port 514 nsew
rlabel metal2 s 6000 48980 6000 48980 4 gnd
port 514 nsew
rlabel metal2 s 6480 49217 6480 49217 4 gnd
port 514 nsew
rlabel metal2 s 5232 47637 5232 47637 4 gnd
port 514 nsew
rlabel metal2 s 7248 47953 7248 47953 4 gnd
port 514 nsew
rlabel metal2 s 6000 50007 6000 50007 4 gnd
port 514 nsew
rlabel metal2 s 7248 49217 7248 49217 4 gnd
port 514 nsew
rlabel metal2 s 5232 48743 5232 48743 4 gnd
port 514 nsew
rlabel metal2 s 6000 48427 6000 48427 4 gnd
port 514 nsew
rlabel metal2 s 6480 48980 6480 48980 4 gnd
port 514 nsew
rlabel metal2 s 6000 48190 6000 48190 4 gnd
port 514 nsew
rlabel metal2 s 5232 49533 5232 49533 4 gnd
port 514 nsew
rlabel metal2 s 7248 50007 7248 50007 4 gnd
port 514 nsew
rlabel metal2 s 6480 49533 6480 49533 4 gnd
port 514 nsew
rlabel metal2 s 7248 48190 7248 48190 4 gnd
port 514 nsew
rlabel metal2 s 5232 50007 5232 50007 4 gnd
port 514 nsew
rlabel metal2 s 6000 47637 6000 47637 4 gnd
port 514 nsew
rlabel metal2 s 7248 48427 7248 48427 4 gnd
port 514 nsew
rlabel metal2 s 7248 48743 7248 48743 4 gnd
port 514 nsew
rlabel metal2 s 5232 48980 5232 48980 4 gnd
port 514 nsew
rlabel metal2 s 6480 48190 6480 48190 4 gnd
port 514 nsew
rlabel metal2 s 7248 47637 7248 47637 4 gnd
port 514 nsew
rlabel metal2 s 6000 49533 6000 49533 4 gnd
port 514 nsew
rlabel metal2 s 5232 49770 5232 49770 4 gnd
port 514 nsew
rlabel metal2 s 6480 50007 6480 50007 4 gnd
port 514 nsew
rlabel metal2 s 6480 48427 6480 48427 4 gnd
port 514 nsew
rlabel metal2 s 6480 50323 6480 50323 4 gnd
port 514 nsew
rlabel metal2 s 5232 48427 5232 48427 4 gnd
port 514 nsew
rlabel metal2 s 6000 49217 6000 49217 4 gnd
port 514 nsew
rlabel metal2 s 5232 50560 5232 50560 4 gnd
port 514 nsew
rlabel metal2 s 7248 50323 7248 50323 4 gnd
port 514 nsew
rlabel metal2 s 6480 48743 6480 48743 4 gnd
port 514 nsew
rlabel metal2 s 7248 49533 7248 49533 4 gnd
port 514 nsew
rlabel metal2 s 5232 50323 5232 50323 4 gnd
port 514 nsew
rlabel metal2 s 6000 49770 6000 49770 4 gnd
port 514 nsew
rlabel metal2 s 6480 47637 6480 47637 4 gnd
port 514 nsew
rlabel metal2 s 6000 50560 6000 50560 4 gnd
port 514 nsew
rlabel metal2 s 5232 46373 5232 46373 4 gnd
port 514 nsew
rlabel metal2 s 6000 47400 6000 47400 4 gnd
port 514 nsew
rlabel metal2 s 7248 45820 7248 45820 4 gnd
port 514 nsew
rlabel metal2 s 7248 44477 7248 44477 4 gnd
port 514 nsew
rlabel metal2 s 6000 45583 6000 45583 4 gnd
port 514 nsew
rlabel metal2 s 6000 46847 6000 46847 4 gnd
port 514 nsew
rlabel metal2 s 5232 45030 5232 45030 4 gnd
port 514 nsew
rlabel metal2 s 6000 46057 6000 46057 4 gnd
port 514 nsew
rlabel metal2 s 6000 47163 6000 47163 4 gnd
port 514 nsew
rlabel metal2 s 7248 47400 7248 47400 4 gnd
port 514 nsew
rlabel metal2 s 6480 46610 6480 46610 4 gnd
port 514 nsew
rlabel metal2 s 7248 47163 7248 47163 4 gnd
port 514 nsew
rlabel metal2 s 7248 45583 7248 45583 4 gnd
port 514 nsew
rlabel metal2 s 5232 45820 5232 45820 4 gnd
port 514 nsew
rlabel metal2 s 6480 46847 6480 46847 4 gnd
port 514 nsew
rlabel metal2 s 6480 44793 6480 44793 4 gnd
port 514 nsew
rlabel metal2 s 6480 45030 6480 45030 4 gnd
port 514 nsew
rlabel metal2 s 6480 45267 6480 45267 4 gnd
port 514 nsew
rlabel metal2 s 6000 45267 6000 45267 4 gnd
port 514 nsew
rlabel metal2 s 5232 46847 5232 46847 4 gnd
port 514 nsew
rlabel metal2 s 6480 47400 6480 47400 4 gnd
port 514 nsew
rlabel metal2 s 6000 45030 6000 45030 4 gnd
port 514 nsew
rlabel metal2 s 6480 45583 6480 45583 4 gnd
port 514 nsew
rlabel metal2 s 6480 46057 6480 46057 4 gnd
port 514 nsew
rlabel metal2 s 5232 46057 5232 46057 4 gnd
port 514 nsew
rlabel metal2 s 6000 45820 6000 45820 4 gnd
port 514 nsew
rlabel metal2 s 5232 45583 5232 45583 4 gnd
port 514 nsew
rlabel metal2 s 5232 44793 5232 44793 4 gnd
port 514 nsew
rlabel metal2 s 5232 46610 5232 46610 4 gnd
port 514 nsew
rlabel metal2 s 7248 46057 7248 46057 4 gnd
port 514 nsew
rlabel metal2 s 6480 45820 6480 45820 4 gnd
port 514 nsew
rlabel metal2 s 6480 44477 6480 44477 4 gnd
port 514 nsew
rlabel metal2 s 5232 44477 5232 44477 4 gnd
port 514 nsew
rlabel metal2 s 5232 47163 5232 47163 4 gnd
port 514 nsew
rlabel metal2 s 5232 45267 5232 45267 4 gnd
port 514 nsew
rlabel metal2 s 7248 45267 7248 45267 4 gnd
port 514 nsew
rlabel metal2 s 6000 46373 6000 46373 4 gnd
port 514 nsew
rlabel metal2 s 6000 46610 6000 46610 4 gnd
port 514 nsew
rlabel metal2 s 7248 44793 7248 44793 4 gnd
port 514 nsew
rlabel metal2 s 7248 46847 7248 46847 4 gnd
port 514 nsew
rlabel metal2 s 5232 47400 5232 47400 4 gnd
port 514 nsew
rlabel metal2 s 7248 45030 7248 45030 4 gnd
port 514 nsew
rlabel metal2 s 6000 44793 6000 44793 4 gnd
port 514 nsew
rlabel metal2 s 6480 46373 6480 46373 4 gnd
port 514 nsew
rlabel metal2 s 6000 44477 6000 44477 4 gnd
port 514 nsew
rlabel metal2 s 7248 46610 7248 46610 4 gnd
port 514 nsew
rlabel metal2 s 7248 46373 7248 46373 4 gnd
port 514 nsew
rlabel metal2 s 6480 47163 6480 47163 4 gnd
port 514 nsew
rlabel metal2 s 8976 45267 8976 45267 4 gnd
port 514 nsew
rlabel metal2 s 8496 46847 8496 46847 4 gnd
port 514 nsew
rlabel metal2 s 8976 46057 8976 46057 4 gnd
port 514 nsew
rlabel metal2 s 7728 45030 7728 45030 4 gnd
port 514 nsew
rlabel metal2 s 8496 44793 8496 44793 4 gnd
port 514 nsew
rlabel metal2 s 8496 46373 8496 46373 4 gnd
port 514 nsew
rlabel metal2 s 7728 44793 7728 44793 4 gnd
port 514 nsew
rlabel metal2 s 7728 45583 7728 45583 4 gnd
port 514 nsew
rlabel metal2 s 8496 47400 8496 47400 4 gnd
port 514 nsew
rlabel metal2 s 8976 46847 8976 46847 4 gnd
port 514 nsew
rlabel metal2 s 9744 44477 9744 44477 4 gnd
port 514 nsew
rlabel metal2 s 9744 47400 9744 47400 4 gnd
port 514 nsew
rlabel metal2 s 8496 45820 8496 45820 4 gnd
port 514 nsew
rlabel metal2 s 8496 47163 8496 47163 4 gnd
port 514 nsew
rlabel metal2 s 8496 45030 8496 45030 4 gnd
port 514 nsew
rlabel metal2 s 8976 46373 8976 46373 4 gnd
port 514 nsew
rlabel metal2 s 7728 45820 7728 45820 4 gnd
port 514 nsew
rlabel metal2 s 8496 46057 8496 46057 4 gnd
port 514 nsew
rlabel metal2 s 7728 47163 7728 47163 4 gnd
port 514 nsew
rlabel metal2 s 8976 47400 8976 47400 4 gnd
port 514 nsew
rlabel metal2 s 8976 45583 8976 45583 4 gnd
port 514 nsew
rlabel metal2 s 7728 45267 7728 45267 4 gnd
port 514 nsew
rlabel metal2 s 7728 46610 7728 46610 4 gnd
port 514 nsew
rlabel metal2 s 8976 46610 8976 46610 4 gnd
port 514 nsew
rlabel metal2 s 9744 45267 9744 45267 4 gnd
port 514 nsew
rlabel metal2 s 7728 46057 7728 46057 4 gnd
port 514 nsew
rlabel metal2 s 8496 46610 8496 46610 4 gnd
port 514 nsew
rlabel metal2 s 9744 46847 9744 46847 4 gnd
port 514 nsew
rlabel metal2 s 8496 44477 8496 44477 4 gnd
port 514 nsew
rlabel metal2 s 7728 46373 7728 46373 4 gnd
port 514 nsew
rlabel metal2 s 9744 45030 9744 45030 4 gnd
port 514 nsew
rlabel metal2 s 9744 45583 9744 45583 4 gnd
port 514 nsew
rlabel metal2 s 9744 47163 9744 47163 4 gnd
port 514 nsew
rlabel metal2 s 9744 46610 9744 46610 4 gnd
port 514 nsew
rlabel metal2 s 9744 44793 9744 44793 4 gnd
port 514 nsew
rlabel metal2 s 7728 47400 7728 47400 4 gnd
port 514 nsew
rlabel metal2 s 9744 46057 9744 46057 4 gnd
port 514 nsew
rlabel metal2 s 8976 44477 8976 44477 4 gnd
port 514 nsew
rlabel metal2 s 8496 45267 8496 45267 4 gnd
port 514 nsew
rlabel metal2 s 9744 46373 9744 46373 4 gnd
port 514 nsew
rlabel metal2 s 8976 45820 8976 45820 4 gnd
port 514 nsew
rlabel metal2 s 9744 45820 9744 45820 4 gnd
port 514 nsew
rlabel metal2 s 8496 45583 8496 45583 4 gnd
port 514 nsew
rlabel metal2 s 8976 47163 8976 47163 4 gnd
port 514 nsew
rlabel metal2 s 7728 44477 7728 44477 4 gnd
port 514 nsew
rlabel metal2 s 7728 46847 7728 46847 4 gnd
port 514 nsew
rlabel metal2 s 8976 45030 8976 45030 4 gnd
port 514 nsew
rlabel metal2 s 8976 44793 8976 44793 4 gnd
port 514 nsew
rlabel metal2 s 3504 47637 3504 47637 4 gnd
port 514 nsew
rlabel metal2 s 3984 49217 3984 49217 4 gnd
port 514 nsew
rlabel metal2 s 2736 48980 2736 48980 4 gnd
port 514 nsew
rlabel metal2 s 3984 48427 3984 48427 4 gnd
port 514 nsew
rlabel metal2 s 4752 50007 4752 50007 4 gnd
port 514 nsew
rlabel metal2 s 4752 49217 4752 49217 4 gnd
port 514 nsew
rlabel metal2 s 3504 49770 3504 49770 4 gnd
port 514 nsew
rlabel metal2 s 3984 49533 3984 49533 4 gnd
port 514 nsew
rlabel metal2 s 3504 48427 3504 48427 4 gnd
port 514 nsew
rlabel metal2 s 2736 50560 2736 50560 4 gnd
port 514 nsew
rlabel metal2 s 3984 49770 3984 49770 4 gnd
port 514 nsew
rlabel metal2 s 3984 48190 3984 48190 4 gnd
port 514 nsew
rlabel metal2 s 4752 47637 4752 47637 4 gnd
port 514 nsew
rlabel metal2 s 2736 47637 2736 47637 4 gnd
port 514 nsew
rlabel metal2 s 3984 50007 3984 50007 4 gnd
port 514 nsew
rlabel metal2 s 3504 48980 3504 48980 4 gnd
port 514 nsew
rlabel metal2 s 4752 48743 4752 48743 4 gnd
port 514 nsew
rlabel metal2 s 4752 50560 4752 50560 4 gnd
port 514 nsew
rlabel metal2 s 3504 50560 3504 50560 4 gnd
port 514 nsew
rlabel metal2 s 4752 50323 4752 50323 4 gnd
port 514 nsew
rlabel metal2 s 3984 50323 3984 50323 4 gnd
port 514 nsew
rlabel metal2 s 2736 50007 2736 50007 4 gnd
port 514 nsew
rlabel metal2 s 4752 49770 4752 49770 4 gnd
port 514 nsew
rlabel metal2 s 3984 47953 3984 47953 4 gnd
port 514 nsew
rlabel metal2 s 2736 49533 2736 49533 4 gnd
port 514 nsew
rlabel metal2 s 3504 47953 3504 47953 4 gnd
port 514 nsew
rlabel metal2 s 3504 49217 3504 49217 4 gnd
port 514 nsew
rlabel metal2 s 2736 50323 2736 50323 4 gnd
port 514 nsew
rlabel metal2 s 4752 48980 4752 48980 4 gnd
port 514 nsew
rlabel metal2 s 3504 50007 3504 50007 4 gnd
port 514 nsew
rlabel metal2 s 3504 48190 3504 48190 4 gnd
port 514 nsew
rlabel metal2 s 2736 48743 2736 48743 4 gnd
port 514 nsew
rlabel metal2 s 4752 48427 4752 48427 4 gnd
port 514 nsew
rlabel metal2 s 3984 48743 3984 48743 4 gnd
port 514 nsew
rlabel metal2 s 3504 49533 3504 49533 4 gnd
port 514 nsew
rlabel metal2 s 3504 50323 3504 50323 4 gnd
port 514 nsew
rlabel metal2 s 2736 47953 2736 47953 4 gnd
port 514 nsew
rlabel metal2 s 2736 48427 2736 48427 4 gnd
port 514 nsew
rlabel metal2 s 4752 49533 4752 49533 4 gnd
port 514 nsew
rlabel metal2 s 3984 47637 3984 47637 4 gnd
port 514 nsew
rlabel metal2 s 4752 48190 4752 48190 4 gnd
port 514 nsew
rlabel metal2 s 3504 48743 3504 48743 4 gnd
port 514 nsew
rlabel metal2 s 2736 48190 2736 48190 4 gnd
port 514 nsew
rlabel metal2 s 2736 49217 2736 49217 4 gnd
port 514 nsew
rlabel metal2 s 4752 47953 4752 47953 4 gnd
port 514 nsew
rlabel metal2 s 3984 50560 3984 50560 4 gnd
port 514 nsew
rlabel metal2 s 2736 49770 2736 49770 4 gnd
port 514 nsew
rlabel metal2 s 3984 48980 3984 48980 4 gnd
port 514 nsew
rlabel metal2 s 240 48743 240 48743 4 gnd
port 514 nsew
rlabel metal2 s 2256 49217 2256 49217 4 gnd
port 514 nsew
rlabel metal2 s 1008 48427 1008 48427 4 gnd
port 514 nsew
rlabel metal2 s 240 48427 240 48427 4 gnd
port 514 nsew
rlabel metal2 s 1488 50323 1488 50323 4 gnd
port 514 nsew
rlabel metal2 s 240 49217 240 49217 4 gnd
port 514 nsew
rlabel metal2 s 1488 48980 1488 48980 4 gnd
port 514 nsew
rlabel metal2 s 1488 48743 1488 48743 4 gnd
port 514 nsew
rlabel metal2 s 1488 49770 1488 49770 4 gnd
port 514 nsew
rlabel metal2 s 240 49533 240 49533 4 gnd
port 514 nsew
rlabel metal2 s 2256 48743 2256 48743 4 gnd
port 514 nsew
rlabel metal2 s 2256 50560 2256 50560 4 gnd
port 514 nsew
rlabel metal2 s 2256 50007 2256 50007 4 gnd
port 514 nsew
rlabel metal2 s 1008 49770 1008 49770 4 gnd
port 514 nsew
rlabel metal2 s 2256 47953 2256 47953 4 gnd
port 514 nsew
rlabel metal2 s 1488 49533 1488 49533 4 gnd
port 514 nsew
rlabel metal2 s 1008 47637 1008 47637 4 gnd
port 514 nsew
rlabel metal2 s 2256 48190 2256 48190 4 gnd
port 514 nsew
rlabel metal2 s 1008 49217 1008 49217 4 gnd
port 514 nsew
rlabel metal2 s 240 49770 240 49770 4 gnd
port 514 nsew
rlabel metal2 s 240 50560 240 50560 4 gnd
port 514 nsew
rlabel metal2 s 1008 48743 1008 48743 4 gnd
port 514 nsew
rlabel metal2 s 2256 47637 2256 47637 4 gnd
port 514 nsew
rlabel metal2 s 2256 48427 2256 48427 4 gnd
port 514 nsew
rlabel metal2 s 2256 50323 2256 50323 4 gnd
port 514 nsew
rlabel metal2 s 240 50007 240 50007 4 gnd
port 514 nsew
rlabel metal2 s 1008 47953 1008 47953 4 gnd
port 514 nsew
rlabel metal2 s 1008 49533 1008 49533 4 gnd
port 514 nsew
rlabel metal2 s 2256 49533 2256 49533 4 gnd
port 514 nsew
rlabel metal2 s 1488 48427 1488 48427 4 gnd
port 514 nsew
rlabel metal2 s 1488 49217 1488 49217 4 gnd
port 514 nsew
rlabel metal2 s 1008 50560 1008 50560 4 gnd
port 514 nsew
rlabel metal2 s 240 47953 240 47953 4 gnd
port 514 nsew
rlabel metal2 s 2256 49770 2256 49770 4 gnd
port 514 nsew
rlabel metal2 s 1488 50007 1488 50007 4 gnd
port 514 nsew
rlabel metal2 s 1008 48980 1008 48980 4 gnd
port 514 nsew
rlabel metal2 s 1488 48190 1488 48190 4 gnd
port 514 nsew
rlabel metal2 s 1488 47637 1488 47637 4 gnd
port 514 nsew
rlabel metal2 s 240 48980 240 48980 4 gnd
port 514 nsew
rlabel metal2 s 1008 50323 1008 50323 4 gnd
port 514 nsew
rlabel metal2 s 1008 50007 1008 50007 4 gnd
port 514 nsew
rlabel metal2 s 2256 48980 2256 48980 4 gnd
port 514 nsew
rlabel metal2 s 1488 50560 1488 50560 4 gnd
port 514 nsew
rlabel metal2 s 240 47637 240 47637 4 gnd
port 514 nsew
rlabel metal2 s 1488 47953 1488 47953 4 gnd
port 514 nsew
rlabel metal2 s 240 50323 240 50323 4 gnd
port 514 nsew
rlabel metal2 s 240 48190 240 48190 4 gnd
port 514 nsew
rlabel metal2 s 1008 48190 1008 48190 4 gnd
port 514 nsew
rlabel metal2 s 1008 46847 1008 46847 4 gnd
port 514 nsew
rlabel metal2 s 1488 44793 1488 44793 4 gnd
port 514 nsew
rlabel metal2 s 2256 46610 2256 46610 4 gnd
port 514 nsew
rlabel metal2 s 2256 44477 2256 44477 4 gnd
port 514 nsew
rlabel metal2 s 1008 45267 1008 45267 4 gnd
port 514 nsew
rlabel metal2 s 1488 46373 1488 46373 4 gnd
port 514 nsew
rlabel metal2 s 1008 47163 1008 47163 4 gnd
port 514 nsew
rlabel metal2 s 2256 45030 2256 45030 4 gnd
port 514 nsew
rlabel metal2 s 2256 44793 2256 44793 4 gnd
port 514 nsew
rlabel metal2 s 1008 46610 1008 46610 4 gnd
port 514 nsew
rlabel metal2 s 1008 46373 1008 46373 4 gnd
port 514 nsew
rlabel metal2 s 240 46847 240 46847 4 gnd
port 514 nsew
rlabel metal2 s 240 46373 240 46373 4 gnd
port 514 nsew
rlabel metal2 s 240 45820 240 45820 4 gnd
port 514 nsew
rlabel metal2 s 1488 45030 1488 45030 4 gnd
port 514 nsew
rlabel metal2 s 1008 44793 1008 44793 4 gnd
port 514 nsew
rlabel metal2 s 1488 46610 1488 46610 4 gnd
port 514 nsew
rlabel metal2 s 1488 45267 1488 45267 4 gnd
port 514 nsew
rlabel metal2 s 2256 46847 2256 46847 4 gnd
port 514 nsew
rlabel metal2 s 240 46057 240 46057 4 gnd
port 514 nsew
rlabel metal2 s 1488 45583 1488 45583 4 gnd
port 514 nsew
rlabel metal2 s 1008 47400 1008 47400 4 gnd
port 514 nsew
rlabel metal2 s 2256 45820 2256 45820 4 gnd
port 514 nsew
rlabel metal2 s 2256 47400 2256 47400 4 gnd
port 514 nsew
rlabel metal2 s 1488 47163 1488 47163 4 gnd
port 514 nsew
rlabel metal2 s 1488 44477 1488 44477 4 gnd
port 514 nsew
rlabel metal2 s 1488 45820 1488 45820 4 gnd
port 514 nsew
rlabel metal2 s 1488 46057 1488 46057 4 gnd
port 514 nsew
rlabel metal2 s 1008 45583 1008 45583 4 gnd
port 514 nsew
rlabel metal2 s 240 45030 240 45030 4 gnd
port 514 nsew
rlabel metal2 s 2256 45267 2256 45267 4 gnd
port 514 nsew
rlabel metal2 s 240 47400 240 47400 4 gnd
port 514 nsew
rlabel metal2 s 1008 45820 1008 45820 4 gnd
port 514 nsew
rlabel metal2 s 240 44477 240 44477 4 gnd
port 514 nsew
rlabel metal2 s 240 47163 240 47163 4 gnd
port 514 nsew
rlabel metal2 s 1008 45030 1008 45030 4 gnd
port 514 nsew
rlabel metal2 s 1008 46057 1008 46057 4 gnd
port 514 nsew
rlabel metal2 s 240 44793 240 44793 4 gnd
port 514 nsew
rlabel metal2 s 240 46610 240 46610 4 gnd
port 514 nsew
rlabel metal2 s 2256 47163 2256 47163 4 gnd
port 514 nsew
rlabel metal2 s 240 45267 240 45267 4 gnd
port 514 nsew
rlabel metal2 s 1488 46847 1488 46847 4 gnd
port 514 nsew
rlabel metal2 s 2256 46373 2256 46373 4 gnd
port 514 nsew
rlabel metal2 s 240 45583 240 45583 4 gnd
port 514 nsew
rlabel metal2 s 1488 47400 1488 47400 4 gnd
port 514 nsew
rlabel metal2 s 1008 44477 1008 44477 4 gnd
port 514 nsew
rlabel metal2 s 2256 45583 2256 45583 4 gnd
port 514 nsew
rlabel metal2 s 2256 46057 2256 46057 4 gnd
port 514 nsew
rlabel metal2 s 2736 46847 2736 46847 4 gnd
port 514 nsew
rlabel metal2 s 3984 44477 3984 44477 4 gnd
port 514 nsew
rlabel metal2 s 3984 45030 3984 45030 4 gnd
port 514 nsew
rlabel metal2 s 4752 44793 4752 44793 4 gnd
port 514 nsew
rlabel metal2 s 3984 47163 3984 47163 4 gnd
port 514 nsew
rlabel metal2 s 4752 45820 4752 45820 4 gnd
port 514 nsew
rlabel metal2 s 3984 45820 3984 45820 4 gnd
port 514 nsew
rlabel metal2 s 4752 45030 4752 45030 4 gnd
port 514 nsew
rlabel metal2 s 3504 46610 3504 46610 4 gnd
port 514 nsew
rlabel metal2 s 3504 45820 3504 45820 4 gnd
port 514 nsew
rlabel metal2 s 4752 45583 4752 45583 4 gnd
port 514 nsew
rlabel metal2 s 3984 46847 3984 46847 4 gnd
port 514 nsew
rlabel metal2 s 2736 47163 2736 47163 4 gnd
port 514 nsew
rlabel metal2 s 3984 44793 3984 44793 4 gnd
port 514 nsew
rlabel metal2 s 3504 47163 3504 47163 4 gnd
port 514 nsew
rlabel metal2 s 3504 44793 3504 44793 4 gnd
port 514 nsew
rlabel metal2 s 2736 45583 2736 45583 4 gnd
port 514 nsew
rlabel metal2 s 3984 46057 3984 46057 4 gnd
port 514 nsew
rlabel metal2 s 2736 45267 2736 45267 4 gnd
port 514 nsew
rlabel metal2 s 3504 46373 3504 46373 4 gnd
port 514 nsew
rlabel metal2 s 3984 47400 3984 47400 4 gnd
port 514 nsew
rlabel metal2 s 3984 46373 3984 46373 4 gnd
port 514 nsew
rlabel metal2 s 2736 46610 2736 46610 4 gnd
port 514 nsew
rlabel metal2 s 2736 44793 2736 44793 4 gnd
port 514 nsew
rlabel metal2 s 3504 45267 3504 45267 4 gnd
port 514 nsew
rlabel metal2 s 4752 46373 4752 46373 4 gnd
port 514 nsew
rlabel metal2 s 4752 46847 4752 46847 4 gnd
port 514 nsew
rlabel metal2 s 2736 45820 2736 45820 4 gnd
port 514 nsew
rlabel metal2 s 2736 46057 2736 46057 4 gnd
port 514 nsew
rlabel metal2 s 4752 44477 4752 44477 4 gnd
port 514 nsew
rlabel metal2 s 3504 46057 3504 46057 4 gnd
port 514 nsew
rlabel metal2 s 3984 46610 3984 46610 4 gnd
port 514 nsew
rlabel metal2 s 4752 46610 4752 46610 4 gnd
port 514 nsew
rlabel metal2 s 4752 47163 4752 47163 4 gnd
port 514 nsew
rlabel metal2 s 3504 46847 3504 46847 4 gnd
port 514 nsew
rlabel metal2 s 3984 45267 3984 45267 4 gnd
port 514 nsew
rlabel metal2 s 2736 46373 2736 46373 4 gnd
port 514 nsew
rlabel metal2 s 3504 45583 3504 45583 4 gnd
port 514 nsew
rlabel metal2 s 3504 44477 3504 44477 4 gnd
port 514 nsew
rlabel metal2 s 2736 44477 2736 44477 4 gnd
port 514 nsew
rlabel metal2 s 4752 46057 4752 46057 4 gnd
port 514 nsew
rlabel metal2 s 3504 47400 3504 47400 4 gnd
port 514 nsew
rlabel metal2 s 3984 45583 3984 45583 4 gnd
port 514 nsew
rlabel metal2 s 3504 45030 3504 45030 4 gnd
port 514 nsew
rlabel metal2 s 4752 47400 4752 47400 4 gnd
port 514 nsew
rlabel metal2 s 2736 45030 2736 45030 4 gnd
port 514 nsew
rlabel metal2 s 2736 47400 2736 47400 4 gnd
port 514 nsew
rlabel metal2 s 4752 45267 4752 45267 4 gnd
port 514 nsew
rlabel metal2 s 3984 42423 3984 42423 4 gnd
port 514 nsew
rlabel metal2 s 3984 42897 3984 42897 4 gnd
port 514 nsew
rlabel metal2 s 4752 42423 4752 42423 4 gnd
port 514 nsew
rlabel metal2 s 4752 41317 4752 41317 4 gnd
port 514 nsew
rlabel metal2 s 2736 41317 2736 41317 4 gnd
port 514 nsew
rlabel metal2 s 4752 44240 4752 44240 4 gnd
port 514 nsew
rlabel metal2 s 2736 41633 2736 41633 4 gnd
port 514 nsew
rlabel metal2 s 3984 43450 3984 43450 4 gnd
port 514 nsew
rlabel metal2 s 3984 43213 3984 43213 4 gnd
port 514 nsew
rlabel metal2 s 3504 41633 3504 41633 4 gnd
port 514 nsew
rlabel metal2 s 2736 42107 2736 42107 4 gnd
port 514 nsew
rlabel metal2 s 3504 41870 3504 41870 4 gnd
port 514 nsew
rlabel metal2 s 3984 41317 3984 41317 4 gnd
port 514 nsew
rlabel metal2 s 3984 44240 3984 44240 4 gnd
port 514 nsew
rlabel metal2 s 3504 42660 3504 42660 4 gnd
port 514 nsew
rlabel metal2 s 3984 41633 3984 41633 4 gnd
port 514 nsew
rlabel metal2 s 2736 41870 2736 41870 4 gnd
port 514 nsew
rlabel metal2 s 4752 43687 4752 43687 4 gnd
port 514 nsew
rlabel metal2 s 3504 41317 3504 41317 4 gnd
port 514 nsew
rlabel metal2 s 2736 44003 2736 44003 4 gnd
port 514 nsew
rlabel metal2 s 3984 44003 3984 44003 4 gnd
port 514 nsew
rlabel metal2 s 4752 41633 4752 41633 4 gnd
port 514 nsew
rlabel metal2 s 3504 43213 3504 43213 4 gnd
port 514 nsew
rlabel metal2 s 2736 42423 2736 42423 4 gnd
port 514 nsew
rlabel metal2 s 3504 42897 3504 42897 4 gnd
port 514 nsew
rlabel metal2 s 3504 42423 3504 42423 4 gnd
port 514 nsew
rlabel metal2 s 4752 41870 4752 41870 4 gnd
port 514 nsew
rlabel metal2 s 3504 44003 3504 44003 4 gnd
port 514 nsew
rlabel metal2 s 3984 43687 3984 43687 4 gnd
port 514 nsew
rlabel metal2 s 3984 42107 3984 42107 4 gnd
port 514 nsew
rlabel metal2 s 3984 41870 3984 41870 4 gnd
port 514 nsew
rlabel metal2 s 4752 42107 4752 42107 4 gnd
port 514 nsew
rlabel metal2 s 2736 43687 2736 43687 4 gnd
port 514 nsew
rlabel metal2 s 4752 43450 4752 43450 4 gnd
port 514 nsew
rlabel metal2 s 4752 42660 4752 42660 4 gnd
port 514 nsew
rlabel metal2 s 2736 42660 2736 42660 4 gnd
port 514 nsew
rlabel metal2 s 4752 42897 4752 42897 4 gnd
port 514 nsew
rlabel metal2 s 2736 43213 2736 43213 4 gnd
port 514 nsew
rlabel metal2 s 3504 44240 3504 44240 4 gnd
port 514 nsew
rlabel metal2 s 3504 43450 3504 43450 4 gnd
port 514 nsew
rlabel metal2 s 2736 43450 2736 43450 4 gnd
port 514 nsew
rlabel metal2 s 2736 44240 2736 44240 4 gnd
port 514 nsew
rlabel metal2 s 2736 42897 2736 42897 4 gnd
port 514 nsew
rlabel metal2 s 3504 43687 3504 43687 4 gnd
port 514 nsew
rlabel metal2 s 4752 43213 4752 43213 4 gnd
port 514 nsew
rlabel metal2 s 3984 42660 3984 42660 4 gnd
port 514 nsew
rlabel metal2 s 4752 44003 4752 44003 4 gnd
port 514 nsew
rlabel metal2 s 3504 42107 3504 42107 4 gnd
port 514 nsew
rlabel metal2 s 2256 44240 2256 44240 4 gnd
port 514 nsew
rlabel metal2 s 1008 41870 1008 41870 4 gnd
port 514 nsew
rlabel metal2 s 1488 41317 1488 41317 4 gnd
port 514 nsew
rlabel metal2 s 1008 42423 1008 42423 4 gnd
port 514 nsew
rlabel metal2 s 1008 43450 1008 43450 4 gnd
port 514 nsew
rlabel metal2 s 1488 44240 1488 44240 4 gnd
port 514 nsew
rlabel metal2 s 1008 42660 1008 42660 4 gnd
port 514 nsew
rlabel metal2 s 2256 43213 2256 43213 4 gnd
port 514 nsew
rlabel metal2 s 1008 43687 1008 43687 4 gnd
port 514 nsew
rlabel metal2 s 2256 41870 2256 41870 4 gnd
port 514 nsew
rlabel metal2 s 2256 42423 2256 42423 4 gnd
port 514 nsew
rlabel metal2 s 1008 44240 1008 44240 4 gnd
port 514 nsew
rlabel metal2 s 2256 41317 2256 41317 4 gnd
port 514 nsew
rlabel metal2 s 1488 42897 1488 42897 4 gnd
port 514 nsew
rlabel metal2 s 2256 42660 2256 42660 4 gnd
port 514 nsew
rlabel metal2 s 2256 44003 2256 44003 4 gnd
port 514 nsew
rlabel metal2 s 240 42660 240 42660 4 gnd
port 514 nsew
rlabel metal2 s 2256 42107 2256 42107 4 gnd
port 514 nsew
rlabel metal2 s 1488 41870 1488 41870 4 gnd
port 514 nsew
rlabel metal2 s 1488 41633 1488 41633 4 gnd
port 514 nsew
rlabel metal2 s 1488 43213 1488 43213 4 gnd
port 514 nsew
rlabel metal2 s 1008 41633 1008 41633 4 gnd
port 514 nsew
rlabel metal2 s 240 41870 240 41870 4 gnd
port 514 nsew
rlabel metal2 s 240 44240 240 44240 4 gnd
port 514 nsew
rlabel metal2 s 1488 43687 1488 43687 4 gnd
port 514 nsew
rlabel metal2 s 240 41633 240 41633 4 gnd
port 514 nsew
rlabel metal2 s 1008 43213 1008 43213 4 gnd
port 514 nsew
rlabel metal2 s 1008 41317 1008 41317 4 gnd
port 514 nsew
rlabel metal2 s 240 44003 240 44003 4 gnd
port 514 nsew
rlabel metal2 s 1008 42897 1008 42897 4 gnd
port 514 nsew
rlabel metal2 s 240 42423 240 42423 4 gnd
port 514 nsew
rlabel metal2 s 2256 42897 2256 42897 4 gnd
port 514 nsew
rlabel metal2 s 1488 42423 1488 42423 4 gnd
port 514 nsew
rlabel metal2 s 2256 43450 2256 43450 4 gnd
port 514 nsew
rlabel metal2 s 240 43213 240 43213 4 gnd
port 514 nsew
rlabel metal2 s 1008 42107 1008 42107 4 gnd
port 514 nsew
rlabel metal2 s 240 43450 240 43450 4 gnd
port 514 nsew
rlabel metal2 s 1008 44003 1008 44003 4 gnd
port 514 nsew
rlabel metal2 s 1488 44003 1488 44003 4 gnd
port 514 nsew
rlabel metal2 s 240 42897 240 42897 4 gnd
port 514 nsew
rlabel metal2 s 1488 42660 1488 42660 4 gnd
port 514 nsew
rlabel metal2 s 240 41317 240 41317 4 gnd
port 514 nsew
rlabel metal2 s 1488 42107 1488 42107 4 gnd
port 514 nsew
rlabel metal2 s 240 42107 240 42107 4 gnd
port 514 nsew
rlabel metal2 s 1488 43450 1488 43450 4 gnd
port 514 nsew
rlabel metal2 s 2256 43687 2256 43687 4 gnd
port 514 nsew
rlabel metal2 s 240 43687 240 43687 4 gnd
port 514 nsew
rlabel metal2 s 2256 41633 2256 41633 4 gnd
port 514 nsew
rlabel metal2 s 1488 39500 1488 39500 4 gnd
port 514 nsew
rlabel metal2 s 1488 38473 1488 38473 4 gnd
port 514 nsew
rlabel metal2 s 240 40527 240 40527 4 gnd
port 514 nsew
rlabel metal2 s 240 38473 240 38473 4 gnd
port 514 nsew
rlabel metal2 s 2256 40053 2256 40053 4 gnd
port 514 nsew
rlabel metal2 s 1008 40053 1008 40053 4 gnd
port 514 nsew
rlabel metal2 s 2256 41080 2256 41080 4 gnd
port 514 nsew
rlabel metal2 s 1488 38947 1488 38947 4 gnd
port 514 nsew
rlabel metal2 s 1488 41080 1488 41080 4 gnd
port 514 nsew
rlabel metal2 s 1008 38157 1008 38157 4 gnd
port 514 nsew
rlabel metal2 s 1008 40290 1008 40290 4 gnd
port 514 nsew
rlabel metal2 s 2256 40527 2256 40527 4 gnd
port 514 nsew
rlabel metal2 s 1488 39737 1488 39737 4 gnd
port 514 nsew
rlabel metal2 s 1008 39500 1008 39500 4 gnd
port 514 nsew
rlabel metal2 s 1488 40843 1488 40843 4 gnd
port 514 nsew
rlabel metal2 s 240 39500 240 39500 4 gnd
port 514 nsew
rlabel metal2 s 1008 41080 1008 41080 4 gnd
port 514 nsew
rlabel metal2 s 2256 38710 2256 38710 4 gnd
port 514 nsew
rlabel metal2 s 1008 38710 1008 38710 4 gnd
port 514 nsew
rlabel metal2 s 1488 38710 1488 38710 4 gnd
port 514 nsew
rlabel metal2 s 1488 39263 1488 39263 4 gnd
port 514 nsew
rlabel metal2 s 240 39263 240 39263 4 gnd
port 514 nsew
rlabel metal2 s 2256 38157 2256 38157 4 gnd
port 514 nsew
rlabel metal2 s 240 40053 240 40053 4 gnd
port 514 nsew
rlabel metal2 s 1008 38947 1008 38947 4 gnd
port 514 nsew
rlabel metal2 s 1008 39737 1008 39737 4 gnd
port 514 nsew
rlabel metal2 s 1008 39263 1008 39263 4 gnd
port 514 nsew
rlabel metal2 s 1488 40527 1488 40527 4 gnd
port 514 nsew
rlabel metal2 s 2256 40843 2256 40843 4 gnd
port 514 nsew
rlabel metal2 s 240 40290 240 40290 4 gnd
port 514 nsew
rlabel metal2 s 240 38710 240 38710 4 gnd
port 514 nsew
rlabel metal2 s 240 40843 240 40843 4 gnd
port 514 nsew
rlabel metal2 s 1488 40290 1488 40290 4 gnd
port 514 nsew
rlabel metal2 s 1008 38473 1008 38473 4 gnd
port 514 nsew
rlabel metal2 s 2256 39500 2256 39500 4 gnd
port 514 nsew
rlabel metal2 s 2256 40290 2256 40290 4 gnd
port 514 nsew
rlabel metal2 s 2256 39263 2256 39263 4 gnd
port 514 nsew
rlabel metal2 s 240 39737 240 39737 4 gnd
port 514 nsew
rlabel metal2 s 1488 38157 1488 38157 4 gnd
port 514 nsew
rlabel metal2 s 240 41080 240 41080 4 gnd
port 514 nsew
rlabel metal2 s 1008 40527 1008 40527 4 gnd
port 514 nsew
rlabel metal2 s 240 38157 240 38157 4 gnd
port 514 nsew
rlabel metal2 s 1488 40053 1488 40053 4 gnd
port 514 nsew
rlabel metal2 s 1008 40843 1008 40843 4 gnd
port 514 nsew
rlabel metal2 s 240 38947 240 38947 4 gnd
port 514 nsew
rlabel metal2 s 2256 38473 2256 38473 4 gnd
port 514 nsew
rlabel metal2 s 2256 39737 2256 39737 4 gnd
port 514 nsew
rlabel metal2 s 2256 38947 2256 38947 4 gnd
port 514 nsew
rlabel metal2 s 2736 40053 2736 40053 4 gnd
port 514 nsew
rlabel metal2 s 3504 38157 3504 38157 4 gnd
port 514 nsew
rlabel metal2 s 3504 40053 3504 40053 4 gnd
port 514 nsew
rlabel metal2 s 2736 38947 2736 38947 4 gnd
port 514 nsew
rlabel metal2 s 4752 40843 4752 40843 4 gnd
port 514 nsew
rlabel metal2 s 3504 38947 3504 38947 4 gnd
port 514 nsew
rlabel metal2 s 3984 38710 3984 38710 4 gnd
port 514 nsew
rlabel metal2 s 2736 40290 2736 40290 4 gnd
port 514 nsew
rlabel metal2 s 2736 39263 2736 39263 4 gnd
port 514 nsew
rlabel metal2 s 3984 40053 3984 40053 4 gnd
port 514 nsew
rlabel metal2 s 2736 40527 2736 40527 4 gnd
port 514 nsew
rlabel metal2 s 2736 40843 2736 40843 4 gnd
port 514 nsew
rlabel metal2 s 3984 39263 3984 39263 4 gnd
port 514 nsew
rlabel metal2 s 4752 38473 4752 38473 4 gnd
port 514 nsew
rlabel metal2 s 3984 40527 3984 40527 4 gnd
port 514 nsew
rlabel metal2 s 3504 39263 3504 39263 4 gnd
port 514 nsew
rlabel metal2 s 4752 38710 4752 38710 4 gnd
port 514 nsew
rlabel metal2 s 4752 39737 4752 39737 4 gnd
port 514 nsew
rlabel metal2 s 3984 39500 3984 39500 4 gnd
port 514 nsew
rlabel metal2 s 3504 40843 3504 40843 4 gnd
port 514 nsew
rlabel metal2 s 2736 39500 2736 39500 4 gnd
port 514 nsew
rlabel metal2 s 3984 38947 3984 38947 4 gnd
port 514 nsew
rlabel metal2 s 3984 39737 3984 39737 4 gnd
port 514 nsew
rlabel metal2 s 4752 38157 4752 38157 4 gnd
port 514 nsew
rlabel metal2 s 3504 38473 3504 38473 4 gnd
port 514 nsew
rlabel metal2 s 3984 38473 3984 38473 4 gnd
port 514 nsew
rlabel metal2 s 3504 39500 3504 39500 4 gnd
port 514 nsew
rlabel metal2 s 2736 38157 2736 38157 4 gnd
port 514 nsew
rlabel metal2 s 3984 41080 3984 41080 4 gnd
port 514 nsew
rlabel metal2 s 2736 38710 2736 38710 4 gnd
port 514 nsew
rlabel metal2 s 4752 38947 4752 38947 4 gnd
port 514 nsew
rlabel metal2 s 3984 38157 3984 38157 4 gnd
port 514 nsew
rlabel metal2 s 4752 39263 4752 39263 4 gnd
port 514 nsew
rlabel metal2 s 3504 40290 3504 40290 4 gnd
port 514 nsew
rlabel metal2 s 2736 41080 2736 41080 4 gnd
port 514 nsew
rlabel metal2 s 4752 41080 4752 41080 4 gnd
port 514 nsew
rlabel metal2 s 2736 39737 2736 39737 4 gnd
port 514 nsew
rlabel metal2 s 2736 38473 2736 38473 4 gnd
port 514 nsew
rlabel metal2 s 3504 40527 3504 40527 4 gnd
port 514 nsew
rlabel metal2 s 3504 39737 3504 39737 4 gnd
port 514 nsew
rlabel metal2 s 4752 40527 4752 40527 4 gnd
port 514 nsew
rlabel metal2 s 3984 40290 3984 40290 4 gnd
port 514 nsew
rlabel metal2 s 4752 39500 4752 39500 4 gnd
port 514 nsew
rlabel metal2 s 3504 41080 3504 41080 4 gnd
port 514 nsew
rlabel metal2 s 3984 40843 3984 40843 4 gnd
port 514 nsew
rlabel metal2 s 3504 38710 3504 38710 4 gnd
port 514 nsew
rlabel metal2 s 4752 40290 4752 40290 4 gnd
port 514 nsew
rlabel metal2 s 4752 40053 4752 40053 4 gnd
port 514 nsew
rlabel metal2 s 9744 42897 9744 42897 4 gnd
port 514 nsew
rlabel metal2 s 8976 42660 8976 42660 4 gnd
port 514 nsew
rlabel metal2 s 9744 42107 9744 42107 4 gnd
port 514 nsew
rlabel metal2 s 9744 41870 9744 41870 4 gnd
port 514 nsew
rlabel metal2 s 8976 41870 8976 41870 4 gnd
port 514 nsew
rlabel metal2 s 7728 42897 7728 42897 4 gnd
port 514 nsew
rlabel metal2 s 9744 44240 9744 44240 4 gnd
port 514 nsew
rlabel metal2 s 9744 44003 9744 44003 4 gnd
port 514 nsew
rlabel metal2 s 9744 42423 9744 42423 4 gnd
port 514 nsew
rlabel metal2 s 7728 41870 7728 41870 4 gnd
port 514 nsew
rlabel metal2 s 8496 41870 8496 41870 4 gnd
port 514 nsew
rlabel metal2 s 8976 44240 8976 44240 4 gnd
port 514 nsew
rlabel metal2 s 8496 41633 8496 41633 4 gnd
port 514 nsew
rlabel metal2 s 8496 43687 8496 43687 4 gnd
port 514 nsew
rlabel metal2 s 8976 43450 8976 43450 4 gnd
port 514 nsew
rlabel metal2 s 7728 42660 7728 42660 4 gnd
port 514 nsew
rlabel metal2 s 7728 43213 7728 43213 4 gnd
port 514 nsew
rlabel metal2 s 8496 42423 8496 42423 4 gnd
port 514 nsew
rlabel metal2 s 8976 44003 8976 44003 4 gnd
port 514 nsew
rlabel metal2 s 9744 42660 9744 42660 4 gnd
port 514 nsew
rlabel metal2 s 8496 42897 8496 42897 4 gnd
port 514 nsew
rlabel metal2 s 8976 41317 8976 41317 4 gnd
port 514 nsew
rlabel metal2 s 8976 43213 8976 43213 4 gnd
port 514 nsew
rlabel metal2 s 8976 42107 8976 42107 4 gnd
port 514 nsew
rlabel metal2 s 7728 44240 7728 44240 4 gnd
port 514 nsew
rlabel metal2 s 7728 44003 7728 44003 4 gnd
port 514 nsew
rlabel metal2 s 7728 42107 7728 42107 4 gnd
port 514 nsew
rlabel metal2 s 7728 41633 7728 41633 4 gnd
port 514 nsew
rlabel metal2 s 9744 43687 9744 43687 4 gnd
port 514 nsew
rlabel metal2 s 7728 42423 7728 42423 4 gnd
port 514 nsew
rlabel metal2 s 9744 43213 9744 43213 4 gnd
port 514 nsew
rlabel metal2 s 8976 42423 8976 42423 4 gnd
port 514 nsew
rlabel metal2 s 8496 43450 8496 43450 4 gnd
port 514 nsew
rlabel metal2 s 9744 41317 9744 41317 4 gnd
port 514 nsew
rlabel metal2 s 7728 41317 7728 41317 4 gnd
port 514 nsew
rlabel metal2 s 8496 42660 8496 42660 4 gnd
port 514 nsew
rlabel metal2 s 9744 41633 9744 41633 4 gnd
port 514 nsew
rlabel metal2 s 8976 41633 8976 41633 4 gnd
port 514 nsew
rlabel metal2 s 8496 44240 8496 44240 4 gnd
port 514 nsew
rlabel metal2 s 8496 43213 8496 43213 4 gnd
port 514 nsew
rlabel metal2 s 7728 43687 7728 43687 4 gnd
port 514 nsew
rlabel metal2 s 7728 43450 7728 43450 4 gnd
port 514 nsew
rlabel metal2 s 8496 41317 8496 41317 4 gnd
port 514 nsew
rlabel metal2 s 9744 43450 9744 43450 4 gnd
port 514 nsew
rlabel metal2 s 8976 43687 8976 43687 4 gnd
port 514 nsew
rlabel metal2 s 8496 42107 8496 42107 4 gnd
port 514 nsew
rlabel metal2 s 8976 42897 8976 42897 4 gnd
port 514 nsew
rlabel metal2 s 8496 44003 8496 44003 4 gnd
port 514 nsew
rlabel metal2 s 6480 42660 6480 42660 4 gnd
port 514 nsew
rlabel metal2 s 5232 42423 5232 42423 4 gnd
port 514 nsew
rlabel metal2 s 7248 41633 7248 41633 4 gnd
port 514 nsew
rlabel metal2 s 7248 42660 7248 42660 4 gnd
port 514 nsew
rlabel metal2 s 7248 42423 7248 42423 4 gnd
port 514 nsew
rlabel metal2 s 5232 42897 5232 42897 4 gnd
port 514 nsew
rlabel metal2 s 6000 42423 6000 42423 4 gnd
port 514 nsew
rlabel metal2 s 6000 41633 6000 41633 4 gnd
port 514 nsew
rlabel metal2 s 6000 41870 6000 41870 4 gnd
port 514 nsew
rlabel metal2 s 7248 42107 7248 42107 4 gnd
port 514 nsew
rlabel metal2 s 6480 44003 6480 44003 4 gnd
port 514 nsew
rlabel metal2 s 7248 41870 7248 41870 4 gnd
port 514 nsew
rlabel metal2 s 6000 42897 6000 42897 4 gnd
port 514 nsew
rlabel metal2 s 5232 43213 5232 43213 4 gnd
port 514 nsew
rlabel metal2 s 7248 43213 7248 43213 4 gnd
port 514 nsew
rlabel metal2 s 6480 44240 6480 44240 4 gnd
port 514 nsew
rlabel metal2 s 6000 43687 6000 43687 4 gnd
port 514 nsew
rlabel metal2 s 7248 44003 7248 44003 4 gnd
port 514 nsew
rlabel metal2 s 5232 44240 5232 44240 4 gnd
port 514 nsew
rlabel metal2 s 6000 44003 6000 44003 4 gnd
port 514 nsew
rlabel metal2 s 7248 43687 7248 43687 4 gnd
port 514 nsew
rlabel metal2 s 7248 44240 7248 44240 4 gnd
port 514 nsew
rlabel metal2 s 5232 42660 5232 42660 4 gnd
port 514 nsew
rlabel metal2 s 6480 43450 6480 43450 4 gnd
port 514 nsew
rlabel metal2 s 5232 43687 5232 43687 4 gnd
port 514 nsew
rlabel metal2 s 6480 41633 6480 41633 4 gnd
port 514 nsew
rlabel metal2 s 6000 42107 6000 42107 4 gnd
port 514 nsew
rlabel metal2 s 5232 41317 5232 41317 4 gnd
port 514 nsew
rlabel metal2 s 6480 42107 6480 42107 4 gnd
port 514 nsew
rlabel metal2 s 5232 41633 5232 41633 4 gnd
port 514 nsew
rlabel metal2 s 6000 42660 6000 42660 4 gnd
port 514 nsew
rlabel metal2 s 6480 42423 6480 42423 4 gnd
port 514 nsew
rlabel metal2 s 6480 43213 6480 43213 4 gnd
port 514 nsew
rlabel metal2 s 5232 42107 5232 42107 4 gnd
port 514 nsew
rlabel metal2 s 7248 41317 7248 41317 4 gnd
port 514 nsew
rlabel metal2 s 5232 43450 5232 43450 4 gnd
port 514 nsew
rlabel metal2 s 6000 44240 6000 44240 4 gnd
port 514 nsew
rlabel metal2 s 6480 42897 6480 42897 4 gnd
port 514 nsew
rlabel metal2 s 6000 43213 6000 43213 4 gnd
port 514 nsew
rlabel metal2 s 6000 41317 6000 41317 4 gnd
port 514 nsew
rlabel metal2 s 5232 41870 5232 41870 4 gnd
port 514 nsew
rlabel metal2 s 6000 43450 6000 43450 4 gnd
port 514 nsew
rlabel metal2 s 6480 43687 6480 43687 4 gnd
port 514 nsew
rlabel metal2 s 7248 42897 7248 42897 4 gnd
port 514 nsew
rlabel metal2 s 6480 41870 6480 41870 4 gnd
port 514 nsew
rlabel metal2 s 5232 44003 5232 44003 4 gnd
port 514 nsew
rlabel metal2 s 7248 43450 7248 43450 4 gnd
port 514 nsew
rlabel metal2 s 6480 41317 6480 41317 4 gnd
port 514 nsew
rlabel metal2 s 7248 41080 7248 41080 4 gnd
port 514 nsew
rlabel metal2 s 6000 39737 6000 39737 4 gnd
port 514 nsew
rlabel metal2 s 6000 40053 6000 40053 4 gnd
port 514 nsew
rlabel metal2 s 7248 38473 7248 38473 4 gnd
port 514 nsew
rlabel metal2 s 5232 39263 5232 39263 4 gnd
port 514 nsew
rlabel metal2 s 6480 41080 6480 41080 4 gnd
port 514 nsew
rlabel metal2 s 7248 40527 7248 40527 4 gnd
port 514 nsew
rlabel metal2 s 6480 40527 6480 40527 4 gnd
port 514 nsew
rlabel metal2 s 6000 38947 6000 38947 4 gnd
port 514 nsew
rlabel metal2 s 5232 40843 5232 40843 4 gnd
port 514 nsew
rlabel metal2 s 6000 39500 6000 39500 4 gnd
port 514 nsew
rlabel metal2 s 5232 40053 5232 40053 4 gnd
port 514 nsew
rlabel metal2 s 6480 38473 6480 38473 4 gnd
port 514 nsew
rlabel metal2 s 7248 40290 7248 40290 4 gnd
port 514 nsew
rlabel metal2 s 6000 38157 6000 38157 4 gnd
port 514 nsew
rlabel metal2 s 6480 39500 6480 39500 4 gnd
port 514 nsew
rlabel metal2 s 5232 41080 5232 41080 4 gnd
port 514 nsew
rlabel metal2 s 7248 40843 7248 40843 4 gnd
port 514 nsew
rlabel metal2 s 5232 40290 5232 40290 4 gnd
port 514 nsew
rlabel metal2 s 5232 38157 5232 38157 4 gnd
port 514 nsew
rlabel metal2 s 7248 39263 7248 39263 4 gnd
port 514 nsew
rlabel metal2 s 6000 41080 6000 41080 4 gnd
port 514 nsew
rlabel metal2 s 6480 38157 6480 38157 4 gnd
port 514 nsew
rlabel metal2 s 6000 38710 6000 38710 4 gnd
port 514 nsew
rlabel metal2 s 6480 38947 6480 38947 4 gnd
port 514 nsew
rlabel metal2 s 6480 39263 6480 39263 4 gnd
port 514 nsew
rlabel metal2 s 6000 40527 6000 40527 4 gnd
port 514 nsew
rlabel metal2 s 7248 38947 7248 38947 4 gnd
port 514 nsew
rlabel metal2 s 7248 40053 7248 40053 4 gnd
port 514 nsew
rlabel metal2 s 5232 38473 5232 38473 4 gnd
port 514 nsew
rlabel metal2 s 6480 40290 6480 40290 4 gnd
port 514 nsew
rlabel metal2 s 5232 39500 5232 39500 4 gnd
port 514 nsew
rlabel metal2 s 5232 40527 5232 40527 4 gnd
port 514 nsew
rlabel metal2 s 7248 39500 7248 39500 4 gnd
port 514 nsew
rlabel metal2 s 6480 38710 6480 38710 4 gnd
port 514 nsew
rlabel metal2 s 6000 40843 6000 40843 4 gnd
port 514 nsew
rlabel metal2 s 6000 39263 6000 39263 4 gnd
port 514 nsew
rlabel metal2 s 5232 39737 5232 39737 4 gnd
port 514 nsew
rlabel metal2 s 6000 40290 6000 40290 4 gnd
port 514 nsew
rlabel metal2 s 6480 39737 6480 39737 4 gnd
port 514 nsew
rlabel metal2 s 7248 38157 7248 38157 4 gnd
port 514 nsew
rlabel metal2 s 5232 38710 5232 38710 4 gnd
port 514 nsew
rlabel metal2 s 7248 38710 7248 38710 4 gnd
port 514 nsew
rlabel metal2 s 6480 40843 6480 40843 4 gnd
port 514 nsew
rlabel metal2 s 7248 39737 7248 39737 4 gnd
port 514 nsew
rlabel metal2 s 6480 40053 6480 40053 4 gnd
port 514 nsew
rlabel metal2 s 5232 38947 5232 38947 4 gnd
port 514 nsew
rlabel metal2 s 6000 38473 6000 38473 4 gnd
port 514 nsew
rlabel metal2 s 8976 38473 8976 38473 4 gnd
port 514 nsew
rlabel metal2 s 7728 40053 7728 40053 4 gnd
port 514 nsew
rlabel metal2 s 8496 39500 8496 39500 4 gnd
port 514 nsew
rlabel metal2 s 9744 40843 9744 40843 4 gnd
port 514 nsew
rlabel metal2 s 8976 38710 8976 38710 4 gnd
port 514 nsew
rlabel metal2 s 9744 38710 9744 38710 4 gnd
port 514 nsew
rlabel metal2 s 9744 38157 9744 38157 4 gnd
port 514 nsew
rlabel metal2 s 8496 38947 8496 38947 4 gnd
port 514 nsew
rlabel metal2 s 8496 38473 8496 38473 4 gnd
port 514 nsew
rlabel metal2 s 8496 39263 8496 39263 4 gnd
port 514 nsew
rlabel metal2 s 9744 38473 9744 38473 4 gnd
port 514 nsew
rlabel metal2 s 8496 40053 8496 40053 4 gnd
port 514 nsew
rlabel metal2 s 7728 39500 7728 39500 4 gnd
port 514 nsew
rlabel metal2 s 7728 41080 7728 41080 4 gnd
port 514 nsew
rlabel metal2 s 8976 39737 8976 39737 4 gnd
port 514 nsew
rlabel metal2 s 8496 41080 8496 41080 4 gnd
port 514 nsew
rlabel metal2 s 9744 40527 9744 40527 4 gnd
port 514 nsew
rlabel metal2 s 9744 41080 9744 41080 4 gnd
port 514 nsew
rlabel metal2 s 8976 40527 8976 40527 4 gnd
port 514 nsew
rlabel metal2 s 8496 40527 8496 40527 4 gnd
port 514 nsew
rlabel metal2 s 9744 39737 9744 39737 4 gnd
port 514 nsew
rlabel metal2 s 8976 38947 8976 38947 4 gnd
port 514 nsew
rlabel metal2 s 8496 38157 8496 38157 4 gnd
port 514 nsew
rlabel metal2 s 7728 38157 7728 38157 4 gnd
port 514 nsew
rlabel metal2 s 7728 39737 7728 39737 4 gnd
port 514 nsew
rlabel metal2 s 8496 39737 8496 39737 4 gnd
port 514 nsew
rlabel metal2 s 8976 40843 8976 40843 4 gnd
port 514 nsew
rlabel metal2 s 8976 40053 8976 40053 4 gnd
port 514 nsew
rlabel metal2 s 7728 38473 7728 38473 4 gnd
port 514 nsew
rlabel metal2 s 7728 40290 7728 40290 4 gnd
port 514 nsew
rlabel metal2 s 9744 39500 9744 39500 4 gnd
port 514 nsew
rlabel metal2 s 8976 39500 8976 39500 4 gnd
port 514 nsew
rlabel metal2 s 8496 40290 8496 40290 4 gnd
port 514 nsew
rlabel metal2 s 7728 38947 7728 38947 4 gnd
port 514 nsew
rlabel metal2 s 8496 40843 8496 40843 4 gnd
port 514 nsew
rlabel metal2 s 9744 38947 9744 38947 4 gnd
port 514 nsew
rlabel metal2 s 7728 40527 7728 40527 4 gnd
port 514 nsew
rlabel metal2 s 8976 39263 8976 39263 4 gnd
port 514 nsew
rlabel metal2 s 8976 41080 8976 41080 4 gnd
port 514 nsew
rlabel metal2 s 9744 39263 9744 39263 4 gnd
port 514 nsew
rlabel metal2 s 8976 38157 8976 38157 4 gnd
port 514 nsew
rlabel metal2 s 8976 40290 8976 40290 4 gnd
port 514 nsew
rlabel metal2 s 7728 38710 7728 38710 4 gnd
port 514 nsew
rlabel metal2 s 9744 40290 9744 40290 4 gnd
port 514 nsew
rlabel metal2 s 7728 40843 7728 40843 4 gnd
port 514 nsew
rlabel metal2 s 8496 38710 8496 38710 4 gnd
port 514 nsew
rlabel metal2 s 9744 40053 9744 40053 4 gnd
port 514 nsew
rlabel metal2 s 7728 39263 7728 39263 4 gnd
port 514 nsew
rlabel metal2 s 9744 36893 9744 36893 4 gnd
port 514 nsew
rlabel metal2 s 7728 36103 7728 36103 4 gnd
port 514 nsew
rlabel metal2 s 8976 37130 8976 37130 4 gnd
port 514 nsew
rlabel metal2 s 9744 36340 9744 36340 4 gnd
port 514 nsew
rlabel metal2 s 7728 37920 7728 37920 4 gnd
port 514 nsew
rlabel metal2 s 7728 36577 7728 36577 4 gnd
port 514 nsew
rlabel metal2 s 8976 36577 8976 36577 4 gnd
port 514 nsew
rlabel metal2 s 9744 35787 9744 35787 4 gnd
port 514 nsew
rlabel metal2 s 8976 37683 8976 37683 4 gnd
port 514 nsew
rlabel metal2 s 8496 37130 8496 37130 4 gnd
port 514 nsew
rlabel metal2 s 8496 36103 8496 36103 4 gnd
port 514 nsew
rlabel metal2 s 9744 37367 9744 37367 4 gnd
port 514 nsew
rlabel metal2 s 9744 36577 9744 36577 4 gnd
port 514 nsew
rlabel metal2 s 8496 35313 8496 35313 4 gnd
port 514 nsew
rlabel metal2 s 8496 36577 8496 36577 4 gnd
port 514 nsew
rlabel metal2 s 8976 37367 8976 37367 4 gnd
port 514 nsew
rlabel metal2 s 9744 35313 9744 35313 4 gnd
port 514 nsew
rlabel metal2 s 8976 35313 8976 35313 4 gnd
port 514 nsew
rlabel metal2 s 8976 35550 8976 35550 4 gnd
port 514 nsew
rlabel metal2 s 9744 37920 9744 37920 4 gnd
port 514 nsew
rlabel metal2 s 8496 36893 8496 36893 4 gnd
port 514 nsew
rlabel metal2 s 7728 36893 7728 36893 4 gnd
port 514 nsew
rlabel metal2 s 7728 37683 7728 37683 4 gnd
port 514 nsew
rlabel metal2 s 8496 37367 8496 37367 4 gnd
port 514 nsew
rlabel metal2 s 7728 34997 7728 34997 4 gnd
port 514 nsew
rlabel metal2 s 8976 36893 8976 36893 4 gnd
port 514 nsew
rlabel metal2 s 9744 37130 9744 37130 4 gnd
port 514 nsew
rlabel metal2 s 9744 34997 9744 34997 4 gnd
port 514 nsew
rlabel metal2 s 7728 37130 7728 37130 4 gnd
port 514 nsew
rlabel metal2 s 8496 35550 8496 35550 4 gnd
port 514 nsew
rlabel metal2 s 9744 35550 9744 35550 4 gnd
port 514 nsew
rlabel metal2 s 8496 34997 8496 34997 4 gnd
port 514 nsew
rlabel metal2 s 7728 35313 7728 35313 4 gnd
port 514 nsew
rlabel metal2 s 8976 36340 8976 36340 4 gnd
port 514 nsew
rlabel metal2 s 8496 35787 8496 35787 4 gnd
port 514 nsew
rlabel metal2 s 8976 37920 8976 37920 4 gnd
port 514 nsew
rlabel metal2 s 7728 35550 7728 35550 4 gnd
port 514 nsew
rlabel metal2 s 9744 37683 9744 37683 4 gnd
port 514 nsew
rlabel metal2 s 8976 36103 8976 36103 4 gnd
port 514 nsew
rlabel metal2 s 8976 35787 8976 35787 4 gnd
port 514 nsew
rlabel metal2 s 8496 37683 8496 37683 4 gnd
port 514 nsew
rlabel metal2 s 7728 35787 7728 35787 4 gnd
port 514 nsew
rlabel metal2 s 7728 37367 7728 37367 4 gnd
port 514 nsew
rlabel metal2 s 8496 37920 8496 37920 4 gnd
port 514 nsew
rlabel metal2 s 8496 36340 8496 36340 4 gnd
port 514 nsew
rlabel metal2 s 7728 36340 7728 36340 4 gnd
port 514 nsew
rlabel metal2 s 9744 36103 9744 36103 4 gnd
port 514 nsew
rlabel metal2 s 8976 34997 8976 34997 4 gnd
port 514 nsew
rlabel metal2 s 5232 36340 5232 36340 4 gnd
port 514 nsew
rlabel metal2 s 5232 37130 5232 37130 4 gnd
port 514 nsew
rlabel metal2 s 6000 36340 6000 36340 4 gnd
port 514 nsew
rlabel metal2 s 6000 35313 6000 35313 4 gnd
port 514 nsew
rlabel metal2 s 7248 36103 7248 36103 4 gnd
port 514 nsew
rlabel metal2 s 7248 37683 7248 37683 4 gnd
port 514 nsew
rlabel metal2 s 5232 36577 5232 36577 4 gnd
port 514 nsew
rlabel metal2 s 7248 37367 7248 37367 4 gnd
port 514 nsew
rlabel metal2 s 5232 36103 5232 36103 4 gnd
port 514 nsew
rlabel metal2 s 5232 37367 5232 37367 4 gnd
port 514 nsew
rlabel metal2 s 6000 36893 6000 36893 4 gnd
port 514 nsew
rlabel metal2 s 6480 35787 6480 35787 4 gnd
port 514 nsew
rlabel metal2 s 7248 34997 7248 34997 4 gnd
port 514 nsew
rlabel metal2 s 6480 37367 6480 37367 4 gnd
port 514 nsew
rlabel metal2 s 7248 36893 7248 36893 4 gnd
port 514 nsew
rlabel metal2 s 5232 35787 5232 35787 4 gnd
port 514 nsew
rlabel metal2 s 6480 36340 6480 36340 4 gnd
port 514 nsew
rlabel metal2 s 6000 37130 6000 37130 4 gnd
port 514 nsew
rlabel metal2 s 6480 34997 6480 34997 4 gnd
port 514 nsew
rlabel metal2 s 7248 35550 7248 35550 4 gnd
port 514 nsew
rlabel metal2 s 6000 37920 6000 37920 4 gnd
port 514 nsew
rlabel metal2 s 5232 35313 5232 35313 4 gnd
port 514 nsew
rlabel metal2 s 6000 36577 6000 36577 4 gnd
port 514 nsew
rlabel metal2 s 7248 35313 7248 35313 4 gnd
port 514 nsew
rlabel metal2 s 6480 36103 6480 36103 4 gnd
port 514 nsew
rlabel metal2 s 6480 36577 6480 36577 4 gnd
port 514 nsew
rlabel metal2 s 7248 36577 7248 36577 4 gnd
port 514 nsew
rlabel metal2 s 6480 37920 6480 37920 4 gnd
port 514 nsew
rlabel metal2 s 5232 34997 5232 34997 4 gnd
port 514 nsew
rlabel metal2 s 7248 35787 7248 35787 4 gnd
port 514 nsew
rlabel metal2 s 6000 36103 6000 36103 4 gnd
port 514 nsew
rlabel metal2 s 5232 37683 5232 37683 4 gnd
port 514 nsew
rlabel metal2 s 6000 37683 6000 37683 4 gnd
port 514 nsew
rlabel metal2 s 6480 35313 6480 35313 4 gnd
port 514 nsew
rlabel metal2 s 6480 36893 6480 36893 4 gnd
port 514 nsew
rlabel metal2 s 6000 37367 6000 37367 4 gnd
port 514 nsew
rlabel metal2 s 6480 37683 6480 37683 4 gnd
port 514 nsew
rlabel metal2 s 5232 35550 5232 35550 4 gnd
port 514 nsew
rlabel metal2 s 6480 35550 6480 35550 4 gnd
port 514 nsew
rlabel metal2 s 7248 37130 7248 37130 4 gnd
port 514 nsew
rlabel metal2 s 6000 35787 6000 35787 4 gnd
port 514 nsew
rlabel metal2 s 6000 35550 6000 35550 4 gnd
port 514 nsew
rlabel metal2 s 6480 37130 6480 37130 4 gnd
port 514 nsew
rlabel metal2 s 7248 36340 7248 36340 4 gnd
port 514 nsew
rlabel metal2 s 6000 34997 6000 34997 4 gnd
port 514 nsew
rlabel metal2 s 5232 37920 5232 37920 4 gnd
port 514 nsew
rlabel metal2 s 7248 37920 7248 37920 4 gnd
port 514 nsew
rlabel metal2 s 5232 36893 5232 36893 4 gnd
port 514 nsew
rlabel metal2 s 5232 31837 5232 31837 4 gnd
port 514 nsew
rlabel metal2 s 6480 33733 6480 33733 4 gnd
port 514 nsew
rlabel metal2 s 6000 33970 6000 33970 4 gnd
port 514 nsew
rlabel metal2 s 6480 32390 6480 32390 4 gnd
port 514 nsew
rlabel metal2 s 6000 33733 6000 33733 4 gnd
port 514 nsew
rlabel metal2 s 6000 34207 6000 34207 4 gnd
port 514 nsew
rlabel metal2 s 7248 34207 7248 34207 4 gnd
port 514 nsew
rlabel metal2 s 7248 32627 7248 32627 4 gnd
port 514 nsew
rlabel metal2 s 6480 32943 6480 32943 4 gnd
port 514 nsew
rlabel metal2 s 5232 32390 5232 32390 4 gnd
port 514 nsew
rlabel metal2 s 6480 33180 6480 33180 4 gnd
port 514 nsew
rlabel metal2 s 6000 33417 6000 33417 4 gnd
port 514 nsew
rlabel metal2 s 7248 32153 7248 32153 4 gnd
port 514 nsew
rlabel metal2 s 5232 33733 5232 33733 4 gnd
port 514 nsew
rlabel metal2 s 7248 33180 7248 33180 4 gnd
port 514 nsew
rlabel metal2 s 5232 32943 5232 32943 4 gnd
port 514 nsew
rlabel metal2 s 6480 32153 6480 32153 4 gnd
port 514 nsew
rlabel metal2 s 6000 32943 6000 32943 4 gnd
port 514 nsew
rlabel metal2 s 5232 32627 5232 32627 4 gnd
port 514 nsew
rlabel metal2 s 6480 34207 6480 34207 4 gnd
port 514 nsew
rlabel metal2 s 5232 34523 5232 34523 4 gnd
port 514 nsew
rlabel metal2 s 6480 34760 6480 34760 4 gnd
port 514 nsew
rlabel metal2 s 5232 33180 5232 33180 4 gnd
port 514 nsew
rlabel metal2 s 5232 34207 5232 34207 4 gnd
port 514 nsew
rlabel metal2 s 7248 34760 7248 34760 4 gnd
port 514 nsew
rlabel metal2 s 6480 33417 6480 33417 4 gnd
port 514 nsew
rlabel metal2 s 5232 33970 5232 33970 4 gnd
port 514 nsew
rlabel metal2 s 7248 33970 7248 33970 4 gnd
port 514 nsew
rlabel metal2 s 7248 31837 7248 31837 4 gnd
port 514 nsew
rlabel metal2 s 7248 32390 7248 32390 4 gnd
port 514 nsew
rlabel metal2 s 6000 34523 6000 34523 4 gnd
port 514 nsew
rlabel metal2 s 6000 32153 6000 32153 4 gnd
port 514 nsew
rlabel metal2 s 7248 32943 7248 32943 4 gnd
port 514 nsew
rlabel metal2 s 6000 33180 6000 33180 4 gnd
port 514 nsew
rlabel metal2 s 7248 34523 7248 34523 4 gnd
port 514 nsew
rlabel metal2 s 6480 32627 6480 32627 4 gnd
port 514 nsew
rlabel metal2 s 6480 31837 6480 31837 4 gnd
port 514 nsew
rlabel metal2 s 6000 32627 6000 32627 4 gnd
port 514 nsew
rlabel metal2 s 5232 34760 5232 34760 4 gnd
port 514 nsew
rlabel metal2 s 5232 33417 5232 33417 4 gnd
port 514 nsew
rlabel metal2 s 6000 34760 6000 34760 4 gnd
port 514 nsew
rlabel metal2 s 6000 31837 6000 31837 4 gnd
port 514 nsew
rlabel metal2 s 7248 33417 7248 33417 4 gnd
port 514 nsew
rlabel metal2 s 6480 34523 6480 34523 4 gnd
port 514 nsew
rlabel metal2 s 6480 33970 6480 33970 4 gnd
port 514 nsew
rlabel metal2 s 7248 33733 7248 33733 4 gnd
port 514 nsew
rlabel metal2 s 6000 32390 6000 32390 4 gnd
port 514 nsew
rlabel metal2 s 5232 32153 5232 32153 4 gnd
port 514 nsew
rlabel metal2 s 7728 32627 7728 32627 4 gnd
port 514 nsew
rlabel metal2 s 8496 34207 8496 34207 4 gnd
port 514 nsew
rlabel metal2 s 9744 34760 9744 34760 4 gnd
port 514 nsew
rlabel metal2 s 8496 32627 8496 32627 4 gnd
port 514 nsew
rlabel metal2 s 8976 33180 8976 33180 4 gnd
port 514 nsew
rlabel metal2 s 7728 32943 7728 32943 4 gnd
port 514 nsew
rlabel metal2 s 8496 34760 8496 34760 4 gnd
port 514 nsew
rlabel metal2 s 8976 33417 8976 33417 4 gnd
port 514 nsew
rlabel metal2 s 8976 34523 8976 34523 4 gnd
port 514 nsew
rlabel metal2 s 8976 34760 8976 34760 4 gnd
port 514 nsew
rlabel metal2 s 9744 33180 9744 33180 4 gnd
port 514 nsew
rlabel metal2 s 9744 32943 9744 32943 4 gnd
port 514 nsew
rlabel metal2 s 9744 31837 9744 31837 4 gnd
port 514 nsew
rlabel metal2 s 8496 32943 8496 32943 4 gnd
port 514 nsew
rlabel metal2 s 8976 34207 8976 34207 4 gnd
port 514 nsew
rlabel metal2 s 8976 32390 8976 32390 4 gnd
port 514 nsew
rlabel metal2 s 9744 33970 9744 33970 4 gnd
port 514 nsew
rlabel metal2 s 8496 32153 8496 32153 4 gnd
port 514 nsew
rlabel metal2 s 7728 33417 7728 33417 4 gnd
port 514 nsew
rlabel metal2 s 7728 32153 7728 32153 4 gnd
port 514 nsew
rlabel metal2 s 8496 33970 8496 33970 4 gnd
port 514 nsew
rlabel metal2 s 9744 33417 9744 33417 4 gnd
port 514 nsew
rlabel metal2 s 8976 33733 8976 33733 4 gnd
port 514 nsew
rlabel metal2 s 8976 32153 8976 32153 4 gnd
port 514 nsew
rlabel metal2 s 7728 33180 7728 33180 4 gnd
port 514 nsew
rlabel metal2 s 7728 34760 7728 34760 4 gnd
port 514 nsew
rlabel metal2 s 9744 34207 9744 34207 4 gnd
port 514 nsew
rlabel metal2 s 8976 32943 8976 32943 4 gnd
port 514 nsew
rlabel metal2 s 7728 33970 7728 33970 4 gnd
port 514 nsew
rlabel metal2 s 8976 31837 8976 31837 4 gnd
port 514 nsew
rlabel metal2 s 9744 33733 9744 33733 4 gnd
port 514 nsew
rlabel metal2 s 8496 33733 8496 33733 4 gnd
port 514 nsew
rlabel metal2 s 7728 32390 7728 32390 4 gnd
port 514 nsew
rlabel metal2 s 7728 34207 7728 34207 4 gnd
port 514 nsew
rlabel metal2 s 9744 32627 9744 32627 4 gnd
port 514 nsew
rlabel metal2 s 8496 32390 8496 32390 4 gnd
port 514 nsew
rlabel metal2 s 9744 32390 9744 32390 4 gnd
port 514 nsew
rlabel metal2 s 8496 34523 8496 34523 4 gnd
port 514 nsew
rlabel metal2 s 8496 33180 8496 33180 4 gnd
port 514 nsew
rlabel metal2 s 7728 31837 7728 31837 4 gnd
port 514 nsew
rlabel metal2 s 8976 32627 8976 32627 4 gnd
port 514 nsew
rlabel metal2 s 9744 32153 9744 32153 4 gnd
port 514 nsew
rlabel metal2 s 9744 34523 9744 34523 4 gnd
port 514 nsew
rlabel metal2 s 7728 34523 7728 34523 4 gnd
port 514 nsew
rlabel metal2 s 8976 33970 8976 33970 4 gnd
port 514 nsew
rlabel metal2 s 8496 33417 8496 33417 4 gnd
port 514 nsew
rlabel metal2 s 8496 31837 8496 31837 4 gnd
port 514 nsew
rlabel metal2 s 7728 33733 7728 33733 4 gnd
port 514 nsew
rlabel metal2 s 3504 35550 3504 35550 4 gnd
port 514 nsew
rlabel metal2 s 4752 37920 4752 37920 4 gnd
port 514 nsew
rlabel metal2 s 3504 36893 3504 36893 4 gnd
port 514 nsew
rlabel metal2 s 4752 37130 4752 37130 4 gnd
port 514 nsew
rlabel metal2 s 2736 35787 2736 35787 4 gnd
port 514 nsew
rlabel metal2 s 3984 37920 3984 37920 4 gnd
port 514 nsew
rlabel metal2 s 3504 36340 3504 36340 4 gnd
port 514 nsew
rlabel metal2 s 2736 37683 2736 37683 4 gnd
port 514 nsew
rlabel metal2 s 3984 34997 3984 34997 4 gnd
port 514 nsew
rlabel metal2 s 3984 35787 3984 35787 4 gnd
port 514 nsew
rlabel metal2 s 4752 36893 4752 36893 4 gnd
port 514 nsew
rlabel metal2 s 3984 36577 3984 36577 4 gnd
port 514 nsew
rlabel metal2 s 4752 36340 4752 36340 4 gnd
port 514 nsew
rlabel metal2 s 2736 35313 2736 35313 4 gnd
port 514 nsew
rlabel metal2 s 3984 37683 3984 37683 4 gnd
port 514 nsew
rlabel metal2 s 3504 35313 3504 35313 4 gnd
port 514 nsew
rlabel metal2 s 2736 36340 2736 36340 4 gnd
port 514 nsew
rlabel metal2 s 3984 37367 3984 37367 4 gnd
port 514 nsew
rlabel metal2 s 3504 37683 3504 37683 4 gnd
port 514 nsew
rlabel metal2 s 3984 36340 3984 36340 4 gnd
port 514 nsew
rlabel metal2 s 3504 36577 3504 36577 4 gnd
port 514 nsew
rlabel metal2 s 4752 35787 4752 35787 4 gnd
port 514 nsew
rlabel metal2 s 3984 37130 3984 37130 4 gnd
port 514 nsew
rlabel metal2 s 2736 37367 2736 37367 4 gnd
port 514 nsew
rlabel metal2 s 4752 34997 4752 34997 4 gnd
port 514 nsew
rlabel metal2 s 4752 35313 4752 35313 4 gnd
port 514 nsew
rlabel metal2 s 2736 36893 2736 36893 4 gnd
port 514 nsew
rlabel metal2 s 4752 37683 4752 37683 4 gnd
port 514 nsew
rlabel metal2 s 2736 35550 2736 35550 4 gnd
port 514 nsew
rlabel metal2 s 3984 36103 3984 36103 4 gnd
port 514 nsew
rlabel metal2 s 3984 36893 3984 36893 4 gnd
port 514 nsew
rlabel metal2 s 4752 35550 4752 35550 4 gnd
port 514 nsew
rlabel metal2 s 3504 37130 3504 37130 4 gnd
port 514 nsew
rlabel metal2 s 3504 36103 3504 36103 4 gnd
port 514 nsew
rlabel metal2 s 2736 34997 2736 34997 4 gnd
port 514 nsew
rlabel metal2 s 3504 34997 3504 34997 4 gnd
port 514 nsew
rlabel metal2 s 2736 36577 2736 36577 4 gnd
port 514 nsew
rlabel metal2 s 3504 35787 3504 35787 4 gnd
port 514 nsew
rlabel metal2 s 2736 36103 2736 36103 4 gnd
port 514 nsew
rlabel metal2 s 4752 36103 4752 36103 4 gnd
port 514 nsew
rlabel metal2 s 4752 36577 4752 36577 4 gnd
port 514 nsew
rlabel metal2 s 3984 35313 3984 35313 4 gnd
port 514 nsew
rlabel metal2 s 4752 37367 4752 37367 4 gnd
port 514 nsew
rlabel metal2 s 3504 37367 3504 37367 4 gnd
port 514 nsew
rlabel metal2 s 3504 37920 3504 37920 4 gnd
port 514 nsew
rlabel metal2 s 2736 37130 2736 37130 4 gnd
port 514 nsew
rlabel metal2 s 2736 37920 2736 37920 4 gnd
port 514 nsew
rlabel metal2 s 3984 35550 3984 35550 4 gnd
port 514 nsew
rlabel metal2 s 2256 36103 2256 36103 4 gnd
port 514 nsew
rlabel metal2 s 1488 37920 1488 37920 4 gnd
port 514 nsew
rlabel metal2 s 2256 36340 2256 36340 4 gnd
port 514 nsew
rlabel metal2 s 1488 35787 1488 35787 4 gnd
port 514 nsew
rlabel metal2 s 1008 36103 1008 36103 4 gnd
port 514 nsew
rlabel metal2 s 2256 36577 2256 36577 4 gnd
port 514 nsew
rlabel metal2 s 1488 36577 1488 36577 4 gnd
port 514 nsew
rlabel metal2 s 1008 36577 1008 36577 4 gnd
port 514 nsew
rlabel metal2 s 1488 36340 1488 36340 4 gnd
port 514 nsew
rlabel metal2 s 2256 37130 2256 37130 4 gnd
port 514 nsew
rlabel metal2 s 1008 35787 1008 35787 4 gnd
port 514 nsew
rlabel metal2 s 1008 36340 1008 36340 4 gnd
port 514 nsew
rlabel metal2 s 2256 35313 2256 35313 4 gnd
port 514 nsew
rlabel metal2 s 240 35787 240 35787 4 gnd
port 514 nsew
rlabel metal2 s 1488 36103 1488 36103 4 gnd
port 514 nsew
rlabel metal2 s 1488 37683 1488 37683 4 gnd
port 514 nsew
rlabel metal2 s 1008 37367 1008 37367 4 gnd
port 514 nsew
rlabel metal2 s 1008 36893 1008 36893 4 gnd
port 514 nsew
rlabel metal2 s 240 37920 240 37920 4 gnd
port 514 nsew
rlabel metal2 s 1008 37683 1008 37683 4 gnd
port 514 nsew
rlabel metal2 s 2256 35787 2256 35787 4 gnd
port 514 nsew
rlabel metal2 s 1008 37920 1008 37920 4 gnd
port 514 nsew
rlabel metal2 s 240 35550 240 35550 4 gnd
port 514 nsew
rlabel metal2 s 240 36340 240 36340 4 gnd
port 514 nsew
rlabel metal2 s 1008 37130 1008 37130 4 gnd
port 514 nsew
rlabel metal2 s 1488 37130 1488 37130 4 gnd
port 514 nsew
rlabel metal2 s 1008 35313 1008 35313 4 gnd
port 514 nsew
rlabel metal2 s 1488 35550 1488 35550 4 gnd
port 514 nsew
rlabel metal2 s 240 36577 240 36577 4 gnd
port 514 nsew
rlabel metal2 s 1488 35313 1488 35313 4 gnd
port 514 nsew
rlabel metal2 s 240 36103 240 36103 4 gnd
port 514 nsew
rlabel metal2 s 2256 37683 2256 37683 4 gnd
port 514 nsew
rlabel metal2 s 1008 34997 1008 34997 4 gnd
port 514 nsew
rlabel metal2 s 1488 36893 1488 36893 4 gnd
port 514 nsew
rlabel metal2 s 2256 37920 2256 37920 4 gnd
port 514 nsew
rlabel metal2 s 240 36893 240 36893 4 gnd
port 514 nsew
rlabel metal2 s 1488 37367 1488 37367 4 gnd
port 514 nsew
rlabel metal2 s 2256 35550 2256 35550 4 gnd
port 514 nsew
rlabel metal2 s 2256 34997 2256 34997 4 gnd
port 514 nsew
rlabel metal2 s 1488 34997 1488 34997 4 gnd
port 514 nsew
rlabel metal2 s 1008 35550 1008 35550 4 gnd
port 514 nsew
rlabel metal2 s 240 37367 240 37367 4 gnd
port 514 nsew
rlabel metal2 s 2256 36893 2256 36893 4 gnd
port 514 nsew
rlabel metal2 s 240 37683 240 37683 4 gnd
port 514 nsew
rlabel metal2 s 240 35313 240 35313 4 gnd
port 514 nsew
rlabel metal2 s 240 37130 240 37130 4 gnd
port 514 nsew
rlabel metal2 s 240 34997 240 34997 4 gnd
port 514 nsew
rlabel metal2 s 2256 37367 2256 37367 4 gnd
port 514 nsew
rlabel metal2 s 2256 31837 2256 31837 4 gnd
port 514 nsew
rlabel metal2 s 2256 33180 2256 33180 4 gnd
port 514 nsew
rlabel metal2 s 1488 33180 1488 33180 4 gnd
port 514 nsew
rlabel metal2 s 240 33733 240 33733 4 gnd
port 514 nsew
rlabel metal2 s 1488 32390 1488 32390 4 gnd
port 514 nsew
rlabel metal2 s 2256 34760 2256 34760 4 gnd
port 514 nsew
rlabel metal2 s 1008 34207 1008 34207 4 gnd
port 514 nsew
rlabel metal2 s 1488 34207 1488 34207 4 gnd
port 514 nsew
rlabel metal2 s 2256 34207 2256 34207 4 gnd
port 514 nsew
rlabel metal2 s 1008 33733 1008 33733 4 gnd
port 514 nsew
rlabel metal2 s 240 34207 240 34207 4 gnd
port 514 nsew
rlabel metal2 s 1488 31837 1488 31837 4 gnd
port 514 nsew
rlabel metal2 s 1488 32943 1488 32943 4 gnd
port 514 nsew
rlabel metal2 s 2256 33970 2256 33970 4 gnd
port 514 nsew
rlabel metal2 s 1008 32390 1008 32390 4 gnd
port 514 nsew
rlabel metal2 s 2256 34523 2256 34523 4 gnd
port 514 nsew
rlabel metal2 s 1008 33970 1008 33970 4 gnd
port 514 nsew
rlabel metal2 s 2256 33733 2256 33733 4 gnd
port 514 nsew
rlabel metal2 s 1488 33970 1488 33970 4 gnd
port 514 nsew
rlabel metal2 s 1488 33417 1488 33417 4 gnd
port 514 nsew
rlabel metal2 s 1488 32627 1488 32627 4 gnd
port 514 nsew
rlabel metal2 s 240 31837 240 31837 4 gnd
port 514 nsew
rlabel metal2 s 240 32943 240 32943 4 gnd
port 514 nsew
rlabel metal2 s 1008 31837 1008 31837 4 gnd
port 514 nsew
rlabel metal2 s 240 34523 240 34523 4 gnd
port 514 nsew
rlabel metal2 s 240 33180 240 33180 4 gnd
port 514 nsew
rlabel metal2 s 240 33970 240 33970 4 gnd
port 514 nsew
rlabel metal2 s 2256 33417 2256 33417 4 gnd
port 514 nsew
rlabel metal2 s 1008 32153 1008 32153 4 gnd
port 514 nsew
rlabel metal2 s 240 32390 240 32390 4 gnd
port 514 nsew
rlabel metal2 s 1008 33417 1008 33417 4 gnd
port 514 nsew
rlabel metal2 s 240 33417 240 33417 4 gnd
port 514 nsew
rlabel metal2 s 1488 34523 1488 34523 4 gnd
port 514 nsew
rlabel metal2 s 1488 33733 1488 33733 4 gnd
port 514 nsew
rlabel metal2 s 1008 32627 1008 32627 4 gnd
port 514 nsew
rlabel metal2 s 2256 32627 2256 32627 4 gnd
port 514 nsew
rlabel metal2 s 2256 32390 2256 32390 4 gnd
port 514 nsew
rlabel metal2 s 1488 32153 1488 32153 4 gnd
port 514 nsew
rlabel metal2 s 1008 33180 1008 33180 4 gnd
port 514 nsew
rlabel metal2 s 1008 34523 1008 34523 4 gnd
port 514 nsew
rlabel metal2 s 1008 32943 1008 32943 4 gnd
port 514 nsew
rlabel metal2 s 2256 32153 2256 32153 4 gnd
port 514 nsew
rlabel metal2 s 2256 32943 2256 32943 4 gnd
port 514 nsew
rlabel metal2 s 240 32627 240 32627 4 gnd
port 514 nsew
rlabel metal2 s 1008 34760 1008 34760 4 gnd
port 514 nsew
rlabel metal2 s 1488 34760 1488 34760 4 gnd
port 514 nsew
rlabel metal2 s 240 32153 240 32153 4 gnd
port 514 nsew
rlabel metal2 s 240 34760 240 34760 4 gnd
port 514 nsew
rlabel metal2 s 3984 33417 3984 33417 4 gnd
port 514 nsew
rlabel metal2 s 4752 33970 4752 33970 4 gnd
port 514 nsew
rlabel metal2 s 2736 32390 2736 32390 4 gnd
port 514 nsew
rlabel metal2 s 2736 31837 2736 31837 4 gnd
port 514 nsew
rlabel metal2 s 2736 33733 2736 33733 4 gnd
port 514 nsew
rlabel metal2 s 3984 32153 3984 32153 4 gnd
port 514 nsew
rlabel metal2 s 3504 33180 3504 33180 4 gnd
port 514 nsew
rlabel metal2 s 3504 32390 3504 32390 4 gnd
port 514 nsew
rlabel metal2 s 2736 32943 2736 32943 4 gnd
port 514 nsew
rlabel metal2 s 3984 34207 3984 34207 4 gnd
port 514 nsew
rlabel metal2 s 3984 33733 3984 33733 4 gnd
port 514 nsew
rlabel metal2 s 3984 32390 3984 32390 4 gnd
port 514 nsew
rlabel metal2 s 3504 31837 3504 31837 4 gnd
port 514 nsew
rlabel metal2 s 3984 33180 3984 33180 4 gnd
port 514 nsew
rlabel metal2 s 4752 32627 4752 32627 4 gnd
port 514 nsew
rlabel metal2 s 4752 31837 4752 31837 4 gnd
port 514 nsew
rlabel metal2 s 3984 33970 3984 33970 4 gnd
port 514 nsew
rlabel metal2 s 3984 34523 3984 34523 4 gnd
port 514 nsew
rlabel metal2 s 4752 33180 4752 33180 4 gnd
port 514 nsew
rlabel metal2 s 3504 33733 3504 33733 4 gnd
port 514 nsew
rlabel metal2 s 3984 32627 3984 32627 4 gnd
port 514 nsew
rlabel metal2 s 3504 32153 3504 32153 4 gnd
port 514 nsew
rlabel metal2 s 3504 34523 3504 34523 4 gnd
port 514 nsew
rlabel metal2 s 4752 32943 4752 32943 4 gnd
port 514 nsew
rlabel metal2 s 4752 34207 4752 34207 4 gnd
port 514 nsew
rlabel metal2 s 3504 32943 3504 32943 4 gnd
port 514 nsew
rlabel metal2 s 4752 32153 4752 32153 4 gnd
port 514 nsew
rlabel metal2 s 2736 33417 2736 33417 4 gnd
port 514 nsew
rlabel metal2 s 2736 32153 2736 32153 4 gnd
port 514 nsew
rlabel metal2 s 3984 32943 3984 32943 4 gnd
port 514 nsew
rlabel metal2 s 2736 34523 2736 34523 4 gnd
port 514 nsew
rlabel metal2 s 2736 33180 2736 33180 4 gnd
port 514 nsew
rlabel metal2 s 3504 34207 3504 34207 4 gnd
port 514 nsew
rlabel metal2 s 3984 34760 3984 34760 4 gnd
port 514 nsew
rlabel metal2 s 3504 33417 3504 33417 4 gnd
port 514 nsew
rlabel metal2 s 3504 32627 3504 32627 4 gnd
port 514 nsew
rlabel metal2 s 4752 34523 4752 34523 4 gnd
port 514 nsew
rlabel metal2 s 2736 34760 2736 34760 4 gnd
port 514 nsew
rlabel metal2 s 3504 34760 3504 34760 4 gnd
port 514 nsew
rlabel metal2 s 2736 34207 2736 34207 4 gnd
port 514 nsew
rlabel metal2 s 4752 33733 4752 33733 4 gnd
port 514 nsew
rlabel metal2 s 3504 33970 3504 33970 4 gnd
port 514 nsew
rlabel metal2 s 2736 32627 2736 32627 4 gnd
port 514 nsew
rlabel metal2 s 4752 34760 4752 34760 4 gnd
port 514 nsew
rlabel metal2 s 2736 33970 2736 33970 4 gnd
port 514 nsew
rlabel metal2 s 4752 33417 4752 33417 4 gnd
port 514 nsew
rlabel metal2 s 3984 31837 3984 31837 4 gnd
port 514 nsew
rlabel metal2 s 4752 32390 4752 32390 4 gnd
port 514 nsew
rlabel metal2 s 4752 30257 4752 30257 4 gnd
port 514 nsew
rlabel metal2 s 3504 31363 3504 31363 4 gnd
port 514 nsew
rlabel metal2 s 3504 31047 3504 31047 4 gnd
port 514 nsew
rlabel metal2 s 3984 30810 3984 30810 4 gnd
port 514 nsew
rlabel metal2 s 4752 30810 4752 30810 4 gnd
port 514 nsew
rlabel metal2 s 2736 30257 2736 30257 4 gnd
port 514 nsew
rlabel metal2 s 3504 28993 3504 28993 4 gnd
port 514 nsew
rlabel metal2 s 3504 30573 3504 30573 4 gnd
port 514 nsew
rlabel metal2 s 3984 28993 3984 28993 4 gnd
port 514 nsew
rlabel metal2 s 3504 28677 3504 28677 4 gnd
port 514 nsew
rlabel metal2 s 2736 30573 2736 30573 4 gnd
port 514 nsew
rlabel metal2 s 3984 31600 3984 31600 4 gnd
port 514 nsew
rlabel metal2 s 3504 29467 3504 29467 4 gnd
port 514 nsew
rlabel metal2 s 4752 30573 4752 30573 4 gnd
port 514 nsew
rlabel metal2 s 3504 30810 3504 30810 4 gnd
port 514 nsew
rlabel metal2 s 3984 31047 3984 31047 4 gnd
port 514 nsew
rlabel metal2 s 4752 28677 4752 28677 4 gnd
port 514 nsew
rlabel metal2 s 4752 31047 4752 31047 4 gnd
port 514 nsew
rlabel metal2 s 3984 30257 3984 30257 4 gnd
port 514 nsew
rlabel metal2 s 4752 28993 4752 28993 4 gnd
port 514 nsew
rlabel metal2 s 3984 29783 3984 29783 4 gnd
port 514 nsew
rlabel metal2 s 3504 30257 3504 30257 4 gnd
port 514 nsew
rlabel metal2 s 2736 29783 2736 29783 4 gnd
port 514 nsew
rlabel metal2 s 3504 29783 3504 29783 4 gnd
port 514 nsew
rlabel metal2 s 3504 30020 3504 30020 4 gnd
port 514 nsew
rlabel metal2 s 2736 31047 2736 31047 4 gnd
port 514 nsew
rlabel metal2 s 2736 31600 2736 31600 4 gnd
port 514 nsew
rlabel metal2 s 4752 30020 4752 30020 4 gnd
port 514 nsew
rlabel metal2 s 3984 29230 3984 29230 4 gnd
port 514 nsew
rlabel metal2 s 2736 30020 2736 30020 4 gnd
port 514 nsew
rlabel metal2 s 3984 28677 3984 28677 4 gnd
port 514 nsew
rlabel metal2 s 4752 31363 4752 31363 4 gnd
port 514 nsew
rlabel metal2 s 3984 30020 3984 30020 4 gnd
port 514 nsew
rlabel metal2 s 3504 29230 3504 29230 4 gnd
port 514 nsew
rlabel metal2 s 4752 29230 4752 29230 4 gnd
port 514 nsew
rlabel metal2 s 2736 28677 2736 28677 4 gnd
port 514 nsew
rlabel metal2 s 2736 28993 2736 28993 4 gnd
port 514 nsew
rlabel metal2 s 3984 30573 3984 30573 4 gnd
port 514 nsew
rlabel metal2 s 2736 29230 2736 29230 4 gnd
port 514 nsew
rlabel metal2 s 4752 31600 4752 31600 4 gnd
port 514 nsew
rlabel metal2 s 4752 29783 4752 29783 4 gnd
port 514 nsew
rlabel metal2 s 2736 30810 2736 30810 4 gnd
port 514 nsew
rlabel metal2 s 2736 31363 2736 31363 4 gnd
port 514 nsew
rlabel metal2 s 3504 31600 3504 31600 4 gnd
port 514 nsew
rlabel metal2 s 3984 31363 3984 31363 4 gnd
port 514 nsew
rlabel metal2 s 2736 29467 2736 29467 4 gnd
port 514 nsew
rlabel metal2 s 3984 29467 3984 29467 4 gnd
port 514 nsew
rlabel metal2 s 4752 29467 4752 29467 4 gnd
port 514 nsew
rlabel metal2 s 240 31363 240 31363 4 gnd
port 514 nsew
rlabel metal2 s 1008 30573 1008 30573 4 gnd
port 514 nsew
rlabel metal2 s 2256 30020 2256 30020 4 gnd
port 514 nsew
rlabel metal2 s 1008 31363 1008 31363 4 gnd
port 514 nsew
rlabel metal2 s 1008 30020 1008 30020 4 gnd
port 514 nsew
rlabel metal2 s 1488 28993 1488 28993 4 gnd
port 514 nsew
rlabel metal2 s 1008 28993 1008 28993 4 gnd
port 514 nsew
rlabel metal2 s 2256 30810 2256 30810 4 gnd
port 514 nsew
rlabel metal2 s 1488 31047 1488 31047 4 gnd
port 514 nsew
rlabel metal2 s 1008 29467 1008 29467 4 gnd
port 514 nsew
rlabel metal2 s 240 28677 240 28677 4 gnd
port 514 nsew
rlabel metal2 s 2256 31600 2256 31600 4 gnd
port 514 nsew
rlabel metal2 s 1008 29783 1008 29783 4 gnd
port 514 nsew
rlabel metal2 s 240 29467 240 29467 4 gnd
port 514 nsew
rlabel metal2 s 240 29783 240 29783 4 gnd
port 514 nsew
rlabel metal2 s 1008 31047 1008 31047 4 gnd
port 514 nsew
rlabel metal2 s 240 30810 240 30810 4 gnd
port 514 nsew
rlabel metal2 s 240 28993 240 28993 4 gnd
port 514 nsew
rlabel metal2 s 240 30573 240 30573 4 gnd
port 514 nsew
rlabel metal2 s 2256 28993 2256 28993 4 gnd
port 514 nsew
rlabel metal2 s 2256 28677 2256 28677 4 gnd
port 514 nsew
rlabel metal2 s 2256 30257 2256 30257 4 gnd
port 514 nsew
rlabel metal2 s 1488 30020 1488 30020 4 gnd
port 514 nsew
rlabel metal2 s 1008 31600 1008 31600 4 gnd
port 514 nsew
rlabel metal2 s 2256 30573 2256 30573 4 gnd
port 514 nsew
rlabel metal2 s 2256 29230 2256 29230 4 gnd
port 514 nsew
rlabel metal2 s 240 31600 240 31600 4 gnd
port 514 nsew
rlabel metal2 s 1488 29230 1488 29230 4 gnd
port 514 nsew
rlabel metal2 s 240 29230 240 29230 4 gnd
port 514 nsew
rlabel metal2 s 1488 31600 1488 31600 4 gnd
port 514 nsew
rlabel metal2 s 1008 30810 1008 30810 4 gnd
port 514 nsew
rlabel metal2 s 1488 29467 1488 29467 4 gnd
port 514 nsew
rlabel metal2 s 1008 30257 1008 30257 4 gnd
port 514 nsew
rlabel metal2 s 1488 30257 1488 30257 4 gnd
port 514 nsew
rlabel metal2 s 240 30257 240 30257 4 gnd
port 514 nsew
rlabel metal2 s 1488 28677 1488 28677 4 gnd
port 514 nsew
rlabel metal2 s 2256 31363 2256 31363 4 gnd
port 514 nsew
rlabel metal2 s 2256 29467 2256 29467 4 gnd
port 514 nsew
rlabel metal2 s 1008 28677 1008 28677 4 gnd
port 514 nsew
rlabel metal2 s 2256 29783 2256 29783 4 gnd
port 514 nsew
rlabel metal2 s 1008 29230 1008 29230 4 gnd
port 514 nsew
rlabel metal2 s 240 31047 240 31047 4 gnd
port 514 nsew
rlabel metal2 s 1488 30810 1488 30810 4 gnd
port 514 nsew
rlabel metal2 s 240 30020 240 30020 4 gnd
port 514 nsew
rlabel metal2 s 1488 29783 1488 29783 4 gnd
port 514 nsew
rlabel metal2 s 1488 30573 1488 30573 4 gnd
port 514 nsew
rlabel metal2 s 1488 31363 1488 31363 4 gnd
port 514 nsew
rlabel metal2 s 2256 31047 2256 31047 4 gnd
port 514 nsew
rlabel metal2 s 1488 27650 1488 27650 4 gnd
port 514 nsew
rlabel metal2 s 1008 28203 1008 28203 4 gnd
port 514 nsew
rlabel metal2 s 240 27887 240 27887 4 gnd
port 514 nsew
rlabel metal2 s 2256 26307 2256 26307 4 gnd
port 514 nsew
rlabel metal2 s 1488 26307 1488 26307 4 gnd
port 514 nsew
rlabel metal2 s 2256 28440 2256 28440 4 gnd
port 514 nsew
rlabel metal2 s 2256 26070 2256 26070 4 gnd
port 514 nsew
rlabel metal2 s 1488 28440 1488 28440 4 gnd
port 514 nsew
rlabel metal2 s 1008 27650 1008 27650 4 gnd
port 514 nsew
rlabel metal2 s 1008 25517 1008 25517 4 gnd
port 514 nsew
rlabel metal2 s 1008 26070 1008 26070 4 gnd
port 514 nsew
rlabel metal2 s 2256 27097 2256 27097 4 gnd
port 514 nsew
rlabel metal2 s 240 27650 240 27650 4 gnd
port 514 nsew
rlabel metal2 s 1488 26070 1488 26070 4 gnd
port 514 nsew
rlabel metal2 s 1488 27887 1488 27887 4 gnd
port 514 nsew
rlabel metal2 s 240 27413 240 27413 4 gnd
port 514 nsew
rlabel metal2 s 240 26860 240 26860 4 gnd
port 514 nsew
rlabel metal2 s 1488 27413 1488 27413 4 gnd
port 514 nsew
rlabel metal2 s 240 25517 240 25517 4 gnd
port 514 nsew
rlabel metal2 s 2256 25833 2256 25833 4 gnd
port 514 nsew
rlabel metal2 s 2256 26860 2256 26860 4 gnd
port 514 nsew
rlabel metal2 s 1008 27097 1008 27097 4 gnd
port 514 nsew
rlabel metal2 s 1008 25833 1008 25833 4 gnd
port 514 nsew
rlabel metal2 s 1488 26860 1488 26860 4 gnd
port 514 nsew
rlabel metal2 s 2256 28203 2256 28203 4 gnd
port 514 nsew
rlabel metal2 s 240 26070 240 26070 4 gnd
port 514 nsew
rlabel metal2 s 240 27097 240 27097 4 gnd
port 514 nsew
rlabel metal2 s 2256 26623 2256 26623 4 gnd
port 514 nsew
rlabel metal2 s 240 26623 240 26623 4 gnd
port 514 nsew
rlabel metal2 s 240 26307 240 26307 4 gnd
port 514 nsew
rlabel metal2 s 2256 27650 2256 27650 4 gnd
port 514 nsew
rlabel metal2 s 1488 28203 1488 28203 4 gnd
port 514 nsew
rlabel metal2 s 1488 25517 1488 25517 4 gnd
port 514 nsew
rlabel metal2 s 240 28440 240 28440 4 gnd
port 514 nsew
rlabel metal2 s 1488 26623 1488 26623 4 gnd
port 514 nsew
rlabel metal2 s 2256 25517 2256 25517 4 gnd
port 514 nsew
rlabel metal2 s 2256 27413 2256 27413 4 gnd
port 514 nsew
rlabel metal2 s 1008 27413 1008 27413 4 gnd
port 514 nsew
rlabel metal2 s 1008 26860 1008 26860 4 gnd
port 514 nsew
rlabel metal2 s 1008 26307 1008 26307 4 gnd
port 514 nsew
rlabel metal2 s 2256 27887 2256 27887 4 gnd
port 514 nsew
rlabel metal2 s 1008 28440 1008 28440 4 gnd
port 514 nsew
rlabel metal2 s 240 25833 240 25833 4 gnd
port 514 nsew
rlabel metal2 s 1488 27097 1488 27097 4 gnd
port 514 nsew
rlabel metal2 s 240 28203 240 28203 4 gnd
port 514 nsew
rlabel metal2 s 1488 25833 1488 25833 4 gnd
port 514 nsew
rlabel metal2 s 1008 26623 1008 26623 4 gnd
port 514 nsew
rlabel metal2 s 1008 27887 1008 27887 4 gnd
port 514 nsew
rlabel metal2 s 3504 26070 3504 26070 4 gnd
port 514 nsew
rlabel metal2 s 3504 26860 3504 26860 4 gnd
port 514 nsew
rlabel metal2 s 3984 27650 3984 27650 4 gnd
port 514 nsew
rlabel metal2 s 3984 26070 3984 26070 4 gnd
port 514 nsew
rlabel metal2 s 4752 26860 4752 26860 4 gnd
port 514 nsew
rlabel metal2 s 3984 27097 3984 27097 4 gnd
port 514 nsew
rlabel metal2 s 2736 26307 2736 26307 4 gnd
port 514 nsew
rlabel metal2 s 2736 27887 2736 27887 4 gnd
port 514 nsew
rlabel metal2 s 2736 27413 2736 27413 4 gnd
port 514 nsew
rlabel metal2 s 2736 25517 2736 25517 4 gnd
port 514 nsew
rlabel metal2 s 2736 27650 2736 27650 4 gnd
port 514 nsew
rlabel metal2 s 2736 26623 2736 26623 4 gnd
port 514 nsew
rlabel metal2 s 2736 27097 2736 27097 4 gnd
port 514 nsew
rlabel metal2 s 3504 26623 3504 26623 4 gnd
port 514 nsew
rlabel metal2 s 3504 27887 3504 27887 4 gnd
port 514 nsew
rlabel metal2 s 3984 28440 3984 28440 4 gnd
port 514 nsew
rlabel metal2 s 4752 26307 4752 26307 4 gnd
port 514 nsew
rlabel metal2 s 2736 26070 2736 26070 4 gnd
port 514 nsew
rlabel metal2 s 4752 27887 4752 27887 4 gnd
port 514 nsew
rlabel metal2 s 3504 25833 3504 25833 4 gnd
port 514 nsew
rlabel metal2 s 4752 28440 4752 28440 4 gnd
port 514 nsew
rlabel metal2 s 4752 26623 4752 26623 4 gnd
port 514 nsew
rlabel metal2 s 2736 28203 2736 28203 4 gnd
port 514 nsew
rlabel metal2 s 4752 25517 4752 25517 4 gnd
port 514 nsew
rlabel metal2 s 3984 25517 3984 25517 4 gnd
port 514 nsew
rlabel metal2 s 4752 27413 4752 27413 4 gnd
port 514 nsew
rlabel metal2 s 2736 26860 2736 26860 4 gnd
port 514 nsew
rlabel metal2 s 3504 27413 3504 27413 4 gnd
port 514 nsew
rlabel metal2 s 3984 25833 3984 25833 4 gnd
port 514 nsew
rlabel metal2 s 3984 26307 3984 26307 4 gnd
port 514 nsew
rlabel metal2 s 4752 26070 4752 26070 4 gnd
port 514 nsew
rlabel metal2 s 2736 25833 2736 25833 4 gnd
port 514 nsew
rlabel metal2 s 3984 26623 3984 26623 4 gnd
port 514 nsew
rlabel metal2 s 3504 28440 3504 28440 4 gnd
port 514 nsew
rlabel metal2 s 4752 28203 4752 28203 4 gnd
port 514 nsew
rlabel metal2 s 3984 26860 3984 26860 4 gnd
port 514 nsew
rlabel metal2 s 3984 27887 3984 27887 4 gnd
port 514 nsew
rlabel metal2 s 4752 27097 4752 27097 4 gnd
port 514 nsew
rlabel metal2 s 3504 27650 3504 27650 4 gnd
port 514 nsew
rlabel metal2 s 3984 27413 3984 27413 4 gnd
port 514 nsew
rlabel metal2 s 3504 26307 3504 26307 4 gnd
port 514 nsew
rlabel metal2 s 3504 28203 3504 28203 4 gnd
port 514 nsew
rlabel metal2 s 3984 28203 3984 28203 4 gnd
port 514 nsew
rlabel metal2 s 4752 27650 4752 27650 4 gnd
port 514 nsew
rlabel metal2 s 3504 27097 3504 27097 4 gnd
port 514 nsew
rlabel metal2 s 3504 25517 3504 25517 4 gnd
port 514 nsew
rlabel metal2 s 4752 25833 4752 25833 4 gnd
port 514 nsew
rlabel metal2 s 2736 28440 2736 28440 4 gnd
port 514 nsew
rlabel metal2 s 9744 29230 9744 29230 4 gnd
port 514 nsew
rlabel metal2 s 8976 29230 8976 29230 4 gnd
port 514 nsew
rlabel metal2 s 8976 30573 8976 30573 4 gnd
port 514 nsew
rlabel metal2 s 7728 30573 7728 30573 4 gnd
port 514 nsew
rlabel metal2 s 9744 30573 9744 30573 4 gnd
port 514 nsew
rlabel metal2 s 8976 31363 8976 31363 4 gnd
port 514 nsew
rlabel metal2 s 7728 31600 7728 31600 4 gnd
port 514 nsew
rlabel metal2 s 7728 30020 7728 30020 4 gnd
port 514 nsew
rlabel metal2 s 8976 29783 8976 29783 4 gnd
port 514 nsew
rlabel metal2 s 7728 28993 7728 28993 4 gnd
port 514 nsew
rlabel metal2 s 8496 29467 8496 29467 4 gnd
port 514 nsew
rlabel metal2 s 9744 30020 9744 30020 4 gnd
port 514 nsew
rlabel metal2 s 8496 30020 8496 30020 4 gnd
port 514 nsew
rlabel metal2 s 8976 31047 8976 31047 4 gnd
port 514 nsew
rlabel metal2 s 7728 29783 7728 29783 4 gnd
port 514 nsew
rlabel metal2 s 7728 31363 7728 31363 4 gnd
port 514 nsew
rlabel metal2 s 7728 31047 7728 31047 4 gnd
port 514 nsew
rlabel metal2 s 9744 28993 9744 28993 4 gnd
port 514 nsew
rlabel metal2 s 7728 28677 7728 28677 4 gnd
port 514 nsew
rlabel metal2 s 8976 31600 8976 31600 4 gnd
port 514 nsew
rlabel metal2 s 8496 28993 8496 28993 4 gnd
port 514 nsew
rlabel metal2 s 8496 28677 8496 28677 4 gnd
port 514 nsew
rlabel metal2 s 8976 30810 8976 30810 4 gnd
port 514 nsew
rlabel metal2 s 9744 30257 9744 30257 4 gnd
port 514 nsew
rlabel metal2 s 8496 30810 8496 30810 4 gnd
port 514 nsew
rlabel metal2 s 8496 31600 8496 31600 4 gnd
port 514 nsew
rlabel metal2 s 9744 30810 9744 30810 4 gnd
port 514 nsew
rlabel metal2 s 8496 29230 8496 29230 4 gnd
port 514 nsew
rlabel metal2 s 8976 30257 8976 30257 4 gnd
port 514 nsew
rlabel metal2 s 8976 28677 8976 28677 4 gnd
port 514 nsew
rlabel metal2 s 8976 29467 8976 29467 4 gnd
port 514 nsew
rlabel metal2 s 9744 28677 9744 28677 4 gnd
port 514 nsew
rlabel metal2 s 8496 31363 8496 31363 4 gnd
port 514 nsew
rlabel metal2 s 8976 30020 8976 30020 4 gnd
port 514 nsew
rlabel metal2 s 7728 29467 7728 29467 4 gnd
port 514 nsew
rlabel metal2 s 7728 30810 7728 30810 4 gnd
port 514 nsew
rlabel metal2 s 9744 31600 9744 31600 4 gnd
port 514 nsew
rlabel metal2 s 8496 30257 8496 30257 4 gnd
port 514 nsew
rlabel metal2 s 9744 29783 9744 29783 4 gnd
port 514 nsew
rlabel metal2 s 8496 30573 8496 30573 4 gnd
port 514 nsew
rlabel metal2 s 9744 31363 9744 31363 4 gnd
port 514 nsew
rlabel metal2 s 8496 29783 8496 29783 4 gnd
port 514 nsew
rlabel metal2 s 9744 29467 9744 29467 4 gnd
port 514 nsew
rlabel metal2 s 8976 28993 8976 28993 4 gnd
port 514 nsew
rlabel metal2 s 7728 29230 7728 29230 4 gnd
port 514 nsew
rlabel metal2 s 7728 30257 7728 30257 4 gnd
port 514 nsew
rlabel metal2 s 9744 31047 9744 31047 4 gnd
port 514 nsew
rlabel metal2 s 8496 31047 8496 31047 4 gnd
port 514 nsew
rlabel metal2 s 6480 31600 6480 31600 4 gnd
port 514 nsew
rlabel metal2 s 5232 31047 5232 31047 4 gnd
port 514 nsew
rlabel metal2 s 6480 29783 6480 29783 4 gnd
port 514 nsew
rlabel metal2 s 6000 31363 6000 31363 4 gnd
port 514 nsew
rlabel metal2 s 5232 28993 5232 28993 4 gnd
port 514 nsew
rlabel metal2 s 6480 30573 6480 30573 4 gnd
port 514 nsew
rlabel metal2 s 7248 29230 7248 29230 4 gnd
port 514 nsew
rlabel metal2 s 5232 31600 5232 31600 4 gnd
port 514 nsew
rlabel metal2 s 6000 30020 6000 30020 4 gnd
port 514 nsew
rlabel metal2 s 6480 29467 6480 29467 4 gnd
port 514 nsew
rlabel metal2 s 6000 29230 6000 29230 4 gnd
port 514 nsew
rlabel metal2 s 6480 31363 6480 31363 4 gnd
port 514 nsew
rlabel metal2 s 7248 30020 7248 30020 4 gnd
port 514 nsew
rlabel metal2 s 6000 28677 6000 28677 4 gnd
port 514 nsew
rlabel metal2 s 5232 29230 5232 29230 4 gnd
port 514 nsew
rlabel metal2 s 6480 29230 6480 29230 4 gnd
port 514 nsew
rlabel metal2 s 6000 30257 6000 30257 4 gnd
port 514 nsew
rlabel metal2 s 6480 28677 6480 28677 4 gnd
port 514 nsew
rlabel metal2 s 6000 31047 6000 31047 4 gnd
port 514 nsew
rlabel metal2 s 7248 29467 7248 29467 4 gnd
port 514 nsew
rlabel metal2 s 6480 30810 6480 30810 4 gnd
port 514 nsew
rlabel metal2 s 5232 29467 5232 29467 4 gnd
port 514 nsew
rlabel metal2 s 6000 30810 6000 30810 4 gnd
port 514 nsew
rlabel metal2 s 5232 30257 5232 30257 4 gnd
port 514 nsew
rlabel metal2 s 7248 30810 7248 30810 4 gnd
port 514 nsew
rlabel metal2 s 6000 29783 6000 29783 4 gnd
port 514 nsew
rlabel metal2 s 5232 30573 5232 30573 4 gnd
port 514 nsew
rlabel metal2 s 6000 29467 6000 29467 4 gnd
port 514 nsew
rlabel metal2 s 5232 31363 5232 31363 4 gnd
port 514 nsew
rlabel metal2 s 6000 30573 6000 30573 4 gnd
port 514 nsew
rlabel metal2 s 7248 30573 7248 30573 4 gnd
port 514 nsew
rlabel metal2 s 7248 30257 7248 30257 4 gnd
port 514 nsew
rlabel metal2 s 7248 29783 7248 29783 4 gnd
port 514 nsew
rlabel metal2 s 7248 28993 7248 28993 4 gnd
port 514 nsew
rlabel metal2 s 6000 28993 6000 28993 4 gnd
port 514 nsew
rlabel metal2 s 5232 30020 5232 30020 4 gnd
port 514 nsew
rlabel metal2 s 5232 28677 5232 28677 4 gnd
port 514 nsew
rlabel metal2 s 6480 30257 6480 30257 4 gnd
port 514 nsew
rlabel metal2 s 6480 30020 6480 30020 4 gnd
port 514 nsew
rlabel metal2 s 7248 31047 7248 31047 4 gnd
port 514 nsew
rlabel metal2 s 6480 31047 6480 31047 4 gnd
port 514 nsew
rlabel metal2 s 5232 29783 5232 29783 4 gnd
port 514 nsew
rlabel metal2 s 7248 31600 7248 31600 4 gnd
port 514 nsew
rlabel metal2 s 6000 31600 6000 31600 4 gnd
port 514 nsew
rlabel metal2 s 7248 28677 7248 28677 4 gnd
port 514 nsew
rlabel metal2 s 5232 30810 5232 30810 4 gnd
port 514 nsew
rlabel metal2 s 6480 28993 6480 28993 4 gnd
port 514 nsew
rlabel metal2 s 7248 31363 7248 31363 4 gnd
port 514 nsew
rlabel metal2 s 7248 28440 7248 28440 4 gnd
port 514 nsew
rlabel metal2 s 7248 28203 7248 28203 4 gnd
port 514 nsew
rlabel metal2 s 7248 27887 7248 27887 4 gnd
port 514 nsew
rlabel metal2 s 6480 27097 6480 27097 4 gnd
port 514 nsew
rlabel metal2 s 6000 27097 6000 27097 4 gnd
port 514 nsew
rlabel metal2 s 6000 26307 6000 26307 4 gnd
port 514 nsew
rlabel metal2 s 6480 26623 6480 26623 4 gnd
port 514 nsew
rlabel metal2 s 5232 28440 5232 28440 4 gnd
port 514 nsew
rlabel metal2 s 5232 26860 5232 26860 4 gnd
port 514 nsew
rlabel metal2 s 7248 27097 7248 27097 4 gnd
port 514 nsew
rlabel metal2 s 5232 26070 5232 26070 4 gnd
port 514 nsew
rlabel metal2 s 5232 27887 5232 27887 4 gnd
port 514 nsew
rlabel metal2 s 5232 25833 5232 25833 4 gnd
port 514 nsew
rlabel metal2 s 7248 26070 7248 26070 4 gnd
port 514 nsew
rlabel metal2 s 7248 26860 7248 26860 4 gnd
port 514 nsew
rlabel metal2 s 6000 26860 6000 26860 4 gnd
port 514 nsew
rlabel metal2 s 6480 26860 6480 26860 4 gnd
port 514 nsew
rlabel metal2 s 6000 25517 6000 25517 4 gnd
port 514 nsew
rlabel metal2 s 6000 27887 6000 27887 4 gnd
port 514 nsew
rlabel metal2 s 6000 27650 6000 27650 4 gnd
port 514 nsew
rlabel metal2 s 7248 27413 7248 27413 4 gnd
port 514 nsew
rlabel metal2 s 5232 26623 5232 26623 4 gnd
port 514 nsew
rlabel metal2 s 6480 27650 6480 27650 4 gnd
port 514 nsew
rlabel metal2 s 7248 25517 7248 25517 4 gnd
port 514 nsew
rlabel metal2 s 6480 26070 6480 26070 4 gnd
port 514 nsew
rlabel metal2 s 7248 27650 7248 27650 4 gnd
port 514 nsew
rlabel metal2 s 7248 26307 7248 26307 4 gnd
port 514 nsew
rlabel metal2 s 6480 28440 6480 28440 4 gnd
port 514 nsew
rlabel metal2 s 6480 25517 6480 25517 4 gnd
port 514 nsew
rlabel metal2 s 5232 27650 5232 27650 4 gnd
port 514 nsew
rlabel metal2 s 6000 28440 6000 28440 4 gnd
port 514 nsew
rlabel metal2 s 6000 26070 6000 26070 4 gnd
port 514 nsew
rlabel metal2 s 6000 27413 6000 27413 4 gnd
port 514 nsew
rlabel metal2 s 5232 26307 5232 26307 4 gnd
port 514 nsew
rlabel metal2 s 5232 27413 5232 27413 4 gnd
port 514 nsew
rlabel metal2 s 5232 28203 5232 28203 4 gnd
port 514 nsew
rlabel metal2 s 6480 26307 6480 26307 4 gnd
port 514 nsew
rlabel metal2 s 5232 27097 5232 27097 4 gnd
port 514 nsew
rlabel metal2 s 6000 28203 6000 28203 4 gnd
port 514 nsew
rlabel metal2 s 6480 28203 6480 28203 4 gnd
port 514 nsew
rlabel metal2 s 6480 25833 6480 25833 4 gnd
port 514 nsew
rlabel metal2 s 7248 26623 7248 26623 4 gnd
port 514 nsew
rlabel metal2 s 5232 25517 5232 25517 4 gnd
port 514 nsew
rlabel metal2 s 6000 26623 6000 26623 4 gnd
port 514 nsew
rlabel metal2 s 6480 27413 6480 27413 4 gnd
port 514 nsew
rlabel metal2 s 6000 25833 6000 25833 4 gnd
port 514 nsew
rlabel metal2 s 6480 27887 6480 27887 4 gnd
port 514 nsew
rlabel metal2 s 7248 25833 7248 25833 4 gnd
port 514 nsew
rlabel metal2 s 9744 28203 9744 28203 4 gnd
port 514 nsew
rlabel metal2 s 8976 25517 8976 25517 4 gnd
port 514 nsew
rlabel metal2 s 9744 26070 9744 26070 4 gnd
port 514 nsew
rlabel metal2 s 7728 25517 7728 25517 4 gnd
port 514 nsew
rlabel metal2 s 7728 26860 7728 26860 4 gnd
port 514 nsew
rlabel metal2 s 9744 25517 9744 25517 4 gnd
port 514 nsew
rlabel metal2 s 8496 27650 8496 27650 4 gnd
port 514 nsew
rlabel metal2 s 8496 27887 8496 27887 4 gnd
port 514 nsew
rlabel metal2 s 8976 27413 8976 27413 4 gnd
port 514 nsew
rlabel metal2 s 8976 26070 8976 26070 4 gnd
port 514 nsew
rlabel metal2 s 8976 28440 8976 28440 4 gnd
port 514 nsew
rlabel metal2 s 9744 26860 9744 26860 4 gnd
port 514 nsew
rlabel metal2 s 9744 25833 9744 25833 4 gnd
port 514 nsew
rlabel metal2 s 7728 27650 7728 27650 4 gnd
port 514 nsew
rlabel metal2 s 8496 28440 8496 28440 4 gnd
port 514 nsew
rlabel metal2 s 8976 26623 8976 26623 4 gnd
port 514 nsew
rlabel metal2 s 9744 26307 9744 26307 4 gnd
port 514 nsew
rlabel metal2 s 7728 26070 7728 26070 4 gnd
port 514 nsew
rlabel metal2 s 8976 25833 8976 25833 4 gnd
port 514 nsew
rlabel metal2 s 8496 26860 8496 26860 4 gnd
port 514 nsew
rlabel metal2 s 8976 26860 8976 26860 4 gnd
port 514 nsew
rlabel metal2 s 8496 25517 8496 25517 4 gnd
port 514 nsew
rlabel metal2 s 7728 28203 7728 28203 4 gnd
port 514 nsew
rlabel metal2 s 8976 27650 8976 27650 4 gnd
port 514 nsew
rlabel metal2 s 9744 27887 9744 27887 4 gnd
port 514 nsew
rlabel metal2 s 8496 27413 8496 27413 4 gnd
port 514 nsew
rlabel metal2 s 8976 28203 8976 28203 4 gnd
port 514 nsew
rlabel metal2 s 9744 27097 9744 27097 4 gnd
port 514 nsew
rlabel metal2 s 7728 26307 7728 26307 4 gnd
port 514 nsew
rlabel metal2 s 8976 27887 8976 27887 4 gnd
port 514 nsew
rlabel metal2 s 7728 25833 7728 25833 4 gnd
port 514 nsew
rlabel metal2 s 7728 28440 7728 28440 4 gnd
port 514 nsew
rlabel metal2 s 9744 26623 9744 26623 4 gnd
port 514 nsew
rlabel metal2 s 8496 26070 8496 26070 4 gnd
port 514 nsew
rlabel metal2 s 9744 27650 9744 27650 4 gnd
port 514 nsew
rlabel metal2 s 8976 27097 8976 27097 4 gnd
port 514 nsew
rlabel metal2 s 7728 27413 7728 27413 4 gnd
port 514 nsew
rlabel metal2 s 9744 28440 9744 28440 4 gnd
port 514 nsew
rlabel metal2 s 8496 27097 8496 27097 4 gnd
port 514 nsew
rlabel metal2 s 8976 26307 8976 26307 4 gnd
port 514 nsew
rlabel metal2 s 8496 26307 8496 26307 4 gnd
port 514 nsew
rlabel metal2 s 7728 27887 7728 27887 4 gnd
port 514 nsew
rlabel metal2 s 8496 28203 8496 28203 4 gnd
port 514 nsew
rlabel metal2 s 8496 26623 8496 26623 4 gnd
port 514 nsew
rlabel metal2 s 7728 27097 7728 27097 4 gnd
port 514 nsew
rlabel metal2 s 7728 26623 7728 26623 4 gnd
port 514 nsew
rlabel metal2 s 8496 25833 8496 25833 4 gnd
port 514 nsew
rlabel metal2 s 9744 27413 9744 27413 4 gnd
port 514 nsew
rlabel metal2 s 17712 36340 17712 36340 4 gnd
port 514 nsew
rlabel metal2 s 18480 36577 18480 36577 4 gnd
port 514 nsew
rlabel metal2 s 19728 35550 19728 35550 4 gnd
port 514 nsew
rlabel metal2 s 18960 35313 18960 35313 4 gnd
port 514 nsew
rlabel metal2 s 17712 36893 17712 36893 4 gnd
port 514 nsew
rlabel metal2 s 18960 34997 18960 34997 4 gnd
port 514 nsew
rlabel metal2 s 17712 35550 17712 35550 4 gnd
port 514 nsew
rlabel metal2 s 19968 36467 19968 36467 4 wl1_92
port 442 nsew
rlabel metal2 s 19968 37003 19968 37003 4 wl1_93
port 444 nsew
rlabel metal2 s 18960 36103 18960 36103 4 gnd
port 514 nsew
rlabel metal2 s 18960 36340 18960 36340 4 gnd
port 514 nsew
rlabel metal2 s 18480 37367 18480 37367 4 gnd
port 514 nsew
rlabel metal2 s 19968 35993 19968 35993 4 wl0_91
port 439 nsew
rlabel metal2 s 18480 36893 18480 36893 4 gnd
port 514 nsew
rlabel metal2 s 18480 34997 18480 34997 4 gnd
port 514 nsew
rlabel metal2 s 19728 37920 19728 37920 4 gnd
port 514 nsew
rlabel metal2 s 17712 34997 17712 34997 4 gnd
port 514 nsew
rlabel metal2 s 18480 36103 18480 36103 4 gnd
port 514 nsew
rlabel metal2 s 19728 36103 19728 36103 4 gnd
port 514 nsew
rlabel metal2 s 17712 36103 17712 36103 4 gnd
port 514 nsew
rlabel metal2 s 18960 37683 18960 37683 4 gnd
port 514 nsew
rlabel metal2 s 19728 36340 19728 36340 4 gnd
port 514 nsew
rlabel metal2 s 18960 35787 18960 35787 4 gnd
port 514 nsew
rlabel metal2 s 19728 35313 19728 35313 4 gnd
port 514 nsew
rlabel metal2 s 19968 37793 19968 37793 4 wl1_95
port 448 nsew
rlabel metal2 s 19728 36577 19728 36577 4 gnd
port 514 nsew
rlabel metal2 s 17712 37683 17712 37683 4 gnd
port 514 nsew
rlabel metal2 s 18960 37130 18960 37130 4 gnd
port 514 nsew
rlabel metal2 s 19968 35677 19968 35677 4 wl1_90
port 438 nsew
rlabel metal2 s 19728 34997 19728 34997 4 gnd
port 514 nsew
rlabel metal2 s 17712 35787 17712 35787 4 gnd
port 514 nsew
rlabel metal2 s 18480 37683 18480 37683 4 gnd
port 514 nsew
rlabel metal2 s 19728 37367 19728 37367 4 gnd
port 514 nsew
rlabel metal2 s 18480 36340 18480 36340 4 gnd
port 514 nsew
rlabel metal2 s 19728 35787 19728 35787 4 gnd
port 514 nsew
rlabel metal2 s 19728 36893 19728 36893 4 gnd
port 514 nsew
rlabel metal2 s 18480 35787 18480 35787 4 gnd
port 514 nsew
rlabel metal2 s 18960 37920 18960 37920 4 gnd
port 514 nsew
rlabel metal2 s 18960 36893 18960 36893 4 gnd
port 514 nsew
rlabel metal2 s 18960 36577 18960 36577 4 gnd
port 514 nsew
rlabel metal2 s 18480 37130 18480 37130 4 gnd
port 514 nsew
rlabel metal2 s 19728 37683 19728 37683 4 gnd
port 514 nsew
rlabel metal2 s 18480 35313 18480 35313 4 gnd
port 514 nsew
rlabel metal2 s 19968 37477 19968 37477 4 wl0_94
port 445 nsew
rlabel metal2 s 17712 37920 17712 37920 4 gnd
port 514 nsew
rlabel metal2 s 18480 37920 18480 37920 4 gnd
port 514 nsew
rlabel metal2 s 19968 35107 19968 35107 4 wl0_88
port 433 nsew
rlabel metal2 s 17712 36577 17712 36577 4 gnd
port 514 nsew
rlabel metal2 s 19728 37130 19728 37130 4 gnd
port 514 nsew
rlabel metal2 s 19968 37257 19968 37257 4 wl1_94
port 446 nsew
rlabel metal2 s 18960 35550 18960 35550 4 gnd
port 514 nsew
rlabel metal2 s 18960 37367 18960 37367 4 gnd
port 514 nsew
rlabel metal2 s 17712 37130 17712 37130 4 gnd
port 514 nsew
rlabel metal2 s 18480 35550 18480 35550 4 gnd
port 514 nsew
rlabel metal2 s 19968 35203 19968 35203 4 wl0_89
port 435 nsew
rlabel metal2 s 19968 37573 19968 37573 4 wl0_95
port 447 nsew
rlabel metal2 s 19968 36783 19968 36783 4 wl0_93
port 443 nsew
rlabel metal2 s 19968 34887 19968 34887 4 wl1_88
port 434 nsew
rlabel metal2 s 17712 37367 17712 37367 4 gnd
port 514 nsew
rlabel metal2 s 19968 36687 19968 36687 4 wl0_92
port 441 nsew
rlabel metal2 s 19968 36213 19968 36213 4 wl1_91
port 440 nsew
rlabel metal2 s 19968 35423 19968 35423 4 wl1_89
port 436 nsew
rlabel metal2 s 19968 35897 19968 35897 4 wl0_90
port 437 nsew
rlabel metal2 s 17712 35313 17712 35313 4 gnd
port 514 nsew
rlabel metal2 s 15216 36577 15216 36577 4 gnd
port 514 nsew
rlabel metal2 s 15216 34997 15216 34997 4 gnd
port 514 nsew
rlabel metal2 s 15216 35550 15216 35550 4 gnd
port 514 nsew
rlabel metal2 s 16464 36893 16464 36893 4 gnd
port 514 nsew
rlabel metal2 s 15984 35787 15984 35787 4 gnd
port 514 nsew
rlabel metal2 s 15216 36893 15216 36893 4 gnd
port 514 nsew
rlabel metal2 s 17232 36103 17232 36103 4 gnd
port 514 nsew
rlabel metal2 s 15984 37130 15984 37130 4 gnd
port 514 nsew
rlabel metal2 s 17232 35313 17232 35313 4 gnd
port 514 nsew
rlabel metal2 s 15984 35313 15984 35313 4 gnd
port 514 nsew
rlabel metal2 s 16464 37683 16464 37683 4 gnd
port 514 nsew
rlabel metal2 s 15216 36103 15216 36103 4 gnd
port 514 nsew
rlabel metal2 s 17232 36340 17232 36340 4 gnd
port 514 nsew
rlabel metal2 s 17232 36577 17232 36577 4 gnd
port 514 nsew
rlabel metal2 s 16464 35313 16464 35313 4 gnd
port 514 nsew
rlabel metal2 s 15216 37130 15216 37130 4 gnd
port 514 nsew
rlabel metal2 s 15984 36893 15984 36893 4 gnd
port 514 nsew
rlabel metal2 s 16464 37920 16464 37920 4 gnd
port 514 nsew
rlabel metal2 s 15216 37920 15216 37920 4 gnd
port 514 nsew
rlabel metal2 s 16464 35550 16464 35550 4 gnd
port 514 nsew
rlabel metal2 s 17232 34997 17232 34997 4 gnd
port 514 nsew
rlabel metal2 s 17232 37130 17232 37130 4 gnd
port 514 nsew
rlabel metal2 s 15984 37920 15984 37920 4 gnd
port 514 nsew
rlabel metal2 s 15984 37683 15984 37683 4 gnd
port 514 nsew
rlabel metal2 s 15216 37683 15216 37683 4 gnd
port 514 nsew
rlabel metal2 s 15984 37367 15984 37367 4 gnd
port 514 nsew
rlabel metal2 s 16464 35787 16464 35787 4 gnd
port 514 nsew
rlabel metal2 s 17232 35787 17232 35787 4 gnd
port 514 nsew
rlabel metal2 s 15216 35313 15216 35313 4 gnd
port 514 nsew
rlabel metal2 s 17232 37367 17232 37367 4 gnd
port 514 nsew
rlabel metal2 s 15984 34997 15984 34997 4 gnd
port 514 nsew
rlabel metal2 s 15216 36340 15216 36340 4 gnd
port 514 nsew
rlabel metal2 s 16464 36577 16464 36577 4 gnd
port 514 nsew
rlabel metal2 s 17232 35550 17232 35550 4 gnd
port 514 nsew
rlabel metal2 s 15984 36103 15984 36103 4 gnd
port 514 nsew
rlabel metal2 s 15984 35550 15984 35550 4 gnd
port 514 nsew
rlabel metal2 s 15984 36577 15984 36577 4 gnd
port 514 nsew
rlabel metal2 s 17232 36893 17232 36893 4 gnd
port 514 nsew
rlabel metal2 s 17232 37920 17232 37920 4 gnd
port 514 nsew
rlabel metal2 s 16464 34997 16464 34997 4 gnd
port 514 nsew
rlabel metal2 s 15984 36340 15984 36340 4 gnd
port 514 nsew
rlabel metal2 s 16464 36340 16464 36340 4 gnd
port 514 nsew
rlabel metal2 s 15216 35787 15216 35787 4 gnd
port 514 nsew
rlabel metal2 s 16464 37367 16464 37367 4 gnd
port 514 nsew
rlabel metal2 s 17232 37683 17232 37683 4 gnd
port 514 nsew
rlabel metal2 s 16464 37130 16464 37130 4 gnd
port 514 nsew
rlabel metal2 s 16464 36103 16464 36103 4 gnd
port 514 nsew
rlabel metal2 s 15216 37367 15216 37367 4 gnd
port 514 nsew
rlabel metal2 s 17232 33733 17232 33733 4 gnd
port 514 nsew
rlabel metal2 s 15984 34207 15984 34207 4 gnd
port 514 nsew
rlabel metal2 s 15984 33417 15984 33417 4 gnd
port 514 nsew
rlabel metal2 s 16464 32390 16464 32390 4 gnd
port 514 nsew
rlabel metal2 s 17232 34523 17232 34523 4 gnd
port 514 nsew
rlabel metal2 s 16464 31837 16464 31837 4 gnd
port 514 nsew
rlabel metal2 s 17232 32943 17232 32943 4 gnd
port 514 nsew
rlabel metal2 s 15216 33180 15216 33180 4 gnd
port 514 nsew
rlabel metal2 s 17232 34760 17232 34760 4 gnd
port 514 nsew
rlabel metal2 s 16464 32627 16464 32627 4 gnd
port 514 nsew
rlabel metal2 s 15216 34523 15216 34523 4 gnd
port 514 nsew
rlabel metal2 s 15984 34523 15984 34523 4 gnd
port 514 nsew
rlabel metal2 s 15984 32390 15984 32390 4 gnd
port 514 nsew
rlabel metal2 s 17232 32390 17232 32390 4 gnd
port 514 nsew
rlabel metal2 s 15216 32943 15216 32943 4 gnd
port 514 nsew
rlabel metal2 s 15216 32153 15216 32153 4 gnd
port 514 nsew
rlabel metal2 s 15216 32627 15216 32627 4 gnd
port 514 nsew
rlabel metal2 s 17232 33417 17232 33417 4 gnd
port 514 nsew
rlabel metal2 s 15984 31837 15984 31837 4 gnd
port 514 nsew
rlabel metal2 s 17232 31837 17232 31837 4 gnd
port 514 nsew
rlabel metal2 s 16464 32153 16464 32153 4 gnd
port 514 nsew
rlabel metal2 s 16464 34207 16464 34207 4 gnd
port 514 nsew
rlabel metal2 s 15984 33733 15984 33733 4 gnd
port 514 nsew
rlabel metal2 s 15216 31837 15216 31837 4 gnd
port 514 nsew
rlabel metal2 s 15984 32153 15984 32153 4 gnd
port 514 nsew
rlabel metal2 s 17232 33180 17232 33180 4 gnd
port 514 nsew
rlabel metal2 s 16464 33180 16464 33180 4 gnd
port 514 nsew
rlabel metal2 s 16464 33970 16464 33970 4 gnd
port 514 nsew
rlabel metal2 s 15216 34760 15216 34760 4 gnd
port 514 nsew
rlabel metal2 s 15216 33733 15216 33733 4 gnd
port 514 nsew
rlabel metal2 s 15216 33970 15216 33970 4 gnd
port 514 nsew
rlabel metal2 s 15216 32390 15216 32390 4 gnd
port 514 nsew
rlabel metal2 s 16464 33417 16464 33417 4 gnd
port 514 nsew
rlabel metal2 s 15984 32943 15984 32943 4 gnd
port 514 nsew
rlabel metal2 s 17232 32627 17232 32627 4 gnd
port 514 nsew
rlabel metal2 s 17232 32153 17232 32153 4 gnd
port 514 nsew
rlabel metal2 s 15216 33417 15216 33417 4 gnd
port 514 nsew
rlabel metal2 s 17232 33970 17232 33970 4 gnd
port 514 nsew
rlabel metal2 s 16464 34760 16464 34760 4 gnd
port 514 nsew
rlabel metal2 s 16464 32943 16464 32943 4 gnd
port 514 nsew
rlabel metal2 s 15984 33180 15984 33180 4 gnd
port 514 nsew
rlabel metal2 s 16464 33733 16464 33733 4 gnd
port 514 nsew
rlabel metal2 s 15984 33970 15984 33970 4 gnd
port 514 nsew
rlabel metal2 s 16464 34523 16464 34523 4 gnd
port 514 nsew
rlabel metal2 s 15984 32627 15984 32627 4 gnd
port 514 nsew
rlabel metal2 s 15216 34207 15216 34207 4 gnd
port 514 nsew
rlabel metal2 s 15984 34760 15984 34760 4 gnd
port 514 nsew
rlabel metal2 s 17232 34207 17232 34207 4 gnd
port 514 nsew
rlabel metal2 s 19728 32153 19728 32153 4 gnd
port 514 nsew
rlabel metal2 s 17712 33970 17712 33970 4 gnd
port 514 nsew
rlabel metal2 s 18960 32390 18960 32390 4 gnd
port 514 nsew
rlabel metal2 s 18960 31837 18960 31837 4 gnd
port 514 nsew
rlabel metal2 s 19728 34523 19728 34523 4 gnd
port 514 nsew
rlabel metal2 s 19968 32833 19968 32833 4 wl0_83
port 423 nsew
rlabel metal2 s 17712 31837 17712 31837 4 gnd
port 514 nsew
rlabel metal2 s 18480 32153 18480 32153 4 gnd
port 514 nsew
rlabel metal2 s 18960 33970 18960 33970 4 gnd
port 514 nsew
rlabel metal2 s 19728 34207 19728 34207 4 gnd
port 514 nsew
rlabel metal2 s 19968 33623 19968 33623 4 wl0_85
port 427 nsew
rlabel metal2 s 18960 32153 18960 32153 4 gnd
port 514 nsew
rlabel metal2 s 19728 33733 19728 33733 4 gnd
port 514 nsew
rlabel metal2 s 17712 34523 17712 34523 4 gnd
port 514 nsew
rlabel metal2 s 18480 34207 18480 34207 4 gnd
port 514 nsew
rlabel metal2 s 17712 32943 17712 32943 4 gnd
port 514 nsew
rlabel metal2 s 18480 32943 18480 32943 4 gnd
port 514 nsew
rlabel metal2 s 19728 32943 19728 32943 4 gnd
port 514 nsew
rlabel metal2 s 18960 34523 18960 34523 4 gnd
port 514 nsew
rlabel metal2 s 19968 34097 19968 34097 4 wl1_86
port 430 nsew
rlabel metal2 s 17712 33180 17712 33180 4 gnd
port 514 nsew
rlabel metal2 s 19728 31837 19728 31837 4 gnd
port 514 nsew
rlabel metal2 s 18480 34523 18480 34523 4 gnd
port 514 nsew
rlabel metal2 s 18480 33970 18480 33970 4 gnd
port 514 nsew
rlabel metal2 s 18960 32627 18960 32627 4 gnd
port 514 nsew
rlabel metal2 s 19728 32390 19728 32390 4 gnd
port 514 nsew
rlabel metal2 s 19728 32627 19728 32627 4 gnd
port 514 nsew
rlabel metal2 s 18960 33733 18960 33733 4 gnd
port 514 nsew
rlabel metal2 s 17712 32390 17712 32390 4 gnd
port 514 nsew
rlabel metal2 s 18480 32627 18480 32627 4 gnd
port 514 nsew
rlabel metal2 s 18480 33417 18480 33417 4 gnd
port 514 nsew
rlabel metal2 s 18480 32390 18480 32390 4 gnd
port 514 nsew
rlabel metal2 s 19728 34760 19728 34760 4 gnd
port 514 nsew
rlabel metal2 s 19968 32263 19968 32263 4 wl1_81
port 420 nsew
rlabel metal2 s 18480 33180 18480 33180 4 gnd
port 514 nsew
rlabel metal2 s 18960 33417 18960 33417 4 gnd
port 514 nsew
rlabel metal2 s 19968 34317 19968 34317 4 wl0_86
port 429 nsew
rlabel metal2 s 19968 33307 19968 33307 4 wl1_84
port 426 nsew
rlabel metal2 s 19968 31947 19968 31947 4 wl0_80
port 417 nsew
rlabel metal2 s 19968 31727 19968 31727 4 wl1_80
port 418 nsew
rlabel metal2 s 19728 33417 19728 33417 4 gnd
port 514 nsew
rlabel metal2 s 17712 33417 17712 33417 4 gnd
port 514 nsew
rlabel metal2 s 17712 32153 17712 32153 4 gnd
port 514 nsew
rlabel metal2 s 19968 32737 19968 32737 4 wl0_82
port 421 nsew
rlabel metal2 s 19968 32043 19968 32043 4 wl0_81
port 419 nsew
rlabel metal2 s 17712 32627 17712 32627 4 gnd
port 514 nsew
rlabel metal2 s 18960 32943 18960 32943 4 gnd
port 514 nsew
rlabel metal2 s 19728 33970 19728 33970 4 gnd
port 514 nsew
rlabel metal2 s 19968 34413 19968 34413 4 wl0_87
port 431 nsew
rlabel metal2 s 17712 33733 17712 33733 4 gnd
port 514 nsew
rlabel metal2 s 18960 34207 18960 34207 4 gnd
port 514 nsew
rlabel metal2 s 18960 33180 18960 33180 4 gnd
port 514 nsew
rlabel metal2 s 17712 34760 17712 34760 4 gnd
port 514 nsew
rlabel metal2 s 18480 34760 18480 34760 4 gnd
port 514 nsew
rlabel metal2 s 19728 33180 19728 33180 4 gnd
port 514 nsew
rlabel metal2 s 19968 32517 19968 32517 4 wl1_82
port 422 nsew
rlabel metal2 s 18480 31837 18480 31837 4 gnd
port 514 nsew
rlabel metal2 s 19968 33843 19968 33843 4 wl1_85
port 428 nsew
rlabel metal2 s 18960 34760 18960 34760 4 gnd
port 514 nsew
rlabel metal2 s 19968 33053 19968 33053 4 wl1_83
port 424 nsew
rlabel metal2 s 17712 34207 17712 34207 4 gnd
port 514 nsew
rlabel metal2 s 19968 33527 19968 33527 4 wl0_84
port 425 nsew
rlabel metal2 s 19968 34633 19968 34633 4 wl1_87
port 432 nsew
rlabel metal2 s 18480 33733 18480 33733 4 gnd
port 514 nsew
rlabel metal2 s 13968 37920 13968 37920 4 gnd
port 514 nsew
rlabel metal2 s 13968 36577 13968 36577 4 gnd
port 514 nsew
rlabel metal2 s 13968 37683 13968 37683 4 gnd
port 514 nsew
rlabel metal2 s 13968 35550 13968 35550 4 gnd
port 514 nsew
rlabel metal2 s 12720 37683 12720 37683 4 gnd
port 514 nsew
rlabel metal2 s 13968 36893 13968 36893 4 gnd
port 514 nsew
rlabel metal2 s 13488 34997 13488 34997 4 gnd
port 514 nsew
rlabel metal2 s 13968 35313 13968 35313 4 gnd
port 514 nsew
rlabel metal2 s 13488 36340 13488 36340 4 gnd
port 514 nsew
rlabel metal2 s 14736 34997 14736 34997 4 gnd
port 514 nsew
rlabel metal2 s 14736 37683 14736 37683 4 gnd
port 514 nsew
rlabel metal2 s 12720 36103 12720 36103 4 gnd
port 514 nsew
rlabel metal2 s 14736 36577 14736 36577 4 gnd
port 514 nsew
rlabel metal2 s 13968 35787 13968 35787 4 gnd
port 514 nsew
rlabel metal2 s 12720 36340 12720 36340 4 gnd
port 514 nsew
rlabel metal2 s 14736 35550 14736 35550 4 gnd
port 514 nsew
rlabel metal2 s 13488 35550 13488 35550 4 gnd
port 514 nsew
rlabel metal2 s 14736 36893 14736 36893 4 gnd
port 514 nsew
rlabel metal2 s 12720 35550 12720 35550 4 gnd
port 514 nsew
rlabel metal2 s 12720 36577 12720 36577 4 gnd
port 514 nsew
rlabel metal2 s 12720 37920 12720 37920 4 gnd
port 514 nsew
rlabel metal2 s 13488 35313 13488 35313 4 gnd
port 514 nsew
rlabel metal2 s 12720 35313 12720 35313 4 gnd
port 514 nsew
rlabel metal2 s 13968 37367 13968 37367 4 gnd
port 514 nsew
rlabel metal2 s 14736 36103 14736 36103 4 gnd
port 514 nsew
rlabel metal2 s 13488 36103 13488 36103 4 gnd
port 514 nsew
rlabel metal2 s 12720 37130 12720 37130 4 gnd
port 514 nsew
rlabel metal2 s 14736 36340 14736 36340 4 gnd
port 514 nsew
rlabel metal2 s 13968 34997 13968 34997 4 gnd
port 514 nsew
rlabel metal2 s 12720 35787 12720 35787 4 gnd
port 514 nsew
rlabel metal2 s 14736 37920 14736 37920 4 gnd
port 514 nsew
rlabel metal2 s 12720 36893 12720 36893 4 gnd
port 514 nsew
rlabel metal2 s 13488 36577 13488 36577 4 gnd
port 514 nsew
rlabel metal2 s 13488 37130 13488 37130 4 gnd
port 514 nsew
rlabel metal2 s 13968 36103 13968 36103 4 gnd
port 514 nsew
rlabel metal2 s 14736 37367 14736 37367 4 gnd
port 514 nsew
rlabel metal2 s 13968 36340 13968 36340 4 gnd
port 514 nsew
rlabel metal2 s 13968 37130 13968 37130 4 gnd
port 514 nsew
rlabel metal2 s 13488 37367 13488 37367 4 gnd
port 514 nsew
rlabel metal2 s 14736 35313 14736 35313 4 gnd
port 514 nsew
rlabel metal2 s 14736 37130 14736 37130 4 gnd
port 514 nsew
rlabel metal2 s 14736 35787 14736 35787 4 gnd
port 514 nsew
rlabel metal2 s 13488 35787 13488 35787 4 gnd
port 514 nsew
rlabel metal2 s 13488 36893 13488 36893 4 gnd
port 514 nsew
rlabel metal2 s 12720 37367 12720 37367 4 gnd
port 514 nsew
rlabel metal2 s 13488 37683 13488 37683 4 gnd
port 514 nsew
rlabel metal2 s 12720 34997 12720 34997 4 gnd
port 514 nsew
rlabel metal2 s 13488 37920 13488 37920 4 gnd
port 514 nsew
rlabel metal2 s 10224 35313 10224 35313 4 gnd
port 514 nsew
rlabel metal2 s 10224 37920 10224 37920 4 gnd
port 514 nsew
rlabel metal2 s 11472 37367 11472 37367 4 gnd
port 514 nsew
rlabel metal2 s 10992 36893 10992 36893 4 gnd
port 514 nsew
rlabel metal2 s 11472 36103 11472 36103 4 gnd
port 514 nsew
rlabel metal2 s 10992 37367 10992 37367 4 gnd
port 514 nsew
rlabel metal2 s 12240 36893 12240 36893 4 gnd
port 514 nsew
rlabel metal2 s 10992 37683 10992 37683 4 gnd
port 514 nsew
rlabel metal2 s 10992 36103 10992 36103 4 gnd
port 514 nsew
rlabel metal2 s 10224 37130 10224 37130 4 gnd
port 514 nsew
rlabel metal2 s 12240 37130 12240 37130 4 gnd
port 514 nsew
rlabel metal2 s 10224 36893 10224 36893 4 gnd
port 514 nsew
rlabel metal2 s 10224 36103 10224 36103 4 gnd
port 514 nsew
rlabel metal2 s 12240 35550 12240 35550 4 gnd
port 514 nsew
rlabel metal2 s 10224 35550 10224 35550 4 gnd
port 514 nsew
rlabel metal2 s 11472 35313 11472 35313 4 gnd
port 514 nsew
rlabel metal2 s 12240 35313 12240 35313 4 gnd
port 514 nsew
rlabel metal2 s 12240 37920 12240 37920 4 gnd
port 514 nsew
rlabel metal2 s 11472 36893 11472 36893 4 gnd
port 514 nsew
rlabel metal2 s 10224 35787 10224 35787 4 gnd
port 514 nsew
rlabel metal2 s 12240 36103 12240 36103 4 gnd
port 514 nsew
rlabel metal2 s 12240 37683 12240 37683 4 gnd
port 514 nsew
rlabel metal2 s 11472 37683 11472 37683 4 gnd
port 514 nsew
rlabel metal2 s 12240 36577 12240 36577 4 gnd
port 514 nsew
rlabel metal2 s 10992 36577 10992 36577 4 gnd
port 514 nsew
rlabel metal2 s 11472 36340 11472 36340 4 gnd
port 514 nsew
rlabel metal2 s 11472 35550 11472 35550 4 gnd
port 514 nsew
rlabel metal2 s 10992 35550 10992 35550 4 gnd
port 514 nsew
rlabel metal2 s 12240 34997 12240 34997 4 gnd
port 514 nsew
rlabel metal2 s 10992 37920 10992 37920 4 gnd
port 514 nsew
rlabel metal2 s 10992 36340 10992 36340 4 gnd
port 514 nsew
rlabel metal2 s 10992 37130 10992 37130 4 gnd
port 514 nsew
rlabel metal2 s 12240 36340 12240 36340 4 gnd
port 514 nsew
rlabel metal2 s 11472 35787 11472 35787 4 gnd
port 514 nsew
rlabel metal2 s 12240 37367 12240 37367 4 gnd
port 514 nsew
rlabel metal2 s 11472 37130 11472 37130 4 gnd
port 514 nsew
rlabel metal2 s 10224 37683 10224 37683 4 gnd
port 514 nsew
rlabel metal2 s 10224 37367 10224 37367 4 gnd
port 514 nsew
rlabel metal2 s 12240 35787 12240 35787 4 gnd
port 514 nsew
rlabel metal2 s 10224 36340 10224 36340 4 gnd
port 514 nsew
rlabel metal2 s 10992 34997 10992 34997 4 gnd
port 514 nsew
rlabel metal2 s 10224 36577 10224 36577 4 gnd
port 514 nsew
rlabel metal2 s 11472 37920 11472 37920 4 gnd
port 514 nsew
rlabel metal2 s 10992 35313 10992 35313 4 gnd
port 514 nsew
rlabel metal2 s 11472 34997 11472 34997 4 gnd
port 514 nsew
rlabel metal2 s 10992 35787 10992 35787 4 gnd
port 514 nsew
rlabel metal2 s 11472 36577 11472 36577 4 gnd
port 514 nsew
rlabel metal2 s 10224 34997 10224 34997 4 gnd
port 514 nsew
rlabel metal2 s 10992 33180 10992 33180 4 gnd
port 514 nsew
rlabel metal2 s 12240 33180 12240 33180 4 gnd
port 514 nsew
rlabel metal2 s 12240 33733 12240 33733 4 gnd
port 514 nsew
rlabel metal2 s 10992 33733 10992 33733 4 gnd
port 514 nsew
rlabel metal2 s 11472 32943 11472 32943 4 gnd
port 514 nsew
rlabel metal2 s 11472 33970 11472 33970 4 gnd
port 514 nsew
rlabel metal2 s 12240 33970 12240 33970 4 gnd
port 514 nsew
rlabel metal2 s 11472 31837 11472 31837 4 gnd
port 514 nsew
rlabel metal2 s 10224 33180 10224 33180 4 gnd
port 514 nsew
rlabel metal2 s 10224 32153 10224 32153 4 gnd
port 514 nsew
rlabel metal2 s 10224 31837 10224 31837 4 gnd
port 514 nsew
rlabel metal2 s 10992 32943 10992 32943 4 gnd
port 514 nsew
rlabel metal2 s 10224 32627 10224 32627 4 gnd
port 514 nsew
rlabel metal2 s 10992 34760 10992 34760 4 gnd
port 514 nsew
rlabel metal2 s 11472 34523 11472 34523 4 gnd
port 514 nsew
rlabel metal2 s 10224 33970 10224 33970 4 gnd
port 514 nsew
rlabel metal2 s 10224 32390 10224 32390 4 gnd
port 514 nsew
rlabel metal2 s 10992 33970 10992 33970 4 gnd
port 514 nsew
rlabel metal2 s 10992 34523 10992 34523 4 gnd
port 514 nsew
rlabel metal2 s 10992 31837 10992 31837 4 gnd
port 514 nsew
rlabel metal2 s 12240 32153 12240 32153 4 gnd
port 514 nsew
rlabel metal2 s 10224 34207 10224 34207 4 gnd
port 514 nsew
rlabel metal2 s 11472 33180 11472 33180 4 gnd
port 514 nsew
rlabel metal2 s 11472 32627 11472 32627 4 gnd
port 514 nsew
rlabel metal2 s 10224 34760 10224 34760 4 gnd
port 514 nsew
rlabel metal2 s 12240 34523 12240 34523 4 gnd
port 514 nsew
rlabel metal2 s 10224 33417 10224 33417 4 gnd
port 514 nsew
rlabel metal2 s 11472 33733 11472 33733 4 gnd
port 514 nsew
rlabel metal2 s 11472 32390 11472 32390 4 gnd
port 514 nsew
rlabel metal2 s 11472 34760 11472 34760 4 gnd
port 514 nsew
rlabel metal2 s 10224 34523 10224 34523 4 gnd
port 514 nsew
rlabel metal2 s 11472 34207 11472 34207 4 gnd
port 514 nsew
rlabel metal2 s 10224 32943 10224 32943 4 gnd
port 514 nsew
rlabel metal2 s 10992 32153 10992 32153 4 gnd
port 514 nsew
rlabel metal2 s 10224 33733 10224 33733 4 gnd
port 514 nsew
rlabel metal2 s 12240 32390 12240 32390 4 gnd
port 514 nsew
rlabel metal2 s 12240 33417 12240 33417 4 gnd
port 514 nsew
rlabel metal2 s 11472 32153 11472 32153 4 gnd
port 514 nsew
rlabel metal2 s 12240 32627 12240 32627 4 gnd
port 514 nsew
rlabel metal2 s 11472 33417 11472 33417 4 gnd
port 514 nsew
rlabel metal2 s 10992 33417 10992 33417 4 gnd
port 514 nsew
rlabel metal2 s 10992 32627 10992 32627 4 gnd
port 514 nsew
rlabel metal2 s 12240 32943 12240 32943 4 gnd
port 514 nsew
rlabel metal2 s 12240 31837 12240 31837 4 gnd
port 514 nsew
rlabel metal2 s 10992 34207 10992 34207 4 gnd
port 514 nsew
rlabel metal2 s 12240 34207 12240 34207 4 gnd
port 514 nsew
rlabel metal2 s 12240 34760 12240 34760 4 gnd
port 514 nsew
rlabel metal2 s 10992 32390 10992 32390 4 gnd
port 514 nsew
rlabel metal2 s 13968 32153 13968 32153 4 gnd
port 514 nsew
rlabel metal2 s 12720 32153 12720 32153 4 gnd
port 514 nsew
rlabel metal2 s 12720 32943 12720 32943 4 gnd
port 514 nsew
rlabel metal2 s 13968 34760 13968 34760 4 gnd
port 514 nsew
rlabel metal2 s 14736 32627 14736 32627 4 gnd
port 514 nsew
rlabel metal2 s 12720 33970 12720 33970 4 gnd
port 514 nsew
rlabel metal2 s 13968 33970 13968 33970 4 gnd
port 514 nsew
rlabel metal2 s 14736 33417 14736 33417 4 gnd
port 514 nsew
rlabel metal2 s 12720 33180 12720 33180 4 gnd
port 514 nsew
rlabel metal2 s 14736 34760 14736 34760 4 gnd
port 514 nsew
rlabel metal2 s 13488 33417 13488 33417 4 gnd
port 514 nsew
rlabel metal2 s 12720 32627 12720 32627 4 gnd
port 514 nsew
rlabel metal2 s 14736 33180 14736 33180 4 gnd
port 514 nsew
rlabel metal2 s 13968 34207 13968 34207 4 gnd
port 514 nsew
rlabel metal2 s 14736 34523 14736 34523 4 gnd
port 514 nsew
rlabel metal2 s 13488 32153 13488 32153 4 gnd
port 514 nsew
rlabel metal2 s 14736 31837 14736 31837 4 gnd
port 514 nsew
rlabel metal2 s 12720 34523 12720 34523 4 gnd
port 514 nsew
rlabel metal2 s 13968 31837 13968 31837 4 gnd
port 514 nsew
rlabel metal2 s 13968 32943 13968 32943 4 gnd
port 514 nsew
rlabel metal2 s 13488 34207 13488 34207 4 gnd
port 514 nsew
rlabel metal2 s 12720 34207 12720 34207 4 gnd
port 514 nsew
rlabel metal2 s 13968 33733 13968 33733 4 gnd
port 514 nsew
rlabel metal2 s 13968 32627 13968 32627 4 gnd
port 514 nsew
rlabel metal2 s 14736 32153 14736 32153 4 gnd
port 514 nsew
rlabel metal2 s 12720 34760 12720 34760 4 gnd
port 514 nsew
rlabel metal2 s 13488 33733 13488 33733 4 gnd
port 514 nsew
rlabel metal2 s 13488 32627 13488 32627 4 gnd
port 514 nsew
rlabel metal2 s 12720 33417 12720 33417 4 gnd
port 514 nsew
rlabel metal2 s 13488 31837 13488 31837 4 gnd
port 514 nsew
rlabel metal2 s 12720 31837 12720 31837 4 gnd
port 514 nsew
rlabel metal2 s 14736 34207 14736 34207 4 gnd
port 514 nsew
rlabel metal2 s 12720 33733 12720 33733 4 gnd
port 514 nsew
rlabel metal2 s 12720 32390 12720 32390 4 gnd
port 514 nsew
rlabel metal2 s 13488 33180 13488 33180 4 gnd
port 514 nsew
rlabel metal2 s 14736 33733 14736 33733 4 gnd
port 514 nsew
rlabel metal2 s 14736 32943 14736 32943 4 gnd
port 514 nsew
rlabel metal2 s 13488 33970 13488 33970 4 gnd
port 514 nsew
rlabel metal2 s 13968 33180 13968 33180 4 gnd
port 514 nsew
rlabel metal2 s 13968 32390 13968 32390 4 gnd
port 514 nsew
rlabel metal2 s 13488 34760 13488 34760 4 gnd
port 514 nsew
rlabel metal2 s 13488 32943 13488 32943 4 gnd
port 514 nsew
rlabel metal2 s 14736 32390 14736 32390 4 gnd
port 514 nsew
rlabel metal2 s 13488 32390 13488 32390 4 gnd
port 514 nsew
rlabel metal2 s 13488 34523 13488 34523 4 gnd
port 514 nsew
rlabel metal2 s 13968 33417 13968 33417 4 gnd
port 514 nsew
rlabel metal2 s 14736 33970 14736 33970 4 gnd
port 514 nsew
rlabel metal2 s 13968 34523 13968 34523 4 gnd
port 514 nsew
rlabel metal2 s 14736 30810 14736 30810 4 gnd
port 514 nsew
rlabel metal2 s 12720 31363 12720 31363 4 gnd
port 514 nsew
rlabel metal2 s 12720 29230 12720 29230 4 gnd
port 514 nsew
rlabel metal2 s 13488 30573 13488 30573 4 gnd
port 514 nsew
rlabel metal2 s 13488 30020 13488 30020 4 gnd
port 514 nsew
rlabel metal2 s 14736 28993 14736 28993 4 gnd
port 514 nsew
rlabel metal2 s 12720 29783 12720 29783 4 gnd
port 514 nsew
rlabel metal2 s 12720 28677 12720 28677 4 gnd
port 514 nsew
rlabel metal2 s 13488 28677 13488 28677 4 gnd
port 514 nsew
rlabel metal2 s 13488 28993 13488 28993 4 gnd
port 514 nsew
rlabel metal2 s 13968 28993 13968 28993 4 gnd
port 514 nsew
rlabel metal2 s 14736 29467 14736 29467 4 gnd
port 514 nsew
rlabel metal2 s 14736 29783 14736 29783 4 gnd
port 514 nsew
rlabel metal2 s 13488 29783 13488 29783 4 gnd
port 514 nsew
rlabel metal2 s 14736 30573 14736 30573 4 gnd
port 514 nsew
rlabel metal2 s 13968 29467 13968 29467 4 gnd
port 514 nsew
rlabel metal2 s 12720 31047 12720 31047 4 gnd
port 514 nsew
rlabel metal2 s 13968 31600 13968 31600 4 gnd
port 514 nsew
rlabel metal2 s 13968 31363 13968 31363 4 gnd
port 514 nsew
rlabel metal2 s 13968 30810 13968 30810 4 gnd
port 514 nsew
rlabel metal2 s 13968 29783 13968 29783 4 gnd
port 514 nsew
rlabel metal2 s 14736 29230 14736 29230 4 gnd
port 514 nsew
rlabel metal2 s 14736 30257 14736 30257 4 gnd
port 514 nsew
rlabel metal2 s 13968 30257 13968 30257 4 gnd
port 514 nsew
rlabel metal2 s 13488 29230 13488 29230 4 gnd
port 514 nsew
rlabel metal2 s 13488 30257 13488 30257 4 gnd
port 514 nsew
rlabel metal2 s 13968 30573 13968 30573 4 gnd
port 514 nsew
rlabel metal2 s 12720 29467 12720 29467 4 gnd
port 514 nsew
rlabel metal2 s 14736 31047 14736 31047 4 gnd
port 514 nsew
rlabel metal2 s 13488 29467 13488 29467 4 gnd
port 514 nsew
rlabel metal2 s 14736 28677 14736 28677 4 gnd
port 514 nsew
rlabel metal2 s 12720 30573 12720 30573 4 gnd
port 514 nsew
rlabel metal2 s 12720 30810 12720 30810 4 gnd
port 514 nsew
rlabel metal2 s 13968 28677 13968 28677 4 gnd
port 514 nsew
rlabel metal2 s 13968 30020 13968 30020 4 gnd
port 514 nsew
rlabel metal2 s 13488 31047 13488 31047 4 gnd
port 514 nsew
rlabel metal2 s 12720 28993 12720 28993 4 gnd
port 514 nsew
rlabel metal2 s 14736 31600 14736 31600 4 gnd
port 514 nsew
rlabel metal2 s 13488 31363 13488 31363 4 gnd
port 514 nsew
rlabel metal2 s 12720 31600 12720 31600 4 gnd
port 514 nsew
rlabel metal2 s 13488 30810 13488 30810 4 gnd
port 514 nsew
rlabel metal2 s 13488 31600 13488 31600 4 gnd
port 514 nsew
rlabel metal2 s 12720 30020 12720 30020 4 gnd
port 514 nsew
rlabel metal2 s 13968 29230 13968 29230 4 gnd
port 514 nsew
rlabel metal2 s 14736 31363 14736 31363 4 gnd
port 514 nsew
rlabel metal2 s 14736 30020 14736 30020 4 gnd
port 514 nsew
rlabel metal2 s 12720 30257 12720 30257 4 gnd
port 514 nsew
rlabel metal2 s 13968 31047 13968 31047 4 gnd
port 514 nsew
rlabel metal2 s 10992 31600 10992 31600 4 gnd
port 514 nsew
rlabel metal2 s 11472 30257 11472 30257 4 gnd
port 514 nsew
rlabel metal2 s 11472 28993 11472 28993 4 gnd
port 514 nsew
rlabel metal2 s 12240 31363 12240 31363 4 gnd
port 514 nsew
rlabel metal2 s 12240 29230 12240 29230 4 gnd
port 514 nsew
rlabel metal2 s 10224 29230 10224 29230 4 gnd
port 514 nsew
rlabel metal2 s 11472 31363 11472 31363 4 gnd
port 514 nsew
rlabel metal2 s 10224 28993 10224 28993 4 gnd
port 514 nsew
rlabel metal2 s 12240 30573 12240 30573 4 gnd
port 514 nsew
rlabel metal2 s 11472 30020 11472 30020 4 gnd
port 514 nsew
rlabel metal2 s 10992 30257 10992 30257 4 gnd
port 514 nsew
rlabel metal2 s 11472 29230 11472 29230 4 gnd
port 514 nsew
rlabel metal2 s 10992 31047 10992 31047 4 gnd
port 514 nsew
rlabel metal2 s 10224 30810 10224 30810 4 gnd
port 514 nsew
rlabel metal2 s 10992 30573 10992 30573 4 gnd
port 514 nsew
rlabel metal2 s 10224 30257 10224 30257 4 gnd
port 514 nsew
rlabel metal2 s 10992 28993 10992 28993 4 gnd
port 514 nsew
rlabel metal2 s 10992 29783 10992 29783 4 gnd
port 514 nsew
rlabel metal2 s 10992 29467 10992 29467 4 gnd
port 514 nsew
rlabel metal2 s 12240 28993 12240 28993 4 gnd
port 514 nsew
rlabel metal2 s 12240 28677 12240 28677 4 gnd
port 514 nsew
rlabel metal2 s 11472 29783 11472 29783 4 gnd
port 514 nsew
rlabel metal2 s 11472 30810 11472 30810 4 gnd
port 514 nsew
rlabel metal2 s 11472 29467 11472 29467 4 gnd
port 514 nsew
rlabel metal2 s 11472 28677 11472 28677 4 gnd
port 514 nsew
rlabel metal2 s 12240 30810 12240 30810 4 gnd
port 514 nsew
rlabel metal2 s 12240 31047 12240 31047 4 gnd
port 514 nsew
rlabel metal2 s 11472 30573 11472 30573 4 gnd
port 514 nsew
rlabel metal2 s 10992 30810 10992 30810 4 gnd
port 514 nsew
rlabel metal2 s 10224 30573 10224 30573 4 gnd
port 514 nsew
rlabel metal2 s 12240 29783 12240 29783 4 gnd
port 514 nsew
rlabel metal2 s 10992 28677 10992 28677 4 gnd
port 514 nsew
rlabel metal2 s 10992 31363 10992 31363 4 gnd
port 514 nsew
rlabel metal2 s 11472 31047 11472 31047 4 gnd
port 514 nsew
rlabel metal2 s 12240 30020 12240 30020 4 gnd
port 514 nsew
rlabel metal2 s 10224 29467 10224 29467 4 gnd
port 514 nsew
rlabel metal2 s 11472 31600 11472 31600 4 gnd
port 514 nsew
rlabel metal2 s 10224 30020 10224 30020 4 gnd
port 514 nsew
rlabel metal2 s 12240 31600 12240 31600 4 gnd
port 514 nsew
rlabel metal2 s 10224 31363 10224 31363 4 gnd
port 514 nsew
rlabel metal2 s 10224 31047 10224 31047 4 gnd
port 514 nsew
rlabel metal2 s 10224 31600 10224 31600 4 gnd
port 514 nsew
rlabel metal2 s 10992 30020 10992 30020 4 gnd
port 514 nsew
rlabel metal2 s 10224 29783 10224 29783 4 gnd
port 514 nsew
rlabel metal2 s 12240 30257 12240 30257 4 gnd
port 514 nsew
rlabel metal2 s 10992 29230 10992 29230 4 gnd
port 514 nsew
rlabel metal2 s 10224 28677 10224 28677 4 gnd
port 514 nsew
rlabel metal2 s 12240 29467 12240 29467 4 gnd
port 514 nsew
rlabel metal2 s 11472 25517 11472 25517 4 gnd
port 514 nsew
rlabel metal2 s 10992 27413 10992 27413 4 gnd
port 514 nsew
rlabel metal2 s 12240 27097 12240 27097 4 gnd
port 514 nsew
rlabel metal2 s 10224 27413 10224 27413 4 gnd
port 514 nsew
rlabel metal2 s 11472 27097 11472 27097 4 gnd
port 514 nsew
rlabel metal2 s 11472 27650 11472 27650 4 gnd
port 514 nsew
rlabel metal2 s 12240 28203 12240 28203 4 gnd
port 514 nsew
rlabel metal2 s 11472 26070 11472 26070 4 gnd
port 514 nsew
rlabel metal2 s 11472 26307 11472 26307 4 gnd
port 514 nsew
rlabel metal2 s 10992 26623 10992 26623 4 gnd
port 514 nsew
rlabel metal2 s 10992 28440 10992 28440 4 gnd
port 514 nsew
rlabel metal2 s 10224 26307 10224 26307 4 gnd
port 514 nsew
rlabel metal2 s 10224 25833 10224 25833 4 gnd
port 514 nsew
rlabel metal2 s 10992 27887 10992 27887 4 gnd
port 514 nsew
rlabel metal2 s 12240 26070 12240 26070 4 gnd
port 514 nsew
rlabel metal2 s 11472 28440 11472 28440 4 gnd
port 514 nsew
rlabel metal2 s 10224 26860 10224 26860 4 gnd
port 514 nsew
rlabel metal2 s 10992 28203 10992 28203 4 gnd
port 514 nsew
rlabel metal2 s 10224 27097 10224 27097 4 gnd
port 514 nsew
rlabel metal2 s 12240 27413 12240 27413 4 gnd
port 514 nsew
rlabel metal2 s 11472 26860 11472 26860 4 gnd
port 514 nsew
rlabel metal2 s 10992 26070 10992 26070 4 gnd
port 514 nsew
rlabel metal2 s 12240 26860 12240 26860 4 gnd
port 514 nsew
rlabel metal2 s 10992 26860 10992 26860 4 gnd
port 514 nsew
rlabel metal2 s 10224 27887 10224 27887 4 gnd
port 514 nsew
rlabel metal2 s 10224 27650 10224 27650 4 gnd
port 514 nsew
rlabel metal2 s 12240 26623 12240 26623 4 gnd
port 514 nsew
rlabel metal2 s 11472 28203 11472 28203 4 gnd
port 514 nsew
rlabel metal2 s 11472 26623 11472 26623 4 gnd
port 514 nsew
rlabel metal2 s 12240 27650 12240 27650 4 gnd
port 514 nsew
rlabel metal2 s 10224 28440 10224 28440 4 gnd
port 514 nsew
rlabel metal2 s 12240 25833 12240 25833 4 gnd
port 514 nsew
rlabel metal2 s 10224 28203 10224 28203 4 gnd
port 514 nsew
rlabel metal2 s 12240 27887 12240 27887 4 gnd
port 514 nsew
rlabel metal2 s 10224 26623 10224 26623 4 gnd
port 514 nsew
rlabel metal2 s 11472 27413 11472 27413 4 gnd
port 514 nsew
rlabel metal2 s 10224 26070 10224 26070 4 gnd
port 514 nsew
rlabel metal2 s 10992 27650 10992 27650 4 gnd
port 514 nsew
rlabel metal2 s 10224 25517 10224 25517 4 gnd
port 514 nsew
rlabel metal2 s 12240 26307 12240 26307 4 gnd
port 514 nsew
rlabel metal2 s 12240 28440 12240 28440 4 gnd
port 514 nsew
rlabel metal2 s 10992 25517 10992 25517 4 gnd
port 514 nsew
rlabel metal2 s 11472 25833 11472 25833 4 gnd
port 514 nsew
rlabel metal2 s 11472 27887 11472 27887 4 gnd
port 514 nsew
rlabel metal2 s 10992 27097 10992 27097 4 gnd
port 514 nsew
rlabel metal2 s 10992 25833 10992 25833 4 gnd
port 514 nsew
rlabel metal2 s 12240 25517 12240 25517 4 gnd
port 514 nsew
rlabel metal2 s 10992 26307 10992 26307 4 gnd
port 514 nsew
rlabel metal2 s 13968 27097 13968 27097 4 gnd
port 514 nsew
rlabel metal2 s 13488 27887 13488 27887 4 gnd
port 514 nsew
rlabel metal2 s 12720 26070 12720 26070 4 gnd
port 514 nsew
rlabel metal2 s 12720 26623 12720 26623 4 gnd
port 514 nsew
rlabel metal2 s 13968 25833 13968 25833 4 gnd
port 514 nsew
rlabel metal2 s 13488 27097 13488 27097 4 gnd
port 514 nsew
rlabel metal2 s 14736 26307 14736 26307 4 gnd
port 514 nsew
rlabel metal2 s 12720 25833 12720 25833 4 gnd
port 514 nsew
rlabel metal2 s 14736 27887 14736 27887 4 gnd
port 514 nsew
rlabel metal2 s 13968 27887 13968 27887 4 gnd
port 514 nsew
rlabel metal2 s 13488 26623 13488 26623 4 gnd
port 514 nsew
rlabel metal2 s 13488 27413 13488 27413 4 gnd
port 514 nsew
rlabel metal2 s 13488 27650 13488 27650 4 gnd
port 514 nsew
rlabel metal2 s 13488 26307 13488 26307 4 gnd
port 514 nsew
rlabel metal2 s 13968 26307 13968 26307 4 gnd
port 514 nsew
rlabel metal2 s 13488 28203 13488 28203 4 gnd
port 514 nsew
rlabel metal2 s 13968 27650 13968 27650 4 gnd
port 514 nsew
rlabel metal2 s 12720 27413 12720 27413 4 gnd
port 514 nsew
rlabel metal2 s 12720 26860 12720 26860 4 gnd
port 514 nsew
rlabel metal2 s 12720 27887 12720 27887 4 gnd
port 514 nsew
rlabel metal2 s 14736 27413 14736 27413 4 gnd
port 514 nsew
rlabel metal2 s 12720 28440 12720 28440 4 gnd
port 514 nsew
rlabel metal2 s 13968 26860 13968 26860 4 gnd
port 514 nsew
rlabel metal2 s 13488 25517 13488 25517 4 gnd
port 514 nsew
rlabel metal2 s 12720 25517 12720 25517 4 gnd
port 514 nsew
rlabel metal2 s 13488 28440 13488 28440 4 gnd
port 514 nsew
rlabel metal2 s 13488 25833 13488 25833 4 gnd
port 514 nsew
rlabel metal2 s 12720 27097 12720 27097 4 gnd
port 514 nsew
rlabel metal2 s 13968 28440 13968 28440 4 gnd
port 514 nsew
rlabel metal2 s 14736 26070 14736 26070 4 gnd
port 514 nsew
rlabel metal2 s 14736 27097 14736 27097 4 gnd
port 514 nsew
rlabel metal2 s 13968 28203 13968 28203 4 gnd
port 514 nsew
rlabel metal2 s 12720 28203 12720 28203 4 gnd
port 514 nsew
rlabel metal2 s 13488 26070 13488 26070 4 gnd
port 514 nsew
rlabel metal2 s 14736 28203 14736 28203 4 gnd
port 514 nsew
rlabel metal2 s 12720 27650 12720 27650 4 gnd
port 514 nsew
rlabel metal2 s 13968 25517 13968 25517 4 gnd
port 514 nsew
rlabel metal2 s 14736 26623 14736 26623 4 gnd
port 514 nsew
rlabel metal2 s 13488 26860 13488 26860 4 gnd
port 514 nsew
rlabel metal2 s 14736 27650 14736 27650 4 gnd
port 514 nsew
rlabel metal2 s 13968 26623 13968 26623 4 gnd
port 514 nsew
rlabel metal2 s 14736 28440 14736 28440 4 gnd
port 514 nsew
rlabel metal2 s 13968 27413 13968 27413 4 gnd
port 514 nsew
rlabel metal2 s 13968 26070 13968 26070 4 gnd
port 514 nsew
rlabel metal2 s 14736 25517 14736 25517 4 gnd
port 514 nsew
rlabel metal2 s 14736 25833 14736 25833 4 gnd
port 514 nsew
rlabel metal2 s 12720 26307 12720 26307 4 gnd
port 514 nsew
rlabel metal2 s 14736 26860 14736 26860 4 gnd
port 514 nsew
rlabel metal2 s 18480 30020 18480 30020 4 gnd
port 514 nsew
rlabel metal2 s 19968 29673 19968 29673 4 wl0_75
port 407 nsew
rlabel metal2 s 19728 30257 19728 30257 4 gnd
port 514 nsew
rlabel metal2 s 19728 30810 19728 30810 4 gnd
port 514 nsew
rlabel metal2 s 18960 29230 18960 29230 4 gnd
port 514 nsew
rlabel metal2 s 19728 29783 19728 29783 4 gnd
port 514 nsew
rlabel metal2 s 17712 30573 17712 30573 4 gnd
port 514 nsew
rlabel metal2 s 17712 29783 17712 29783 4 gnd
port 514 nsew
rlabel metal2 s 18960 30810 18960 30810 4 gnd
port 514 nsew
rlabel metal2 s 18480 31363 18480 31363 4 gnd
port 514 nsew
rlabel metal2 s 18960 30257 18960 30257 4 gnd
port 514 nsew
rlabel metal2 s 18480 30257 18480 30257 4 gnd
port 514 nsew
rlabel metal2 s 17712 31363 17712 31363 4 gnd
port 514 nsew
rlabel metal2 s 18960 28993 18960 28993 4 gnd
port 514 nsew
rlabel metal2 s 18480 31047 18480 31047 4 gnd
port 514 nsew
rlabel metal2 s 18960 28677 18960 28677 4 gnd
port 514 nsew
rlabel metal2 s 17712 31600 17712 31600 4 gnd
port 514 nsew
rlabel metal2 s 19728 31363 19728 31363 4 gnd
port 514 nsew
rlabel metal2 s 18480 30573 18480 30573 4 gnd
port 514 nsew
rlabel metal2 s 17712 30810 17712 30810 4 gnd
port 514 nsew
rlabel metal2 s 17712 28677 17712 28677 4 gnd
port 514 nsew
rlabel metal2 s 17712 30257 17712 30257 4 gnd
port 514 nsew
rlabel metal2 s 17712 29230 17712 29230 4 gnd
port 514 nsew
rlabel metal2 s 19728 29467 19728 29467 4 gnd
port 514 nsew
rlabel metal2 s 19728 28677 19728 28677 4 gnd
port 514 nsew
rlabel metal2 s 18960 31047 18960 31047 4 gnd
port 514 nsew
rlabel metal2 s 18960 30020 18960 30020 4 gnd
port 514 nsew
rlabel metal2 s 19728 30020 19728 30020 4 gnd
port 514 nsew
rlabel metal2 s 18480 28993 18480 28993 4 gnd
port 514 nsew
rlabel metal2 s 18480 28677 18480 28677 4 gnd
port 514 nsew
rlabel metal2 s 19968 30463 19968 30463 4 wl0_77
port 411 nsew
rlabel metal2 s 19968 30683 19968 30683 4 wl1_77
port 412 nsew
rlabel metal2 s 19968 29103 19968 29103 4 wl1_73
port 404 nsew
rlabel metal2 s 18480 29230 18480 29230 4 gnd
port 514 nsew
rlabel metal2 s 18960 30573 18960 30573 4 gnd
port 514 nsew
rlabel metal2 s 19968 28787 19968 28787 4 wl0_72
port 401 nsew
rlabel metal2 s 17712 28993 17712 28993 4 gnd
port 514 nsew
rlabel metal2 s 17712 30020 17712 30020 4 gnd
port 514 nsew
rlabel metal2 s 19968 31157 19968 31157 4 wl0_78
port 413 nsew
rlabel metal2 s 19968 30367 19968 30367 4 wl0_76
port 409 nsew
rlabel metal2 s 19728 31600 19728 31600 4 gnd
port 514 nsew
rlabel metal2 s 18480 29783 18480 29783 4 gnd
port 514 nsew
rlabel metal2 s 19968 28883 19968 28883 4 wl0_73
port 403 nsew
rlabel metal2 s 19968 28567 19968 28567 4 wl1_72
port 402 nsew
rlabel metal2 s 19968 29577 19968 29577 4 wl0_74
port 405 nsew
rlabel metal2 s 18960 31363 18960 31363 4 gnd
port 514 nsew
rlabel metal2 s 18960 29467 18960 29467 4 gnd
port 514 nsew
rlabel metal2 s 19968 31473 19968 31473 4 wl1_79
port 416 nsew
rlabel metal2 s 19728 28993 19728 28993 4 gnd
port 514 nsew
rlabel metal2 s 19968 29357 19968 29357 4 wl1_74
port 406 nsew
rlabel metal2 s 19968 31253 19968 31253 4 wl0_79
port 415 nsew
rlabel metal2 s 18960 31600 18960 31600 4 gnd
port 514 nsew
rlabel metal2 s 17712 31047 17712 31047 4 gnd
port 514 nsew
rlabel metal2 s 17712 29467 17712 29467 4 gnd
port 514 nsew
rlabel metal2 s 19968 30147 19968 30147 4 wl1_76
port 410 nsew
rlabel metal2 s 19728 29230 19728 29230 4 gnd
port 514 nsew
rlabel metal2 s 19968 30937 19968 30937 4 wl1_78
port 414 nsew
rlabel metal2 s 18480 30810 18480 30810 4 gnd
port 514 nsew
rlabel metal2 s 19728 30573 19728 30573 4 gnd
port 514 nsew
rlabel metal2 s 18480 29467 18480 29467 4 gnd
port 514 nsew
rlabel metal2 s 18480 31600 18480 31600 4 gnd
port 514 nsew
rlabel metal2 s 19728 31047 19728 31047 4 gnd
port 514 nsew
rlabel metal2 s 18960 29783 18960 29783 4 gnd
port 514 nsew
rlabel metal2 s 19968 29893 19968 29893 4 wl1_75
port 408 nsew
rlabel metal2 s 15216 30573 15216 30573 4 gnd
port 514 nsew
rlabel metal2 s 17232 28993 17232 28993 4 gnd
port 514 nsew
rlabel metal2 s 15984 31600 15984 31600 4 gnd
port 514 nsew
rlabel metal2 s 16464 30257 16464 30257 4 gnd
port 514 nsew
rlabel metal2 s 16464 30573 16464 30573 4 gnd
port 514 nsew
rlabel metal2 s 15216 28677 15216 28677 4 gnd
port 514 nsew
rlabel metal2 s 15216 31047 15216 31047 4 gnd
port 514 nsew
rlabel metal2 s 15216 30020 15216 30020 4 gnd
port 514 nsew
rlabel metal2 s 16464 29783 16464 29783 4 gnd
port 514 nsew
rlabel metal2 s 15216 29783 15216 29783 4 gnd
port 514 nsew
rlabel metal2 s 15984 30257 15984 30257 4 gnd
port 514 nsew
rlabel metal2 s 16464 31047 16464 31047 4 gnd
port 514 nsew
rlabel metal2 s 16464 29230 16464 29230 4 gnd
port 514 nsew
rlabel metal2 s 16464 31363 16464 31363 4 gnd
port 514 nsew
rlabel metal2 s 15216 28993 15216 28993 4 gnd
port 514 nsew
rlabel metal2 s 15984 29230 15984 29230 4 gnd
port 514 nsew
rlabel metal2 s 15216 31600 15216 31600 4 gnd
port 514 nsew
rlabel metal2 s 17232 30810 17232 30810 4 gnd
port 514 nsew
rlabel metal2 s 17232 31600 17232 31600 4 gnd
port 514 nsew
rlabel metal2 s 17232 28677 17232 28677 4 gnd
port 514 nsew
rlabel metal2 s 15984 30573 15984 30573 4 gnd
port 514 nsew
rlabel metal2 s 15216 30810 15216 30810 4 gnd
port 514 nsew
rlabel metal2 s 17232 29467 17232 29467 4 gnd
port 514 nsew
rlabel metal2 s 15984 29467 15984 29467 4 gnd
port 514 nsew
rlabel metal2 s 17232 29783 17232 29783 4 gnd
port 514 nsew
rlabel metal2 s 16464 30810 16464 30810 4 gnd
port 514 nsew
rlabel metal2 s 17232 31363 17232 31363 4 gnd
port 514 nsew
rlabel metal2 s 16464 30020 16464 30020 4 gnd
port 514 nsew
rlabel metal2 s 16464 31600 16464 31600 4 gnd
port 514 nsew
rlabel metal2 s 15984 28677 15984 28677 4 gnd
port 514 nsew
rlabel metal2 s 15984 31047 15984 31047 4 gnd
port 514 nsew
rlabel metal2 s 15984 29783 15984 29783 4 gnd
port 514 nsew
rlabel metal2 s 15984 31363 15984 31363 4 gnd
port 514 nsew
rlabel metal2 s 15216 31363 15216 31363 4 gnd
port 514 nsew
rlabel metal2 s 17232 29230 17232 29230 4 gnd
port 514 nsew
rlabel metal2 s 17232 30573 17232 30573 4 gnd
port 514 nsew
rlabel metal2 s 15216 29467 15216 29467 4 gnd
port 514 nsew
rlabel metal2 s 17232 30020 17232 30020 4 gnd
port 514 nsew
rlabel metal2 s 17232 30257 17232 30257 4 gnd
port 514 nsew
rlabel metal2 s 15216 29230 15216 29230 4 gnd
port 514 nsew
rlabel metal2 s 15984 30810 15984 30810 4 gnd
port 514 nsew
rlabel metal2 s 16464 28993 16464 28993 4 gnd
port 514 nsew
rlabel metal2 s 17232 31047 17232 31047 4 gnd
port 514 nsew
rlabel metal2 s 15984 30020 15984 30020 4 gnd
port 514 nsew
rlabel metal2 s 15216 30257 15216 30257 4 gnd
port 514 nsew
rlabel metal2 s 16464 28677 16464 28677 4 gnd
port 514 nsew
rlabel metal2 s 15984 28993 15984 28993 4 gnd
port 514 nsew
rlabel metal2 s 16464 29467 16464 29467 4 gnd
port 514 nsew
rlabel metal2 s 16464 27650 16464 27650 4 gnd
port 514 nsew
rlabel metal2 s 17232 26860 17232 26860 4 gnd
port 514 nsew
rlabel metal2 s 15216 27650 15216 27650 4 gnd
port 514 nsew
rlabel metal2 s 17232 27887 17232 27887 4 gnd
port 514 nsew
rlabel metal2 s 15216 26623 15216 26623 4 gnd
port 514 nsew
rlabel metal2 s 15216 27097 15216 27097 4 gnd
port 514 nsew
rlabel metal2 s 15216 25833 15216 25833 4 gnd
port 514 nsew
rlabel metal2 s 15216 27413 15216 27413 4 gnd
port 514 nsew
rlabel metal2 s 16464 26307 16464 26307 4 gnd
port 514 nsew
rlabel metal2 s 17232 27650 17232 27650 4 gnd
port 514 nsew
rlabel metal2 s 17232 25517 17232 25517 4 gnd
port 514 nsew
rlabel metal2 s 17232 28203 17232 28203 4 gnd
port 514 nsew
rlabel metal2 s 16464 26623 16464 26623 4 gnd
port 514 nsew
rlabel metal2 s 15984 27650 15984 27650 4 gnd
port 514 nsew
rlabel metal2 s 17232 26307 17232 26307 4 gnd
port 514 nsew
rlabel metal2 s 15216 26860 15216 26860 4 gnd
port 514 nsew
rlabel metal2 s 17232 27097 17232 27097 4 gnd
port 514 nsew
rlabel metal2 s 15984 25833 15984 25833 4 gnd
port 514 nsew
rlabel metal2 s 15216 28203 15216 28203 4 gnd
port 514 nsew
rlabel metal2 s 17232 26070 17232 26070 4 gnd
port 514 nsew
rlabel metal2 s 16464 26860 16464 26860 4 gnd
port 514 nsew
rlabel metal2 s 15984 25517 15984 25517 4 gnd
port 514 nsew
rlabel metal2 s 15216 28440 15216 28440 4 gnd
port 514 nsew
rlabel metal2 s 15984 28440 15984 28440 4 gnd
port 514 nsew
rlabel metal2 s 15216 25517 15216 25517 4 gnd
port 514 nsew
rlabel metal2 s 17232 26623 17232 26623 4 gnd
port 514 nsew
rlabel metal2 s 17232 28440 17232 28440 4 gnd
port 514 nsew
rlabel metal2 s 16464 27413 16464 27413 4 gnd
port 514 nsew
rlabel metal2 s 15984 26860 15984 26860 4 gnd
port 514 nsew
rlabel metal2 s 15984 26307 15984 26307 4 gnd
port 514 nsew
rlabel metal2 s 16464 25833 16464 25833 4 gnd
port 514 nsew
rlabel metal2 s 15216 27887 15216 27887 4 gnd
port 514 nsew
rlabel metal2 s 17232 25833 17232 25833 4 gnd
port 514 nsew
rlabel metal2 s 16464 28440 16464 28440 4 gnd
port 514 nsew
rlabel metal2 s 16464 26070 16464 26070 4 gnd
port 514 nsew
rlabel metal2 s 15216 26070 15216 26070 4 gnd
port 514 nsew
rlabel metal2 s 15984 26623 15984 26623 4 gnd
port 514 nsew
rlabel metal2 s 16464 28203 16464 28203 4 gnd
port 514 nsew
rlabel metal2 s 16464 25517 16464 25517 4 gnd
port 514 nsew
rlabel metal2 s 16464 27887 16464 27887 4 gnd
port 514 nsew
rlabel metal2 s 15216 26307 15216 26307 4 gnd
port 514 nsew
rlabel metal2 s 16464 27097 16464 27097 4 gnd
port 514 nsew
rlabel metal2 s 15984 27887 15984 27887 4 gnd
port 514 nsew
rlabel metal2 s 15984 27097 15984 27097 4 gnd
port 514 nsew
rlabel metal2 s 15984 26070 15984 26070 4 gnd
port 514 nsew
rlabel metal2 s 15984 28203 15984 28203 4 gnd
port 514 nsew
rlabel metal2 s 15984 27413 15984 27413 4 gnd
port 514 nsew
rlabel metal2 s 17232 27413 17232 27413 4 gnd
port 514 nsew
rlabel metal2 s 19968 26197 19968 26197 4 wl1_66
port 390 nsew
rlabel metal2 s 19968 26513 19968 26513 4 wl0_67
port 391 nsew
rlabel metal2 s 19968 27997 19968 27997 4 wl0_70
port 397 nsew
rlabel metal2 s 18960 25517 18960 25517 4 gnd
port 514 nsew
rlabel metal2 s 19968 25627 19968 25627 4 wl0_64
port 385 nsew
rlabel metal2 s 18480 26070 18480 26070 4 gnd
port 514 nsew
rlabel metal2 s 19728 26307 19728 26307 4 gnd
port 514 nsew
rlabel metal2 s 17712 28440 17712 28440 4 gnd
port 514 nsew
rlabel metal2 s 19728 25517 19728 25517 4 gnd
port 514 nsew
rlabel metal2 s 18960 26623 18960 26623 4 gnd
port 514 nsew
rlabel metal2 s 18480 28203 18480 28203 4 gnd
port 514 nsew
rlabel metal2 s 19728 28440 19728 28440 4 gnd
port 514 nsew
rlabel metal2 s 17712 27650 17712 27650 4 gnd
port 514 nsew
rlabel metal2 s 18960 28203 18960 28203 4 gnd
port 514 nsew
rlabel metal2 s 18960 25833 18960 25833 4 gnd
port 514 nsew
rlabel metal2 s 17712 25833 17712 25833 4 gnd
port 514 nsew
rlabel metal2 s 18960 27650 18960 27650 4 gnd
port 514 nsew
rlabel metal2 s 18960 28440 18960 28440 4 gnd
port 514 nsew
rlabel metal2 s 18480 27413 18480 27413 4 gnd
port 514 nsew
rlabel metal2 s 17712 28203 17712 28203 4 gnd
port 514 nsew
rlabel metal2 s 19968 26733 19968 26733 4 wl1_67
port 392 nsew
rlabel metal2 s 18480 27650 18480 27650 4 gnd
port 514 nsew
rlabel metal2 s 19728 26860 19728 26860 4 gnd
port 514 nsew
rlabel metal2 s 19968 26417 19968 26417 4 wl0_66
port 389 nsew
rlabel metal2 s 19728 27887 19728 27887 4 gnd
port 514 nsew
rlabel metal2 s 17712 26307 17712 26307 4 gnd
port 514 nsew
rlabel metal2 s 18960 27413 18960 27413 4 gnd
port 514 nsew
rlabel metal2 s 19968 25943 19968 25943 4 wl1_65
port 388 nsew
rlabel metal2 s 17712 25517 17712 25517 4 gnd
port 514 nsew
rlabel metal2 s 18480 26623 18480 26623 4 gnd
port 514 nsew
rlabel metal2 s 18480 25517 18480 25517 4 gnd
port 514 nsew
rlabel metal2 s 19968 27207 19968 27207 4 wl0_68
port 393 nsew
rlabel metal2 s 19728 25833 19728 25833 4 gnd
port 514 nsew
rlabel metal2 s 17712 26623 17712 26623 4 gnd
port 514 nsew
rlabel metal2 s 19968 25723 19968 25723 4 wl0_65
port 387 nsew
rlabel metal2 s 18480 28440 18480 28440 4 gnd
port 514 nsew
rlabel metal2 s 18960 27097 18960 27097 4 gnd
port 514 nsew
rlabel metal2 s 19968 27777 19968 27777 4 wl1_70
port 398 nsew
rlabel metal2 s 18480 25833 18480 25833 4 gnd
port 514 nsew
rlabel metal2 s 18480 26860 18480 26860 4 gnd
port 514 nsew
rlabel metal2 s 19968 26987 19968 26987 4 wl1_68
port 394 nsew
rlabel metal2 s 17712 27097 17712 27097 4 gnd
port 514 nsew
rlabel metal2 s 19728 26623 19728 26623 4 gnd
port 514 nsew
rlabel metal2 s 18960 26860 18960 26860 4 gnd
port 514 nsew
rlabel metal2 s 17712 26860 17712 26860 4 gnd
port 514 nsew
rlabel metal2 s 17712 27413 17712 27413 4 gnd
port 514 nsew
rlabel metal2 s 19968 27303 19968 27303 4 wl0_69
port 395 nsew
rlabel metal2 s 19728 27413 19728 27413 4 gnd
port 514 nsew
rlabel metal2 s 17712 26070 17712 26070 4 gnd
port 514 nsew
rlabel metal2 s 19968 28313 19968 28313 4 wl1_71
port 400 nsew
rlabel metal2 s 18960 26307 18960 26307 4 gnd
port 514 nsew
rlabel metal2 s 18960 26070 18960 26070 4 gnd
port 514 nsew
rlabel metal2 s 19968 28093 19968 28093 4 wl0_71
port 399 nsew
rlabel metal2 s 18480 27887 18480 27887 4 gnd
port 514 nsew
rlabel metal2 s 17712 27887 17712 27887 4 gnd
port 514 nsew
rlabel metal2 s 19728 27650 19728 27650 4 gnd
port 514 nsew
rlabel metal2 s 19728 26070 19728 26070 4 gnd
port 514 nsew
rlabel metal2 s 18480 27097 18480 27097 4 gnd
port 514 nsew
rlabel metal2 s 19728 28203 19728 28203 4 gnd
port 514 nsew
rlabel metal2 s 19728 27097 19728 27097 4 gnd
port 514 nsew
rlabel metal2 s 19968 27523 19968 27523 4 wl1_69
port 396 nsew
rlabel metal2 s 18480 26307 18480 26307 4 gnd
port 514 nsew
rlabel metal2 s 18960 27887 18960 27887 4 gnd
port 514 nsew
rlabel metal2 s 19968 25407 19968 25407 4 wl1_64
port 386 nsew
rlabel metal2 s 18960 23463 18960 23463 4 gnd
port 514 nsew
rlabel metal2 s 19728 25043 19728 25043 4 gnd
port 514 nsew
rlabel metal2 s 19728 24490 19728 24490 4 gnd
port 514 nsew
rlabel metal2 s 19728 24727 19728 24727 4 gnd
port 514 nsew
rlabel metal2 s 17712 23700 17712 23700 4 gnd
port 514 nsew
rlabel metal2 s 18480 24253 18480 24253 4 gnd
port 514 nsew
rlabel metal2 s 19968 23037 19968 23037 4 wl1_58
port 374 nsew
rlabel metal2 s 18480 22673 18480 22673 4 gnd
port 514 nsew
rlabel metal2 s 18960 22673 18960 22673 4 gnd
port 514 nsew
rlabel metal2 s 19968 24047 19968 24047 4 wl0_60
port 377 nsew
rlabel metal2 s 17712 22673 17712 22673 4 gnd
port 514 nsew
rlabel metal2 s 19728 25280 19728 25280 4 gnd
port 514 nsew
rlabel metal2 s 18960 24253 18960 24253 4 gnd
port 514 nsew
rlabel metal2 s 18960 23700 18960 23700 4 gnd
port 514 nsew
rlabel metal2 s 17712 25043 17712 25043 4 gnd
port 514 nsew
rlabel metal2 s 17712 22910 17712 22910 4 gnd
port 514 nsew
rlabel metal2 s 19728 24253 19728 24253 4 gnd
port 514 nsew
rlabel metal2 s 19968 25153 19968 25153 4 wl1_63
port 384 nsew
rlabel metal2 s 17712 22357 17712 22357 4 gnd
port 514 nsew
rlabel metal2 s 18480 24727 18480 24727 4 gnd
port 514 nsew
rlabel metal2 s 19968 24617 19968 24617 4 wl1_62
port 382 nsew
rlabel metal2 s 18960 25043 18960 25043 4 gnd
port 514 nsew
rlabel metal2 s 17712 25280 17712 25280 4 gnd
port 514 nsew
rlabel metal2 s 18960 25280 18960 25280 4 gnd
port 514 nsew
rlabel metal2 s 17712 23147 17712 23147 4 gnd
port 514 nsew
rlabel metal2 s 18480 23700 18480 23700 4 gnd
port 514 nsew
rlabel metal2 s 19968 24933 19968 24933 4 wl0_63
port 383 nsew
rlabel metal2 s 18960 22910 18960 22910 4 gnd
port 514 nsew
rlabel metal2 s 17712 24253 17712 24253 4 gnd
port 514 nsew
rlabel metal2 s 18480 25043 18480 25043 4 gnd
port 514 nsew
rlabel metal2 s 18480 23937 18480 23937 4 gnd
port 514 nsew
rlabel metal2 s 19728 23700 19728 23700 4 gnd
port 514 nsew
rlabel metal2 s 19728 23463 19728 23463 4 gnd
port 514 nsew
rlabel metal2 s 18480 22357 18480 22357 4 gnd
port 514 nsew
rlabel metal2 s 18960 24727 18960 24727 4 gnd
port 514 nsew
rlabel metal2 s 19968 23257 19968 23257 4 wl0_58
port 373 nsew
rlabel metal2 s 18960 22357 18960 22357 4 gnd
port 514 nsew
rlabel metal2 s 18480 22910 18480 22910 4 gnd
port 514 nsew
rlabel metal2 s 19728 23147 19728 23147 4 gnd
port 514 nsew
rlabel metal2 s 17712 24490 17712 24490 4 gnd
port 514 nsew
rlabel metal2 s 18480 24490 18480 24490 4 gnd
port 514 nsew
rlabel metal2 s 18480 25280 18480 25280 4 gnd
port 514 nsew
rlabel metal2 s 19728 22910 19728 22910 4 gnd
port 514 nsew
rlabel metal2 s 19728 23937 19728 23937 4 gnd
port 514 nsew
rlabel metal2 s 18960 23937 18960 23937 4 gnd
port 514 nsew
rlabel metal2 s 19728 22357 19728 22357 4 gnd
port 514 nsew
rlabel metal2 s 18480 23147 18480 23147 4 gnd
port 514 nsew
rlabel metal2 s 18960 24490 18960 24490 4 gnd
port 514 nsew
rlabel metal2 s 17712 23937 17712 23937 4 gnd
port 514 nsew
rlabel metal2 s 17712 23463 17712 23463 4 gnd
port 514 nsew
rlabel metal2 s 19728 22673 19728 22673 4 gnd
port 514 nsew
rlabel metal2 s 17712 24727 17712 24727 4 gnd
port 514 nsew
rlabel metal2 s 18960 23147 18960 23147 4 gnd
port 514 nsew
rlabel metal2 s 18480 23463 18480 23463 4 gnd
port 514 nsew
rlabel metal2 s 19968 22467 19968 22467 4 wl0_56
port 369 nsew
rlabel metal2 s 19968 23827 19968 23827 4 wl1_60
port 378 nsew
rlabel metal2 s 19968 24837 19968 24837 4 wl0_62
port 381 nsew
rlabel metal2 s 19968 22563 19968 22563 4 wl0_57
port 371 nsew
rlabel metal2 s 19968 24363 19968 24363 4 wl1_61
port 380 nsew
rlabel metal2 s 19968 23353 19968 23353 4 wl0_59
port 375 nsew
rlabel metal2 s 19968 23573 19968 23573 4 wl1_59
port 376 nsew
rlabel metal2 s 19968 22783 19968 22783 4 wl1_57
port 372 nsew
rlabel metal2 s 19968 22247 19968 22247 4 wl1_56
port 370 nsew
rlabel metal2 s 19968 24143 19968 24143 4 wl0_61
port 379 nsew
rlabel metal2 s 15984 25280 15984 25280 4 gnd
port 514 nsew
rlabel metal2 s 17232 23147 17232 23147 4 gnd
port 514 nsew
rlabel metal2 s 15216 22910 15216 22910 4 gnd
port 514 nsew
rlabel metal2 s 15216 25280 15216 25280 4 gnd
port 514 nsew
rlabel metal2 s 16464 22673 16464 22673 4 gnd
port 514 nsew
rlabel metal2 s 15984 22673 15984 22673 4 gnd
port 514 nsew
rlabel metal2 s 15984 25043 15984 25043 4 gnd
port 514 nsew
rlabel metal2 s 16464 23463 16464 23463 4 gnd
port 514 nsew
rlabel metal2 s 16464 22910 16464 22910 4 gnd
port 514 nsew
rlabel metal2 s 16464 23700 16464 23700 4 gnd
port 514 nsew
rlabel metal2 s 15216 22673 15216 22673 4 gnd
port 514 nsew
rlabel metal2 s 16464 24253 16464 24253 4 gnd
port 514 nsew
rlabel metal2 s 16464 23937 16464 23937 4 gnd
port 514 nsew
rlabel metal2 s 15984 22910 15984 22910 4 gnd
port 514 nsew
rlabel metal2 s 15216 23700 15216 23700 4 gnd
port 514 nsew
rlabel metal2 s 15984 23700 15984 23700 4 gnd
port 514 nsew
rlabel metal2 s 17232 25043 17232 25043 4 gnd
port 514 nsew
rlabel metal2 s 15984 23937 15984 23937 4 gnd
port 514 nsew
rlabel metal2 s 17232 24727 17232 24727 4 gnd
port 514 nsew
rlabel metal2 s 17232 24490 17232 24490 4 gnd
port 514 nsew
rlabel metal2 s 15984 23147 15984 23147 4 gnd
port 514 nsew
rlabel metal2 s 16464 25043 16464 25043 4 gnd
port 514 nsew
rlabel metal2 s 17232 24253 17232 24253 4 gnd
port 514 nsew
rlabel metal2 s 15984 23463 15984 23463 4 gnd
port 514 nsew
rlabel metal2 s 17232 22910 17232 22910 4 gnd
port 514 nsew
rlabel metal2 s 16464 22357 16464 22357 4 gnd
port 514 nsew
rlabel metal2 s 17232 25280 17232 25280 4 gnd
port 514 nsew
rlabel metal2 s 15216 23463 15216 23463 4 gnd
port 514 nsew
rlabel metal2 s 15216 24490 15216 24490 4 gnd
port 514 nsew
rlabel metal2 s 15216 24727 15216 24727 4 gnd
port 514 nsew
rlabel metal2 s 16464 24490 16464 24490 4 gnd
port 514 nsew
rlabel metal2 s 15984 24253 15984 24253 4 gnd
port 514 nsew
rlabel metal2 s 17232 23937 17232 23937 4 gnd
port 514 nsew
rlabel metal2 s 15984 24727 15984 24727 4 gnd
port 514 nsew
rlabel metal2 s 15984 24490 15984 24490 4 gnd
port 514 nsew
rlabel metal2 s 17232 22673 17232 22673 4 gnd
port 514 nsew
rlabel metal2 s 15216 24253 15216 24253 4 gnd
port 514 nsew
rlabel metal2 s 15216 25043 15216 25043 4 gnd
port 514 nsew
rlabel metal2 s 17232 23700 17232 23700 4 gnd
port 514 nsew
rlabel metal2 s 15216 23937 15216 23937 4 gnd
port 514 nsew
rlabel metal2 s 16464 25280 16464 25280 4 gnd
port 514 nsew
rlabel metal2 s 15984 22357 15984 22357 4 gnd
port 514 nsew
rlabel metal2 s 16464 23147 16464 23147 4 gnd
port 514 nsew
rlabel metal2 s 17232 23463 17232 23463 4 gnd
port 514 nsew
rlabel metal2 s 17232 22357 17232 22357 4 gnd
port 514 nsew
rlabel metal2 s 15216 22357 15216 22357 4 gnd
port 514 nsew
rlabel metal2 s 16464 24727 16464 24727 4 gnd
port 514 nsew
rlabel metal2 s 15216 23147 15216 23147 4 gnd
port 514 nsew
rlabel metal2 s 15216 21330 15216 21330 4 gnd
port 514 nsew
rlabel metal2 s 17232 22120 17232 22120 4 gnd
port 514 nsew
rlabel metal2 s 17232 19197 17232 19197 4 gnd
port 514 nsew
rlabel metal2 s 15216 21093 15216 21093 4 gnd
port 514 nsew
rlabel metal2 s 15984 19513 15984 19513 4 gnd
port 514 nsew
rlabel metal2 s 17232 20303 17232 20303 4 gnd
port 514 nsew
rlabel metal2 s 16464 19513 16464 19513 4 gnd
port 514 nsew
rlabel metal2 s 17232 21567 17232 21567 4 gnd
port 514 nsew
rlabel metal2 s 17232 20540 17232 20540 4 gnd
port 514 nsew
rlabel metal2 s 15216 21883 15216 21883 4 gnd
port 514 nsew
rlabel metal2 s 15216 22120 15216 22120 4 gnd
port 514 nsew
rlabel metal2 s 16464 21330 16464 21330 4 gnd
port 514 nsew
rlabel metal2 s 16464 21883 16464 21883 4 gnd
port 514 nsew
rlabel metal2 s 15216 21567 15216 21567 4 gnd
port 514 nsew
rlabel metal2 s 16464 20303 16464 20303 4 gnd
port 514 nsew
rlabel metal2 s 15984 20540 15984 20540 4 gnd
port 514 nsew
rlabel metal2 s 15216 19513 15216 19513 4 gnd
port 514 nsew
rlabel metal2 s 15984 19197 15984 19197 4 gnd
port 514 nsew
rlabel metal2 s 17232 21883 17232 21883 4 gnd
port 514 nsew
rlabel metal2 s 15984 21567 15984 21567 4 gnd
port 514 nsew
rlabel metal2 s 15216 19987 15216 19987 4 gnd
port 514 nsew
rlabel metal2 s 16464 19750 16464 19750 4 gnd
port 514 nsew
rlabel metal2 s 16464 22120 16464 22120 4 gnd
port 514 nsew
rlabel metal2 s 15984 21330 15984 21330 4 gnd
port 514 nsew
rlabel metal2 s 16464 20777 16464 20777 4 gnd
port 514 nsew
rlabel metal2 s 15984 21093 15984 21093 4 gnd
port 514 nsew
rlabel metal2 s 17232 20777 17232 20777 4 gnd
port 514 nsew
rlabel metal2 s 17232 21330 17232 21330 4 gnd
port 514 nsew
rlabel metal2 s 15216 20777 15216 20777 4 gnd
port 514 nsew
rlabel metal2 s 16464 19987 16464 19987 4 gnd
port 514 nsew
rlabel metal2 s 15216 20540 15216 20540 4 gnd
port 514 nsew
rlabel metal2 s 15216 19750 15216 19750 4 gnd
port 514 nsew
rlabel metal2 s 15216 20303 15216 20303 4 gnd
port 514 nsew
rlabel metal2 s 15984 21883 15984 21883 4 gnd
port 514 nsew
rlabel metal2 s 15216 19197 15216 19197 4 gnd
port 514 nsew
rlabel metal2 s 15984 20777 15984 20777 4 gnd
port 514 nsew
rlabel metal2 s 17232 19513 17232 19513 4 gnd
port 514 nsew
rlabel metal2 s 17232 21093 17232 21093 4 gnd
port 514 nsew
rlabel metal2 s 16464 20540 16464 20540 4 gnd
port 514 nsew
rlabel metal2 s 16464 19197 16464 19197 4 gnd
port 514 nsew
rlabel metal2 s 15984 19987 15984 19987 4 gnd
port 514 nsew
rlabel metal2 s 15984 19750 15984 19750 4 gnd
port 514 nsew
rlabel metal2 s 17232 19750 17232 19750 4 gnd
port 514 nsew
rlabel metal2 s 16464 21093 16464 21093 4 gnd
port 514 nsew
rlabel metal2 s 15984 22120 15984 22120 4 gnd
port 514 nsew
rlabel metal2 s 15984 20303 15984 20303 4 gnd
port 514 nsew
rlabel metal2 s 16464 21567 16464 21567 4 gnd
port 514 nsew
rlabel metal2 s 17232 19987 17232 19987 4 gnd
port 514 nsew
rlabel metal2 s 17712 21567 17712 21567 4 gnd
port 514 nsew
rlabel metal2 s 18480 19987 18480 19987 4 gnd
port 514 nsew
rlabel metal2 s 19728 20303 19728 20303 4 gnd
port 514 nsew
rlabel metal2 s 18480 22120 18480 22120 4 gnd
port 514 nsew
rlabel metal2 s 18960 21093 18960 21093 4 gnd
port 514 nsew
rlabel metal2 s 19728 19750 19728 19750 4 gnd
port 514 nsew
rlabel metal2 s 18960 21567 18960 21567 4 gnd
port 514 nsew
rlabel metal2 s 18960 19197 18960 19197 4 gnd
port 514 nsew
rlabel metal2 s 19728 19197 19728 19197 4 gnd
port 514 nsew
rlabel metal2 s 19728 20777 19728 20777 4 gnd
port 514 nsew
rlabel metal2 s 18960 19750 18960 19750 4 gnd
port 514 nsew
rlabel metal2 s 17712 21330 17712 21330 4 gnd
port 514 nsew
rlabel metal2 s 18480 19750 18480 19750 4 gnd
port 514 nsew
rlabel metal2 s 19728 21567 19728 21567 4 gnd
port 514 nsew
rlabel metal2 s 18480 21883 18480 21883 4 gnd
port 514 nsew
rlabel metal2 s 18480 21330 18480 21330 4 gnd
port 514 nsew
rlabel metal2 s 19728 19987 19728 19987 4 gnd
port 514 nsew
rlabel metal2 s 19728 20540 19728 20540 4 gnd
port 514 nsew
rlabel metal2 s 18480 20540 18480 20540 4 gnd
port 514 nsew
rlabel metal2 s 17712 19513 17712 19513 4 gnd
port 514 nsew
rlabel metal2 s 18480 20777 18480 20777 4 gnd
port 514 nsew
rlabel metal2 s 19728 21330 19728 21330 4 gnd
port 514 nsew
rlabel metal2 s 19728 21093 19728 21093 4 gnd
port 514 nsew
rlabel metal2 s 18480 21093 18480 21093 4 gnd
port 514 nsew
rlabel metal2 s 18960 21883 18960 21883 4 gnd
port 514 nsew
rlabel metal2 s 18960 19987 18960 19987 4 gnd
port 514 nsew
rlabel metal2 s 19728 22120 19728 22120 4 gnd
port 514 nsew
rlabel metal2 s 18960 20303 18960 20303 4 gnd
port 514 nsew
rlabel metal2 s 17712 20540 17712 20540 4 gnd
port 514 nsew
rlabel metal2 s 17712 21883 17712 21883 4 gnd
port 514 nsew
rlabel metal2 s 17712 22120 17712 22120 4 gnd
port 514 nsew
rlabel metal2 s 18480 21567 18480 21567 4 gnd
port 514 nsew
rlabel metal2 s 19728 19513 19728 19513 4 gnd
port 514 nsew
rlabel metal2 s 19968 20667 19968 20667 4 wl1_52
port 362 nsew
rlabel metal2 s 19968 19877 19968 19877 4 wl1_50
port 358 nsew
rlabel metal2 s 18960 21330 18960 21330 4 gnd
port 514 nsew
rlabel metal2 s 17712 19197 17712 19197 4 gnd
port 514 nsew
rlabel metal2 s 19968 20413 19968 20413 4 wl1_51
port 360 nsew
rlabel metal2 s 18960 20777 18960 20777 4 gnd
port 514 nsew
rlabel metal2 s 18480 19197 18480 19197 4 gnd
port 514 nsew
rlabel metal2 s 19968 20887 19968 20887 4 wl0_52
port 361 nsew
rlabel metal2 s 19968 20097 19968 20097 4 wl0_50
port 357 nsew
rlabel metal2 s 19968 19087 19968 19087 4 wl1_48
port 354 nsew
rlabel metal2 s 19968 19403 19968 19403 4 wl0_49
port 355 nsew
rlabel metal2 s 18960 19513 18960 19513 4 gnd
port 514 nsew
rlabel metal2 s 19968 21203 19968 21203 4 wl1_53
port 364 nsew
rlabel metal2 s 18960 20540 18960 20540 4 gnd
port 514 nsew
rlabel metal2 s 19968 21457 19968 21457 4 wl1_54
port 366 nsew
rlabel metal2 s 19968 19623 19968 19623 4 wl1_49
port 356 nsew
rlabel metal2 s 19968 20193 19968 20193 4 wl0_51
port 359 nsew
rlabel metal2 s 19968 21677 19968 21677 4 wl0_54
port 365 nsew
rlabel metal2 s 19968 21773 19968 21773 4 wl0_55
port 367 nsew
rlabel metal2 s 18480 19513 18480 19513 4 gnd
port 514 nsew
rlabel metal2 s 17712 20777 17712 20777 4 gnd
port 514 nsew
rlabel metal2 s 19968 19307 19968 19307 4 wl0_48
port 353 nsew
rlabel metal2 s 19968 21993 19968 21993 4 wl1_55
port 368 nsew
rlabel metal2 s 17712 19987 17712 19987 4 gnd
port 514 nsew
rlabel metal2 s 17712 19750 17712 19750 4 gnd
port 514 nsew
rlabel metal2 s 17712 21093 17712 21093 4 gnd
port 514 nsew
rlabel metal2 s 18480 20303 18480 20303 4 gnd
port 514 nsew
rlabel metal2 s 18960 22120 18960 22120 4 gnd
port 514 nsew
rlabel metal2 s 19728 21883 19728 21883 4 gnd
port 514 nsew
rlabel metal2 s 17712 20303 17712 20303 4 gnd
port 514 nsew
rlabel metal2 s 19968 20983 19968 20983 4 wl0_53
port 363 nsew
rlabel metal2 s 13968 22673 13968 22673 4 gnd
port 514 nsew
rlabel metal2 s 13968 22357 13968 22357 4 gnd
port 514 nsew
rlabel metal2 s 12720 25043 12720 25043 4 gnd
port 514 nsew
rlabel metal2 s 14736 22357 14736 22357 4 gnd
port 514 nsew
rlabel metal2 s 13488 24253 13488 24253 4 gnd
port 514 nsew
rlabel metal2 s 12720 25280 12720 25280 4 gnd
port 514 nsew
rlabel metal2 s 12720 24490 12720 24490 4 gnd
port 514 nsew
rlabel metal2 s 14736 24253 14736 24253 4 gnd
port 514 nsew
rlabel metal2 s 14736 25280 14736 25280 4 gnd
port 514 nsew
rlabel metal2 s 14736 23147 14736 23147 4 gnd
port 514 nsew
rlabel metal2 s 13488 24727 13488 24727 4 gnd
port 514 nsew
rlabel metal2 s 13488 23700 13488 23700 4 gnd
port 514 nsew
rlabel metal2 s 13968 25043 13968 25043 4 gnd
port 514 nsew
rlabel metal2 s 13488 22357 13488 22357 4 gnd
port 514 nsew
rlabel metal2 s 14736 23700 14736 23700 4 gnd
port 514 nsew
rlabel metal2 s 13968 23937 13968 23937 4 gnd
port 514 nsew
rlabel metal2 s 13968 24490 13968 24490 4 gnd
port 514 nsew
rlabel metal2 s 14736 24490 14736 24490 4 gnd
port 514 nsew
rlabel metal2 s 13488 24490 13488 24490 4 gnd
port 514 nsew
rlabel metal2 s 13968 23147 13968 23147 4 gnd
port 514 nsew
rlabel metal2 s 14736 22673 14736 22673 4 gnd
port 514 nsew
rlabel metal2 s 13968 24727 13968 24727 4 gnd
port 514 nsew
rlabel metal2 s 13488 25043 13488 25043 4 gnd
port 514 nsew
rlabel metal2 s 13488 25280 13488 25280 4 gnd
port 514 nsew
rlabel metal2 s 12720 23700 12720 23700 4 gnd
port 514 nsew
rlabel metal2 s 12720 22673 12720 22673 4 gnd
port 514 nsew
rlabel metal2 s 12720 24253 12720 24253 4 gnd
port 514 nsew
rlabel metal2 s 13968 24253 13968 24253 4 gnd
port 514 nsew
rlabel metal2 s 13968 25280 13968 25280 4 gnd
port 514 nsew
rlabel metal2 s 13968 23700 13968 23700 4 gnd
port 514 nsew
rlabel metal2 s 14736 24727 14736 24727 4 gnd
port 514 nsew
rlabel metal2 s 12720 23463 12720 23463 4 gnd
port 514 nsew
rlabel metal2 s 14736 22910 14736 22910 4 gnd
port 514 nsew
rlabel metal2 s 13488 23147 13488 23147 4 gnd
port 514 nsew
rlabel metal2 s 13968 22910 13968 22910 4 gnd
port 514 nsew
rlabel metal2 s 12720 22357 12720 22357 4 gnd
port 514 nsew
rlabel metal2 s 12720 23937 12720 23937 4 gnd
port 514 nsew
rlabel metal2 s 14736 23937 14736 23937 4 gnd
port 514 nsew
rlabel metal2 s 12720 24727 12720 24727 4 gnd
port 514 nsew
rlabel metal2 s 12720 23147 12720 23147 4 gnd
port 514 nsew
rlabel metal2 s 13488 22910 13488 22910 4 gnd
port 514 nsew
rlabel metal2 s 13488 23937 13488 23937 4 gnd
port 514 nsew
rlabel metal2 s 12720 22910 12720 22910 4 gnd
port 514 nsew
rlabel metal2 s 13488 22673 13488 22673 4 gnd
port 514 nsew
rlabel metal2 s 14736 25043 14736 25043 4 gnd
port 514 nsew
rlabel metal2 s 14736 23463 14736 23463 4 gnd
port 514 nsew
rlabel metal2 s 13968 23463 13968 23463 4 gnd
port 514 nsew
rlabel metal2 s 13488 23463 13488 23463 4 gnd
port 514 nsew
rlabel metal2 s 12240 24253 12240 24253 4 gnd
port 514 nsew
rlabel metal2 s 10224 24490 10224 24490 4 gnd
port 514 nsew
rlabel metal2 s 11472 24490 11472 24490 4 gnd
port 514 nsew
rlabel metal2 s 10224 23937 10224 23937 4 gnd
port 514 nsew
rlabel metal2 s 11472 22673 11472 22673 4 gnd
port 514 nsew
rlabel metal2 s 10224 22357 10224 22357 4 gnd
port 514 nsew
rlabel metal2 s 10224 23463 10224 23463 4 gnd
port 514 nsew
rlabel metal2 s 11472 25280 11472 25280 4 gnd
port 514 nsew
rlabel metal2 s 11472 22910 11472 22910 4 gnd
port 514 nsew
rlabel metal2 s 10992 24253 10992 24253 4 gnd
port 514 nsew
rlabel metal2 s 10224 22673 10224 22673 4 gnd
port 514 nsew
rlabel metal2 s 12240 23700 12240 23700 4 gnd
port 514 nsew
rlabel metal2 s 12240 22910 12240 22910 4 gnd
port 514 nsew
rlabel metal2 s 10224 23147 10224 23147 4 gnd
port 514 nsew
rlabel metal2 s 10992 23147 10992 23147 4 gnd
port 514 nsew
rlabel metal2 s 10224 24253 10224 24253 4 gnd
port 514 nsew
rlabel metal2 s 12240 23463 12240 23463 4 gnd
port 514 nsew
rlabel metal2 s 10992 25043 10992 25043 4 gnd
port 514 nsew
rlabel metal2 s 10992 22910 10992 22910 4 gnd
port 514 nsew
rlabel metal2 s 11472 22357 11472 22357 4 gnd
port 514 nsew
rlabel metal2 s 11472 23463 11472 23463 4 gnd
port 514 nsew
rlabel metal2 s 12240 22357 12240 22357 4 gnd
port 514 nsew
rlabel metal2 s 10992 25280 10992 25280 4 gnd
port 514 nsew
rlabel metal2 s 11472 23937 11472 23937 4 gnd
port 514 nsew
rlabel metal2 s 10992 24490 10992 24490 4 gnd
port 514 nsew
rlabel metal2 s 11472 25043 11472 25043 4 gnd
port 514 nsew
rlabel metal2 s 10224 24727 10224 24727 4 gnd
port 514 nsew
rlabel metal2 s 12240 24727 12240 24727 4 gnd
port 514 nsew
rlabel metal2 s 12240 23147 12240 23147 4 gnd
port 514 nsew
rlabel metal2 s 10992 22357 10992 22357 4 gnd
port 514 nsew
rlabel metal2 s 11472 24727 11472 24727 4 gnd
port 514 nsew
rlabel metal2 s 10992 24727 10992 24727 4 gnd
port 514 nsew
rlabel metal2 s 11472 23700 11472 23700 4 gnd
port 514 nsew
rlabel metal2 s 10224 25280 10224 25280 4 gnd
port 514 nsew
rlabel metal2 s 10224 25043 10224 25043 4 gnd
port 514 nsew
rlabel metal2 s 10224 22910 10224 22910 4 gnd
port 514 nsew
rlabel metal2 s 12240 23937 12240 23937 4 gnd
port 514 nsew
rlabel metal2 s 11472 24253 11472 24253 4 gnd
port 514 nsew
rlabel metal2 s 10224 23700 10224 23700 4 gnd
port 514 nsew
rlabel metal2 s 11472 23147 11472 23147 4 gnd
port 514 nsew
rlabel metal2 s 10992 23463 10992 23463 4 gnd
port 514 nsew
rlabel metal2 s 10992 23700 10992 23700 4 gnd
port 514 nsew
rlabel metal2 s 10992 22673 10992 22673 4 gnd
port 514 nsew
rlabel metal2 s 12240 25043 12240 25043 4 gnd
port 514 nsew
rlabel metal2 s 12240 24490 12240 24490 4 gnd
port 514 nsew
rlabel metal2 s 12240 22673 12240 22673 4 gnd
port 514 nsew
rlabel metal2 s 12240 25280 12240 25280 4 gnd
port 514 nsew
rlabel metal2 s 10992 23937 10992 23937 4 gnd
port 514 nsew
rlabel metal2 s 10224 21093 10224 21093 4 gnd
port 514 nsew
rlabel metal2 s 10992 19513 10992 19513 4 gnd
port 514 nsew
rlabel metal2 s 10992 19750 10992 19750 4 gnd
port 514 nsew
rlabel metal2 s 10992 20777 10992 20777 4 gnd
port 514 nsew
rlabel metal2 s 10224 19750 10224 19750 4 gnd
port 514 nsew
rlabel metal2 s 11472 20303 11472 20303 4 gnd
port 514 nsew
rlabel metal2 s 12240 20777 12240 20777 4 gnd
port 514 nsew
rlabel metal2 s 11472 21330 11472 21330 4 gnd
port 514 nsew
rlabel metal2 s 10992 21567 10992 21567 4 gnd
port 514 nsew
rlabel metal2 s 10224 19513 10224 19513 4 gnd
port 514 nsew
rlabel metal2 s 10224 21883 10224 21883 4 gnd
port 514 nsew
rlabel metal2 s 10992 20303 10992 20303 4 gnd
port 514 nsew
rlabel metal2 s 12240 19513 12240 19513 4 gnd
port 514 nsew
rlabel metal2 s 11472 22120 11472 22120 4 gnd
port 514 nsew
rlabel metal2 s 10224 20303 10224 20303 4 gnd
port 514 nsew
rlabel metal2 s 12240 19197 12240 19197 4 gnd
port 514 nsew
rlabel metal2 s 10992 20540 10992 20540 4 gnd
port 514 nsew
rlabel metal2 s 10992 19197 10992 19197 4 gnd
port 514 nsew
rlabel metal2 s 12240 21093 12240 21093 4 gnd
port 514 nsew
rlabel metal2 s 11472 21093 11472 21093 4 gnd
port 514 nsew
rlabel metal2 s 10224 19987 10224 19987 4 gnd
port 514 nsew
rlabel metal2 s 12240 21883 12240 21883 4 gnd
port 514 nsew
rlabel metal2 s 11472 20540 11472 20540 4 gnd
port 514 nsew
rlabel metal2 s 11472 19513 11472 19513 4 gnd
port 514 nsew
rlabel metal2 s 11472 21883 11472 21883 4 gnd
port 514 nsew
rlabel metal2 s 10224 21567 10224 21567 4 gnd
port 514 nsew
rlabel metal2 s 10224 19197 10224 19197 4 gnd
port 514 nsew
rlabel metal2 s 10224 21330 10224 21330 4 gnd
port 514 nsew
rlabel metal2 s 10224 22120 10224 22120 4 gnd
port 514 nsew
rlabel metal2 s 12240 22120 12240 22120 4 gnd
port 514 nsew
rlabel metal2 s 10992 22120 10992 22120 4 gnd
port 514 nsew
rlabel metal2 s 11472 21567 11472 21567 4 gnd
port 514 nsew
rlabel metal2 s 12240 19987 12240 19987 4 gnd
port 514 nsew
rlabel metal2 s 11472 19987 11472 19987 4 gnd
port 514 nsew
rlabel metal2 s 12240 20303 12240 20303 4 gnd
port 514 nsew
rlabel metal2 s 11472 19750 11472 19750 4 gnd
port 514 nsew
rlabel metal2 s 11472 19197 11472 19197 4 gnd
port 514 nsew
rlabel metal2 s 12240 21567 12240 21567 4 gnd
port 514 nsew
rlabel metal2 s 10224 20540 10224 20540 4 gnd
port 514 nsew
rlabel metal2 s 12240 20540 12240 20540 4 gnd
port 514 nsew
rlabel metal2 s 10992 21093 10992 21093 4 gnd
port 514 nsew
rlabel metal2 s 11472 20777 11472 20777 4 gnd
port 514 nsew
rlabel metal2 s 12240 19750 12240 19750 4 gnd
port 514 nsew
rlabel metal2 s 10992 21883 10992 21883 4 gnd
port 514 nsew
rlabel metal2 s 12240 21330 12240 21330 4 gnd
port 514 nsew
rlabel metal2 s 10992 19987 10992 19987 4 gnd
port 514 nsew
rlabel metal2 s 10224 20777 10224 20777 4 gnd
port 514 nsew
rlabel metal2 s 10992 21330 10992 21330 4 gnd
port 514 nsew
rlabel metal2 s 14736 21567 14736 21567 4 gnd
port 514 nsew
rlabel metal2 s 14736 19987 14736 19987 4 gnd
port 514 nsew
rlabel metal2 s 13488 20540 13488 20540 4 gnd
port 514 nsew
rlabel metal2 s 14736 19513 14736 19513 4 gnd
port 514 nsew
rlabel metal2 s 12720 20777 12720 20777 4 gnd
port 514 nsew
rlabel metal2 s 13488 19987 13488 19987 4 gnd
port 514 nsew
rlabel metal2 s 12720 22120 12720 22120 4 gnd
port 514 nsew
rlabel metal2 s 12720 21330 12720 21330 4 gnd
port 514 nsew
rlabel metal2 s 12720 19750 12720 19750 4 gnd
port 514 nsew
rlabel metal2 s 14736 22120 14736 22120 4 gnd
port 514 nsew
rlabel metal2 s 13488 19750 13488 19750 4 gnd
port 514 nsew
rlabel metal2 s 13488 21330 13488 21330 4 gnd
port 514 nsew
rlabel metal2 s 12720 21567 12720 21567 4 gnd
port 514 nsew
rlabel metal2 s 13968 20777 13968 20777 4 gnd
port 514 nsew
rlabel metal2 s 14736 20777 14736 20777 4 gnd
port 514 nsew
rlabel metal2 s 14736 21883 14736 21883 4 gnd
port 514 nsew
rlabel metal2 s 12720 19197 12720 19197 4 gnd
port 514 nsew
rlabel metal2 s 13488 20303 13488 20303 4 gnd
port 514 nsew
rlabel metal2 s 12720 20540 12720 20540 4 gnd
port 514 nsew
rlabel metal2 s 13968 21330 13968 21330 4 gnd
port 514 nsew
rlabel metal2 s 13968 21567 13968 21567 4 gnd
port 514 nsew
rlabel metal2 s 13968 19513 13968 19513 4 gnd
port 514 nsew
rlabel metal2 s 14736 21330 14736 21330 4 gnd
port 514 nsew
rlabel metal2 s 12720 19513 12720 19513 4 gnd
port 514 nsew
rlabel metal2 s 12720 20303 12720 20303 4 gnd
port 514 nsew
rlabel metal2 s 12720 21093 12720 21093 4 gnd
port 514 nsew
rlabel metal2 s 13488 20777 13488 20777 4 gnd
port 514 nsew
rlabel metal2 s 14736 20540 14736 20540 4 gnd
port 514 nsew
rlabel metal2 s 13968 21093 13968 21093 4 gnd
port 514 nsew
rlabel metal2 s 13968 22120 13968 22120 4 gnd
port 514 nsew
rlabel metal2 s 13968 19197 13968 19197 4 gnd
port 514 nsew
rlabel metal2 s 12720 19987 12720 19987 4 gnd
port 514 nsew
rlabel metal2 s 13968 20540 13968 20540 4 gnd
port 514 nsew
rlabel metal2 s 13488 21567 13488 21567 4 gnd
port 514 nsew
rlabel metal2 s 13968 19987 13968 19987 4 gnd
port 514 nsew
rlabel metal2 s 13488 19513 13488 19513 4 gnd
port 514 nsew
rlabel metal2 s 13488 19197 13488 19197 4 gnd
port 514 nsew
rlabel metal2 s 13968 20303 13968 20303 4 gnd
port 514 nsew
rlabel metal2 s 12720 21883 12720 21883 4 gnd
port 514 nsew
rlabel metal2 s 13968 21883 13968 21883 4 gnd
port 514 nsew
rlabel metal2 s 14736 20303 14736 20303 4 gnd
port 514 nsew
rlabel metal2 s 13488 21883 13488 21883 4 gnd
port 514 nsew
rlabel metal2 s 14736 19750 14736 19750 4 gnd
port 514 nsew
rlabel metal2 s 14736 21093 14736 21093 4 gnd
port 514 nsew
rlabel metal2 s 13488 22120 13488 22120 4 gnd
port 514 nsew
rlabel metal2 s 13968 19750 13968 19750 4 gnd
port 514 nsew
rlabel metal2 s 14736 19197 14736 19197 4 gnd
port 514 nsew
rlabel metal2 s 13488 21093 13488 21093 4 gnd
port 514 nsew
rlabel metal2 s 12720 17933 12720 17933 4 gnd
port 514 nsew
rlabel metal2 s 12720 18960 12720 18960 4 gnd
port 514 nsew
rlabel metal2 s 13488 18723 13488 18723 4 gnd
port 514 nsew
rlabel metal2 s 13968 17143 13968 17143 4 gnd
port 514 nsew
rlabel metal2 s 14736 16827 14736 16827 4 gnd
port 514 nsew
rlabel metal2 s 13968 18723 13968 18723 4 gnd
port 514 nsew
rlabel metal2 s 12720 16590 12720 16590 4 gnd
port 514 nsew
rlabel metal2 s 14736 16590 14736 16590 4 gnd
port 514 nsew
rlabel metal2 s 13968 18960 13968 18960 4 gnd
port 514 nsew
rlabel metal2 s 13968 16590 13968 16590 4 gnd
port 514 nsew
rlabel metal2 s 14736 17143 14736 17143 4 gnd
port 514 nsew
rlabel metal2 s 14736 16353 14736 16353 4 gnd
port 514 nsew
rlabel metal2 s 12720 18407 12720 18407 4 gnd
port 514 nsew
rlabel metal2 s 13968 16827 13968 16827 4 gnd
port 514 nsew
rlabel metal2 s 12720 18723 12720 18723 4 gnd
port 514 nsew
rlabel metal2 s 14736 16037 14736 16037 4 gnd
port 514 nsew
rlabel metal2 s 13968 18170 13968 18170 4 gnd
port 514 nsew
rlabel metal2 s 13968 16037 13968 16037 4 gnd
port 514 nsew
rlabel metal2 s 13488 18170 13488 18170 4 gnd
port 514 nsew
rlabel metal2 s 13488 17143 13488 17143 4 gnd
port 514 nsew
rlabel metal2 s 13968 18407 13968 18407 4 gnd
port 514 nsew
rlabel metal2 s 12720 17143 12720 17143 4 gnd
port 514 nsew
rlabel metal2 s 12720 17380 12720 17380 4 gnd
port 514 nsew
rlabel metal2 s 14736 18170 14736 18170 4 gnd
port 514 nsew
rlabel metal2 s 12720 16037 12720 16037 4 gnd
port 514 nsew
rlabel metal2 s 14736 17380 14736 17380 4 gnd
port 514 nsew
rlabel metal2 s 14736 18723 14736 18723 4 gnd
port 514 nsew
rlabel metal2 s 13488 16353 13488 16353 4 gnd
port 514 nsew
rlabel metal2 s 13488 17933 13488 17933 4 gnd
port 514 nsew
rlabel metal2 s 12720 18170 12720 18170 4 gnd
port 514 nsew
rlabel metal2 s 14736 17617 14736 17617 4 gnd
port 514 nsew
rlabel metal2 s 14736 17933 14736 17933 4 gnd
port 514 nsew
rlabel metal2 s 13488 16590 13488 16590 4 gnd
port 514 nsew
rlabel metal2 s 12720 17617 12720 17617 4 gnd
port 514 nsew
rlabel metal2 s 12720 16827 12720 16827 4 gnd
port 514 nsew
rlabel metal2 s 13488 17380 13488 17380 4 gnd
port 514 nsew
rlabel metal2 s 14736 18960 14736 18960 4 gnd
port 514 nsew
rlabel metal2 s 12720 16353 12720 16353 4 gnd
port 514 nsew
rlabel metal2 s 13488 18960 13488 18960 4 gnd
port 514 nsew
rlabel metal2 s 13488 18407 13488 18407 4 gnd
port 514 nsew
rlabel metal2 s 13968 17617 13968 17617 4 gnd
port 514 nsew
rlabel metal2 s 13488 16037 13488 16037 4 gnd
port 514 nsew
rlabel metal2 s 13968 16353 13968 16353 4 gnd
port 514 nsew
rlabel metal2 s 13488 16827 13488 16827 4 gnd
port 514 nsew
rlabel metal2 s 14736 18407 14736 18407 4 gnd
port 514 nsew
rlabel metal2 s 13968 17933 13968 17933 4 gnd
port 514 nsew
rlabel metal2 s 13968 17380 13968 17380 4 gnd
port 514 nsew
rlabel metal2 s 13488 17617 13488 17617 4 gnd
port 514 nsew
rlabel metal2 s 12240 18960 12240 18960 4 gnd
port 514 nsew
rlabel metal2 s 12240 17933 12240 17933 4 gnd
port 514 nsew
rlabel metal2 s 11472 17933 11472 17933 4 gnd
port 514 nsew
rlabel metal2 s 12240 18723 12240 18723 4 gnd
port 514 nsew
rlabel metal2 s 12240 16827 12240 16827 4 gnd
port 514 nsew
rlabel metal2 s 10224 17933 10224 17933 4 gnd
port 514 nsew
rlabel metal2 s 10992 16353 10992 16353 4 gnd
port 514 nsew
rlabel metal2 s 10992 17380 10992 17380 4 gnd
port 514 nsew
rlabel metal2 s 10224 18170 10224 18170 4 gnd
port 514 nsew
rlabel metal2 s 11472 17617 11472 17617 4 gnd
port 514 nsew
rlabel metal2 s 10224 17617 10224 17617 4 gnd
port 514 nsew
rlabel metal2 s 10992 16590 10992 16590 4 gnd
port 514 nsew
rlabel metal2 s 11472 16590 11472 16590 4 gnd
port 514 nsew
rlabel metal2 s 10992 16827 10992 16827 4 gnd
port 514 nsew
rlabel metal2 s 10224 18960 10224 18960 4 gnd
port 514 nsew
rlabel metal2 s 10992 18170 10992 18170 4 gnd
port 514 nsew
rlabel metal2 s 11472 17143 11472 17143 4 gnd
port 514 nsew
rlabel metal2 s 10224 18723 10224 18723 4 gnd
port 514 nsew
rlabel metal2 s 10992 17617 10992 17617 4 gnd
port 514 nsew
rlabel metal2 s 12240 17143 12240 17143 4 gnd
port 514 nsew
rlabel metal2 s 10224 16037 10224 16037 4 gnd
port 514 nsew
rlabel metal2 s 11472 18723 11472 18723 4 gnd
port 514 nsew
rlabel metal2 s 12240 16590 12240 16590 4 gnd
port 514 nsew
rlabel metal2 s 10224 16353 10224 16353 4 gnd
port 514 nsew
rlabel metal2 s 10224 18407 10224 18407 4 gnd
port 514 nsew
rlabel metal2 s 10992 18723 10992 18723 4 gnd
port 514 nsew
rlabel metal2 s 12240 17380 12240 17380 4 gnd
port 514 nsew
rlabel metal2 s 12240 17617 12240 17617 4 gnd
port 514 nsew
rlabel metal2 s 10992 17143 10992 17143 4 gnd
port 514 nsew
rlabel metal2 s 12240 16037 12240 16037 4 gnd
port 514 nsew
rlabel metal2 s 10224 17143 10224 17143 4 gnd
port 514 nsew
rlabel metal2 s 11472 16827 11472 16827 4 gnd
port 514 nsew
rlabel metal2 s 12240 18170 12240 18170 4 gnd
port 514 nsew
rlabel metal2 s 11472 17380 11472 17380 4 gnd
port 514 nsew
rlabel metal2 s 11472 16037 11472 16037 4 gnd
port 514 nsew
rlabel metal2 s 11472 18407 11472 18407 4 gnd
port 514 nsew
rlabel metal2 s 11472 18960 11472 18960 4 gnd
port 514 nsew
rlabel metal2 s 10992 18960 10992 18960 4 gnd
port 514 nsew
rlabel metal2 s 11472 16353 11472 16353 4 gnd
port 514 nsew
rlabel metal2 s 10992 17933 10992 17933 4 gnd
port 514 nsew
rlabel metal2 s 10224 16590 10224 16590 4 gnd
port 514 nsew
rlabel metal2 s 12240 18407 12240 18407 4 gnd
port 514 nsew
rlabel metal2 s 11472 18170 11472 18170 4 gnd
port 514 nsew
rlabel metal2 s 12240 16353 12240 16353 4 gnd
port 514 nsew
rlabel metal2 s 10224 16827 10224 16827 4 gnd
port 514 nsew
rlabel metal2 s 10992 18407 10992 18407 4 gnd
port 514 nsew
rlabel metal2 s 10224 17380 10224 17380 4 gnd
port 514 nsew
rlabel metal2 s 10992 16037 10992 16037 4 gnd
port 514 nsew
rlabel metal2 s 12240 15010 12240 15010 4 gnd
port 514 nsew
rlabel metal2 s 11472 13193 11472 13193 4 gnd
port 514 nsew
rlabel metal2 s 12240 15247 12240 15247 4 gnd
port 514 nsew
rlabel metal2 s 10224 14773 10224 14773 4 gnd
port 514 nsew
rlabel metal2 s 12240 14457 12240 14457 4 gnd
port 514 nsew
rlabel metal2 s 10992 13430 10992 13430 4 gnd
port 514 nsew
rlabel metal2 s 10224 13193 10224 13193 4 gnd
port 514 nsew
rlabel metal2 s 12240 15800 12240 15800 4 gnd
port 514 nsew
rlabel metal2 s 12240 13430 12240 13430 4 gnd
port 514 nsew
rlabel metal2 s 11472 12877 11472 12877 4 gnd
port 514 nsew
rlabel metal2 s 10992 14457 10992 14457 4 gnd
port 514 nsew
rlabel metal2 s 10224 15247 10224 15247 4 gnd
port 514 nsew
rlabel metal2 s 11472 13667 11472 13667 4 gnd
port 514 nsew
rlabel metal2 s 11472 14220 11472 14220 4 gnd
port 514 nsew
rlabel metal2 s 10992 14220 10992 14220 4 gnd
port 514 nsew
rlabel metal2 s 10224 15010 10224 15010 4 gnd
port 514 nsew
rlabel metal2 s 10992 14773 10992 14773 4 gnd
port 514 nsew
rlabel metal2 s 12240 14773 12240 14773 4 gnd
port 514 nsew
rlabel metal2 s 11472 15800 11472 15800 4 gnd
port 514 nsew
rlabel metal2 s 10224 13430 10224 13430 4 gnd
port 514 nsew
rlabel metal2 s 10224 12877 10224 12877 4 gnd
port 514 nsew
rlabel metal2 s 12240 15563 12240 15563 4 gnd
port 514 nsew
rlabel metal2 s 12240 13667 12240 13667 4 gnd
port 514 nsew
rlabel metal2 s 10224 15800 10224 15800 4 gnd
port 514 nsew
rlabel metal2 s 11472 15563 11472 15563 4 gnd
port 514 nsew
rlabel metal2 s 11472 15247 11472 15247 4 gnd
port 514 nsew
rlabel metal2 s 10992 15247 10992 15247 4 gnd
port 514 nsew
rlabel metal2 s 10992 15563 10992 15563 4 gnd
port 514 nsew
rlabel metal2 s 10224 14220 10224 14220 4 gnd
port 514 nsew
rlabel metal2 s 11472 14773 11472 14773 4 gnd
port 514 nsew
rlabel metal2 s 10992 12877 10992 12877 4 gnd
port 514 nsew
rlabel metal2 s 11472 13983 11472 13983 4 gnd
port 514 nsew
rlabel metal2 s 12240 14220 12240 14220 4 gnd
port 514 nsew
rlabel metal2 s 10992 15800 10992 15800 4 gnd
port 514 nsew
rlabel metal2 s 10992 15010 10992 15010 4 gnd
port 514 nsew
rlabel metal2 s 11472 14457 11472 14457 4 gnd
port 514 nsew
rlabel metal2 s 10992 13193 10992 13193 4 gnd
port 514 nsew
rlabel metal2 s 11472 15010 11472 15010 4 gnd
port 514 nsew
rlabel metal2 s 12240 13193 12240 13193 4 gnd
port 514 nsew
rlabel metal2 s 10224 13667 10224 13667 4 gnd
port 514 nsew
rlabel metal2 s 10992 13667 10992 13667 4 gnd
port 514 nsew
rlabel metal2 s 10224 15563 10224 15563 4 gnd
port 514 nsew
rlabel metal2 s 12240 13983 12240 13983 4 gnd
port 514 nsew
rlabel metal2 s 10224 13983 10224 13983 4 gnd
port 514 nsew
rlabel metal2 s 11472 13430 11472 13430 4 gnd
port 514 nsew
rlabel metal2 s 10224 14457 10224 14457 4 gnd
port 514 nsew
rlabel metal2 s 12240 12877 12240 12877 4 gnd
port 514 nsew
rlabel metal2 s 10992 13983 10992 13983 4 gnd
port 514 nsew
rlabel metal2 s 14736 13193 14736 13193 4 gnd
port 514 nsew
rlabel metal2 s 13488 13667 13488 13667 4 gnd
port 514 nsew
rlabel metal2 s 12720 12877 12720 12877 4 gnd
port 514 nsew
rlabel metal2 s 13968 12877 13968 12877 4 gnd
port 514 nsew
rlabel metal2 s 13968 15563 13968 15563 4 gnd
port 514 nsew
rlabel metal2 s 14736 15010 14736 15010 4 gnd
port 514 nsew
rlabel metal2 s 14736 15247 14736 15247 4 gnd
port 514 nsew
rlabel metal2 s 12720 14457 12720 14457 4 gnd
port 514 nsew
rlabel metal2 s 13488 13983 13488 13983 4 gnd
port 514 nsew
rlabel metal2 s 13968 13430 13968 13430 4 gnd
port 514 nsew
rlabel metal2 s 12720 14220 12720 14220 4 gnd
port 514 nsew
rlabel metal2 s 12720 15247 12720 15247 4 gnd
port 514 nsew
rlabel metal2 s 14736 14773 14736 14773 4 gnd
port 514 nsew
rlabel metal2 s 14736 14457 14736 14457 4 gnd
port 514 nsew
rlabel metal2 s 14736 12877 14736 12877 4 gnd
port 514 nsew
rlabel metal2 s 14736 13983 14736 13983 4 gnd
port 514 nsew
rlabel metal2 s 13968 15010 13968 15010 4 gnd
port 514 nsew
rlabel metal2 s 12720 15563 12720 15563 4 gnd
port 514 nsew
rlabel metal2 s 13968 14457 13968 14457 4 gnd
port 514 nsew
rlabel metal2 s 12720 13430 12720 13430 4 gnd
port 514 nsew
rlabel metal2 s 13488 15010 13488 15010 4 gnd
port 514 nsew
rlabel metal2 s 12720 14773 12720 14773 4 gnd
port 514 nsew
rlabel metal2 s 13488 15563 13488 15563 4 gnd
port 514 nsew
rlabel metal2 s 13488 13430 13488 13430 4 gnd
port 514 nsew
rlabel metal2 s 13968 15247 13968 15247 4 gnd
port 514 nsew
rlabel metal2 s 13488 14220 13488 14220 4 gnd
port 514 nsew
rlabel metal2 s 12720 15800 12720 15800 4 gnd
port 514 nsew
rlabel metal2 s 13488 14773 13488 14773 4 gnd
port 514 nsew
rlabel metal2 s 13488 12877 13488 12877 4 gnd
port 514 nsew
rlabel metal2 s 13488 15800 13488 15800 4 gnd
port 514 nsew
rlabel metal2 s 14736 15800 14736 15800 4 gnd
port 514 nsew
rlabel metal2 s 12720 13983 12720 13983 4 gnd
port 514 nsew
rlabel metal2 s 12720 13667 12720 13667 4 gnd
port 514 nsew
rlabel metal2 s 13968 13667 13968 13667 4 gnd
port 514 nsew
rlabel metal2 s 13968 14220 13968 14220 4 gnd
port 514 nsew
rlabel metal2 s 13968 13193 13968 13193 4 gnd
port 514 nsew
rlabel metal2 s 13488 15247 13488 15247 4 gnd
port 514 nsew
rlabel metal2 s 14736 13667 14736 13667 4 gnd
port 514 nsew
rlabel metal2 s 13968 14773 13968 14773 4 gnd
port 514 nsew
rlabel metal2 s 13488 14457 13488 14457 4 gnd
port 514 nsew
rlabel metal2 s 14736 14220 14736 14220 4 gnd
port 514 nsew
rlabel metal2 s 14736 15563 14736 15563 4 gnd
port 514 nsew
rlabel metal2 s 13968 13983 13968 13983 4 gnd
port 514 nsew
rlabel metal2 s 12720 13193 12720 13193 4 gnd
port 514 nsew
rlabel metal2 s 14736 13430 14736 13430 4 gnd
port 514 nsew
rlabel metal2 s 13488 13193 13488 13193 4 gnd
port 514 nsew
rlabel metal2 s 13968 15800 13968 15800 4 gnd
port 514 nsew
rlabel metal2 s 12720 15010 12720 15010 4 gnd
port 514 nsew
rlabel metal2 s 17712 16590 17712 16590 4 gnd
port 514 nsew
rlabel metal2 s 19728 16037 19728 16037 4 gnd
port 514 nsew
rlabel metal2 s 19728 18407 19728 18407 4 gnd
port 514 nsew
rlabel metal2 s 17712 17617 17712 17617 4 gnd
port 514 nsew
rlabel metal2 s 18960 17933 18960 17933 4 gnd
port 514 nsew
rlabel metal2 s 18960 16590 18960 16590 4 gnd
port 514 nsew
rlabel metal2 s 19728 18960 19728 18960 4 gnd
port 514 nsew
rlabel metal2 s 18480 18723 18480 18723 4 gnd
port 514 nsew
rlabel metal2 s 18960 18407 18960 18407 4 gnd
port 514 nsew
rlabel metal2 s 19728 17617 19728 17617 4 gnd
port 514 nsew
rlabel metal2 s 19728 16590 19728 16590 4 gnd
port 514 nsew
rlabel metal2 s 17712 18170 17712 18170 4 gnd
port 514 nsew
rlabel metal2 s 19728 18723 19728 18723 4 gnd
port 514 nsew
rlabel metal2 s 18960 17617 18960 17617 4 gnd
port 514 nsew
rlabel metal2 s 17712 17380 17712 17380 4 gnd
port 514 nsew
rlabel metal2 s 18480 16590 18480 16590 4 gnd
port 514 nsew
rlabel metal2 s 17712 18723 17712 18723 4 gnd
port 514 nsew
rlabel metal2 s 19728 17143 19728 17143 4 gnd
port 514 nsew
rlabel metal2 s 17712 16353 17712 16353 4 gnd
port 514 nsew
rlabel metal2 s 19728 16353 19728 16353 4 gnd
port 514 nsew
rlabel metal2 s 17712 17933 17712 17933 4 gnd
port 514 nsew
rlabel metal2 s 18480 18170 18480 18170 4 gnd
port 514 nsew
rlabel metal2 s 18480 18960 18480 18960 4 gnd
port 514 nsew
rlabel metal2 s 18960 16827 18960 16827 4 gnd
port 514 nsew
rlabel metal2 s 18480 17933 18480 17933 4 gnd
port 514 nsew
rlabel metal2 s 17712 16037 17712 16037 4 gnd
port 514 nsew
rlabel metal2 s 17712 16827 17712 16827 4 gnd
port 514 nsew
rlabel metal2 s 19728 17380 19728 17380 4 gnd
port 514 nsew
rlabel metal2 s 17712 17143 17712 17143 4 gnd
port 514 nsew
rlabel metal2 s 18480 17380 18480 17380 4 gnd
port 514 nsew
rlabel metal2 s 18480 16827 18480 16827 4 gnd
port 514 nsew
rlabel metal2 s 18480 17617 18480 17617 4 gnd
port 514 nsew
rlabel metal2 s 17712 18407 17712 18407 4 gnd
port 514 nsew
rlabel metal2 s 18480 17143 18480 17143 4 gnd
port 514 nsew
rlabel metal2 s 18960 18170 18960 18170 4 gnd
port 514 nsew
rlabel metal2 s 18960 18723 18960 18723 4 gnd
port 514 nsew
rlabel metal2 s 18480 16353 18480 16353 4 gnd
port 514 nsew
rlabel metal2 s 18480 16037 18480 16037 4 gnd
port 514 nsew
rlabel metal2 s 19728 17933 19728 17933 4 gnd
port 514 nsew
rlabel metal2 s 19728 18170 19728 18170 4 gnd
port 514 nsew
rlabel metal2 s 19968 15927 19968 15927 4 wl1_40
port 338 nsew
rlabel metal2 s 19968 17253 19968 17253 4 wl1_43
port 344 nsew
rlabel metal2 s 19968 18613 19968 18613 4 wl0_47
port 351 nsew
rlabel metal2 s 19728 16827 19728 16827 4 gnd
port 514 nsew
rlabel metal2 s 18960 17143 18960 17143 4 gnd
port 514 nsew
rlabel metal2 s 19968 17823 19968 17823 4 wl0_45
port 347 nsew
rlabel metal2 s 18480 18407 18480 18407 4 gnd
port 514 nsew
rlabel metal2 s 19968 18297 19968 18297 4 wl1_46
port 350 nsew
rlabel metal2 s 19968 16937 19968 16937 4 wl0_42
port 341 nsew
rlabel metal2 s 18960 17380 18960 17380 4 gnd
port 514 nsew
rlabel metal2 s 19968 18043 19968 18043 4 wl1_45
port 348 nsew
rlabel metal2 s 18960 16353 18960 16353 4 gnd
port 514 nsew
rlabel metal2 s 18960 16037 18960 16037 4 gnd
port 514 nsew
rlabel metal2 s 19968 16463 19968 16463 4 wl1_41
port 340 nsew
rlabel metal2 s 19968 18517 19968 18517 4 wl0_46
port 349 nsew
rlabel metal2 s 19968 17727 19968 17727 4 wl0_44
port 345 nsew
rlabel metal2 s 19968 16717 19968 16717 4 wl1_42
port 342 nsew
rlabel metal2 s 19968 17033 19968 17033 4 wl0_43
port 343 nsew
rlabel metal2 s 19968 18833 19968 18833 4 wl1_47
port 352 nsew
rlabel metal2 s 18960 18960 18960 18960 4 gnd
port 514 nsew
rlabel metal2 s 17712 18960 17712 18960 4 gnd
port 514 nsew
rlabel metal2 s 19968 16147 19968 16147 4 wl0_40
port 337 nsew
rlabel metal2 s 19968 16243 19968 16243 4 wl0_41
port 339 nsew
rlabel metal2 s 19968 17507 19968 17507 4 wl1_44
port 346 nsew
rlabel metal2 s 15984 16590 15984 16590 4 gnd
port 514 nsew
rlabel metal2 s 15216 16590 15216 16590 4 gnd
port 514 nsew
rlabel metal2 s 15216 17617 15216 17617 4 gnd
port 514 nsew
rlabel metal2 s 17232 17617 17232 17617 4 gnd
port 514 nsew
rlabel metal2 s 16464 17617 16464 17617 4 gnd
port 514 nsew
rlabel metal2 s 15984 17143 15984 17143 4 gnd
port 514 nsew
rlabel metal2 s 15216 16827 15216 16827 4 gnd
port 514 nsew
rlabel metal2 s 17232 17933 17232 17933 4 gnd
port 514 nsew
rlabel metal2 s 15216 17933 15216 17933 4 gnd
port 514 nsew
rlabel metal2 s 16464 16037 16464 16037 4 gnd
port 514 nsew
rlabel metal2 s 16464 18407 16464 18407 4 gnd
port 514 nsew
rlabel metal2 s 17232 18170 17232 18170 4 gnd
port 514 nsew
rlabel metal2 s 15216 17380 15216 17380 4 gnd
port 514 nsew
rlabel metal2 s 17232 18960 17232 18960 4 gnd
port 514 nsew
rlabel metal2 s 17232 17380 17232 17380 4 gnd
port 514 nsew
rlabel metal2 s 15216 18407 15216 18407 4 gnd
port 514 nsew
rlabel metal2 s 16464 18960 16464 18960 4 gnd
port 514 nsew
rlabel metal2 s 15984 17380 15984 17380 4 gnd
port 514 nsew
rlabel metal2 s 17232 18407 17232 18407 4 gnd
port 514 nsew
rlabel metal2 s 16464 17933 16464 17933 4 gnd
port 514 nsew
rlabel metal2 s 16464 16590 16464 16590 4 gnd
port 514 nsew
rlabel metal2 s 16464 16353 16464 16353 4 gnd
port 514 nsew
rlabel metal2 s 17232 17143 17232 17143 4 gnd
port 514 nsew
rlabel metal2 s 15984 18723 15984 18723 4 gnd
port 514 nsew
rlabel metal2 s 15984 16353 15984 16353 4 gnd
port 514 nsew
rlabel metal2 s 15984 16037 15984 16037 4 gnd
port 514 nsew
rlabel metal2 s 15984 18170 15984 18170 4 gnd
port 514 nsew
rlabel metal2 s 17232 16037 17232 16037 4 gnd
port 514 nsew
rlabel metal2 s 17232 16827 17232 16827 4 gnd
port 514 nsew
rlabel metal2 s 17232 16353 17232 16353 4 gnd
port 514 nsew
rlabel metal2 s 15984 17933 15984 17933 4 gnd
port 514 nsew
rlabel metal2 s 16464 18170 16464 18170 4 gnd
port 514 nsew
rlabel metal2 s 15984 16827 15984 16827 4 gnd
port 514 nsew
rlabel metal2 s 15216 16037 15216 16037 4 gnd
port 514 nsew
rlabel metal2 s 15216 16353 15216 16353 4 gnd
port 514 nsew
rlabel metal2 s 15984 18407 15984 18407 4 gnd
port 514 nsew
rlabel metal2 s 15216 18723 15216 18723 4 gnd
port 514 nsew
rlabel metal2 s 16464 18723 16464 18723 4 gnd
port 514 nsew
rlabel metal2 s 15216 18170 15216 18170 4 gnd
port 514 nsew
rlabel metal2 s 15216 18960 15216 18960 4 gnd
port 514 nsew
rlabel metal2 s 17232 18723 17232 18723 4 gnd
port 514 nsew
rlabel metal2 s 16464 17380 16464 17380 4 gnd
port 514 nsew
rlabel metal2 s 15984 17617 15984 17617 4 gnd
port 514 nsew
rlabel metal2 s 16464 17143 16464 17143 4 gnd
port 514 nsew
rlabel metal2 s 16464 16827 16464 16827 4 gnd
port 514 nsew
rlabel metal2 s 15984 18960 15984 18960 4 gnd
port 514 nsew
rlabel metal2 s 15216 17143 15216 17143 4 gnd
port 514 nsew
rlabel metal2 s 17232 16590 17232 16590 4 gnd
port 514 nsew
rlabel metal2 s 16464 13983 16464 13983 4 gnd
port 514 nsew
rlabel metal2 s 15984 13667 15984 13667 4 gnd
port 514 nsew
rlabel metal2 s 15216 14457 15216 14457 4 gnd
port 514 nsew
rlabel metal2 s 17232 13667 17232 13667 4 gnd
port 514 nsew
rlabel metal2 s 15216 15010 15216 15010 4 gnd
port 514 nsew
rlabel metal2 s 15984 15563 15984 15563 4 gnd
port 514 nsew
rlabel metal2 s 16464 15563 16464 15563 4 gnd
port 514 nsew
rlabel metal2 s 16464 14457 16464 14457 4 gnd
port 514 nsew
rlabel metal2 s 15216 15563 15216 15563 4 gnd
port 514 nsew
rlabel metal2 s 17232 14457 17232 14457 4 gnd
port 514 nsew
rlabel metal2 s 16464 14220 16464 14220 4 gnd
port 514 nsew
rlabel metal2 s 16464 15800 16464 15800 4 gnd
port 514 nsew
rlabel metal2 s 16464 13667 16464 13667 4 gnd
port 514 nsew
rlabel metal2 s 16464 13430 16464 13430 4 gnd
port 514 nsew
rlabel metal2 s 17232 13983 17232 13983 4 gnd
port 514 nsew
rlabel metal2 s 15216 13667 15216 13667 4 gnd
port 514 nsew
rlabel metal2 s 17232 14773 17232 14773 4 gnd
port 514 nsew
rlabel metal2 s 16464 14773 16464 14773 4 gnd
port 514 nsew
rlabel metal2 s 16464 15010 16464 15010 4 gnd
port 514 nsew
rlabel metal2 s 17232 15010 17232 15010 4 gnd
port 514 nsew
rlabel metal2 s 16464 13193 16464 13193 4 gnd
port 514 nsew
rlabel metal2 s 15984 13430 15984 13430 4 gnd
port 514 nsew
rlabel metal2 s 15216 12877 15216 12877 4 gnd
port 514 nsew
rlabel metal2 s 15216 15247 15216 15247 4 gnd
port 514 nsew
rlabel metal2 s 16464 15247 16464 15247 4 gnd
port 514 nsew
rlabel metal2 s 15216 14220 15216 14220 4 gnd
port 514 nsew
rlabel metal2 s 15984 12877 15984 12877 4 gnd
port 514 nsew
rlabel metal2 s 15984 15247 15984 15247 4 gnd
port 514 nsew
rlabel metal2 s 16464 12877 16464 12877 4 gnd
port 514 nsew
rlabel metal2 s 15984 15800 15984 15800 4 gnd
port 514 nsew
rlabel metal2 s 17232 12877 17232 12877 4 gnd
port 514 nsew
rlabel metal2 s 15216 13983 15216 13983 4 gnd
port 514 nsew
rlabel metal2 s 17232 14220 17232 14220 4 gnd
port 514 nsew
rlabel metal2 s 15216 13430 15216 13430 4 gnd
port 514 nsew
rlabel metal2 s 15984 13193 15984 13193 4 gnd
port 514 nsew
rlabel metal2 s 17232 13430 17232 13430 4 gnd
port 514 nsew
rlabel metal2 s 15984 13983 15984 13983 4 gnd
port 514 nsew
rlabel metal2 s 15984 15010 15984 15010 4 gnd
port 514 nsew
rlabel metal2 s 17232 15800 17232 15800 4 gnd
port 514 nsew
rlabel metal2 s 15984 14220 15984 14220 4 gnd
port 514 nsew
rlabel metal2 s 15216 13193 15216 13193 4 gnd
port 514 nsew
rlabel metal2 s 15984 14773 15984 14773 4 gnd
port 514 nsew
rlabel metal2 s 17232 13193 17232 13193 4 gnd
port 514 nsew
rlabel metal2 s 17232 15563 17232 15563 4 gnd
port 514 nsew
rlabel metal2 s 15984 14457 15984 14457 4 gnd
port 514 nsew
rlabel metal2 s 15216 14773 15216 14773 4 gnd
port 514 nsew
rlabel metal2 s 17232 15247 17232 15247 4 gnd
port 514 nsew
rlabel metal2 s 15216 15800 15216 15800 4 gnd
port 514 nsew
rlabel metal2 s 19968 13303 19968 13303 4 wl1_33
port 324 nsew
rlabel metal2 s 18960 13430 18960 13430 4 gnd
port 514 nsew
rlabel metal2 s 19968 13083 19968 13083 4 wl0_33
port 323 nsew
rlabel metal2 s 18480 15800 18480 15800 4 gnd
port 514 nsew
rlabel metal2 s 18480 15247 18480 15247 4 gnd
port 514 nsew
rlabel metal2 s 19968 15453 19968 15453 4 wl0_39
port 335 nsew
rlabel metal2 s 17712 15010 17712 15010 4 gnd
port 514 nsew
rlabel metal2 s 17712 13667 17712 13667 4 gnd
port 514 nsew
rlabel metal2 s 17712 15563 17712 15563 4 gnd
port 514 nsew
rlabel metal2 s 19968 15357 19968 15357 4 wl0_38
port 333 nsew
rlabel metal2 s 19968 14347 19968 14347 4 wl1_36
port 330 nsew
rlabel metal2 s 17712 13430 17712 13430 4 gnd
port 514 nsew
rlabel metal2 s 18960 14773 18960 14773 4 gnd
port 514 nsew
rlabel metal2 s 19968 13557 19968 13557 4 wl1_34
port 326 nsew
rlabel metal2 s 18480 13430 18480 13430 4 gnd
port 514 nsew
rlabel metal2 s 19728 15247 19728 15247 4 gnd
port 514 nsew
rlabel metal2 s 19728 13983 19728 13983 4 gnd
port 514 nsew
rlabel metal2 s 17712 14220 17712 14220 4 gnd
port 514 nsew
rlabel metal2 s 18480 14220 18480 14220 4 gnd
port 514 nsew
rlabel metal2 s 19728 15010 19728 15010 4 gnd
port 514 nsew
rlabel metal2 s 19728 14457 19728 14457 4 gnd
port 514 nsew
rlabel metal2 s 19968 14567 19968 14567 4 wl0_36
port 329 nsew
rlabel metal2 s 18960 13667 18960 13667 4 gnd
port 514 nsew
rlabel metal2 s 18960 14220 18960 14220 4 gnd
port 514 nsew
rlabel metal2 s 18960 14457 18960 14457 4 gnd
port 514 nsew
rlabel metal2 s 18960 12877 18960 12877 4 gnd
port 514 nsew
rlabel metal2 s 18480 15563 18480 15563 4 gnd
port 514 nsew
rlabel metal2 s 19968 14883 19968 14883 4 wl1_37
port 332 nsew
rlabel metal2 s 19968 13873 19968 13873 4 wl0_35
port 327 nsew
rlabel metal2 s 19968 15137 19968 15137 4 wl1_38
port 334 nsew
rlabel metal2 s 18960 15010 18960 15010 4 gnd
port 514 nsew
rlabel metal2 s 19728 14220 19728 14220 4 gnd
port 514 nsew
rlabel metal2 s 18480 13983 18480 13983 4 gnd
port 514 nsew
rlabel metal2 s 17712 14773 17712 14773 4 gnd
port 514 nsew
rlabel metal2 s 19728 15563 19728 15563 4 gnd
port 514 nsew
rlabel metal2 s 17712 13983 17712 13983 4 gnd
port 514 nsew
rlabel metal2 s 18480 15010 18480 15010 4 gnd
port 514 nsew
rlabel metal2 s 18960 15800 18960 15800 4 gnd
port 514 nsew
rlabel metal2 s 18480 14773 18480 14773 4 gnd
port 514 nsew
rlabel metal2 s 19728 12877 19728 12877 4 gnd
port 514 nsew
rlabel metal2 s 17712 12877 17712 12877 4 gnd
port 514 nsew
rlabel metal2 s 19728 13430 19728 13430 4 gnd
port 514 nsew
rlabel metal2 s 17712 13193 17712 13193 4 gnd
port 514 nsew
rlabel metal2 s 17712 15247 17712 15247 4 gnd
port 514 nsew
rlabel metal2 s 18960 13983 18960 13983 4 gnd
port 514 nsew
rlabel metal2 s 19968 14663 19968 14663 4 wl0_37
port 331 nsew
rlabel metal2 s 18480 14457 18480 14457 4 gnd
port 514 nsew
rlabel metal2 s 18960 13193 18960 13193 4 gnd
port 514 nsew
rlabel metal2 s 19968 12767 19968 12767 4 wl1_32
port 322 nsew
rlabel metal2 s 19968 15673 19968 15673 4 wl1_39
port 336 nsew
rlabel metal2 s 19728 13667 19728 13667 4 gnd
port 514 nsew
rlabel metal2 s 18960 15563 18960 15563 4 gnd
port 514 nsew
rlabel metal2 s 19728 13193 19728 13193 4 gnd
port 514 nsew
rlabel metal2 s 17712 14457 17712 14457 4 gnd
port 514 nsew
rlabel metal2 s 18480 13193 18480 13193 4 gnd
port 514 nsew
rlabel metal2 s 19728 14773 19728 14773 4 gnd
port 514 nsew
rlabel metal2 s 19728 15800 19728 15800 4 gnd
port 514 nsew
rlabel metal2 s 18480 13667 18480 13667 4 gnd
port 514 nsew
rlabel metal2 s 18960 15247 18960 15247 4 gnd
port 514 nsew
rlabel metal2 s 18480 12877 18480 12877 4 gnd
port 514 nsew
rlabel metal2 s 19968 12987 19968 12987 4 wl0_32
port 321 nsew
rlabel metal2 s 17712 15800 17712 15800 4 gnd
port 514 nsew
rlabel metal2 s 19968 14093 19968 14093 4 wl1_35
port 328 nsew
rlabel metal2 s 19968 13777 19968 13777 4 wl0_34
port 325 nsew
rlabel metal2 s 7728 24253 7728 24253 4 gnd
port 514 nsew
rlabel metal2 s 9744 25280 9744 25280 4 gnd
port 514 nsew
rlabel metal2 s 7728 22910 7728 22910 4 gnd
port 514 nsew
rlabel metal2 s 8976 25280 8976 25280 4 gnd
port 514 nsew
rlabel metal2 s 9744 23463 9744 23463 4 gnd
port 514 nsew
rlabel metal2 s 8496 22910 8496 22910 4 gnd
port 514 nsew
rlabel metal2 s 8976 23463 8976 23463 4 gnd
port 514 nsew
rlabel metal2 s 9744 24253 9744 24253 4 gnd
port 514 nsew
rlabel metal2 s 7728 23147 7728 23147 4 gnd
port 514 nsew
rlabel metal2 s 8976 23147 8976 23147 4 gnd
port 514 nsew
rlabel metal2 s 8496 23463 8496 23463 4 gnd
port 514 nsew
rlabel metal2 s 7728 24727 7728 24727 4 gnd
port 514 nsew
rlabel metal2 s 8976 25043 8976 25043 4 gnd
port 514 nsew
rlabel metal2 s 9744 23700 9744 23700 4 gnd
port 514 nsew
rlabel metal2 s 9744 23937 9744 23937 4 gnd
port 514 nsew
rlabel metal2 s 8496 24253 8496 24253 4 gnd
port 514 nsew
rlabel metal2 s 8496 24490 8496 24490 4 gnd
port 514 nsew
rlabel metal2 s 8496 23700 8496 23700 4 gnd
port 514 nsew
rlabel metal2 s 7728 24490 7728 24490 4 gnd
port 514 nsew
rlabel metal2 s 7728 25280 7728 25280 4 gnd
port 514 nsew
rlabel metal2 s 8976 23937 8976 23937 4 gnd
port 514 nsew
rlabel metal2 s 8976 24727 8976 24727 4 gnd
port 514 nsew
rlabel metal2 s 8496 22357 8496 22357 4 gnd
port 514 nsew
rlabel metal2 s 8976 22357 8976 22357 4 gnd
port 514 nsew
rlabel metal2 s 7728 23463 7728 23463 4 gnd
port 514 nsew
rlabel metal2 s 7728 25043 7728 25043 4 gnd
port 514 nsew
rlabel metal2 s 9744 25043 9744 25043 4 gnd
port 514 nsew
rlabel metal2 s 9744 24727 9744 24727 4 gnd
port 514 nsew
rlabel metal2 s 7728 22673 7728 22673 4 gnd
port 514 nsew
rlabel metal2 s 9744 22357 9744 22357 4 gnd
port 514 nsew
rlabel metal2 s 8976 24253 8976 24253 4 gnd
port 514 nsew
rlabel metal2 s 8496 25043 8496 25043 4 gnd
port 514 nsew
rlabel metal2 s 8496 23147 8496 23147 4 gnd
port 514 nsew
rlabel metal2 s 7728 22357 7728 22357 4 gnd
port 514 nsew
rlabel metal2 s 8976 22673 8976 22673 4 gnd
port 514 nsew
rlabel metal2 s 8496 25280 8496 25280 4 gnd
port 514 nsew
rlabel metal2 s 8496 22673 8496 22673 4 gnd
port 514 nsew
rlabel metal2 s 9744 24490 9744 24490 4 gnd
port 514 nsew
rlabel metal2 s 8976 23700 8976 23700 4 gnd
port 514 nsew
rlabel metal2 s 8976 22910 8976 22910 4 gnd
port 514 nsew
rlabel metal2 s 7728 23700 7728 23700 4 gnd
port 514 nsew
rlabel metal2 s 8496 23937 8496 23937 4 gnd
port 514 nsew
rlabel metal2 s 9744 23147 9744 23147 4 gnd
port 514 nsew
rlabel metal2 s 8496 24727 8496 24727 4 gnd
port 514 nsew
rlabel metal2 s 9744 22910 9744 22910 4 gnd
port 514 nsew
rlabel metal2 s 7728 23937 7728 23937 4 gnd
port 514 nsew
rlabel metal2 s 9744 22673 9744 22673 4 gnd
port 514 nsew
rlabel metal2 s 8976 24490 8976 24490 4 gnd
port 514 nsew
rlabel metal2 s 6000 25280 6000 25280 4 gnd
port 514 nsew
rlabel metal2 s 7248 24253 7248 24253 4 gnd
port 514 nsew
rlabel metal2 s 7248 22910 7248 22910 4 gnd
port 514 nsew
rlabel metal2 s 5232 23463 5232 23463 4 gnd
port 514 nsew
rlabel metal2 s 6480 24490 6480 24490 4 gnd
port 514 nsew
rlabel metal2 s 6480 23700 6480 23700 4 gnd
port 514 nsew
rlabel metal2 s 5232 25280 5232 25280 4 gnd
port 514 nsew
rlabel metal2 s 6480 23147 6480 23147 4 gnd
port 514 nsew
rlabel metal2 s 7248 24727 7248 24727 4 gnd
port 514 nsew
rlabel metal2 s 5232 23700 5232 23700 4 gnd
port 514 nsew
rlabel metal2 s 5232 25043 5232 25043 4 gnd
port 514 nsew
rlabel metal2 s 6000 22673 6000 22673 4 gnd
port 514 nsew
rlabel metal2 s 6000 24727 6000 24727 4 gnd
port 514 nsew
rlabel metal2 s 6000 22357 6000 22357 4 gnd
port 514 nsew
rlabel metal2 s 6480 25280 6480 25280 4 gnd
port 514 nsew
rlabel metal2 s 5232 24253 5232 24253 4 gnd
port 514 nsew
rlabel metal2 s 5232 23147 5232 23147 4 gnd
port 514 nsew
rlabel metal2 s 6000 24253 6000 24253 4 gnd
port 514 nsew
rlabel metal2 s 7248 22357 7248 22357 4 gnd
port 514 nsew
rlabel metal2 s 6480 22357 6480 22357 4 gnd
port 514 nsew
rlabel metal2 s 7248 22673 7248 22673 4 gnd
port 514 nsew
rlabel metal2 s 5232 23937 5232 23937 4 gnd
port 514 nsew
rlabel metal2 s 6480 23463 6480 23463 4 gnd
port 514 nsew
rlabel metal2 s 5232 24727 5232 24727 4 gnd
port 514 nsew
rlabel metal2 s 6000 25043 6000 25043 4 gnd
port 514 nsew
rlabel metal2 s 6000 23937 6000 23937 4 gnd
port 514 nsew
rlabel metal2 s 5232 22910 5232 22910 4 gnd
port 514 nsew
rlabel metal2 s 7248 25043 7248 25043 4 gnd
port 514 nsew
rlabel metal2 s 6480 22673 6480 22673 4 gnd
port 514 nsew
rlabel metal2 s 6000 23463 6000 23463 4 gnd
port 514 nsew
rlabel metal2 s 7248 23147 7248 23147 4 gnd
port 514 nsew
rlabel metal2 s 6480 22910 6480 22910 4 gnd
port 514 nsew
rlabel metal2 s 5232 24490 5232 24490 4 gnd
port 514 nsew
rlabel metal2 s 6000 24490 6000 24490 4 gnd
port 514 nsew
rlabel metal2 s 6480 24727 6480 24727 4 gnd
port 514 nsew
rlabel metal2 s 6480 24253 6480 24253 4 gnd
port 514 nsew
rlabel metal2 s 7248 25280 7248 25280 4 gnd
port 514 nsew
rlabel metal2 s 7248 23937 7248 23937 4 gnd
port 514 nsew
rlabel metal2 s 6000 23700 6000 23700 4 gnd
port 514 nsew
rlabel metal2 s 5232 22357 5232 22357 4 gnd
port 514 nsew
rlabel metal2 s 6480 25043 6480 25043 4 gnd
port 514 nsew
rlabel metal2 s 6480 23937 6480 23937 4 gnd
port 514 nsew
rlabel metal2 s 6000 22910 6000 22910 4 gnd
port 514 nsew
rlabel metal2 s 5232 22673 5232 22673 4 gnd
port 514 nsew
rlabel metal2 s 7248 23700 7248 23700 4 gnd
port 514 nsew
rlabel metal2 s 7248 24490 7248 24490 4 gnd
port 514 nsew
rlabel metal2 s 7248 23463 7248 23463 4 gnd
port 514 nsew
rlabel metal2 s 6000 23147 6000 23147 4 gnd
port 514 nsew
rlabel metal2 s 6000 20777 6000 20777 4 gnd
port 514 nsew
rlabel metal2 s 5232 19197 5232 19197 4 gnd
port 514 nsew
rlabel metal2 s 5232 20777 5232 20777 4 gnd
port 514 nsew
rlabel metal2 s 5232 19750 5232 19750 4 gnd
port 514 nsew
rlabel metal2 s 5232 21567 5232 21567 4 gnd
port 514 nsew
rlabel metal2 s 7248 19750 7248 19750 4 gnd
port 514 nsew
rlabel metal2 s 7248 22120 7248 22120 4 gnd
port 514 nsew
rlabel metal2 s 6000 21883 6000 21883 4 gnd
port 514 nsew
rlabel metal2 s 5232 19987 5232 19987 4 gnd
port 514 nsew
rlabel metal2 s 6000 19513 6000 19513 4 gnd
port 514 nsew
rlabel metal2 s 6480 22120 6480 22120 4 gnd
port 514 nsew
rlabel metal2 s 6480 19197 6480 19197 4 gnd
port 514 nsew
rlabel metal2 s 6480 21093 6480 21093 4 gnd
port 514 nsew
rlabel metal2 s 6000 19987 6000 19987 4 gnd
port 514 nsew
rlabel metal2 s 6480 21883 6480 21883 4 gnd
port 514 nsew
rlabel metal2 s 5232 22120 5232 22120 4 gnd
port 514 nsew
rlabel metal2 s 7248 19513 7248 19513 4 gnd
port 514 nsew
rlabel metal2 s 7248 19987 7248 19987 4 gnd
port 514 nsew
rlabel metal2 s 6000 21567 6000 21567 4 gnd
port 514 nsew
rlabel metal2 s 6480 19750 6480 19750 4 gnd
port 514 nsew
rlabel metal2 s 5232 21883 5232 21883 4 gnd
port 514 nsew
rlabel metal2 s 5232 21093 5232 21093 4 gnd
port 514 nsew
rlabel metal2 s 6480 20777 6480 20777 4 gnd
port 514 nsew
rlabel metal2 s 6480 21567 6480 21567 4 gnd
port 514 nsew
rlabel metal2 s 6480 19513 6480 19513 4 gnd
port 514 nsew
rlabel metal2 s 5232 19513 5232 19513 4 gnd
port 514 nsew
rlabel metal2 s 6000 22120 6000 22120 4 gnd
port 514 nsew
rlabel metal2 s 6480 20540 6480 20540 4 gnd
port 514 nsew
rlabel metal2 s 5232 21330 5232 21330 4 gnd
port 514 nsew
rlabel metal2 s 7248 21093 7248 21093 4 gnd
port 514 nsew
rlabel metal2 s 7248 21883 7248 21883 4 gnd
port 514 nsew
rlabel metal2 s 6000 19750 6000 19750 4 gnd
port 514 nsew
rlabel metal2 s 6000 20303 6000 20303 4 gnd
port 514 nsew
rlabel metal2 s 6000 20540 6000 20540 4 gnd
port 514 nsew
rlabel metal2 s 6000 19197 6000 19197 4 gnd
port 514 nsew
rlabel metal2 s 7248 20540 7248 20540 4 gnd
port 514 nsew
rlabel metal2 s 7248 20777 7248 20777 4 gnd
port 514 nsew
rlabel metal2 s 6480 20303 6480 20303 4 gnd
port 514 nsew
rlabel metal2 s 7248 21330 7248 21330 4 gnd
port 514 nsew
rlabel metal2 s 5232 20540 5232 20540 4 gnd
port 514 nsew
rlabel metal2 s 6480 19987 6480 19987 4 gnd
port 514 nsew
rlabel metal2 s 7248 21567 7248 21567 4 gnd
port 514 nsew
rlabel metal2 s 6000 21330 6000 21330 4 gnd
port 514 nsew
rlabel metal2 s 5232 20303 5232 20303 4 gnd
port 514 nsew
rlabel metal2 s 7248 20303 7248 20303 4 gnd
port 514 nsew
rlabel metal2 s 6480 21330 6480 21330 4 gnd
port 514 nsew
rlabel metal2 s 7248 19197 7248 19197 4 gnd
port 514 nsew
rlabel metal2 s 6000 21093 6000 21093 4 gnd
port 514 nsew
rlabel metal2 s 8976 19513 8976 19513 4 gnd
port 514 nsew
rlabel metal2 s 8976 21883 8976 21883 4 gnd
port 514 nsew
rlabel metal2 s 8496 21567 8496 21567 4 gnd
port 514 nsew
rlabel metal2 s 8976 21093 8976 21093 4 gnd
port 514 nsew
rlabel metal2 s 8976 20540 8976 20540 4 gnd
port 514 nsew
rlabel metal2 s 9744 22120 9744 22120 4 gnd
port 514 nsew
rlabel metal2 s 9744 21093 9744 21093 4 gnd
port 514 nsew
rlabel metal2 s 8496 19513 8496 19513 4 gnd
port 514 nsew
rlabel metal2 s 9744 20303 9744 20303 4 gnd
port 514 nsew
rlabel metal2 s 9744 20540 9744 20540 4 gnd
port 514 nsew
rlabel metal2 s 7728 20777 7728 20777 4 gnd
port 514 nsew
rlabel metal2 s 8496 19197 8496 19197 4 gnd
port 514 nsew
rlabel metal2 s 8976 19987 8976 19987 4 gnd
port 514 nsew
rlabel metal2 s 7728 20540 7728 20540 4 gnd
port 514 nsew
rlabel metal2 s 8496 20303 8496 20303 4 gnd
port 514 nsew
rlabel metal2 s 7728 19987 7728 19987 4 gnd
port 514 nsew
rlabel metal2 s 9744 21330 9744 21330 4 gnd
port 514 nsew
rlabel metal2 s 7728 20303 7728 20303 4 gnd
port 514 nsew
rlabel metal2 s 7728 21330 7728 21330 4 gnd
port 514 nsew
rlabel metal2 s 9744 19750 9744 19750 4 gnd
port 514 nsew
rlabel metal2 s 7728 21093 7728 21093 4 gnd
port 514 nsew
rlabel metal2 s 8496 21093 8496 21093 4 gnd
port 514 nsew
rlabel metal2 s 9744 19987 9744 19987 4 gnd
port 514 nsew
rlabel metal2 s 8496 20540 8496 20540 4 gnd
port 514 nsew
rlabel metal2 s 8496 19987 8496 19987 4 gnd
port 514 nsew
rlabel metal2 s 9744 21567 9744 21567 4 gnd
port 514 nsew
rlabel metal2 s 7728 19197 7728 19197 4 gnd
port 514 nsew
rlabel metal2 s 8976 20303 8976 20303 4 gnd
port 514 nsew
rlabel metal2 s 7728 21883 7728 21883 4 gnd
port 514 nsew
rlabel metal2 s 8976 19750 8976 19750 4 gnd
port 514 nsew
rlabel metal2 s 8976 21567 8976 21567 4 gnd
port 514 nsew
rlabel metal2 s 7728 19513 7728 19513 4 gnd
port 514 nsew
rlabel metal2 s 7728 19750 7728 19750 4 gnd
port 514 nsew
rlabel metal2 s 8496 21330 8496 21330 4 gnd
port 514 nsew
rlabel metal2 s 7728 21567 7728 21567 4 gnd
port 514 nsew
rlabel metal2 s 9744 19197 9744 19197 4 gnd
port 514 nsew
rlabel metal2 s 8496 22120 8496 22120 4 gnd
port 514 nsew
rlabel metal2 s 8976 20777 8976 20777 4 gnd
port 514 nsew
rlabel metal2 s 8496 19750 8496 19750 4 gnd
port 514 nsew
rlabel metal2 s 8496 20777 8496 20777 4 gnd
port 514 nsew
rlabel metal2 s 7728 22120 7728 22120 4 gnd
port 514 nsew
rlabel metal2 s 8496 21883 8496 21883 4 gnd
port 514 nsew
rlabel metal2 s 9744 19513 9744 19513 4 gnd
port 514 nsew
rlabel metal2 s 8976 21330 8976 21330 4 gnd
port 514 nsew
rlabel metal2 s 8976 22120 8976 22120 4 gnd
port 514 nsew
rlabel metal2 s 9744 20777 9744 20777 4 gnd
port 514 nsew
rlabel metal2 s 9744 21883 9744 21883 4 gnd
port 514 nsew
rlabel metal2 s 8976 19197 8976 19197 4 gnd
port 514 nsew
rlabel metal2 s 3984 23463 3984 23463 4 gnd
port 514 nsew
rlabel metal2 s 2736 23937 2736 23937 4 gnd
port 514 nsew
rlabel metal2 s 2736 22357 2736 22357 4 gnd
port 514 nsew
rlabel metal2 s 2736 24490 2736 24490 4 gnd
port 514 nsew
rlabel metal2 s 3504 23700 3504 23700 4 gnd
port 514 nsew
rlabel metal2 s 4752 24490 4752 24490 4 gnd
port 514 nsew
rlabel metal2 s 4752 23463 4752 23463 4 gnd
port 514 nsew
rlabel metal2 s 2736 24253 2736 24253 4 gnd
port 514 nsew
rlabel metal2 s 3984 22673 3984 22673 4 gnd
port 514 nsew
rlabel metal2 s 4752 25043 4752 25043 4 gnd
port 514 nsew
rlabel metal2 s 4752 23147 4752 23147 4 gnd
port 514 nsew
rlabel metal2 s 3984 23700 3984 23700 4 gnd
port 514 nsew
rlabel metal2 s 4752 23937 4752 23937 4 gnd
port 514 nsew
rlabel metal2 s 2736 25043 2736 25043 4 gnd
port 514 nsew
rlabel metal2 s 4752 22673 4752 22673 4 gnd
port 514 nsew
rlabel metal2 s 3984 22910 3984 22910 4 gnd
port 514 nsew
rlabel metal2 s 3984 25280 3984 25280 4 gnd
port 514 nsew
rlabel metal2 s 4752 24253 4752 24253 4 gnd
port 514 nsew
rlabel metal2 s 3984 23147 3984 23147 4 gnd
port 514 nsew
rlabel metal2 s 2736 22910 2736 22910 4 gnd
port 514 nsew
rlabel metal2 s 3984 24253 3984 24253 4 gnd
port 514 nsew
rlabel metal2 s 3504 23147 3504 23147 4 gnd
port 514 nsew
rlabel metal2 s 3504 24253 3504 24253 4 gnd
port 514 nsew
rlabel metal2 s 3504 22673 3504 22673 4 gnd
port 514 nsew
rlabel metal2 s 3504 23463 3504 23463 4 gnd
port 514 nsew
rlabel metal2 s 3504 23937 3504 23937 4 gnd
port 514 nsew
rlabel metal2 s 3504 22357 3504 22357 4 gnd
port 514 nsew
rlabel metal2 s 2736 25280 2736 25280 4 gnd
port 514 nsew
rlabel metal2 s 3504 22910 3504 22910 4 gnd
port 514 nsew
rlabel metal2 s 3984 24727 3984 24727 4 gnd
port 514 nsew
rlabel metal2 s 3984 23937 3984 23937 4 gnd
port 514 nsew
rlabel metal2 s 3984 22357 3984 22357 4 gnd
port 514 nsew
rlabel metal2 s 3504 25043 3504 25043 4 gnd
port 514 nsew
rlabel metal2 s 3504 24490 3504 24490 4 gnd
port 514 nsew
rlabel metal2 s 4752 24727 4752 24727 4 gnd
port 514 nsew
rlabel metal2 s 2736 23463 2736 23463 4 gnd
port 514 nsew
rlabel metal2 s 3504 24727 3504 24727 4 gnd
port 514 nsew
rlabel metal2 s 4752 22357 4752 22357 4 gnd
port 514 nsew
rlabel metal2 s 4752 25280 4752 25280 4 gnd
port 514 nsew
rlabel metal2 s 3504 25280 3504 25280 4 gnd
port 514 nsew
rlabel metal2 s 3984 25043 3984 25043 4 gnd
port 514 nsew
rlabel metal2 s 4752 23700 4752 23700 4 gnd
port 514 nsew
rlabel metal2 s 2736 23147 2736 23147 4 gnd
port 514 nsew
rlabel metal2 s 2736 23700 2736 23700 4 gnd
port 514 nsew
rlabel metal2 s 2736 24727 2736 24727 4 gnd
port 514 nsew
rlabel metal2 s 2736 22673 2736 22673 4 gnd
port 514 nsew
rlabel metal2 s 3984 24490 3984 24490 4 gnd
port 514 nsew
rlabel metal2 s 4752 22910 4752 22910 4 gnd
port 514 nsew
rlabel metal2 s 2256 23937 2256 23937 4 gnd
port 514 nsew
rlabel metal2 s 1008 23147 1008 23147 4 gnd
port 514 nsew
rlabel metal2 s 240 23463 240 23463 4 gnd
port 514 nsew
rlabel metal2 s 1008 25043 1008 25043 4 gnd
port 514 nsew
rlabel metal2 s 1008 22673 1008 22673 4 gnd
port 514 nsew
rlabel metal2 s 1488 23147 1488 23147 4 gnd
port 514 nsew
rlabel metal2 s 1008 23937 1008 23937 4 gnd
port 514 nsew
rlabel metal2 s 2256 24253 2256 24253 4 gnd
port 514 nsew
rlabel metal2 s 1488 24727 1488 24727 4 gnd
port 514 nsew
rlabel metal2 s 2256 23700 2256 23700 4 gnd
port 514 nsew
rlabel metal2 s 2256 24727 2256 24727 4 gnd
port 514 nsew
rlabel metal2 s 1488 25280 1488 25280 4 gnd
port 514 nsew
rlabel metal2 s 1488 25043 1488 25043 4 gnd
port 514 nsew
rlabel metal2 s 2256 23463 2256 23463 4 gnd
port 514 nsew
rlabel metal2 s 1008 23463 1008 23463 4 gnd
port 514 nsew
rlabel metal2 s 240 23700 240 23700 4 gnd
port 514 nsew
rlabel metal2 s 240 25043 240 25043 4 gnd
port 514 nsew
rlabel metal2 s 2256 25043 2256 25043 4 gnd
port 514 nsew
rlabel metal2 s 1008 25280 1008 25280 4 gnd
port 514 nsew
rlabel metal2 s 2256 22357 2256 22357 4 gnd
port 514 nsew
rlabel metal2 s 1008 24727 1008 24727 4 gnd
port 514 nsew
rlabel metal2 s 2256 24490 2256 24490 4 gnd
port 514 nsew
rlabel metal2 s 240 22910 240 22910 4 gnd
port 514 nsew
rlabel metal2 s 1488 22673 1488 22673 4 gnd
port 514 nsew
rlabel metal2 s 240 23147 240 23147 4 gnd
port 514 nsew
rlabel metal2 s 1488 23700 1488 23700 4 gnd
port 514 nsew
rlabel metal2 s 1008 22357 1008 22357 4 gnd
port 514 nsew
rlabel metal2 s 2256 22910 2256 22910 4 gnd
port 514 nsew
rlabel metal2 s 240 24727 240 24727 4 gnd
port 514 nsew
rlabel metal2 s 1008 24253 1008 24253 4 gnd
port 514 nsew
rlabel metal2 s 240 25280 240 25280 4 gnd
port 514 nsew
rlabel metal2 s 1488 23937 1488 23937 4 gnd
port 514 nsew
rlabel metal2 s 1008 22910 1008 22910 4 gnd
port 514 nsew
rlabel metal2 s 2256 23147 2256 23147 4 gnd
port 514 nsew
rlabel metal2 s 1008 24490 1008 24490 4 gnd
port 514 nsew
rlabel metal2 s 240 24490 240 24490 4 gnd
port 514 nsew
rlabel metal2 s 1488 24490 1488 24490 4 gnd
port 514 nsew
rlabel metal2 s 240 22673 240 22673 4 gnd
port 514 nsew
rlabel metal2 s 2256 25280 2256 25280 4 gnd
port 514 nsew
rlabel metal2 s 240 24253 240 24253 4 gnd
port 514 nsew
rlabel metal2 s 1488 23463 1488 23463 4 gnd
port 514 nsew
rlabel metal2 s 1488 22357 1488 22357 4 gnd
port 514 nsew
rlabel metal2 s 2256 22673 2256 22673 4 gnd
port 514 nsew
rlabel metal2 s 1008 23700 1008 23700 4 gnd
port 514 nsew
rlabel metal2 s 240 22357 240 22357 4 gnd
port 514 nsew
rlabel metal2 s 1488 24253 1488 24253 4 gnd
port 514 nsew
rlabel metal2 s 240 23937 240 23937 4 gnd
port 514 nsew
rlabel metal2 s 1488 22910 1488 22910 4 gnd
port 514 nsew
rlabel metal2 s 2256 19197 2256 19197 4 gnd
port 514 nsew
rlabel metal2 s 240 20777 240 20777 4 gnd
port 514 nsew
rlabel metal2 s 1488 19750 1488 19750 4 gnd
port 514 nsew
rlabel metal2 s 240 21883 240 21883 4 gnd
port 514 nsew
rlabel metal2 s 2256 19513 2256 19513 4 gnd
port 514 nsew
rlabel metal2 s 1008 20303 1008 20303 4 gnd
port 514 nsew
rlabel metal2 s 2256 19987 2256 19987 4 gnd
port 514 nsew
rlabel metal2 s 1008 22120 1008 22120 4 gnd
port 514 nsew
rlabel metal2 s 1488 21883 1488 21883 4 gnd
port 514 nsew
rlabel metal2 s 1008 19750 1008 19750 4 gnd
port 514 nsew
rlabel metal2 s 240 21330 240 21330 4 gnd
port 514 nsew
rlabel metal2 s 1008 20777 1008 20777 4 gnd
port 514 nsew
rlabel metal2 s 240 20540 240 20540 4 gnd
port 514 nsew
rlabel metal2 s 2256 21567 2256 21567 4 gnd
port 514 nsew
rlabel metal2 s 2256 20303 2256 20303 4 gnd
port 514 nsew
rlabel metal2 s 1488 21567 1488 21567 4 gnd
port 514 nsew
rlabel metal2 s 1488 21093 1488 21093 4 gnd
port 514 nsew
rlabel metal2 s 1488 20777 1488 20777 4 gnd
port 514 nsew
rlabel metal2 s 1488 21330 1488 21330 4 gnd
port 514 nsew
rlabel metal2 s 1008 21567 1008 21567 4 gnd
port 514 nsew
rlabel metal2 s 240 21093 240 21093 4 gnd
port 514 nsew
rlabel metal2 s 1008 19513 1008 19513 4 gnd
port 514 nsew
rlabel metal2 s 2256 20540 2256 20540 4 gnd
port 514 nsew
rlabel metal2 s 1008 20540 1008 20540 4 gnd
port 514 nsew
rlabel metal2 s 240 19750 240 19750 4 gnd
port 514 nsew
rlabel metal2 s 2256 19750 2256 19750 4 gnd
port 514 nsew
rlabel metal2 s 1488 19197 1488 19197 4 gnd
port 514 nsew
rlabel metal2 s 1488 20303 1488 20303 4 gnd
port 514 nsew
rlabel metal2 s 240 19197 240 19197 4 gnd
port 514 nsew
rlabel metal2 s 2256 21093 2256 21093 4 gnd
port 514 nsew
rlabel metal2 s 240 21567 240 21567 4 gnd
port 514 nsew
rlabel metal2 s 1488 20540 1488 20540 4 gnd
port 514 nsew
rlabel metal2 s 1008 21883 1008 21883 4 gnd
port 514 nsew
rlabel metal2 s 1008 19987 1008 19987 4 gnd
port 514 nsew
rlabel metal2 s 1488 19987 1488 19987 4 gnd
port 514 nsew
rlabel metal2 s 240 22120 240 22120 4 gnd
port 514 nsew
rlabel metal2 s 2256 21883 2256 21883 4 gnd
port 514 nsew
rlabel metal2 s 1488 19513 1488 19513 4 gnd
port 514 nsew
rlabel metal2 s 2256 21330 2256 21330 4 gnd
port 514 nsew
rlabel metal2 s 240 20303 240 20303 4 gnd
port 514 nsew
rlabel metal2 s 2256 22120 2256 22120 4 gnd
port 514 nsew
rlabel metal2 s 1008 21330 1008 21330 4 gnd
port 514 nsew
rlabel metal2 s 240 19987 240 19987 4 gnd
port 514 nsew
rlabel metal2 s 1008 19197 1008 19197 4 gnd
port 514 nsew
rlabel metal2 s 240 19513 240 19513 4 gnd
port 514 nsew
rlabel metal2 s 2256 20777 2256 20777 4 gnd
port 514 nsew
rlabel metal2 s 1488 22120 1488 22120 4 gnd
port 514 nsew
rlabel metal2 s 1008 21093 1008 21093 4 gnd
port 514 nsew
rlabel metal2 s 2736 19197 2736 19197 4 gnd
port 514 nsew
rlabel metal2 s 3504 19197 3504 19197 4 gnd
port 514 nsew
rlabel metal2 s 4752 22120 4752 22120 4 gnd
port 514 nsew
rlabel metal2 s 3984 20540 3984 20540 4 gnd
port 514 nsew
rlabel metal2 s 4752 20540 4752 20540 4 gnd
port 514 nsew
rlabel metal2 s 3504 19750 3504 19750 4 gnd
port 514 nsew
rlabel metal2 s 2736 22120 2736 22120 4 gnd
port 514 nsew
rlabel metal2 s 4752 21093 4752 21093 4 gnd
port 514 nsew
rlabel metal2 s 3984 19513 3984 19513 4 gnd
port 514 nsew
rlabel metal2 s 2736 21883 2736 21883 4 gnd
port 514 nsew
rlabel metal2 s 3504 22120 3504 22120 4 gnd
port 514 nsew
rlabel metal2 s 2736 19987 2736 19987 4 gnd
port 514 nsew
rlabel metal2 s 3984 21567 3984 21567 4 gnd
port 514 nsew
rlabel metal2 s 2736 19513 2736 19513 4 gnd
port 514 nsew
rlabel metal2 s 3984 19197 3984 19197 4 gnd
port 514 nsew
rlabel metal2 s 3504 21883 3504 21883 4 gnd
port 514 nsew
rlabel metal2 s 3984 21330 3984 21330 4 gnd
port 514 nsew
rlabel metal2 s 2736 20777 2736 20777 4 gnd
port 514 nsew
rlabel metal2 s 3504 21093 3504 21093 4 gnd
port 514 nsew
rlabel metal2 s 4752 21567 4752 21567 4 gnd
port 514 nsew
rlabel metal2 s 4752 19197 4752 19197 4 gnd
port 514 nsew
rlabel metal2 s 4752 21330 4752 21330 4 gnd
port 514 nsew
rlabel metal2 s 2736 21330 2736 21330 4 gnd
port 514 nsew
rlabel metal2 s 3504 20303 3504 20303 4 gnd
port 514 nsew
rlabel metal2 s 3504 19513 3504 19513 4 gnd
port 514 nsew
rlabel metal2 s 3504 20777 3504 20777 4 gnd
port 514 nsew
rlabel metal2 s 2736 19750 2736 19750 4 gnd
port 514 nsew
rlabel metal2 s 3984 19750 3984 19750 4 gnd
port 514 nsew
rlabel metal2 s 4752 21883 4752 21883 4 gnd
port 514 nsew
rlabel metal2 s 2736 21567 2736 21567 4 gnd
port 514 nsew
rlabel metal2 s 3984 20303 3984 20303 4 gnd
port 514 nsew
rlabel metal2 s 3504 20540 3504 20540 4 gnd
port 514 nsew
rlabel metal2 s 4752 20303 4752 20303 4 gnd
port 514 nsew
rlabel metal2 s 4752 19750 4752 19750 4 gnd
port 514 nsew
rlabel metal2 s 3984 20777 3984 20777 4 gnd
port 514 nsew
rlabel metal2 s 3504 19987 3504 19987 4 gnd
port 514 nsew
rlabel metal2 s 3984 19987 3984 19987 4 gnd
port 514 nsew
rlabel metal2 s 3504 21567 3504 21567 4 gnd
port 514 nsew
rlabel metal2 s 4752 20777 4752 20777 4 gnd
port 514 nsew
rlabel metal2 s 2736 21093 2736 21093 4 gnd
port 514 nsew
rlabel metal2 s 4752 19987 4752 19987 4 gnd
port 514 nsew
rlabel metal2 s 3504 21330 3504 21330 4 gnd
port 514 nsew
rlabel metal2 s 3984 21093 3984 21093 4 gnd
port 514 nsew
rlabel metal2 s 4752 19513 4752 19513 4 gnd
port 514 nsew
rlabel metal2 s 3984 21883 3984 21883 4 gnd
port 514 nsew
rlabel metal2 s 2736 20303 2736 20303 4 gnd
port 514 nsew
rlabel metal2 s 2736 20540 2736 20540 4 gnd
port 514 nsew
rlabel metal2 s 3984 22120 3984 22120 4 gnd
port 514 nsew
rlabel metal2 s 3504 17143 3504 17143 4 gnd
port 514 nsew
rlabel metal2 s 3504 17933 3504 17933 4 gnd
port 514 nsew
rlabel metal2 s 2736 17933 2736 17933 4 gnd
port 514 nsew
rlabel metal2 s 3984 16590 3984 16590 4 gnd
port 514 nsew
rlabel metal2 s 3984 18407 3984 18407 4 gnd
port 514 nsew
rlabel metal2 s 3504 17617 3504 17617 4 gnd
port 514 nsew
rlabel metal2 s 4752 17933 4752 17933 4 gnd
port 514 nsew
rlabel metal2 s 3984 18723 3984 18723 4 gnd
port 514 nsew
rlabel metal2 s 2736 18170 2736 18170 4 gnd
port 514 nsew
rlabel metal2 s 2736 17143 2736 17143 4 gnd
port 514 nsew
rlabel metal2 s 4752 18407 4752 18407 4 gnd
port 514 nsew
rlabel metal2 s 2736 16827 2736 16827 4 gnd
port 514 nsew
rlabel metal2 s 2736 16353 2736 16353 4 gnd
port 514 nsew
rlabel metal2 s 2736 18960 2736 18960 4 gnd
port 514 nsew
rlabel metal2 s 3984 17617 3984 17617 4 gnd
port 514 nsew
rlabel metal2 s 3504 17380 3504 17380 4 gnd
port 514 nsew
rlabel metal2 s 4752 16037 4752 16037 4 gnd
port 514 nsew
rlabel metal2 s 4752 18723 4752 18723 4 gnd
port 514 nsew
rlabel metal2 s 3504 16590 3504 16590 4 gnd
port 514 nsew
rlabel metal2 s 4752 16827 4752 16827 4 gnd
port 514 nsew
rlabel metal2 s 3504 18170 3504 18170 4 gnd
port 514 nsew
rlabel metal2 s 3504 18407 3504 18407 4 gnd
port 514 nsew
rlabel metal2 s 4752 16353 4752 16353 4 gnd
port 514 nsew
rlabel metal2 s 2736 16590 2736 16590 4 gnd
port 514 nsew
rlabel metal2 s 3504 16827 3504 16827 4 gnd
port 514 nsew
rlabel metal2 s 3984 17380 3984 17380 4 gnd
port 514 nsew
rlabel metal2 s 3504 18723 3504 18723 4 gnd
port 514 nsew
rlabel metal2 s 4752 18960 4752 18960 4 gnd
port 514 nsew
rlabel metal2 s 3984 16353 3984 16353 4 gnd
port 514 nsew
rlabel metal2 s 2736 18723 2736 18723 4 gnd
port 514 nsew
rlabel metal2 s 3504 16353 3504 16353 4 gnd
port 514 nsew
rlabel metal2 s 2736 16037 2736 16037 4 gnd
port 514 nsew
rlabel metal2 s 3984 18960 3984 18960 4 gnd
port 514 nsew
rlabel metal2 s 3504 16037 3504 16037 4 gnd
port 514 nsew
rlabel metal2 s 4752 16590 4752 16590 4 gnd
port 514 nsew
rlabel metal2 s 4752 18170 4752 18170 4 gnd
port 514 nsew
rlabel metal2 s 3984 16827 3984 16827 4 gnd
port 514 nsew
rlabel metal2 s 3984 16037 3984 16037 4 gnd
port 514 nsew
rlabel metal2 s 4752 17380 4752 17380 4 gnd
port 514 nsew
rlabel metal2 s 2736 18407 2736 18407 4 gnd
port 514 nsew
rlabel metal2 s 3984 18170 3984 18170 4 gnd
port 514 nsew
rlabel metal2 s 2736 17617 2736 17617 4 gnd
port 514 nsew
rlabel metal2 s 4752 17143 4752 17143 4 gnd
port 514 nsew
rlabel metal2 s 3984 17143 3984 17143 4 gnd
port 514 nsew
rlabel metal2 s 4752 17617 4752 17617 4 gnd
port 514 nsew
rlabel metal2 s 3984 17933 3984 17933 4 gnd
port 514 nsew
rlabel metal2 s 3504 18960 3504 18960 4 gnd
port 514 nsew
rlabel metal2 s 2736 17380 2736 17380 4 gnd
port 514 nsew
rlabel metal2 s 1008 16353 1008 16353 4 gnd
port 514 nsew
rlabel metal2 s 2256 17933 2256 17933 4 gnd
port 514 nsew
rlabel metal2 s 2256 16590 2256 16590 4 gnd
port 514 nsew
rlabel metal2 s 240 17617 240 17617 4 gnd
port 514 nsew
rlabel metal2 s 240 18407 240 18407 4 gnd
port 514 nsew
rlabel metal2 s 2256 17143 2256 17143 4 gnd
port 514 nsew
rlabel metal2 s 1008 17933 1008 17933 4 gnd
port 514 nsew
rlabel metal2 s 240 18723 240 18723 4 gnd
port 514 nsew
rlabel metal2 s 1008 16827 1008 16827 4 gnd
port 514 nsew
rlabel metal2 s 240 16590 240 16590 4 gnd
port 514 nsew
rlabel metal2 s 2256 18407 2256 18407 4 gnd
port 514 nsew
rlabel metal2 s 1008 17143 1008 17143 4 gnd
port 514 nsew
rlabel metal2 s 1488 17380 1488 17380 4 gnd
port 514 nsew
rlabel metal2 s 1488 17143 1488 17143 4 gnd
port 514 nsew
rlabel metal2 s 1008 16037 1008 16037 4 gnd
port 514 nsew
rlabel metal2 s 2256 18960 2256 18960 4 gnd
port 514 nsew
rlabel metal2 s 2256 18170 2256 18170 4 gnd
port 514 nsew
rlabel metal2 s 1488 16037 1488 16037 4 gnd
port 514 nsew
rlabel metal2 s 2256 16037 2256 16037 4 gnd
port 514 nsew
rlabel metal2 s 2256 17617 2256 17617 4 gnd
port 514 nsew
rlabel metal2 s 1488 18170 1488 18170 4 gnd
port 514 nsew
rlabel metal2 s 1488 16827 1488 16827 4 gnd
port 514 nsew
rlabel metal2 s 1008 18170 1008 18170 4 gnd
port 514 nsew
rlabel metal2 s 1008 17380 1008 17380 4 gnd
port 514 nsew
rlabel metal2 s 1008 16590 1008 16590 4 gnd
port 514 nsew
rlabel metal2 s 1008 18723 1008 18723 4 gnd
port 514 nsew
rlabel metal2 s 1488 17617 1488 17617 4 gnd
port 514 nsew
rlabel metal2 s 2256 16827 2256 16827 4 gnd
port 514 nsew
rlabel metal2 s 2256 16353 2256 16353 4 gnd
port 514 nsew
rlabel metal2 s 2256 18723 2256 18723 4 gnd
port 514 nsew
rlabel metal2 s 240 17380 240 17380 4 gnd
port 514 nsew
rlabel metal2 s 240 17143 240 17143 4 gnd
port 514 nsew
rlabel metal2 s 240 16353 240 16353 4 gnd
port 514 nsew
rlabel metal2 s 240 17933 240 17933 4 gnd
port 514 nsew
rlabel metal2 s 1008 18407 1008 18407 4 gnd
port 514 nsew
rlabel metal2 s 1488 18407 1488 18407 4 gnd
port 514 nsew
rlabel metal2 s 1488 18723 1488 18723 4 gnd
port 514 nsew
rlabel metal2 s 1008 17617 1008 17617 4 gnd
port 514 nsew
rlabel metal2 s 1488 18960 1488 18960 4 gnd
port 514 nsew
rlabel metal2 s 240 16827 240 16827 4 gnd
port 514 nsew
rlabel metal2 s 1488 16353 1488 16353 4 gnd
port 514 nsew
rlabel metal2 s 240 18960 240 18960 4 gnd
port 514 nsew
rlabel metal2 s 1008 18960 1008 18960 4 gnd
port 514 nsew
rlabel metal2 s 240 18170 240 18170 4 gnd
port 514 nsew
rlabel metal2 s 1488 16590 1488 16590 4 gnd
port 514 nsew
rlabel metal2 s 2256 17380 2256 17380 4 gnd
port 514 nsew
rlabel metal2 s 240 16037 240 16037 4 gnd
port 514 nsew
rlabel metal2 s 1488 17933 1488 17933 4 gnd
port 514 nsew
rlabel metal2 s 2256 15010 2256 15010 4 gnd
port 514 nsew
rlabel metal2 s 1008 12877 1008 12877 4 gnd
port 514 nsew
rlabel metal2 s 1008 13430 1008 13430 4 gnd
port 514 nsew
rlabel metal2 s 1008 15563 1008 15563 4 gnd
port 514 nsew
rlabel metal2 s 1008 13983 1008 13983 4 gnd
port 514 nsew
rlabel metal2 s 2256 12877 2256 12877 4 gnd
port 514 nsew
rlabel metal2 s 1488 15563 1488 15563 4 gnd
port 514 nsew
rlabel metal2 s 1008 15247 1008 15247 4 gnd
port 514 nsew
rlabel metal2 s 1488 13667 1488 13667 4 gnd
port 514 nsew
rlabel metal2 s 240 13667 240 13667 4 gnd
port 514 nsew
rlabel metal2 s 2256 14457 2256 14457 4 gnd
port 514 nsew
rlabel metal2 s 1488 15247 1488 15247 4 gnd
port 514 nsew
rlabel metal2 s 240 15563 240 15563 4 gnd
port 514 nsew
rlabel metal2 s 1008 13193 1008 13193 4 gnd
port 514 nsew
rlabel metal2 s 240 13430 240 13430 4 gnd
port 514 nsew
rlabel metal2 s 1488 15800 1488 15800 4 gnd
port 514 nsew
rlabel metal2 s 1008 14220 1008 14220 4 gnd
port 514 nsew
rlabel metal2 s 1488 12877 1488 12877 4 gnd
port 514 nsew
rlabel metal2 s 2256 13667 2256 13667 4 gnd
port 514 nsew
rlabel metal2 s 1008 14457 1008 14457 4 gnd
port 514 nsew
rlabel metal2 s 240 14457 240 14457 4 gnd
port 514 nsew
rlabel metal2 s 1488 13430 1488 13430 4 gnd
port 514 nsew
rlabel metal2 s 1488 14773 1488 14773 4 gnd
port 514 nsew
rlabel metal2 s 240 13193 240 13193 4 gnd
port 514 nsew
rlabel metal2 s 240 14773 240 14773 4 gnd
port 514 nsew
rlabel metal2 s 1488 13983 1488 13983 4 gnd
port 514 nsew
rlabel metal2 s 1488 13193 1488 13193 4 gnd
port 514 nsew
rlabel metal2 s 240 13983 240 13983 4 gnd
port 514 nsew
rlabel metal2 s 2256 14220 2256 14220 4 gnd
port 514 nsew
rlabel metal2 s 1488 15010 1488 15010 4 gnd
port 514 nsew
rlabel metal2 s 2256 13430 2256 13430 4 gnd
port 514 nsew
rlabel metal2 s 240 12877 240 12877 4 gnd
port 514 nsew
rlabel metal2 s 240 14220 240 14220 4 gnd
port 514 nsew
rlabel metal2 s 240 15247 240 15247 4 gnd
port 514 nsew
rlabel metal2 s 240 15010 240 15010 4 gnd
port 514 nsew
rlabel metal2 s 240 15800 240 15800 4 gnd
port 514 nsew
rlabel metal2 s 2256 15563 2256 15563 4 gnd
port 514 nsew
rlabel metal2 s 1008 13667 1008 13667 4 gnd
port 514 nsew
rlabel metal2 s 1008 15010 1008 15010 4 gnd
port 514 nsew
rlabel metal2 s 1488 14220 1488 14220 4 gnd
port 514 nsew
rlabel metal2 s 1008 15800 1008 15800 4 gnd
port 514 nsew
rlabel metal2 s 1008 14773 1008 14773 4 gnd
port 514 nsew
rlabel metal2 s 2256 13983 2256 13983 4 gnd
port 514 nsew
rlabel metal2 s 1488 14457 1488 14457 4 gnd
port 514 nsew
rlabel metal2 s 2256 15800 2256 15800 4 gnd
port 514 nsew
rlabel metal2 s 2256 15247 2256 15247 4 gnd
port 514 nsew
rlabel metal2 s 2256 14773 2256 14773 4 gnd
port 514 nsew
rlabel metal2 s 2256 13193 2256 13193 4 gnd
port 514 nsew
rlabel metal2 s 3984 13983 3984 13983 4 gnd
port 514 nsew
rlabel metal2 s 3984 14457 3984 14457 4 gnd
port 514 nsew
rlabel metal2 s 2736 15800 2736 15800 4 gnd
port 514 nsew
rlabel metal2 s 2736 15563 2736 15563 4 gnd
port 514 nsew
rlabel metal2 s 3504 15247 3504 15247 4 gnd
port 514 nsew
rlabel metal2 s 4752 13983 4752 13983 4 gnd
port 514 nsew
rlabel metal2 s 2736 13430 2736 13430 4 gnd
port 514 nsew
rlabel metal2 s 3984 15563 3984 15563 4 gnd
port 514 nsew
rlabel metal2 s 3504 13430 3504 13430 4 gnd
port 514 nsew
rlabel metal2 s 3504 12877 3504 12877 4 gnd
port 514 nsew
rlabel metal2 s 3504 15800 3504 15800 4 gnd
port 514 nsew
rlabel metal2 s 4752 14773 4752 14773 4 gnd
port 514 nsew
rlabel metal2 s 4752 15800 4752 15800 4 gnd
port 514 nsew
rlabel metal2 s 3984 14773 3984 14773 4 gnd
port 514 nsew
rlabel metal2 s 4752 15247 4752 15247 4 gnd
port 514 nsew
rlabel metal2 s 3504 14457 3504 14457 4 gnd
port 514 nsew
rlabel metal2 s 3504 15010 3504 15010 4 gnd
port 514 nsew
rlabel metal2 s 3984 13193 3984 13193 4 gnd
port 514 nsew
rlabel metal2 s 3504 13193 3504 13193 4 gnd
port 514 nsew
rlabel metal2 s 2736 15010 2736 15010 4 gnd
port 514 nsew
rlabel metal2 s 2736 14457 2736 14457 4 gnd
port 514 nsew
rlabel metal2 s 2736 13983 2736 13983 4 gnd
port 514 nsew
rlabel metal2 s 3984 15247 3984 15247 4 gnd
port 514 nsew
rlabel metal2 s 3984 12877 3984 12877 4 gnd
port 514 nsew
rlabel metal2 s 4752 15010 4752 15010 4 gnd
port 514 nsew
rlabel metal2 s 3504 13983 3504 13983 4 gnd
port 514 nsew
rlabel metal2 s 2736 14220 2736 14220 4 gnd
port 514 nsew
rlabel metal2 s 2736 13667 2736 13667 4 gnd
port 514 nsew
rlabel metal2 s 4752 13193 4752 13193 4 gnd
port 514 nsew
rlabel metal2 s 2736 14773 2736 14773 4 gnd
port 514 nsew
rlabel metal2 s 2736 13193 2736 13193 4 gnd
port 514 nsew
rlabel metal2 s 4752 14457 4752 14457 4 gnd
port 514 nsew
rlabel metal2 s 2736 15247 2736 15247 4 gnd
port 514 nsew
rlabel metal2 s 3984 13430 3984 13430 4 gnd
port 514 nsew
rlabel metal2 s 2736 12877 2736 12877 4 gnd
port 514 nsew
rlabel metal2 s 4752 15563 4752 15563 4 gnd
port 514 nsew
rlabel metal2 s 3504 13667 3504 13667 4 gnd
port 514 nsew
rlabel metal2 s 4752 13667 4752 13667 4 gnd
port 514 nsew
rlabel metal2 s 4752 13430 4752 13430 4 gnd
port 514 nsew
rlabel metal2 s 4752 14220 4752 14220 4 gnd
port 514 nsew
rlabel metal2 s 3504 14220 3504 14220 4 gnd
port 514 nsew
rlabel metal2 s 3984 13667 3984 13667 4 gnd
port 514 nsew
rlabel metal2 s 3984 15010 3984 15010 4 gnd
port 514 nsew
rlabel metal2 s 4752 12877 4752 12877 4 gnd
port 514 nsew
rlabel metal2 s 3504 14773 3504 14773 4 gnd
port 514 nsew
rlabel metal2 s 3984 15800 3984 15800 4 gnd
port 514 nsew
rlabel metal2 s 3984 14220 3984 14220 4 gnd
port 514 nsew
rlabel metal2 s 3504 15563 3504 15563 4 gnd
port 514 nsew
rlabel metal2 s 9744 17143 9744 17143 4 gnd
port 514 nsew
rlabel metal2 s 7728 17380 7728 17380 4 gnd
port 514 nsew
rlabel metal2 s 8976 17617 8976 17617 4 gnd
port 514 nsew
rlabel metal2 s 9744 17380 9744 17380 4 gnd
port 514 nsew
rlabel metal2 s 9744 16353 9744 16353 4 gnd
port 514 nsew
rlabel metal2 s 9744 18723 9744 18723 4 gnd
port 514 nsew
rlabel metal2 s 7728 18723 7728 18723 4 gnd
port 514 nsew
rlabel metal2 s 8976 18170 8976 18170 4 gnd
port 514 nsew
rlabel metal2 s 8496 18723 8496 18723 4 gnd
port 514 nsew
rlabel metal2 s 8976 18407 8976 18407 4 gnd
port 514 nsew
rlabel metal2 s 7728 16590 7728 16590 4 gnd
port 514 nsew
rlabel metal2 s 7728 16037 7728 16037 4 gnd
port 514 nsew
rlabel metal2 s 9744 18170 9744 18170 4 gnd
port 514 nsew
rlabel metal2 s 7728 18407 7728 18407 4 gnd
port 514 nsew
rlabel metal2 s 7728 18170 7728 18170 4 gnd
port 514 nsew
rlabel metal2 s 8976 18960 8976 18960 4 gnd
port 514 nsew
rlabel metal2 s 7728 17143 7728 17143 4 gnd
port 514 nsew
rlabel metal2 s 8976 17380 8976 17380 4 gnd
port 514 nsew
rlabel metal2 s 8496 17143 8496 17143 4 gnd
port 514 nsew
rlabel metal2 s 7728 18960 7728 18960 4 gnd
port 514 nsew
rlabel metal2 s 8976 17933 8976 17933 4 gnd
port 514 nsew
rlabel metal2 s 8496 16353 8496 16353 4 gnd
port 514 nsew
rlabel metal2 s 8496 17617 8496 17617 4 gnd
port 514 nsew
rlabel metal2 s 9744 17617 9744 17617 4 gnd
port 514 nsew
rlabel metal2 s 8496 16590 8496 16590 4 gnd
port 514 nsew
rlabel metal2 s 8496 18407 8496 18407 4 gnd
port 514 nsew
rlabel metal2 s 8976 16590 8976 16590 4 gnd
port 514 nsew
rlabel metal2 s 9744 16037 9744 16037 4 gnd
port 514 nsew
rlabel metal2 s 8976 16037 8976 16037 4 gnd
port 514 nsew
rlabel metal2 s 8496 17380 8496 17380 4 gnd
port 514 nsew
rlabel metal2 s 8496 18960 8496 18960 4 gnd
port 514 nsew
rlabel metal2 s 8976 16827 8976 16827 4 gnd
port 514 nsew
rlabel metal2 s 7728 16827 7728 16827 4 gnd
port 514 nsew
rlabel metal2 s 9744 16827 9744 16827 4 gnd
port 514 nsew
rlabel metal2 s 8976 16353 8976 16353 4 gnd
port 514 nsew
rlabel metal2 s 7728 17933 7728 17933 4 gnd
port 514 nsew
rlabel metal2 s 9744 18407 9744 18407 4 gnd
port 514 nsew
rlabel metal2 s 8496 16037 8496 16037 4 gnd
port 514 nsew
rlabel metal2 s 7728 17617 7728 17617 4 gnd
port 514 nsew
rlabel metal2 s 8496 16827 8496 16827 4 gnd
port 514 nsew
rlabel metal2 s 9744 18960 9744 18960 4 gnd
port 514 nsew
rlabel metal2 s 7728 16353 7728 16353 4 gnd
port 514 nsew
rlabel metal2 s 9744 16590 9744 16590 4 gnd
port 514 nsew
rlabel metal2 s 8496 17933 8496 17933 4 gnd
port 514 nsew
rlabel metal2 s 8976 18723 8976 18723 4 gnd
port 514 nsew
rlabel metal2 s 8976 17143 8976 17143 4 gnd
port 514 nsew
rlabel metal2 s 9744 17933 9744 17933 4 gnd
port 514 nsew
rlabel metal2 s 8496 18170 8496 18170 4 gnd
port 514 nsew
rlabel metal2 s 7248 18960 7248 18960 4 gnd
port 514 nsew
rlabel metal2 s 6000 17380 6000 17380 4 gnd
port 514 nsew
rlabel metal2 s 6000 18960 6000 18960 4 gnd
port 514 nsew
rlabel metal2 s 6480 17143 6480 17143 4 gnd
port 514 nsew
rlabel metal2 s 7248 16037 7248 16037 4 gnd
port 514 nsew
rlabel metal2 s 5232 16590 5232 16590 4 gnd
port 514 nsew
rlabel metal2 s 6480 16037 6480 16037 4 gnd
port 514 nsew
rlabel metal2 s 7248 18723 7248 18723 4 gnd
port 514 nsew
rlabel metal2 s 6480 17617 6480 17617 4 gnd
port 514 nsew
rlabel metal2 s 6480 17933 6480 17933 4 gnd
port 514 nsew
rlabel metal2 s 5232 16353 5232 16353 4 gnd
port 514 nsew
rlabel metal2 s 6000 16590 6000 16590 4 gnd
port 514 nsew
rlabel metal2 s 7248 18170 7248 18170 4 gnd
port 514 nsew
rlabel metal2 s 7248 16827 7248 16827 4 gnd
port 514 nsew
rlabel metal2 s 5232 17143 5232 17143 4 gnd
port 514 nsew
rlabel metal2 s 5232 18723 5232 18723 4 gnd
port 514 nsew
rlabel metal2 s 7248 18407 7248 18407 4 gnd
port 514 nsew
rlabel metal2 s 6000 16827 6000 16827 4 gnd
port 514 nsew
rlabel metal2 s 7248 17933 7248 17933 4 gnd
port 514 nsew
rlabel metal2 s 7248 17617 7248 17617 4 gnd
port 514 nsew
rlabel metal2 s 5232 16037 5232 16037 4 gnd
port 514 nsew
rlabel metal2 s 6000 16037 6000 16037 4 gnd
port 514 nsew
rlabel metal2 s 6480 16590 6480 16590 4 gnd
port 514 nsew
rlabel metal2 s 5232 18407 5232 18407 4 gnd
port 514 nsew
rlabel metal2 s 6480 16353 6480 16353 4 gnd
port 514 nsew
rlabel metal2 s 7248 17380 7248 17380 4 gnd
port 514 nsew
rlabel metal2 s 6480 18407 6480 18407 4 gnd
port 514 nsew
rlabel metal2 s 7248 17143 7248 17143 4 gnd
port 514 nsew
rlabel metal2 s 6480 16827 6480 16827 4 gnd
port 514 nsew
rlabel metal2 s 5232 17380 5232 17380 4 gnd
port 514 nsew
rlabel metal2 s 6480 18960 6480 18960 4 gnd
port 514 nsew
rlabel metal2 s 5232 18170 5232 18170 4 gnd
port 514 nsew
rlabel metal2 s 6480 17380 6480 17380 4 gnd
port 514 nsew
rlabel metal2 s 6000 18723 6000 18723 4 gnd
port 514 nsew
rlabel metal2 s 6000 17143 6000 17143 4 gnd
port 514 nsew
rlabel metal2 s 6000 16353 6000 16353 4 gnd
port 514 nsew
rlabel metal2 s 6000 18407 6000 18407 4 gnd
port 514 nsew
rlabel metal2 s 6480 18170 6480 18170 4 gnd
port 514 nsew
rlabel metal2 s 6480 18723 6480 18723 4 gnd
port 514 nsew
rlabel metal2 s 5232 16827 5232 16827 4 gnd
port 514 nsew
rlabel metal2 s 6000 18170 6000 18170 4 gnd
port 514 nsew
rlabel metal2 s 5232 18960 5232 18960 4 gnd
port 514 nsew
rlabel metal2 s 6000 17933 6000 17933 4 gnd
port 514 nsew
rlabel metal2 s 5232 17617 5232 17617 4 gnd
port 514 nsew
rlabel metal2 s 6000 17617 6000 17617 4 gnd
port 514 nsew
rlabel metal2 s 5232 17933 5232 17933 4 gnd
port 514 nsew
rlabel metal2 s 7248 16353 7248 16353 4 gnd
port 514 nsew
rlabel metal2 s 7248 16590 7248 16590 4 gnd
port 514 nsew
rlabel metal2 s 6000 14220 6000 14220 4 gnd
port 514 nsew
rlabel metal2 s 5232 15247 5232 15247 4 gnd
port 514 nsew
rlabel metal2 s 6000 13983 6000 13983 4 gnd
port 514 nsew
rlabel metal2 s 5232 13430 5232 13430 4 gnd
port 514 nsew
rlabel metal2 s 5232 14457 5232 14457 4 gnd
port 514 nsew
rlabel metal2 s 6000 13667 6000 13667 4 gnd
port 514 nsew
rlabel metal2 s 5232 12877 5232 12877 4 gnd
port 514 nsew
rlabel metal2 s 6000 13430 6000 13430 4 gnd
port 514 nsew
rlabel metal2 s 7248 13193 7248 13193 4 gnd
port 514 nsew
rlabel metal2 s 5232 13983 5232 13983 4 gnd
port 514 nsew
rlabel metal2 s 6480 13667 6480 13667 4 gnd
port 514 nsew
rlabel metal2 s 7248 14220 7248 14220 4 gnd
port 514 nsew
rlabel metal2 s 7248 14457 7248 14457 4 gnd
port 514 nsew
rlabel metal2 s 5232 13193 5232 13193 4 gnd
port 514 nsew
rlabel metal2 s 7248 14773 7248 14773 4 gnd
port 514 nsew
rlabel metal2 s 6480 15800 6480 15800 4 gnd
port 514 nsew
rlabel metal2 s 7248 13983 7248 13983 4 gnd
port 514 nsew
rlabel metal2 s 6000 15800 6000 15800 4 gnd
port 514 nsew
rlabel metal2 s 5232 14220 5232 14220 4 gnd
port 514 nsew
rlabel metal2 s 6480 13430 6480 13430 4 gnd
port 514 nsew
rlabel metal2 s 5232 13667 5232 13667 4 gnd
port 514 nsew
rlabel metal2 s 5232 14773 5232 14773 4 gnd
port 514 nsew
rlabel metal2 s 6480 14457 6480 14457 4 gnd
port 514 nsew
rlabel metal2 s 7248 12877 7248 12877 4 gnd
port 514 nsew
rlabel metal2 s 6480 15563 6480 15563 4 gnd
port 514 nsew
rlabel metal2 s 6480 13193 6480 13193 4 gnd
port 514 nsew
rlabel metal2 s 7248 15563 7248 15563 4 gnd
port 514 nsew
rlabel metal2 s 6480 14220 6480 14220 4 gnd
port 514 nsew
rlabel metal2 s 6000 12877 6000 12877 4 gnd
port 514 nsew
rlabel metal2 s 6480 15010 6480 15010 4 gnd
port 514 nsew
rlabel metal2 s 6000 15247 6000 15247 4 gnd
port 514 nsew
rlabel metal2 s 6000 14457 6000 14457 4 gnd
port 514 nsew
rlabel metal2 s 6000 13193 6000 13193 4 gnd
port 514 nsew
rlabel metal2 s 7248 15010 7248 15010 4 gnd
port 514 nsew
rlabel metal2 s 7248 15800 7248 15800 4 gnd
port 514 nsew
rlabel metal2 s 7248 15247 7248 15247 4 gnd
port 514 nsew
rlabel metal2 s 6000 15010 6000 15010 4 gnd
port 514 nsew
rlabel metal2 s 6480 13983 6480 13983 4 gnd
port 514 nsew
rlabel metal2 s 5232 15010 5232 15010 4 gnd
port 514 nsew
rlabel metal2 s 7248 13430 7248 13430 4 gnd
port 514 nsew
rlabel metal2 s 5232 15563 5232 15563 4 gnd
port 514 nsew
rlabel metal2 s 5232 15800 5232 15800 4 gnd
port 514 nsew
rlabel metal2 s 7248 13667 7248 13667 4 gnd
port 514 nsew
rlabel metal2 s 6000 15563 6000 15563 4 gnd
port 514 nsew
rlabel metal2 s 6000 14773 6000 14773 4 gnd
port 514 nsew
rlabel metal2 s 6480 15247 6480 15247 4 gnd
port 514 nsew
rlabel metal2 s 6480 12877 6480 12877 4 gnd
port 514 nsew
rlabel metal2 s 6480 14773 6480 14773 4 gnd
port 514 nsew
rlabel metal2 s 8496 12877 8496 12877 4 gnd
port 514 nsew
rlabel metal2 s 7728 12877 7728 12877 4 gnd
port 514 nsew
rlabel metal2 s 7728 14220 7728 14220 4 gnd
port 514 nsew
rlabel metal2 s 7728 13667 7728 13667 4 gnd
port 514 nsew
rlabel metal2 s 9744 13667 9744 13667 4 gnd
port 514 nsew
rlabel metal2 s 9744 12877 9744 12877 4 gnd
port 514 nsew
rlabel metal2 s 8496 13193 8496 13193 4 gnd
port 514 nsew
rlabel metal2 s 9744 14220 9744 14220 4 gnd
port 514 nsew
rlabel metal2 s 7728 14457 7728 14457 4 gnd
port 514 nsew
rlabel metal2 s 9744 15247 9744 15247 4 gnd
port 514 nsew
rlabel metal2 s 9744 13983 9744 13983 4 gnd
port 514 nsew
rlabel metal2 s 8976 13983 8976 13983 4 gnd
port 514 nsew
rlabel metal2 s 7728 13193 7728 13193 4 gnd
port 514 nsew
rlabel metal2 s 7728 14773 7728 14773 4 gnd
port 514 nsew
rlabel metal2 s 8976 14457 8976 14457 4 gnd
port 514 nsew
rlabel metal2 s 8976 14220 8976 14220 4 gnd
port 514 nsew
rlabel metal2 s 8976 13430 8976 13430 4 gnd
port 514 nsew
rlabel metal2 s 8976 13667 8976 13667 4 gnd
port 514 nsew
rlabel metal2 s 9744 13430 9744 13430 4 gnd
port 514 nsew
rlabel metal2 s 7728 15563 7728 15563 4 gnd
port 514 nsew
rlabel metal2 s 8496 15563 8496 15563 4 gnd
port 514 nsew
rlabel metal2 s 7728 15010 7728 15010 4 gnd
port 514 nsew
rlabel metal2 s 7728 15800 7728 15800 4 gnd
port 514 nsew
rlabel metal2 s 8496 14220 8496 14220 4 gnd
port 514 nsew
rlabel metal2 s 8496 13983 8496 13983 4 gnd
port 514 nsew
rlabel metal2 s 8496 14773 8496 14773 4 gnd
port 514 nsew
rlabel metal2 s 8976 14773 8976 14773 4 gnd
port 514 nsew
rlabel metal2 s 8976 15563 8976 15563 4 gnd
port 514 nsew
rlabel metal2 s 8496 15800 8496 15800 4 gnd
port 514 nsew
rlabel metal2 s 8976 12877 8976 12877 4 gnd
port 514 nsew
rlabel metal2 s 8496 13430 8496 13430 4 gnd
port 514 nsew
rlabel metal2 s 8496 15010 8496 15010 4 gnd
port 514 nsew
rlabel metal2 s 8496 14457 8496 14457 4 gnd
port 514 nsew
rlabel metal2 s 8496 13667 8496 13667 4 gnd
port 514 nsew
rlabel metal2 s 9744 14773 9744 14773 4 gnd
port 514 nsew
rlabel metal2 s 7728 15247 7728 15247 4 gnd
port 514 nsew
rlabel metal2 s 9744 14457 9744 14457 4 gnd
port 514 nsew
rlabel metal2 s 8976 15247 8976 15247 4 gnd
port 514 nsew
rlabel metal2 s 7728 13983 7728 13983 4 gnd
port 514 nsew
rlabel metal2 s 8976 15010 8976 15010 4 gnd
port 514 nsew
rlabel metal2 s 9744 13193 9744 13193 4 gnd
port 514 nsew
rlabel metal2 s 8976 15800 8976 15800 4 gnd
port 514 nsew
rlabel metal2 s 7728 13430 7728 13430 4 gnd
port 514 nsew
rlabel metal2 s 9744 15563 9744 15563 4 gnd
port 514 nsew
rlabel metal2 s 8976 13193 8976 13193 4 gnd
port 514 nsew
rlabel metal2 s 9744 15010 9744 15010 4 gnd
port 514 nsew
rlabel metal2 s 8496 15247 8496 15247 4 gnd
port 514 nsew
rlabel metal2 s 9744 15800 9744 15800 4 gnd
port 514 nsew
rlabel metal2 s 8976 10823 8976 10823 4 gnd
port 514 nsew
rlabel metal2 s 7728 12403 7728 12403 4 gnd
port 514 nsew
rlabel metal2 s 8496 12640 8496 12640 4 gnd
port 514 nsew
rlabel metal2 s 7728 10823 7728 10823 4 gnd
port 514 nsew
rlabel metal2 s 8976 11060 8976 11060 4 gnd
port 514 nsew
rlabel metal2 s 9744 10270 9744 10270 4 gnd
port 514 nsew
rlabel metal2 s 8496 10033 8496 10033 4 gnd
port 514 nsew
rlabel metal2 s 9744 11850 9744 11850 4 gnd
port 514 nsew
rlabel metal2 s 9744 12087 9744 12087 4 gnd
port 514 nsew
rlabel metal2 s 8976 10033 8976 10033 4 gnd
port 514 nsew
rlabel metal2 s 7728 11060 7728 11060 4 gnd
port 514 nsew
rlabel metal2 s 7728 11297 7728 11297 4 gnd
port 514 nsew
rlabel metal2 s 9744 12403 9744 12403 4 gnd
port 514 nsew
rlabel metal2 s 9744 11613 9744 11613 4 gnd
port 514 nsew
rlabel metal2 s 8976 11297 8976 11297 4 gnd
port 514 nsew
rlabel metal2 s 8496 11613 8496 11613 4 gnd
port 514 nsew
rlabel metal2 s 7728 11850 7728 11850 4 gnd
port 514 nsew
rlabel metal2 s 8976 10507 8976 10507 4 gnd
port 514 nsew
rlabel metal2 s 8496 12403 8496 12403 4 gnd
port 514 nsew
rlabel metal2 s 8976 11850 8976 11850 4 gnd
port 514 nsew
rlabel metal2 s 8496 10507 8496 10507 4 gnd
port 514 nsew
rlabel metal2 s 8496 11850 8496 11850 4 gnd
port 514 nsew
rlabel metal2 s 8976 12087 8976 12087 4 gnd
port 514 nsew
rlabel metal2 s 8976 9717 8976 9717 4 gnd
port 514 nsew
rlabel metal2 s 9744 9717 9744 9717 4 gnd
port 514 nsew
rlabel metal2 s 8496 10823 8496 10823 4 gnd
port 514 nsew
rlabel metal2 s 7728 12087 7728 12087 4 gnd
port 514 nsew
rlabel metal2 s 8496 9717 8496 9717 4 gnd
port 514 nsew
rlabel metal2 s 7728 11613 7728 11613 4 gnd
port 514 nsew
rlabel metal2 s 8976 11613 8976 11613 4 gnd
port 514 nsew
rlabel metal2 s 9744 11297 9744 11297 4 gnd
port 514 nsew
rlabel metal2 s 9744 12640 9744 12640 4 gnd
port 514 nsew
rlabel metal2 s 8976 12640 8976 12640 4 gnd
port 514 nsew
rlabel metal2 s 8496 10270 8496 10270 4 gnd
port 514 nsew
rlabel metal2 s 7728 10033 7728 10033 4 gnd
port 514 nsew
rlabel metal2 s 9744 10507 9744 10507 4 gnd
port 514 nsew
rlabel metal2 s 7728 9717 7728 9717 4 gnd
port 514 nsew
rlabel metal2 s 9744 11060 9744 11060 4 gnd
port 514 nsew
rlabel metal2 s 8496 11297 8496 11297 4 gnd
port 514 nsew
rlabel metal2 s 9744 10033 9744 10033 4 gnd
port 514 nsew
rlabel metal2 s 8496 11060 8496 11060 4 gnd
port 514 nsew
rlabel metal2 s 8496 12087 8496 12087 4 gnd
port 514 nsew
rlabel metal2 s 8976 10270 8976 10270 4 gnd
port 514 nsew
rlabel metal2 s 9744 10823 9744 10823 4 gnd
port 514 nsew
rlabel metal2 s 7728 10507 7728 10507 4 gnd
port 514 nsew
rlabel metal2 s 8976 12403 8976 12403 4 gnd
port 514 nsew
rlabel metal2 s 7728 10270 7728 10270 4 gnd
port 514 nsew
rlabel metal2 s 7728 12640 7728 12640 4 gnd
port 514 nsew
rlabel metal2 s 6480 12087 6480 12087 4 gnd
port 514 nsew
rlabel metal2 s 6000 10033 6000 10033 4 gnd
port 514 nsew
rlabel metal2 s 5232 10507 5232 10507 4 gnd
port 514 nsew
rlabel metal2 s 5232 10270 5232 10270 4 gnd
port 514 nsew
rlabel metal2 s 7248 12640 7248 12640 4 gnd
port 514 nsew
rlabel metal2 s 6000 10823 6000 10823 4 gnd
port 514 nsew
rlabel metal2 s 7248 10270 7248 10270 4 gnd
port 514 nsew
rlabel metal2 s 5232 10033 5232 10033 4 gnd
port 514 nsew
rlabel metal2 s 5232 11297 5232 11297 4 gnd
port 514 nsew
rlabel metal2 s 7248 11060 7248 11060 4 gnd
port 514 nsew
rlabel metal2 s 5232 12403 5232 12403 4 gnd
port 514 nsew
rlabel metal2 s 6000 11297 6000 11297 4 gnd
port 514 nsew
rlabel metal2 s 6480 11060 6480 11060 4 gnd
port 514 nsew
rlabel metal2 s 6480 12640 6480 12640 4 gnd
port 514 nsew
rlabel metal2 s 6480 10270 6480 10270 4 gnd
port 514 nsew
rlabel metal2 s 7248 11850 7248 11850 4 gnd
port 514 nsew
rlabel metal2 s 7248 11613 7248 11613 4 gnd
port 514 nsew
rlabel metal2 s 5232 12087 5232 12087 4 gnd
port 514 nsew
rlabel metal2 s 6000 9717 6000 9717 4 gnd
port 514 nsew
rlabel metal2 s 7248 12087 7248 12087 4 gnd
port 514 nsew
rlabel metal2 s 7248 11297 7248 11297 4 gnd
port 514 nsew
rlabel metal2 s 6000 12640 6000 12640 4 gnd
port 514 nsew
rlabel metal2 s 6000 10507 6000 10507 4 gnd
port 514 nsew
rlabel metal2 s 6480 11297 6480 11297 4 gnd
port 514 nsew
rlabel metal2 s 5232 11850 5232 11850 4 gnd
port 514 nsew
rlabel metal2 s 5232 9717 5232 9717 4 gnd
port 514 nsew
rlabel metal2 s 5232 11613 5232 11613 4 gnd
port 514 nsew
rlabel metal2 s 7248 12403 7248 12403 4 gnd
port 514 nsew
rlabel metal2 s 7248 10823 7248 10823 4 gnd
port 514 nsew
rlabel metal2 s 6480 10823 6480 10823 4 gnd
port 514 nsew
rlabel metal2 s 6480 12403 6480 12403 4 gnd
port 514 nsew
rlabel metal2 s 6000 11060 6000 11060 4 gnd
port 514 nsew
rlabel metal2 s 6480 10033 6480 10033 4 gnd
port 514 nsew
rlabel metal2 s 6000 12087 6000 12087 4 gnd
port 514 nsew
rlabel metal2 s 6480 10507 6480 10507 4 gnd
port 514 nsew
rlabel metal2 s 6000 11613 6000 11613 4 gnd
port 514 nsew
rlabel metal2 s 5232 10823 5232 10823 4 gnd
port 514 nsew
rlabel metal2 s 6480 11613 6480 11613 4 gnd
port 514 nsew
rlabel metal2 s 5232 11060 5232 11060 4 gnd
port 514 nsew
rlabel metal2 s 6480 11850 6480 11850 4 gnd
port 514 nsew
rlabel metal2 s 5232 12640 5232 12640 4 gnd
port 514 nsew
rlabel metal2 s 6000 10270 6000 10270 4 gnd
port 514 nsew
rlabel metal2 s 6000 12403 6000 12403 4 gnd
port 514 nsew
rlabel metal2 s 7248 10033 7248 10033 4 gnd
port 514 nsew
rlabel metal2 s 6480 9717 6480 9717 4 gnd
port 514 nsew
rlabel metal2 s 6000 11850 6000 11850 4 gnd
port 514 nsew
rlabel metal2 s 7248 9717 7248 9717 4 gnd
port 514 nsew
rlabel metal2 s 7248 10507 7248 10507 4 gnd
port 514 nsew
rlabel metal2 s 7248 7110 7248 7110 4 gnd
port 514 nsew
rlabel metal2 s 5232 8453 5232 8453 4 gnd
port 514 nsew
rlabel metal2 s 6480 8690 6480 8690 4 gnd
port 514 nsew
rlabel metal2 s 7248 8690 7248 8690 4 gnd
port 514 nsew
rlabel metal2 s 5232 7347 5232 7347 4 gnd
port 514 nsew
rlabel metal2 s 6480 7347 6480 7347 4 gnd
port 514 nsew
rlabel metal2 s 7248 7663 7248 7663 4 gnd
port 514 nsew
rlabel metal2 s 5232 6873 5232 6873 4 gnd
port 514 nsew
rlabel metal2 s 6480 7663 6480 7663 4 gnd
port 514 nsew
rlabel metal2 s 6000 8690 6000 8690 4 gnd
port 514 nsew
rlabel metal2 s 7248 9480 7248 9480 4 gnd
port 514 nsew
rlabel metal2 s 6000 7900 6000 7900 4 gnd
port 514 nsew
rlabel metal2 s 6000 7347 6000 7347 4 gnd
port 514 nsew
rlabel metal2 s 7248 7347 7248 7347 4 gnd
port 514 nsew
rlabel metal2 s 5232 9480 5232 9480 4 gnd
port 514 nsew
rlabel metal2 s 5232 8927 5232 8927 4 gnd
port 514 nsew
rlabel metal2 s 6480 6873 6480 6873 4 gnd
port 514 nsew
rlabel metal2 s 6480 9243 6480 9243 4 gnd
port 514 nsew
rlabel metal2 s 7248 9243 7248 9243 4 gnd
port 514 nsew
rlabel metal2 s 5232 6557 5232 6557 4 gnd
port 514 nsew
rlabel metal2 s 6000 6557 6000 6557 4 gnd
port 514 nsew
rlabel metal2 s 6000 7663 6000 7663 4 gnd
port 514 nsew
rlabel metal2 s 6480 9480 6480 9480 4 gnd
port 514 nsew
rlabel metal2 s 5232 8690 5232 8690 4 gnd
port 514 nsew
rlabel metal2 s 7248 6557 7248 6557 4 gnd
port 514 nsew
rlabel metal2 s 6000 9480 6000 9480 4 gnd
port 514 nsew
rlabel metal2 s 5232 7663 5232 7663 4 gnd
port 514 nsew
rlabel metal2 s 6000 9243 6000 9243 4 gnd
port 514 nsew
rlabel metal2 s 5232 7110 5232 7110 4 gnd
port 514 nsew
rlabel metal2 s 6000 7110 6000 7110 4 gnd
port 514 nsew
rlabel metal2 s 7248 7900 7248 7900 4 gnd
port 514 nsew
rlabel metal2 s 7248 8453 7248 8453 4 gnd
port 514 nsew
rlabel metal2 s 7248 8927 7248 8927 4 gnd
port 514 nsew
rlabel metal2 s 6480 7900 6480 7900 4 gnd
port 514 nsew
rlabel metal2 s 6000 8137 6000 8137 4 gnd
port 514 nsew
rlabel metal2 s 7248 8137 7248 8137 4 gnd
port 514 nsew
rlabel metal2 s 6480 8453 6480 8453 4 gnd
port 514 nsew
rlabel metal2 s 6000 8927 6000 8927 4 gnd
port 514 nsew
rlabel metal2 s 6480 7110 6480 7110 4 gnd
port 514 nsew
rlabel metal2 s 5232 9243 5232 9243 4 gnd
port 514 nsew
rlabel metal2 s 5232 7900 5232 7900 4 gnd
port 514 nsew
rlabel metal2 s 5232 8137 5232 8137 4 gnd
port 514 nsew
rlabel metal2 s 6000 6873 6000 6873 4 gnd
port 514 nsew
rlabel metal2 s 6480 8137 6480 8137 4 gnd
port 514 nsew
rlabel metal2 s 7248 6873 7248 6873 4 gnd
port 514 nsew
rlabel metal2 s 6000 8453 6000 8453 4 gnd
port 514 nsew
rlabel metal2 s 6480 6557 6480 6557 4 gnd
port 514 nsew
rlabel metal2 s 6480 8927 6480 8927 4 gnd
port 514 nsew
rlabel metal2 s 8976 6557 8976 6557 4 gnd
port 514 nsew
rlabel metal2 s 8976 8137 8976 8137 4 gnd
port 514 nsew
rlabel metal2 s 8496 6873 8496 6873 4 gnd
port 514 nsew
rlabel metal2 s 8976 9243 8976 9243 4 gnd
port 514 nsew
rlabel metal2 s 8976 8453 8976 8453 4 gnd
port 514 nsew
rlabel metal2 s 8976 7663 8976 7663 4 gnd
port 514 nsew
rlabel metal2 s 9744 9243 9744 9243 4 gnd
port 514 nsew
rlabel metal2 s 8976 7110 8976 7110 4 gnd
port 514 nsew
rlabel metal2 s 8496 7663 8496 7663 4 gnd
port 514 nsew
rlabel metal2 s 9744 8927 9744 8927 4 gnd
port 514 nsew
rlabel metal2 s 7728 8690 7728 8690 4 gnd
port 514 nsew
rlabel metal2 s 7728 8927 7728 8927 4 gnd
port 514 nsew
rlabel metal2 s 7728 9480 7728 9480 4 gnd
port 514 nsew
rlabel metal2 s 7728 8453 7728 8453 4 gnd
port 514 nsew
rlabel metal2 s 9744 8137 9744 8137 4 gnd
port 514 nsew
rlabel metal2 s 8976 7900 8976 7900 4 gnd
port 514 nsew
rlabel metal2 s 8976 7347 8976 7347 4 gnd
port 514 nsew
rlabel metal2 s 7728 9243 7728 9243 4 gnd
port 514 nsew
rlabel metal2 s 8496 8137 8496 8137 4 gnd
port 514 nsew
rlabel metal2 s 8496 8927 8496 8927 4 gnd
port 514 nsew
rlabel metal2 s 8976 6873 8976 6873 4 gnd
port 514 nsew
rlabel metal2 s 9744 7110 9744 7110 4 gnd
port 514 nsew
rlabel metal2 s 9744 7900 9744 7900 4 gnd
port 514 nsew
rlabel metal2 s 9744 6873 9744 6873 4 gnd
port 514 nsew
rlabel metal2 s 7728 7663 7728 7663 4 gnd
port 514 nsew
rlabel metal2 s 8496 8690 8496 8690 4 gnd
port 514 nsew
rlabel metal2 s 9744 7663 9744 7663 4 gnd
port 514 nsew
rlabel metal2 s 9744 8453 9744 8453 4 gnd
port 514 nsew
rlabel metal2 s 8496 6557 8496 6557 4 gnd
port 514 nsew
rlabel metal2 s 9744 8690 9744 8690 4 gnd
port 514 nsew
rlabel metal2 s 8496 7900 8496 7900 4 gnd
port 514 nsew
rlabel metal2 s 8496 9480 8496 9480 4 gnd
port 514 nsew
rlabel metal2 s 7728 6873 7728 6873 4 gnd
port 514 nsew
rlabel metal2 s 9744 9480 9744 9480 4 gnd
port 514 nsew
rlabel metal2 s 9744 7347 9744 7347 4 gnd
port 514 nsew
rlabel metal2 s 8496 7347 8496 7347 4 gnd
port 514 nsew
rlabel metal2 s 8496 7110 8496 7110 4 gnd
port 514 nsew
rlabel metal2 s 7728 8137 7728 8137 4 gnd
port 514 nsew
rlabel metal2 s 7728 7900 7728 7900 4 gnd
port 514 nsew
rlabel metal2 s 7728 7347 7728 7347 4 gnd
port 514 nsew
rlabel metal2 s 8496 9243 8496 9243 4 gnd
port 514 nsew
rlabel metal2 s 8496 8453 8496 8453 4 gnd
port 514 nsew
rlabel metal2 s 8976 8927 8976 8927 4 gnd
port 514 nsew
rlabel metal2 s 9744 6557 9744 6557 4 gnd
port 514 nsew
rlabel metal2 s 7728 6557 7728 6557 4 gnd
port 514 nsew
rlabel metal2 s 8976 9480 8976 9480 4 gnd
port 514 nsew
rlabel metal2 s 8976 8690 8976 8690 4 gnd
port 514 nsew
rlabel metal2 s 7728 7110 7728 7110 4 gnd
port 514 nsew
rlabel metal2 s 4752 10823 4752 10823 4 gnd
port 514 nsew
rlabel metal2 s 4752 10033 4752 10033 4 gnd
port 514 nsew
rlabel metal2 s 3504 11850 3504 11850 4 gnd
port 514 nsew
rlabel metal2 s 4752 11297 4752 11297 4 gnd
port 514 nsew
rlabel metal2 s 4752 12087 4752 12087 4 gnd
port 514 nsew
rlabel metal2 s 3504 12640 3504 12640 4 gnd
port 514 nsew
rlabel metal2 s 3984 11060 3984 11060 4 gnd
port 514 nsew
rlabel metal2 s 3984 12403 3984 12403 4 gnd
port 514 nsew
rlabel metal2 s 2736 10507 2736 10507 4 gnd
port 514 nsew
rlabel metal2 s 2736 11060 2736 11060 4 gnd
port 514 nsew
rlabel metal2 s 3504 11060 3504 11060 4 gnd
port 514 nsew
rlabel metal2 s 4752 11613 4752 11613 4 gnd
port 514 nsew
rlabel metal2 s 2736 11850 2736 11850 4 gnd
port 514 nsew
rlabel metal2 s 4752 11060 4752 11060 4 gnd
port 514 nsew
rlabel metal2 s 2736 10823 2736 10823 4 gnd
port 514 nsew
rlabel metal2 s 3504 10270 3504 10270 4 gnd
port 514 nsew
rlabel metal2 s 3984 12087 3984 12087 4 gnd
port 514 nsew
rlabel metal2 s 3504 10033 3504 10033 4 gnd
port 514 nsew
rlabel metal2 s 3984 11850 3984 11850 4 gnd
port 514 nsew
rlabel metal2 s 4752 11850 4752 11850 4 gnd
port 514 nsew
rlabel metal2 s 2736 12640 2736 12640 4 gnd
port 514 nsew
rlabel metal2 s 2736 10270 2736 10270 4 gnd
port 514 nsew
rlabel metal2 s 2736 11297 2736 11297 4 gnd
port 514 nsew
rlabel metal2 s 2736 9717 2736 9717 4 gnd
port 514 nsew
rlabel metal2 s 4752 12403 4752 12403 4 gnd
port 514 nsew
rlabel metal2 s 3984 10507 3984 10507 4 gnd
port 514 nsew
rlabel metal2 s 3504 9717 3504 9717 4 gnd
port 514 nsew
rlabel metal2 s 3984 11297 3984 11297 4 gnd
port 514 nsew
rlabel metal2 s 2736 11613 2736 11613 4 gnd
port 514 nsew
rlabel metal2 s 4752 9717 4752 9717 4 gnd
port 514 nsew
rlabel metal2 s 4752 10507 4752 10507 4 gnd
port 514 nsew
rlabel metal2 s 3984 9717 3984 9717 4 gnd
port 514 nsew
rlabel metal2 s 3504 11613 3504 11613 4 gnd
port 514 nsew
rlabel metal2 s 2736 12087 2736 12087 4 gnd
port 514 nsew
rlabel metal2 s 3504 10823 3504 10823 4 gnd
port 514 nsew
rlabel metal2 s 2736 10033 2736 10033 4 gnd
port 514 nsew
rlabel metal2 s 3984 10823 3984 10823 4 gnd
port 514 nsew
rlabel metal2 s 3984 12640 3984 12640 4 gnd
port 514 nsew
rlabel metal2 s 3984 11613 3984 11613 4 gnd
port 514 nsew
rlabel metal2 s 3504 12087 3504 12087 4 gnd
port 514 nsew
rlabel metal2 s 3984 10033 3984 10033 4 gnd
port 514 nsew
rlabel metal2 s 3504 11297 3504 11297 4 gnd
port 514 nsew
rlabel metal2 s 3504 12403 3504 12403 4 gnd
port 514 nsew
rlabel metal2 s 4752 10270 4752 10270 4 gnd
port 514 nsew
rlabel metal2 s 3984 10270 3984 10270 4 gnd
port 514 nsew
rlabel metal2 s 4752 12640 4752 12640 4 gnd
port 514 nsew
rlabel metal2 s 2736 12403 2736 12403 4 gnd
port 514 nsew
rlabel metal2 s 3504 10507 3504 10507 4 gnd
port 514 nsew
rlabel metal2 s 240 12640 240 12640 4 gnd
port 514 nsew
rlabel metal2 s 2256 11060 2256 11060 4 gnd
port 514 nsew
rlabel metal2 s 1488 12087 1488 12087 4 gnd
port 514 nsew
rlabel metal2 s 1488 12640 1488 12640 4 gnd
port 514 nsew
rlabel metal2 s 1488 11613 1488 11613 4 gnd
port 514 nsew
rlabel metal2 s 1488 12403 1488 12403 4 gnd
port 514 nsew
rlabel metal2 s 240 12403 240 12403 4 gnd
port 514 nsew
rlabel metal2 s 2256 10033 2256 10033 4 gnd
port 514 nsew
rlabel metal2 s 1488 10033 1488 10033 4 gnd
port 514 nsew
rlabel metal2 s 240 11060 240 11060 4 gnd
port 514 nsew
rlabel metal2 s 240 12087 240 12087 4 gnd
port 514 nsew
rlabel metal2 s 2256 12087 2256 12087 4 gnd
port 514 nsew
rlabel metal2 s 1488 11060 1488 11060 4 gnd
port 514 nsew
rlabel metal2 s 2256 11850 2256 11850 4 gnd
port 514 nsew
rlabel metal2 s 2256 10823 2256 10823 4 gnd
port 514 nsew
rlabel metal2 s 240 10823 240 10823 4 gnd
port 514 nsew
rlabel metal2 s 1488 11297 1488 11297 4 gnd
port 514 nsew
rlabel metal2 s 2256 11297 2256 11297 4 gnd
port 514 nsew
rlabel metal2 s 2256 11613 2256 11613 4 gnd
port 514 nsew
rlabel metal2 s 1008 12403 1008 12403 4 gnd
port 514 nsew
rlabel metal2 s 240 10270 240 10270 4 gnd
port 514 nsew
rlabel metal2 s 240 11297 240 11297 4 gnd
port 514 nsew
rlabel metal2 s 1008 10823 1008 10823 4 gnd
port 514 nsew
rlabel metal2 s 1008 12640 1008 12640 4 gnd
port 514 nsew
rlabel metal2 s 1008 11850 1008 11850 4 gnd
port 514 nsew
rlabel metal2 s 2256 12640 2256 12640 4 gnd
port 514 nsew
rlabel metal2 s 1008 11297 1008 11297 4 gnd
port 514 nsew
rlabel metal2 s 1008 10507 1008 10507 4 gnd
port 514 nsew
rlabel metal2 s 240 10507 240 10507 4 gnd
port 514 nsew
rlabel metal2 s 2256 10507 2256 10507 4 gnd
port 514 nsew
rlabel metal2 s 1008 9717 1008 9717 4 gnd
port 514 nsew
rlabel metal2 s 1008 10033 1008 10033 4 gnd
port 514 nsew
rlabel metal2 s 1488 10270 1488 10270 4 gnd
port 514 nsew
rlabel metal2 s 1008 11613 1008 11613 4 gnd
port 514 nsew
rlabel metal2 s 2256 9717 2256 9717 4 gnd
port 514 nsew
rlabel metal2 s 240 11850 240 11850 4 gnd
port 514 nsew
rlabel metal2 s 240 11613 240 11613 4 gnd
port 514 nsew
rlabel metal2 s 240 9717 240 9717 4 gnd
port 514 nsew
rlabel metal2 s 1488 11850 1488 11850 4 gnd
port 514 nsew
rlabel metal2 s 2256 12403 2256 12403 4 gnd
port 514 nsew
rlabel metal2 s 1488 10507 1488 10507 4 gnd
port 514 nsew
rlabel metal2 s 240 10033 240 10033 4 gnd
port 514 nsew
rlabel metal2 s 1008 12087 1008 12087 4 gnd
port 514 nsew
rlabel metal2 s 1008 11060 1008 11060 4 gnd
port 514 nsew
rlabel metal2 s 2256 10270 2256 10270 4 gnd
port 514 nsew
rlabel metal2 s 1488 10823 1488 10823 4 gnd
port 514 nsew
rlabel metal2 s 1008 10270 1008 10270 4 gnd
port 514 nsew
rlabel metal2 s 1488 9717 1488 9717 4 gnd
port 514 nsew
rlabel metal2 s 2256 7900 2256 7900 4 gnd
port 514 nsew
rlabel metal2 s 1008 6557 1008 6557 4 gnd
port 514 nsew
rlabel metal2 s 240 8927 240 8927 4 gnd
port 514 nsew
rlabel metal2 s 1488 9243 1488 9243 4 gnd
port 514 nsew
rlabel metal2 s 2256 6557 2256 6557 4 gnd
port 514 nsew
rlabel metal2 s 1008 7347 1008 7347 4 gnd
port 514 nsew
rlabel metal2 s 1008 7663 1008 7663 4 gnd
port 514 nsew
rlabel metal2 s 240 6873 240 6873 4 gnd
port 514 nsew
rlabel metal2 s 1008 8453 1008 8453 4 gnd
port 514 nsew
rlabel metal2 s 1488 7110 1488 7110 4 gnd
port 514 nsew
rlabel metal2 s 1488 8137 1488 8137 4 gnd
port 514 nsew
rlabel metal2 s 1488 7347 1488 7347 4 gnd
port 514 nsew
rlabel metal2 s 1008 9480 1008 9480 4 gnd
port 514 nsew
rlabel metal2 s 1488 6557 1488 6557 4 gnd
port 514 nsew
rlabel metal2 s 240 6557 240 6557 4 gnd
port 514 nsew
rlabel metal2 s 240 7347 240 7347 4 gnd
port 514 nsew
rlabel metal2 s 2256 8137 2256 8137 4 gnd
port 514 nsew
rlabel metal2 s 2256 9243 2256 9243 4 gnd
port 514 nsew
rlabel metal2 s 1008 7110 1008 7110 4 gnd
port 514 nsew
rlabel metal2 s 1008 8927 1008 8927 4 gnd
port 514 nsew
rlabel metal2 s 1488 7663 1488 7663 4 gnd
port 514 nsew
rlabel metal2 s 1008 8137 1008 8137 4 gnd
port 514 nsew
rlabel metal2 s 240 8453 240 8453 4 gnd
port 514 nsew
rlabel metal2 s 1488 6873 1488 6873 4 gnd
port 514 nsew
rlabel metal2 s 2256 8690 2256 8690 4 gnd
port 514 nsew
rlabel metal2 s 240 7110 240 7110 4 gnd
port 514 nsew
rlabel metal2 s 1488 9480 1488 9480 4 gnd
port 514 nsew
rlabel metal2 s 1008 8690 1008 8690 4 gnd
port 514 nsew
rlabel metal2 s 1488 8690 1488 8690 4 gnd
port 514 nsew
rlabel metal2 s 1008 9243 1008 9243 4 gnd
port 514 nsew
rlabel metal2 s 1488 8453 1488 8453 4 gnd
port 514 nsew
rlabel metal2 s 2256 8927 2256 8927 4 gnd
port 514 nsew
rlabel metal2 s 2256 7347 2256 7347 4 gnd
port 514 nsew
rlabel metal2 s 240 9243 240 9243 4 gnd
port 514 nsew
rlabel metal2 s 1488 8927 1488 8927 4 gnd
port 514 nsew
rlabel metal2 s 2256 8453 2256 8453 4 gnd
port 514 nsew
rlabel metal2 s 2256 9480 2256 9480 4 gnd
port 514 nsew
rlabel metal2 s 2256 7110 2256 7110 4 gnd
port 514 nsew
rlabel metal2 s 2256 6873 2256 6873 4 gnd
port 514 nsew
rlabel metal2 s 240 8690 240 8690 4 gnd
port 514 nsew
rlabel metal2 s 240 7663 240 7663 4 gnd
port 514 nsew
rlabel metal2 s 2256 7663 2256 7663 4 gnd
port 514 nsew
rlabel metal2 s 240 7900 240 7900 4 gnd
port 514 nsew
rlabel metal2 s 240 9480 240 9480 4 gnd
port 514 nsew
rlabel metal2 s 240 8137 240 8137 4 gnd
port 514 nsew
rlabel metal2 s 1008 7900 1008 7900 4 gnd
port 514 nsew
rlabel metal2 s 1488 7900 1488 7900 4 gnd
port 514 nsew
rlabel metal2 s 1008 6873 1008 6873 4 gnd
port 514 nsew
rlabel metal2 s 3984 9243 3984 9243 4 gnd
port 514 nsew
rlabel metal2 s 2736 6557 2736 6557 4 gnd
port 514 nsew
rlabel metal2 s 2736 7900 2736 7900 4 gnd
port 514 nsew
rlabel metal2 s 3984 6557 3984 6557 4 gnd
port 514 nsew
rlabel metal2 s 3504 7347 3504 7347 4 gnd
port 514 nsew
rlabel metal2 s 3504 7110 3504 7110 4 gnd
port 514 nsew
rlabel metal2 s 3984 6873 3984 6873 4 gnd
port 514 nsew
rlabel metal2 s 2736 6873 2736 6873 4 gnd
port 514 nsew
rlabel metal2 s 4752 8690 4752 8690 4 gnd
port 514 nsew
rlabel metal2 s 2736 7110 2736 7110 4 gnd
port 514 nsew
rlabel metal2 s 4752 8927 4752 8927 4 gnd
port 514 nsew
rlabel metal2 s 4752 7663 4752 7663 4 gnd
port 514 nsew
rlabel metal2 s 3504 7663 3504 7663 4 gnd
port 514 nsew
rlabel metal2 s 2736 9243 2736 9243 4 gnd
port 514 nsew
rlabel metal2 s 3504 8927 3504 8927 4 gnd
port 514 nsew
rlabel metal2 s 3504 8453 3504 8453 4 gnd
port 514 nsew
rlabel metal2 s 3504 8690 3504 8690 4 gnd
port 514 nsew
rlabel metal2 s 3504 9243 3504 9243 4 gnd
port 514 nsew
rlabel metal2 s 3984 7347 3984 7347 4 gnd
port 514 nsew
rlabel metal2 s 3984 9480 3984 9480 4 gnd
port 514 nsew
rlabel metal2 s 3984 8453 3984 8453 4 gnd
port 514 nsew
rlabel metal2 s 4752 7347 4752 7347 4 gnd
port 514 nsew
rlabel metal2 s 2736 7663 2736 7663 4 gnd
port 514 nsew
rlabel metal2 s 4752 7110 4752 7110 4 gnd
port 514 nsew
rlabel metal2 s 3984 8927 3984 8927 4 gnd
port 514 nsew
rlabel metal2 s 3504 7900 3504 7900 4 gnd
port 514 nsew
rlabel metal2 s 2736 8927 2736 8927 4 gnd
port 514 nsew
rlabel metal2 s 4752 7900 4752 7900 4 gnd
port 514 nsew
rlabel metal2 s 3984 7900 3984 7900 4 gnd
port 514 nsew
rlabel metal2 s 2736 9480 2736 9480 4 gnd
port 514 nsew
rlabel metal2 s 4752 9480 4752 9480 4 gnd
port 514 nsew
rlabel metal2 s 4752 6557 4752 6557 4 gnd
port 514 nsew
rlabel metal2 s 2736 7347 2736 7347 4 gnd
port 514 nsew
rlabel metal2 s 4752 6873 4752 6873 4 gnd
port 514 nsew
rlabel metal2 s 3984 7110 3984 7110 4 gnd
port 514 nsew
rlabel metal2 s 3504 6557 3504 6557 4 gnd
port 514 nsew
rlabel metal2 s 4752 9243 4752 9243 4 gnd
port 514 nsew
rlabel metal2 s 3984 8137 3984 8137 4 gnd
port 514 nsew
rlabel metal2 s 4752 8137 4752 8137 4 gnd
port 514 nsew
rlabel metal2 s 3984 8690 3984 8690 4 gnd
port 514 nsew
rlabel metal2 s 2736 8137 2736 8137 4 gnd
port 514 nsew
rlabel metal2 s 2736 8690 2736 8690 4 gnd
port 514 nsew
rlabel metal2 s 4752 8453 4752 8453 4 gnd
port 514 nsew
rlabel metal2 s 3504 8137 3504 8137 4 gnd
port 514 nsew
rlabel metal2 s 3504 9480 3504 9480 4 gnd
port 514 nsew
rlabel metal2 s 3504 6873 3504 6873 4 gnd
port 514 nsew
rlabel metal2 s 2736 8453 2736 8453 4 gnd
port 514 nsew
rlabel metal2 s 3984 7663 3984 7663 4 gnd
port 514 nsew
rlabel metal2 s 2736 3950 2736 3950 4 gnd
port 514 nsew
rlabel metal2 s 4752 3713 4752 3713 4 gnd
port 514 nsew
rlabel metal2 s 3504 3713 3504 3713 4 gnd
port 514 nsew
rlabel metal2 s 4752 4503 4752 4503 4 gnd
port 514 nsew
rlabel metal2 s 3984 4187 3984 4187 4 gnd
port 514 nsew
rlabel metal2 s 4752 3397 4752 3397 4 gnd
port 514 nsew
rlabel metal2 s 3984 5530 3984 5530 4 gnd
port 514 nsew
rlabel metal2 s 3504 4977 3504 4977 4 gnd
port 514 nsew
rlabel metal2 s 4752 4187 4752 4187 4 gnd
port 514 nsew
rlabel metal2 s 3504 5767 3504 5767 4 gnd
port 514 nsew
rlabel metal2 s 4752 6083 4752 6083 4 gnd
port 514 nsew
rlabel metal2 s 2736 5293 2736 5293 4 gnd
port 514 nsew
rlabel metal2 s 2736 4977 2736 4977 4 gnd
port 514 nsew
rlabel metal2 s 4752 5530 4752 5530 4 gnd
port 514 nsew
rlabel metal2 s 4752 5293 4752 5293 4 gnd
port 514 nsew
rlabel metal2 s 3984 3950 3984 3950 4 gnd
port 514 nsew
rlabel metal2 s 2736 4187 2736 4187 4 gnd
port 514 nsew
rlabel metal2 s 2736 3397 2736 3397 4 gnd
port 514 nsew
rlabel metal2 s 2736 4503 2736 4503 4 gnd
port 514 nsew
rlabel metal2 s 4752 6320 4752 6320 4 gnd
port 514 nsew
rlabel metal2 s 3504 4503 3504 4503 4 gnd
port 514 nsew
rlabel metal2 s 3984 4503 3984 4503 4 gnd
port 514 nsew
rlabel metal2 s 3504 4740 3504 4740 4 gnd
port 514 nsew
rlabel metal2 s 2736 5767 2736 5767 4 gnd
port 514 nsew
rlabel metal2 s 3984 5293 3984 5293 4 gnd
port 514 nsew
rlabel metal2 s 2736 5530 2736 5530 4 gnd
port 514 nsew
rlabel metal2 s 2736 6083 2736 6083 4 gnd
port 514 nsew
rlabel metal2 s 2736 6320 2736 6320 4 gnd
port 514 nsew
rlabel metal2 s 3984 4977 3984 4977 4 gnd
port 514 nsew
rlabel metal2 s 4752 4740 4752 4740 4 gnd
port 514 nsew
rlabel metal2 s 3504 4187 3504 4187 4 gnd
port 514 nsew
rlabel metal2 s 3984 3713 3984 3713 4 gnd
port 514 nsew
rlabel metal2 s 3504 3950 3504 3950 4 gnd
port 514 nsew
rlabel metal2 s 4752 3950 4752 3950 4 gnd
port 514 nsew
rlabel metal2 s 2736 4740 2736 4740 4 gnd
port 514 nsew
rlabel metal2 s 2736 3713 2736 3713 4 gnd
port 514 nsew
rlabel metal2 s 3984 3397 3984 3397 4 gnd
port 514 nsew
rlabel metal2 s 3984 5767 3984 5767 4 gnd
port 514 nsew
rlabel metal2 s 3984 6320 3984 6320 4 gnd
port 514 nsew
rlabel metal2 s 3984 6083 3984 6083 4 gnd
port 514 nsew
rlabel metal2 s 3984 4740 3984 4740 4 gnd
port 514 nsew
rlabel metal2 s 4752 5767 4752 5767 4 gnd
port 514 nsew
rlabel metal2 s 3504 5293 3504 5293 4 gnd
port 514 nsew
rlabel metal2 s 3504 6083 3504 6083 4 gnd
port 514 nsew
rlabel metal2 s 3504 3397 3504 3397 4 gnd
port 514 nsew
rlabel metal2 s 4752 4977 4752 4977 4 gnd
port 514 nsew
rlabel metal2 s 3504 5530 3504 5530 4 gnd
port 514 nsew
rlabel metal2 s 3504 6320 3504 6320 4 gnd
port 514 nsew
rlabel metal2 s 2256 6083 2256 6083 4 gnd
port 514 nsew
rlabel metal2 s 240 4977 240 4977 4 gnd
port 514 nsew
rlabel metal2 s 240 5767 240 5767 4 gnd
port 514 nsew
rlabel metal2 s 1008 3950 1008 3950 4 gnd
port 514 nsew
rlabel metal2 s 2256 6320 2256 6320 4 gnd
port 514 nsew
rlabel metal2 s 240 6083 240 6083 4 gnd
port 514 nsew
rlabel metal2 s 1008 5530 1008 5530 4 gnd
port 514 nsew
rlabel metal2 s 1008 5293 1008 5293 4 gnd
port 514 nsew
rlabel metal2 s 1488 4740 1488 4740 4 gnd
port 514 nsew
rlabel metal2 s 240 5530 240 5530 4 gnd
port 514 nsew
rlabel metal2 s 2256 4740 2256 4740 4 gnd
port 514 nsew
rlabel metal2 s 2256 5767 2256 5767 4 gnd
port 514 nsew
rlabel metal2 s 1488 4977 1488 4977 4 gnd
port 514 nsew
rlabel metal2 s 2256 4187 2256 4187 4 gnd
port 514 nsew
rlabel metal2 s 2256 3950 2256 3950 4 gnd
port 514 nsew
rlabel metal2 s 240 3950 240 3950 4 gnd
port 514 nsew
rlabel metal2 s 240 4503 240 4503 4 gnd
port 514 nsew
rlabel metal2 s 1008 3397 1008 3397 4 gnd
port 514 nsew
rlabel metal2 s 1008 4503 1008 4503 4 gnd
port 514 nsew
rlabel metal2 s 1488 3950 1488 3950 4 gnd
port 514 nsew
rlabel metal2 s 1488 5293 1488 5293 4 gnd
port 514 nsew
rlabel metal2 s 1488 3397 1488 3397 4 gnd
port 514 nsew
rlabel metal2 s 2256 4503 2256 4503 4 gnd
port 514 nsew
rlabel metal2 s 1488 5530 1488 5530 4 gnd
port 514 nsew
rlabel metal2 s 240 3713 240 3713 4 gnd
port 514 nsew
rlabel metal2 s 2256 5293 2256 5293 4 gnd
port 514 nsew
rlabel metal2 s 240 4740 240 4740 4 gnd
port 514 nsew
rlabel metal2 s 240 3397 240 3397 4 gnd
port 514 nsew
rlabel metal2 s 240 4187 240 4187 4 gnd
port 514 nsew
rlabel metal2 s 1008 6320 1008 6320 4 gnd
port 514 nsew
rlabel metal2 s 1008 4977 1008 4977 4 gnd
port 514 nsew
rlabel metal2 s 1488 4503 1488 4503 4 gnd
port 514 nsew
rlabel metal2 s 1008 6083 1008 6083 4 gnd
port 514 nsew
rlabel metal2 s 1488 5767 1488 5767 4 gnd
port 514 nsew
rlabel metal2 s 240 6320 240 6320 4 gnd
port 514 nsew
rlabel metal2 s 1488 3713 1488 3713 4 gnd
port 514 nsew
rlabel metal2 s 1008 4187 1008 4187 4 gnd
port 514 nsew
rlabel metal2 s 1008 5767 1008 5767 4 gnd
port 514 nsew
rlabel metal2 s 1488 6320 1488 6320 4 gnd
port 514 nsew
rlabel metal2 s 1488 6083 1488 6083 4 gnd
port 514 nsew
rlabel metal2 s 2256 3397 2256 3397 4 gnd
port 514 nsew
rlabel metal2 s 2256 3713 2256 3713 4 gnd
port 514 nsew
rlabel metal2 s 2256 5530 2256 5530 4 gnd
port 514 nsew
rlabel metal2 s 240 5293 240 5293 4 gnd
port 514 nsew
rlabel metal2 s 2256 4977 2256 4977 4 gnd
port 514 nsew
rlabel metal2 s 1488 4187 1488 4187 4 gnd
port 514 nsew
rlabel metal2 s 1008 4740 1008 4740 4 gnd
port 514 nsew
rlabel metal2 s 1008 3713 1008 3713 4 gnd
port 514 nsew
rlabel metal2 s 1008 2370 1008 2370 4 gnd
port 514 nsew
rlabel metal2 s 1008 237 1008 237 4 gnd
port 514 nsew
rlabel metal2 s 240 1027 240 1027 4 gnd
port 514 nsew
rlabel metal2 s 1488 1027 1488 1027 4 gnd
port 514 nsew
rlabel metal2 s 1488 2923 1488 2923 4 gnd
port 514 nsew
rlabel metal2 s 1488 2133 1488 2133 4 gnd
port 514 nsew
rlabel metal2 s 1488 553 1488 553 4 gnd
port 514 nsew
rlabel metal2 s 2256 2607 2256 2607 4 gnd
port 514 nsew
rlabel metal2 s 1488 1817 1488 1817 4 gnd
port 514 nsew
rlabel metal2 s 1488 237 1488 237 4 gnd
port 514 nsew
rlabel metal2 s 2256 237 2256 237 4 gnd
port 514 nsew
rlabel metal2 s 1488 1343 1488 1343 4 gnd
port 514 nsew
rlabel metal2 s 1008 1343 1008 1343 4 gnd
port 514 nsew
rlabel metal2 s 1488 2607 1488 2607 4 gnd
port 514 nsew
rlabel metal2 s 2256 0 2256 0 4 gnd
port 514 nsew
rlabel metal2 s 2256 790 2256 790 4 gnd
port 514 nsew
rlabel metal2 s 2256 2133 2256 2133 4 gnd
port 514 nsew
rlabel metal2 s 1488 1580 1488 1580 4 gnd
port 514 nsew
rlabel metal2 s 1008 1027 1008 1027 4 gnd
port 514 nsew
rlabel metal2 s 240 0 240 0 4 gnd
port 514 nsew
rlabel metal2 s 1008 1817 1008 1817 4 gnd
port 514 nsew
rlabel metal2 s 2256 553 2256 553 4 gnd
port 514 nsew
rlabel metal2 s 2256 1027 2256 1027 4 gnd
port 514 nsew
rlabel metal2 s 240 2923 240 2923 4 gnd
port 514 nsew
rlabel metal2 s 2256 2923 2256 2923 4 gnd
port 514 nsew
rlabel metal2 s 2256 1343 2256 1343 4 gnd
port 514 nsew
rlabel metal2 s 240 790 240 790 4 gnd
port 514 nsew
rlabel metal2 s 240 2607 240 2607 4 gnd
port 514 nsew
rlabel metal2 s 240 553 240 553 4 gnd
port 514 nsew
rlabel metal2 s 240 237 240 237 4 gnd
port 514 nsew
rlabel metal2 s 1008 2607 1008 2607 4 gnd
port 514 nsew
rlabel metal2 s 1488 0 1488 0 4 gnd
port 514 nsew
rlabel metal2 s 1008 790 1008 790 4 gnd
port 514 nsew
rlabel metal2 s 240 1580 240 1580 4 gnd
port 514 nsew
rlabel metal2 s 2256 2370 2256 2370 4 gnd
port 514 nsew
rlabel metal2 s 1488 3160 1488 3160 4 gnd
port 514 nsew
rlabel metal2 s 1008 2133 1008 2133 4 gnd
port 514 nsew
rlabel metal2 s 1008 553 1008 553 4 gnd
port 514 nsew
rlabel metal2 s 240 2370 240 2370 4 gnd
port 514 nsew
rlabel metal2 s 2256 1817 2256 1817 4 gnd
port 514 nsew
rlabel metal2 s 240 1343 240 1343 4 gnd
port 514 nsew
rlabel metal2 s 1008 3160 1008 3160 4 gnd
port 514 nsew
rlabel metal2 s 1008 1580 1008 1580 4 gnd
port 514 nsew
rlabel metal2 s 1488 2370 1488 2370 4 gnd
port 514 nsew
rlabel metal2 s 2256 1580 2256 1580 4 gnd
port 514 nsew
rlabel metal2 s 240 2133 240 2133 4 gnd
port 514 nsew
rlabel metal2 s 1008 2923 1008 2923 4 gnd
port 514 nsew
rlabel metal2 s 240 1817 240 1817 4 gnd
port 514 nsew
rlabel metal2 s 2256 3160 2256 3160 4 gnd
port 514 nsew
rlabel metal2 s 1008 0 1008 0 4 gnd
port 514 nsew
rlabel metal2 s 1488 790 1488 790 4 gnd
port 514 nsew
rlabel metal2 s 240 3160 240 3160 4 gnd
port 514 nsew
rlabel metal2 s 3984 1343 3984 1343 4 gnd
port 514 nsew
rlabel metal2 s 2736 790 2736 790 4 gnd
port 514 nsew
rlabel metal2 s 3504 2607 3504 2607 4 gnd
port 514 nsew
rlabel metal2 s 3504 553 3504 553 4 gnd
port 514 nsew
rlabel metal2 s 3504 1343 3504 1343 4 gnd
port 514 nsew
rlabel metal2 s 3504 3160 3504 3160 4 gnd
port 514 nsew
rlabel metal2 s 4752 1817 4752 1817 4 gnd
port 514 nsew
rlabel metal2 s 3504 1580 3504 1580 4 gnd
port 514 nsew
rlabel metal2 s 3984 2923 3984 2923 4 gnd
port 514 nsew
rlabel metal2 s 4752 2607 4752 2607 4 gnd
port 514 nsew
rlabel metal2 s 4752 553 4752 553 4 gnd
port 514 nsew
rlabel metal2 s 2736 0 2736 0 4 gnd
port 514 nsew
rlabel metal2 s 4752 1027 4752 1027 4 gnd
port 514 nsew
rlabel metal2 s 3984 2133 3984 2133 4 gnd
port 514 nsew
rlabel metal2 s 2736 2133 2736 2133 4 gnd
port 514 nsew
rlabel metal2 s 3984 2607 3984 2607 4 gnd
port 514 nsew
rlabel metal2 s 4752 2133 4752 2133 4 gnd
port 514 nsew
rlabel metal2 s 4752 237 4752 237 4 gnd
port 514 nsew
rlabel metal2 s 3984 1817 3984 1817 4 gnd
port 514 nsew
rlabel metal2 s 4752 3160 4752 3160 4 gnd
port 514 nsew
rlabel metal2 s 3984 0 3984 0 4 gnd
port 514 nsew
rlabel metal2 s 3984 1580 3984 1580 4 gnd
port 514 nsew
rlabel metal2 s 3504 2923 3504 2923 4 gnd
port 514 nsew
rlabel metal2 s 3984 790 3984 790 4 gnd
port 514 nsew
rlabel metal2 s 2736 2923 2736 2923 4 gnd
port 514 nsew
rlabel metal2 s 4752 2923 4752 2923 4 gnd
port 514 nsew
rlabel metal2 s 2736 1580 2736 1580 4 gnd
port 514 nsew
rlabel metal2 s 4752 2370 4752 2370 4 gnd
port 514 nsew
rlabel metal2 s 4752 790 4752 790 4 gnd
port 514 nsew
rlabel metal2 s 4752 1343 4752 1343 4 gnd
port 514 nsew
rlabel metal2 s 4752 1580 4752 1580 4 gnd
port 514 nsew
rlabel metal2 s 3504 237 3504 237 4 gnd
port 514 nsew
rlabel metal2 s 3504 2370 3504 2370 4 gnd
port 514 nsew
rlabel metal2 s 2736 1343 2736 1343 4 gnd
port 514 nsew
rlabel metal2 s 3504 790 3504 790 4 gnd
port 514 nsew
rlabel metal2 s 3984 1027 3984 1027 4 gnd
port 514 nsew
rlabel metal2 s 2736 2607 2736 2607 4 gnd
port 514 nsew
rlabel metal2 s 3984 3160 3984 3160 4 gnd
port 514 nsew
rlabel metal2 s 3504 0 3504 0 4 gnd
port 514 nsew
rlabel metal2 s 3984 2370 3984 2370 4 gnd
port 514 nsew
rlabel metal2 s 3504 1027 3504 1027 4 gnd
port 514 nsew
rlabel metal2 s 3984 237 3984 237 4 gnd
port 514 nsew
rlabel metal2 s 3984 553 3984 553 4 gnd
port 514 nsew
rlabel metal2 s 2736 1027 2736 1027 4 gnd
port 514 nsew
rlabel metal2 s 4752 0 4752 0 4 gnd
port 514 nsew
rlabel metal2 s 2736 237 2736 237 4 gnd
port 514 nsew
rlabel metal2 s 3504 2133 3504 2133 4 gnd
port 514 nsew
rlabel metal2 s 2736 1817 2736 1817 4 gnd
port 514 nsew
rlabel metal2 s 2736 553 2736 553 4 gnd
port 514 nsew
rlabel metal2 s 2736 2370 2736 2370 4 gnd
port 514 nsew
rlabel metal2 s 2736 3160 2736 3160 4 gnd
port 514 nsew
rlabel metal2 s 3504 1817 3504 1817 4 gnd
port 514 nsew
rlabel metal2 s 8496 4187 8496 4187 4 gnd
port 514 nsew
rlabel metal2 s 7728 3950 7728 3950 4 gnd
port 514 nsew
rlabel metal2 s 8976 4187 8976 4187 4 gnd
port 514 nsew
rlabel metal2 s 7728 4977 7728 4977 4 gnd
port 514 nsew
rlabel metal2 s 9744 6320 9744 6320 4 gnd
port 514 nsew
rlabel metal2 s 9744 5293 9744 5293 4 gnd
port 514 nsew
rlabel metal2 s 8976 5767 8976 5767 4 gnd
port 514 nsew
rlabel metal2 s 8976 5293 8976 5293 4 gnd
port 514 nsew
rlabel metal2 s 8496 5530 8496 5530 4 gnd
port 514 nsew
rlabel metal2 s 8976 4503 8976 4503 4 gnd
port 514 nsew
rlabel metal2 s 8976 3713 8976 3713 4 gnd
port 514 nsew
rlabel metal2 s 9744 4503 9744 4503 4 gnd
port 514 nsew
rlabel metal2 s 9744 5530 9744 5530 4 gnd
port 514 nsew
rlabel metal2 s 8976 6083 8976 6083 4 gnd
port 514 nsew
rlabel metal2 s 7728 3713 7728 3713 4 gnd
port 514 nsew
rlabel metal2 s 7728 5293 7728 5293 4 gnd
port 514 nsew
rlabel metal2 s 8496 5767 8496 5767 4 gnd
port 514 nsew
rlabel metal2 s 7728 6083 7728 6083 4 gnd
port 514 nsew
rlabel metal2 s 8496 5293 8496 5293 4 gnd
port 514 nsew
rlabel metal2 s 8976 6320 8976 6320 4 gnd
port 514 nsew
rlabel metal2 s 8496 3397 8496 3397 4 gnd
port 514 nsew
rlabel metal2 s 7728 6320 7728 6320 4 gnd
port 514 nsew
rlabel metal2 s 8976 3397 8976 3397 4 gnd
port 514 nsew
rlabel metal2 s 9744 3397 9744 3397 4 gnd
port 514 nsew
rlabel metal2 s 8976 3950 8976 3950 4 gnd
port 514 nsew
rlabel metal2 s 9744 3950 9744 3950 4 gnd
port 514 nsew
rlabel metal2 s 7728 4503 7728 4503 4 gnd
port 514 nsew
rlabel metal2 s 8976 4740 8976 4740 4 gnd
port 514 nsew
rlabel metal2 s 7728 5530 7728 5530 4 gnd
port 514 nsew
rlabel metal2 s 8976 4977 8976 4977 4 gnd
port 514 nsew
rlabel metal2 s 8496 4740 8496 4740 4 gnd
port 514 nsew
rlabel metal2 s 8496 6083 8496 6083 4 gnd
port 514 nsew
rlabel metal2 s 9744 3713 9744 3713 4 gnd
port 514 nsew
rlabel metal2 s 9744 4187 9744 4187 4 gnd
port 514 nsew
rlabel metal2 s 8496 6320 8496 6320 4 gnd
port 514 nsew
rlabel metal2 s 7728 4740 7728 4740 4 gnd
port 514 nsew
rlabel metal2 s 7728 5767 7728 5767 4 gnd
port 514 nsew
rlabel metal2 s 7728 3397 7728 3397 4 gnd
port 514 nsew
rlabel metal2 s 8496 3713 8496 3713 4 gnd
port 514 nsew
rlabel metal2 s 9744 4977 9744 4977 4 gnd
port 514 nsew
rlabel metal2 s 9744 5767 9744 5767 4 gnd
port 514 nsew
rlabel metal2 s 8496 4977 8496 4977 4 gnd
port 514 nsew
rlabel metal2 s 8496 4503 8496 4503 4 gnd
port 514 nsew
rlabel metal2 s 9744 4740 9744 4740 4 gnd
port 514 nsew
rlabel metal2 s 7728 4187 7728 4187 4 gnd
port 514 nsew
rlabel metal2 s 9744 6083 9744 6083 4 gnd
port 514 nsew
rlabel metal2 s 8976 5530 8976 5530 4 gnd
port 514 nsew
rlabel metal2 s 8496 3950 8496 3950 4 gnd
port 514 nsew
rlabel metal2 s 6000 3713 6000 3713 4 gnd
port 514 nsew
rlabel metal2 s 7248 4503 7248 4503 4 gnd
port 514 nsew
rlabel metal2 s 6000 6083 6000 6083 4 gnd
port 514 nsew
rlabel metal2 s 6480 4187 6480 4187 4 gnd
port 514 nsew
rlabel metal2 s 5232 3397 5232 3397 4 gnd
port 514 nsew
rlabel metal2 s 6000 3950 6000 3950 4 gnd
port 514 nsew
rlabel metal2 s 7248 6083 7248 6083 4 gnd
port 514 nsew
rlabel metal2 s 5232 3713 5232 3713 4 gnd
port 514 nsew
rlabel metal2 s 5232 5530 5232 5530 4 gnd
port 514 nsew
rlabel metal2 s 5232 6320 5232 6320 4 gnd
port 514 nsew
rlabel metal2 s 7248 5767 7248 5767 4 gnd
port 514 nsew
rlabel metal2 s 7248 3713 7248 3713 4 gnd
port 514 nsew
rlabel metal2 s 7248 4977 7248 4977 4 gnd
port 514 nsew
rlabel metal2 s 7248 5530 7248 5530 4 gnd
port 514 nsew
rlabel metal2 s 6480 3950 6480 3950 4 gnd
port 514 nsew
rlabel metal2 s 6000 6320 6000 6320 4 gnd
port 514 nsew
rlabel metal2 s 6000 4187 6000 4187 4 gnd
port 514 nsew
rlabel metal2 s 6480 3397 6480 3397 4 gnd
port 514 nsew
rlabel metal2 s 7248 4740 7248 4740 4 gnd
port 514 nsew
rlabel metal2 s 6480 6320 6480 6320 4 gnd
port 514 nsew
rlabel metal2 s 5232 4977 5232 4977 4 gnd
port 514 nsew
rlabel metal2 s 6480 5293 6480 5293 4 gnd
port 514 nsew
rlabel metal2 s 6000 5293 6000 5293 4 gnd
port 514 nsew
rlabel metal2 s 5232 4187 5232 4187 4 gnd
port 514 nsew
rlabel metal2 s 7248 5293 7248 5293 4 gnd
port 514 nsew
rlabel metal2 s 6000 4977 6000 4977 4 gnd
port 514 nsew
rlabel metal2 s 6480 5530 6480 5530 4 gnd
port 514 nsew
rlabel metal2 s 6000 5530 6000 5530 4 gnd
port 514 nsew
rlabel metal2 s 6480 3713 6480 3713 4 gnd
port 514 nsew
rlabel metal2 s 6480 4503 6480 4503 4 gnd
port 514 nsew
rlabel metal2 s 5232 5767 5232 5767 4 gnd
port 514 nsew
rlabel metal2 s 5232 6083 5232 6083 4 gnd
port 514 nsew
rlabel metal2 s 5232 5293 5232 5293 4 gnd
port 514 nsew
rlabel metal2 s 6480 5767 6480 5767 4 gnd
port 514 nsew
rlabel metal2 s 5232 3950 5232 3950 4 gnd
port 514 nsew
rlabel metal2 s 6000 5767 6000 5767 4 gnd
port 514 nsew
rlabel metal2 s 7248 4187 7248 4187 4 gnd
port 514 nsew
rlabel metal2 s 6000 3397 6000 3397 4 gnd
port 514 nsew
rlabel metal2 s 5232 4503 5232 4503 4 gnd
port 514 nsew
rlabel metal2 s 6000 4740 6000 4740 4 gnd
port 514 nsew
rlabel metal2 s 5232 4740 5232 4740 4 gnd
port 514 nsew
rlabel metal2 s 7248 6320 7248 6320 4 gnd
port 514 nsew
rlabel metal2 s 6480 4977 6480 4977 4 gnd
port 514 nsew
rlabel metal2 s 7248 3397 7248 3397 4 gnd
port 514 nsew
rlabel metal2 s 6480 4740 6480 4740 4 gnd
port 514 nsew
rlabel metal2 s 7248 3950 7248 3950 4 gnd
port 514 nsew
rlabel metal2 s 6000 4503 6000 4503 4 gnd
port 514 nsew
rlabel metal2 s 6480 6083 6480 6083 4 gnd
port 514 nsew
rlabel metal2 s 6480 790 6480 790 4 gnd
port 514 nsew
rlabel metal2 s 6480 553 6480 553 4 gnd
port 514 nsew
rlabel metal2 s 7248 1580 7248 1580 4 gnd
port 514 nsew
rlabel metal2 s 6000 2607 6000 2607 4 gnd
port 514 nsew
rlabel metal2 s 6480 237 6480 237 4 gnd
port 514 nsew
rlabel metal2 s 7248 2370 7248 2370 4 gnd
port 514 nsew
rlabel metal2 s 5232 0 5232 0 4 gnd
port 514 nsew
rlabel metal2 s 6000 1580 6000 1580 4 gnd
port 514 nsew
rlabel metal2 s 5232 553 5232 553 4 gnd
port 514 nsew
rlabel metal2 s 5232 2133 5232 2133 4 gnd
port 514 nsew
rlabel metal2 s 7248 1343 7248 1343 4 gnd
port 514 nsew
rlabel metal2 s 6480 0 6480 0 4 gnd
port 514 nsew
rlabel metal2 s 6000 3160 6000 3160 4 gnd
port 514 nsew
rlabel metal2 s 6480 2923 6480 2923 4 gnd
port 514 nsew
rlabel metal2 s 5232 2370 5232 2370 4 gnd
port 514 nsew
rlabel metal2 s 7248 790 7248 790 4 gnd
port 514 nsew
rlabel metal2 s 5232 2607 5232 2607 4 gnd
port 514 nsew
rlabel metal2 s 6480 1343 6480 1343 4 gnd
port 514 nsew
rlabel metal2 s 6000 237 6000 237 4 gnd
port 514 nsew
rlabel metal2 s 6480 2607 6480 2607 4 gnd
port 514 nsew
rlabel metal2 s 7248 1817 7248 1817 4 gnd
port 514 nsew
rlabel metal2 s 5232 1027 5232 1027 4 gnd
port 514 nsew
rlabel metal2 s 7248 2607 7248 2607 4 gnd
port 514 nsew
rlabel metal2 s 6480 2133 6480 2133 4 gnd
port 514 nsew
rlabel metal2 s 7248 2133 7248 2133 4 gnd
port 514 nsew
rlabel metal2 s 7248 3160 7248 3160 4 gnd
port 514 nsew
rlabel metal2 s 7248 1027 7248 1027 4 gnd
port 514 nsew
rlabel metal2 s 6000 553 6000 553 4 gnd
port 514 nsew
rlabel metal2 s 5232 1580 5232 1580 4 gnd
port 514 nsew
rlabel metal2 s 7248 237 7248 237 4 gnd
port 514 nsew
rlabel metal2 s 6480 2370 6480 2370 4 gnd
port 514 nsew
rlabel metal2 s 6000 2370 6000 2370 4 gnd
port 514 nsew
rlabel metal2 s 6000 1343 6000 1343 4 gnd
port 514 nsew
rlabel metal2 s 5232 1343 5232 1343 4 gnd
port 514 nsew
rlabel metal2 s 5232 3160 5232 3160 4 gnd
port 514 nsew
rlabel metal2 s 7248 553 7248 553 4 gnd
port 514 nsew
rlabel metal2 s 6480 1580 6480 1580 4 gnd
port 514 nsew
rlabel metal2 s 6480 1027 6480 1027 4 gnd
port 514 nsew
rlabel metal2 s 6480 3160 6480 3160 4 gnd
port 514 nsew
rlabel metal2 s 6480 1817 6480 1817 4 gnd
port 514 nsew
rlabel metal2 s 5232 237 5232 237 4 gnd
port 514 nsew
rlabel metal2 s 6000 2923 6000 2923 4 gnd
port 514 nsew
rlabel metal2 s 6000 1027 6000 1027 4 gnd
port 514 nsew
rlabel metal2 s 7248 2923 7248 2923 4 gnd
port 514 nsew
rlabel metal2 s 6000 2133 6000 2133 4 gnd
port 514 nsew
rlabel metal2 s 5232 1817 5232 1817 4 gnd
port 514 nsew
rlabel metal2 s 7248 0 7248 0 4 gnd
port 514 nsew
rlabel metal2 s 6000 1817 6000 1817 4 gnd
port 514 nsew
rlabel metal2 s 5232 2923 5232 2923 4 gnd
port 514 nsew
rlabel metal2 s 5232 790 5232 790 4 gnd
port 514 nsew
rlabel metal2 s 6000 0 6000 0 4 gnd
port 514 nsew
rlabel metal2 s 6000 790 6000 790 4 gnd
port 514 nsew
rlabel metal2 s 9744 790 9744 790 4 gnd
port 514 nsew
rlabel metal2 s 8976 2133 8976 2133 4 gnd
port 514 nsew
rlabel metal2 s 7728 790 7728 790 4 gnd
port 514 nsew
rlabel metal2 s 8496 1027 8496 1027 4 gnd
port 514 nsew
rlabel metal2 s 9744 2607 9744 2607 4 gnd
port 514 nsew
rlabel metal2 s 8976 2607 8976 2607 4 gnd
port 514 nsew
rlabel metal2 s 8976 3160 8976 3160 4 gnd
port 514 nsew
rlabel metal2 s 8976 2370 8976 2370 4 gnd
port 514 nsew
rlabel metal2 s 9744 2370 9744 2370 4 gnd
port 514 nsew
rlabel metal2 s 9744 1580 9744 1580 4 gnd
port 514 nsew
rlabel metal2 s 7728 1580 7728 1580 4 gnd
port 514 nsew
rlabel metal2 s 7728 1027 7728 1027 4 gnd
port 514 nsew
rlabel metal2 s 9744 2923 9744 2923 4 gnd
port 514 nsew
rlabel metal2 s 9744 3160 9744 3160 4 gnd
port 514 nsew
rlabel metal2 s 9744 237 9744 237 4 gnd
port 514 nsew
rlabel metal2 s 8496 1580 8496 1580 4 gnd
port 514 nsew
rlabel metal2 s 8496 1343 8496 1343 4 gnd
port 514 nsew
rlabel metal2 s 7728 3160 7728 3160 4 gnd
port 514 nsew
rlabel metal2 s 7728 2607 7728 2607 4 gnd
port 514 nsew
rlabel metal2 s 7728 0 7728 0 4 gnd
port 514 nsew
rlabel metal2 s 8496 3160 8496 3160 4 gnd
port 514 nsew
rlabel metal2 s 8976 237 8976 237 4 gnd
port 514 nsew
rlabel metal2 s 9744 553 9744 553 4 gnd
port 514 nsew
rlabel metal2 s 9744 2133 9744 2133 4 gnd
port 514 nsew
rlabel metal2 s 7728 1817 7728 1817 4 gnd
port 514 nsew
rlabel metal2 s 7728 1343 7728 1343 4 gnd
port 514 nsew
rlabel metal2 s 7728 2133 7728 2133 4 gnd
port 514 nsew
rlabel metal2 s 8976 1580 8976 1580 4 gnd
port 514 nsew
rlabel metal2 s 9744 0 9744 0 4 gnd
port 514 nsew
rlabel metal2 s 8496 790 8496 790 4 gnd
port 514 nsew
rlabel metal2 s 8976 1817 8976 1817 4 gnd
port 514 nsew
rlabel metal2 s 8496 2133 8496 2133 4 gnd
port 514 nsew
rlabel metal2 s 8976 1343 8976 1343 4 gnd
port 514 nsew
rlabel metal2 s 7728 2923 7728 2923 4 gnd
port 514 nsew
rlabel metal2 s 8496 2607 8496 2607 4 gnd
port 514 nsew
rlabel metal2 s 8976 0 8976 0 4 gnd
port 514 nsew
rlabel metal2 s 9744 1817 9744 1817 4 gnd
port 514 nsew
rlabel metal2 s 8976 2923 8976 2923 4 gnd
port 514 nsew
rlabel metal2 s 8976 553 8976 553 4 gnd
port 514 nsew
rlabel metal2 s 8976 1027 8976 1027 4 gnd
port 514 nsew
rlabel metal2 s 8496 0 8496 0 4 gnd
port 514 nsew
rlabel metal2 s 7728 2370 7728 2370 4 gnd
port 514 nsew
rlabel metal2 s 8496 553 8496 553 4 gnd
port 514 nsew
rlabel metal2 s 9744 1343 9744 1343 4 gnd
port 514 nsew
rlabel metal2 s 7728 237 7728 237 4 gnd
port 514 nsew
rlabel metal2 s 8496 2923 8496 2923 4 gnd
port 514 nsew
rlabel metal2 s 8496 1817 8496 1817 4 gnd
port 514 nsew
rlabel metal2 s 8976 790 8976 790 4 gnd
port 514 nsew
rlabel metal2 s 8496 2370 8496 2370 4 gnd
port 514 nsew
rlabel metal2 s 9744 1027 9744 1027 4 gnd
port 514 nsew
rlabel metal2 s 7728 553 7728 553 4 gnd
port 514 nsew
rlabel metal2 s 8496 237 8496 237 4 gnd
port 514 nsew
rlabel metal2 s 18960 10270 18960 10270 4 gnd
port 514 nsew
rlabel metal2 s 18480 12403 18480 12403 4 gnd
port 514 nsew
rlabel metal2 s 19968 12293 19968 12293 4 wl0_31
port 319 nsew
rlabel metal2 s 18480 10033 18480 10033 4 gnd
port 514 nsew
rlabel metal2 s 19728 11060 19728 11060 4 gnd
port 514 nsew
rlabel metal2 s 18480 9717 18480 9717 4 gnd
port 514 nsew
rlabel metal2 s 18480 11060 18480 11060 4 gnd
port 514 nsew
rlabel metal2 s 19728 10033 19728 10033 4 gnd
port 514 nsew
rlabel metal2 s 19968 11723 19968 11723 4 wl1_29
port 316 nsew
rlabel metal2 s 17712 12640 17712 12640 4 gnd
port 514 nsew
rlabel metal2 s 19728 11613 19728 11613 4 gnd
port 514 nsew
rlabel metal2 s 18480 10823 18480 10823 4 gnd
port 514 nsew
rlabel metal2 s 17712 11297 17712 11297 4 gnd
port 514 nsew
rlabel metal2 s 19728 11850 19728 11850 4 gnd
port 514 nsew
rlabel metal2 s 18960 11297 18960 11297 4 gnd
port 514 nsew
rlabel metal2 s 17712 11850 17712 11850 4 gnd
port 514 nsew
rlabel metal2 s 19728 12403 19728 12403 4 gnd
port 514 nsew
rlabel metal2 s 19728 11297 19728 11297 4 gnd
port 514 nsew
rlabel metal2 s 18480 12087 18480 12087 4 gnd
port 514 nsew
rlabel metal2 s 18960 11850 18960 11850 4 gnd
port 514 nsew
rlabel metal2 s 19728 9717 19728 9717 4 gnd
port 514 nsew
rlabel metal2 s 17712 10507 17712 10507 4 gnd
port 514 nsew
rlabel metal2 s 19728 10270 19728 10270 4 gnd
port 514 nsew
rlabel metal2 s 19968 10713 19968 10713 4 wl0_27
port 311 nsew
rlabel metal2 s 19968 10397 19968 10397 4 wl1_26
port 310 nsew
rlabel metal2 s 18480 10270 18480 10270 4 gnd
port 514 nsew
rlabel metal2 s 18960 9717 18960 9717 4 gnd
port 514 nsew
rlabel metal2 s 17712 10270 17712 10270 4 gnd
port 514 nsew
rlabel metal2 s 19968 10617 19968 10617 4 wl0_26
port 309 nsew
rlabel metal2 s 18960 10033 18960 10033 4 gnd
port 514 nsew
rlabel metal2 s 18960 11613 18960 11613 4 gnd
port 514 nsew
rlabel metal2 s 18480 10507 18480 10507 4 gnd
port 514 nsew
rlabel metal2 s 18960 10507 18960 10507 4 gnd
port 514 nsew
rlabel metal2 s 19968 10143 19968 10143 4 wl1_25
port 308 nsew
rlabel metal2 s 18480 11850 18480 11850 4 gnd
port 514 nsew
rlabel metal2 s 17712 9717 17712 9717 4 gnd
port 514 nsew
rlabel metal2 s 18480 12640 18480 12640 4 gnd
port 514 nsew
rlabel metal2 s 18960 12087 18960 12087 4 gnd
port 514 nsew
rlabel metal2 s 18960 12640 18960 12640 4 gnd
port 514 nsew
rlabel metal2 s 18960 11060 18960 11060 4 gnd
port 514 nsew
rlabel metal2 s 17712 10033 17712 10033 4 gnd
port 514 nsew
rlabel metal2 s 19968 12197 19968 12197 4 wl0_30
port 317 nsew
rlabel metal2 s 17712 10823 17712 10823 4 gnd
port 514 nsew
rlabel metal2 s 19728 12640 19728 12640 4 gnd
port 514 nsew
rlabel metal2 s 17712 12403 17712 12403 4 gnd
port 514 nsew
rlabel metal2 s 19728 12087 19728 12087 4 gnd
port 514 nsew
rlabel metal2 s 18960 12403 18960 12403 4 gnd
port 514 nsew
rlabel metal2 s 18960 10823 18960 10823 4 gnd
port 514 nsew
rlabel metal2 s 17712 11613 17712 11613 4 gnd
port 514 nsew
rlabel metal2 s 19968 9607 19968 9607 4 wl1_24
port 306 nsew
rlabel metal2 s 19968 9923 19968 9923 4 wl0_25
port 307 nsew
rlabel metal2 s 17712 12087 17712 12087 4 gnd
port 514 nsew
rlabel metal2 s 17712 11060 17712 11060 4 gnd
port 514 nsew
rlabel metal2 s 19968 11977 19968 11977 4 wl1_30
port 318 nsew
rlabel metal2 s 18480 11613 18480 11613 4 gnd
port 514 nsew
rlabel metal2 s 19968 12513 19968 12513 4 wl1_31
port 320 nsew
rlabel metal2 s 19968 10933 19968 10933 4 wl1_27
port 312 nsew
rlabel metal2 s 19728 10823 19728 10823 4 gnd
port 514 nsew
rlabel metal2 s 19968 9827 19968 9827 4 wl0_24
port 305 nsew
rlabel metal2 s 19728 10507 19728 10507 4 gnd
port 514 nsew
rlabel metal2 s 19968 11187 19968 11187 4 wl1_28
port 314 nsew
rlabel metal2 s 19968 11503 19968 11503 4 wl0_29
port 315 nsew
rlabel metal2 s 19968 11407 19968 11407 4 wl0_28
port 313 nsew
rlabel metal2 s 18480 11297 18480 11297 4 gnd
port 514 nsew
rlabel metal2 s 15984 11060 15984 11060 4 gnd
port 514 nsew
rlabel metal2 s 15216 10507 15216 10507 4 gnd
port 514 nsew
rlabel metal2 s 15216 12403 15216 12403 4 gnd
port 514 nsew
rlabel metal2 s 16464 12403 16464 12403 4 gnd
port 514 nsew
rlabel metal2 s 16464 10507 16464 10507 4 gnd
port 514 nsew
rlabel metal2 s 17232 11613 17232 11613 4 gnd
port 514 nsew
rlabel metal2 s 16464 11850 16464 11850 4 gnd
port 514 nsew
rlabel metal2 s 15216 11297 15216 11297 4 gnd
port 514 nsew
rlabel metal2 s 17232 12640 17232 12640 4 gnd
port 514 nsew
rlabel metal2 s 16464 10270 16464 10270 4 gnd
port 514 nsew
rlabel metal2 s 17232 10033 17232 10033 4 gnd
port 514 nsew
rlabel metal2 s 15216 12640 15216 12640 4 gnd
port 514 nsew
rlabel metal2 s 15984 10033 15984 10033 4 gnd
port 514 nsew
rlabel metal2 s 16464 9717 16464 9717 4 gnd
port 514 nsew
rlabel metal2 s 16464 12087 16464 12087 4 gnd
port 514 nsew
rlabel metal2 s 17232 12403 17232 12403 4 gnd
port 514 nsew
rlabel metal2 s 17232 11060 17232 11060 4 gnd
port 514 nsew
rlabel metal2 s 17232 10507 17232 10507 4 gnd
port 514 nsew
rlabel metal2 s 16464 10823 16464 10823 4 gnd
port 514 nsew
rlabel metal2 s 15216 11613 15216 11613 4 gnd
port 514 nsew
rlabel metal2 s 17232 11850 17232 11850 4 gnd
port 514 nsew
rlabel metal2 s 15984 10507 15984 10507 4 gnd
port 514 nsew
rlabel metal2 s 17232 10270 17232 10270 4 gnd
port 514 nsew
rlabel metal2 s 16464 10033 16464 10033 4 gnd
port 514 nsew
rlabel metal2 s 15984 11850 15984 11850 4 gnd
port 514 nsew
rlabel metal2 s 15984 12403 15984 12403 4 gnd
port 514 nsew
rlabel metal2 s 15216 10270 15216 10270 4 gnd
port 514 nsew
rlabel metal2 s 15216 10823 15216 10823 4 gnd
port 514 nsew
rlabel metal2 s 15984 10823 15984 10823 4 gnd
port 514 nsew
rlabel metal2 s 15984 10270 15984 10270 4 gnd
port 514 nsew
rlabel metal2 s 15216 11060 15216 11060 4 gnd
port 514 nsew
rlabel metal2 s 17232 9717 17232 9717 4 gnd
port 514 nsew
rlabel metal2 s 17232 10823 17232 10823 4 gnd
port 514 nsew
rlabel metal2 s 15216 9717 15216 9717 4 gnd
port 514 nsew
rlabel metal2 s 15984 12087 15984 12087 4 gnd
port 514 nsew
rlabel metal2 s 15216 12087 15216 12087 4 gnd
port 514 nsew
rlabel metal2 s 16464 11613 16464 11613 4 gnd
port 514 nsew
rlabel metal2 s 15984 12640 15984 12640 4 gnd
port 514 nsew
rlabel metal2 s 15216 11850 15216 11850 4 gnd
port 514 nsew
rlabel metal2 s 16464 11297 16464 11297 4 gnd
port 514 nsew
rlabel metal2 s 15216 10033 15216 10033 4 gnd
port 514 nsew
rlabel metal2 s 17232 12087 17232 12087 4 gnd
port 514 nsew
rlabel metal2 s 17232 11297 17232 11297 4 gnd
port 514 nsew
rlabel metal2 s 15984 11613 15984 11613 4 gnd
port 514 nsew
rlabel metal2 s 16464 11060 16464 11060 4 gnd
port 514 nsew
rlabel metal2 s 16464 12640 16464 12640 4 gnd
port 514 nsew
rlabel metal2 s 15984 11297 15984 11297 4 gnd
port 514 nsew
rlabel metal2 s 15984 9717 15984 9717 4 gnd
port 514 nsew
rlabel metal2 s 16464 7663 16464 7663 4 gnd
port 514 nsew
rlabel metal2 s 16464 9243 16464 9243 4 gnd
port 514 nsew
rlabel metal2 s 15984 7347 15984 7347 4 gnd
port 514 nsew
rlabel metal2 s 15216 8927 15216 8927 4 gnd
port 514 nsew
rlabel metal2 s 17232 9480 17232 9480 4 gnd
port 514 nsew
rlabel metal2 s 15216 7900 15216 7900 4 gnd
port 514 nsew
rlabel metal2 s 15984 7110 15984 7110 4 gnd
port 514 nsew
rlabel metal2 s 15984 9243 15984 9243 4 gnd
port 514 nsew
rlabel metal2 s 16464 6557 16464 6557 4 gnd
port 514 nsew
rlabel metal2 s 16464 9480 16464 9480 4 gnd
port 514 nsew
rlabel metal2 s 16464 8453 16464 8453 4 gnd
port 514 nsew
rlabel metal2 s 17232 8927 17232 8927 4 gnd
port 514 nsew
rlabel metal2 s 15216 9243 15216 9243 4 gnd
port 514 nsew
rlabel metal2 s 16464 8927 16464 8927 4 gnd
port 514 nsew
rlabel metal2 s 15216 8690 15216 8690 4 gnd
port 514 nsew
rlabel metal2 s 16464 8690 16464 8690 4 gnd
port 514 nsew
rlabel metal2 s 15216 6873 15216 6873 4 gnd
port 514 nsew
rlabel metal2 s 16464 6873 16464 6873 4 gnd
port 514 nsew
rlabel metal2 s 15984 8453 15984 8453 4 gnd
port 514 nsew
rlabel metal2 s 15984 6873 15984 6873 4 gnd
port 514 nsew
rlabel metal2 s 15216 7347 15216 7347 4 gnd
port 514 nsew
rlabel metal2 s 17232 7900 17232 7900 4 gnd
port 514 nsew
rlabel metal2 s 17232 9243 17232 9243 4 gnd
port 514 nsew
rlabel metal2 s 17232 6557 17232 6557 4 gnd
port 514 nsew
rlabel metal2 s 15984 6557 15984 6557 4 gnd
port 514 nsew
rlabel metal2 s 16464 7110 16464 7110 4 gnd
port 514 nsew
rlabel metal2 s 15216 9480 15216 9480 4 gnd
port 514 nsew
rlabel metal2 s 15984 8690 15984 8690 4 gnd
port 514 nsew
rlabel metal2 s 16464 7900 16464 7900 4 gnd
port 514 nsew
rlabel metal2 s 15216 8453 15216 8453 4 gnd
port 514 nsew
rlabel metal2 s 17232 8137 17232 8137 4 gnd
port 514 nsew
rlabel metal2 s 15984 9480 15984 9480 4 gnd
port 514 nsew
rlabel metal2 s 15984 7900 15984 7900 4 gnd
port 514 nsew
rlabel metal2 s 15216 7110 15216 7110 4 gnd
port 514 nsew
rlabel metal2 s 16464 7347 16464 7347 4 gnd
port 514 nsew
rlabel metal2 s 15984 8927 15984 8927 4 gnd
port 514 nsew
rlabel metal2 s 17232 8690 17232 8690 4 gnd
port 514 nsew
rlabel metal2 s 15216 7663 15216 7663 4 gnd
port 514 nsew
rlabel metal2 s 17232 7347 17232 7347 4 gnd
port 514 nsew
rlabel metal2 s 17232 7663 17232 7663 4 gnd
port 514 nsew
rlabel metal2 s 17232 7110 17232 7110 4 gnd
port 514 nsew
rlabel metal2 s 17232 8453 17232 8453 4 gnd
port 514 nsew
rlabel metal2 s 16464 8137 16464 8137 4 gnd
port 514 nsew
rlabel metal2 s 15984 7663 15984 7663 4 gnd
port 514 nsew
rlabel metal2 s 15984 8137 15984 8137 4 gnd
port 514 nsew
rlabel metal2 s 17232 6873 17232 6873 4 gnd
port 514 nsew
rlabel metal2 s 15216 8137 15216 8137 4 gnd
port 514 nsew
rlabel metal2 s 15216 6557 15216 6557 4 gnd
port 514 nsew
rlabel metal2 s 17712 8690 17712 8690 4 gnd
port 514 nsew
rlabel metal2 s 19728 6873 19728 6873 4 gnd
port 514 nsew
rlabel metal2 s 17712 7347 17712 7347 4 gnd
port 514 nsew
rlabel metal2 s 18960 7110 18960 7110 4 gnd
port 514 nsew
rlabel metal2 s 18960 9480 18960 9480 4 gnd
port 514 nsew
rlabel metal2 s 17712 7110 17712 7110 4 gnd
port 514 nsew
rlabel metal2 s 17712 9243 17712 9243 4 gnd
port 514 nsew
rlabel metal2 s 18960 8453 18960 8453 4 gnd
port 514 nsew
rlabel metal2 s 18480 7110 18480 7110 4 gnd
port 514 nsew
rlabel metal2 s 19968 9037 19968 9037 4 wl0_22
port 301 nsew
rlabel metal2 s 17712 8137 17712 8137 4 gnd
port 514 nsew
rlabel metal2 s 19728 7110 19728 7110 4 gnd
port 514 nsew
rlabel metal2 s 19968 8247 19968 8247 4 wl0_20
port 297 nsew
rlabel metal2 s 18480 7900 18480 7900 4 gnd
port 514 nsew
rlabel metal2 s 19728 9480 19728 9480 4 gnd
port 514 nsew
rlabel metal2 s 17712 9480 17712 9480 4 gnd
port 514 nsew
rlabel metal2 s 17712 7663 17712 7663 4 gnd
port 514 nsew
rlabel metal2 s 18480 7663 18480 7663 4 gnd
port 514 nsew
rlabel metal2 s 19968 6447 19968 6447 4 wl1_16
port 290 nsew
rlabel metal2 s 18960 9243 18960 9243 4 gnd
port 514 nsew
rlabel metal2 s 18960 7900 18960 7900 4 gnd
port 514 nsew
rlabel metal2 s 17712 7900 17712 7900 4 gnd
port 514 nsew
rlabel metal2 s 17712 8927 17712 8927 4 gnd
port 514 nsew
rlabel metal2 s 19968 8343 19968 8343 4 wl0_21
port 299 nsew
rlabel metal2 s 18960 6873 18960 6873 4 gnd
port 514 nsew
rlabel metal2 s 19968 8563 19968 8563 4 wl1_21
port 300 nsew
rlabel metal2 s 17712 6557 17712 6557 4 gnd
port 514 nsew
rlabel metal2 s 19728 8453 19728 8453 4 gnd
port 514 nsew
rlabel metal2 s 19968 7237 19968 7237 4 wl1_18
port 294 nsew
rlabel metal2 s 19968 7457 19968 7457 4 wl0_18
port 293 nsew
rlabel metal2 s 19968 8817 19968 8817 4 wl1_22
port 302 nsew
rlabel metal2 s 19728 7347 19728 7347 4 gnd
port 514 nsew
rlabel metal2 s 19728 6557 19728 6557 4 gnd
port 514 nsew
rlabel metal2 s 19728 8690 19728 8690 4 gnd
port 514 nsew
rlabel metal2 s 18960 8927 18960 8927 4 gnd
port 514 nsew
rlabel metal2 s 18480 7347 18480 7347 4 gnd
port 514 nsew
rlabel metal2 s 18480 6873 18480 6873 4 gnd
port 514 nsew
rlabel metal2 s 18960 8137 18960 8137 4 gnd
port 514 nsew
rlabel metal2 s 19968 9133 19968 9133 4 wl0_23
port 303 nsew
rlabel metal2 s 17712 8453 17712 8453 4 gnd
port 514 nsew
rlabel metal2 s 18960 8690 18960 8690 4 gnd
port 514 nsew
rlabel metal2 s 19968 6983 19968 6983 4 wl1_17
port 292 nsew
rlabel metal2 s 19968 8027 19968 8027 4 wl1_20
port 298 nsew
rlabel metal2 s 18960 6557 18960 6557 4 gnd
port 514 nsew
rlabel metal2 s 19968 9353 19968 9353 4 wl1_23
port 304 nsew
rlabel metal2 s 19728 7900 19728 7900 4 gnd
port 514 nsew
rlabel metal2 s 18480 6557 18480 6557 4 gnd
port 514 nsew
rlabel metal2 s 18960 7663 18960 7663 4 gnd
port 514 nsew
rlabel metal2 s 18480 8927 18480 8927 4 gnd
port 514 nsew
rlabel metal2 s 18480 9480 18480 9480 4 gnd
port 514 nsew
rlabel metal2 s 19728 7663 19728 7663 4 gnd
port 514 nsew
rlabel metal2 s 18960 7347 18960 7347 4 gnd
port 514 nsew
rlabel metal2 s 19728 9243 19728 9243 4 gnd
port 514 nsew
rlabel metal2 s 19728 8927 19728 8927 4 gnd
port 514 nsew
rlabel metal2 s 19968 7773 19968 7773 4 wl1_19
port 296 nsew
rlabel metal2 s 19968 6763 19968 6763 4 wl0_17
port 291 nsew
rlabel metal2 s 18480 9243 18480 9243 4 gnd
port 514 nsew
rlabel metal2 s 18480 8453 18480 8453 4 gnd
port 514 nsew
rlabel metal2 s 18480 8690 18480 8690 4 gnd
port 514 nsew
rlabel metal2 s 19728 8137 19728 8137 4 gnd
port 514 nsew
rlabel metal2 s 19968 7553 19968 7553 4 wl0_19
port 295 nsew
rlabel metal2 s 17712 6873 17712 6873 4 gnd
port 514 nsew
rlabel metal2 s 19968 6667 19968 6667 4 wl0_16
port 289 nsew
rlabel metal2 s 18480 8137 18480 8137 4 gnd
port 514 nsew
rlabel metal2 s 12720 10270 12720 10270 4 gnd
port 514 nsew
rlabel metal2 s 13968 11060 13968 11060 4 gnd
port 514 nsew
rlabel metal2 s 14736 11297 14736 11297 4 gnd
port 514 nsew
rlabel metal2 s 13488 12640 13488 12640 4 gnd
port 514 nsew
rlabel metal2 s 14736 11850 14736 11850 4 gnd
port 514 nsew
rlabel metal2 s 14736 10033 14736 10033 4 gnd
port 514 nsew
rlabel metal2 s 13968 11850 13968 11850 4 gnd
port 514 nsew
rlabel metal2 s 14736 10270 14736 10270 4 gnd
port 514 nsew
rlabel metal2 s 13968 10033 13968 10033 4 gnd
port 514 nsew
rlabel metal2 s 13488 11850 13488 11850 4 gnd
port 514 nsew
rlabel metal2 s 12720 11613 12720 11613 4 gnd
port 514 nsew
rlabel metal2 s 13488 10507 13488 10507 4 gnd
port 514 nsew
rlabel metal2 s 13488 12403 13488 12403 4 gnd
port 514 nsew
rlabel metal2 s 13488 11297 13488 11297 4 gnd
port 514 nsew
rlabel metal2 s 13488 10823 13488 10823 4 gnd
port 514 nsew
rlabel metal2 s 12720 10823 12720 10823 4 gnd
port 514 nsew
rlabel metal2 s 12720 10033 12720 10033 4 gnd
port 514 nsew
rlabel metal2 s 13968 11297 13968 11297 4 gnd
port 514 nsew
rlabel metal2 s 13488 10270 13488 10270 4 gnd
port 514 nsew
rlabel metal2 s 13488 11613 13488 11613 4 gnd
port 514 nsew
rlabel metal2 s 14736 10823 14736 10823 4 gnd
port 514 nsew
rlabel metal2 s 12720 11297 12720 11297 4 gnd
port 514 nsew
rlabel metal2 s 12720 11060 12720 11060 4 gnd
port 514 nsew
rlabel metal2 s 12720 12087 12720 12087 4 gnd
port 514 nsew
rlabel metal2 s 13968 10270 13968 10270 4 gnd
port 514 nsew
rlabel metal2 s 14736 9717 14736 9717 4 gnd
port 514 nsew
rlabel metal2 s 13488 10033 13488 10033 4 gnd
port 514 nsew
rlabel metal2 s 14736 11613 14736 11613 4 gnd
port 514 nsew
rlabel metal2 s 13968 12087 13968 12087 4 gnd
port 514 nsew
rlabel metal2 s 14736 12087 14736 12087 4 gnd
port 514 nsew
rlabel metal2 s 12720 9717 12720 9717 4 gnd
port 514 nsew
rlabel metal2 s 12720 12403 12720 12403 4 gnd
port 514 nsew
rlabel metal2 s 14736 12640 14736 12640 4 gnd
port 514 nsew
rlabel metal2 s 14736 12403 14736 12403 4 gnd
port 514 nsew
rlabel metal2 s 13968 12403 13968 12403 4 gnd
port 514 nsew
rlabel metal2 s 13488 11060 13488 11060 4 gnd
port 514 nsew
rlabel metal2 s 13968 11613 13968 11613 4 gnd
port 514 nsew
rlabel metal2 s 13968 12640 13968 12640 4 gnd
port 514 nsew
rlabel metal2 s 13488 12087 13488 12087 4 gnd
port 514 nsew
rlabel metal2 s 12720 12640 12720 12640 4 gnd
port 514 nsew
rlabel metal2 s 13968 10507 13968 10507 4 gnd
port 514 nsew
rlabel metal2 s 14736 10507 14736 10507 4 gnd
port 514 nsew
rlabel metal2 s 12720 11850 12720 11850 4 gnd
port 514 nsew
rlabel metal2 s 13968 9717 13968 9717 4 gnd
port 514 nsew
rlabel metal2 s 13968 10823 13968 10823 4 gnd
port 514 nsew
rlabel metal2 s 14736 11060 14736 11060 4 gnd
port 514 nsew
rlabel metal2 s 13488 9717 13488 9717 4 gnd
port 514 nsew
rlabel metal2 s 12720 10507 12720 10507 4 gnd
port 514 nsew
rlabel metal2 s 12240 11850 12240 11850 4 gnd
port 514 nsew
rlabel metal2 s 11472 10033 11472 10033 4 gnd
port 514 nsew
rlabel metal2 s 11472 12087 11472 12087 4 gnd
port 514 nsew
rlabel metal2 s 10224 11297 10224 11297 4 gnd
port 514 nsew
rlabel metal2 s 10992 10270 10992 10270 4 gnd
port 514 nsew
rlabel metal2 s 11472 9717 11472 9717 4 gnd
port 514 nsew
rlabel metal2 s 10992 9717 10992 9717 4 gnd
port 514 nsew
rlabel metal2 s 11472 12403 11472 12403 4 gnd
port 514 nsew
rlabel metal2 s 10992 12640 10992 12640 4 gnd
port 514 nsew
rlabel metal2 s 10224 11613 10224 11613 4 gnd
port 514 nsew
rlabel metal2 s 12240 11613 12240 11613 4 gnd
port 514 nsew
rlabel metal2 s 10224 12640 10224 12640 4 gnd
port 514 nsew
rlabel metal2 s 11472 11613 11472 11613 4 gnd
port 514 nsew
rlabel metal2 s 10992 12087 10992 12087 4 gnd
port 514 nsew
rlabel metal2 s 12240 10507 12240 10507 4 gnd
port 514 nsew
rlabel metal2 s 10992 11613 10992 11613 4 gnd
port 514 nsew
rlabel metal2 s 10992 10823 10992 10823 4 gnd
port 514 nsew
rlabel metal2 s 11472 10507 11472 10507 4 gnd
port 514 nsew
rlabel metal2 s 12240 12640 12240 12640 4 gnd
port 514 nsew
rlabel metal2 s 10224 11850 10224 11850 4 gnd
port 514 nsew
rlabel metal2 s 12240 11060 12240 11060 4 gnd
port 514 nsew
rlabel metal2 s 11472 10270 11472 10270 4 gnd
port 514 nsew
rlabel metal2 s 12240 10033 12240 10033 4 gnd
port 514 nsew
rlabel metal2 s 11472 11297 11472 11297 4 gnd
port 514 nsew
rlabel metal2 s 10224 9717 10224 9717 4 gnd
port 514 nsew
rlabel metal2 s 10992 11297 10992 11297 4 gnd
port 514 nsew
rlabel metal2 s 10224 10507 10224 10507 4 gnd
port 514 nsew
rlabel metal2 s 10224 12087 10224 12087 4 gnd
port 514 nsew
rlabel metal2 s 12240 9717 12240 9717 4 gnd
port 514 nsew
rlabel metal2 s 10992 11850 10992 11850 4 gnd
port 514 nsew
rlabel metal2 s 10224 11060 10224 11060 4 gnd
port 514 nsew
rlabel metal2 s 10224 10823 10224 10823 4 gnd
port 514 nsew
rlabel metal2 s 12240 12087 12240 12087 4 gnd
port 514 nsew
rlabel metal2 s 10224 10270 10224 10270 4 gnd
port 514 nsew
rlabel metal2 s 12240 12403 12240 12403 4 gnd
port 514 nsew
rlabel metal2 s 12240 11297 12240 11297 4 gnd
port 514 nsew
rlabel metal2 s 10992 10033 10992 10033 4 gnd
port 514 nsew
rlabel metal2 s 12240 10823 12240 10823 4 gnd
port 514 nsew
rlabel metal2 s 10224 10033 10224 10033 4 gnd
port 514 nsew
rlabel metal2 s 11472 12640 11472 12640 4 gnd
port 514 nsew
rlabel metal2 s 11472 11850 11472 11850 4 gnd
port 514 nsew
rlabel metal2 s 10992 10507 10992 10507 4 gnd
port 514 nsew
rlabel metal2 s 10992 11060 10992 11060 4 gnd
port 514 nsew
rlabel metal2 s 10992 12403 10992 12403 4 gnd
port 514 nsew
rlabel metal2 s 12240 10270 12240 10270 4 gnd
port 514 nsew
rlabel metal2 s 11472 11060 11472 11060 4 gnd
port 514 nsew
rlabel metal2 s 11472 10823 11472 10823 4 gnd
port 514 nsew
rlabel metal2 s 10224 12403 10224 12403 4 gnd
port 514 nsew
rlabel metal2 s 10992 9243 10992 9243 4 gnd
port 514 nsew
rlabel metal2 s 11472 8690 11472 8690 4 gnd
port 514 nsew
rlabel metal2 s 12240 8927 12240 8927 4 gnd
port 514 nsew
rlabel metal2 s 12240 9243 12240 9243 4 gnd
port 514 nsew
rlabel metal2 s 11472 6873 11472 6873 4 gnd
port 514 nsew
rlabel metal2 s 10992 9480 10992 9480 4 gnd
port 514 nsew
rlabel metal2 s 12240 9480 12240 9480 4 gnd
port 514 nsew
rlabel metal2 s 10224 9243 10224 9243 4 gnd
port 514 nsew
rlabel metal2 s 12240 7110 12240 7110 4 gnd
port 514 nsew
rlabel metal2 s 10224 8137 10224 8137 4 gnd
port 514 nsew
rlabel metal2 s 11472 8137 11472 8137 4 gnd
port 514 nsew
rlabel metal2 s 10992 6557 10992 6557 4 gnd
port 514 nsew
rlabel metal2 s 11472 7900 11472 7900 4 gnd
port 514 nsew
rlabel metal2 s 10992 8927 10992 8927 4 gnd
port 514 nsew
rlabel metal2 s 10992 8690 10992 8690 4 gnd
port 514 nsew
rlabel metal2 s 11472 7663 11472 7663 4 gnd
port 514 nsew
rlabel metal2 s 12240 7663 12240 7663 4 gnd
port 514 nsew
rlabel metal2 s 11472 9243 11472 9243 4 gnd
port 514 nsew
rlabel metal2 s 12240 8690 12240 8690 4 gnd
port 514 nsew
rlabel metal2 s 10992 7900 10992 7900 4 gnd
port 514 nsew
rlabel metal2 s 12240 8137 12240 8137 4 gnd
port 514 nsew
rlabel metal2 s 12240 6873 12240 6873 4 gnd
port 514 nsew
rlabel metal2 s 10224 8927 10224 8927 4 gnd
port 514 nsew
rlabel metal2 s 10224 6873 10224 6873 4 gnd
port 514 nsew
rlabel metal2 s 10224 8453 10224 8453 4 gnd
port 514 nsew
rlabel metal2 s 12240 7900 12240 7900 4 gnd
port 514 nsew
rlabel metal2 s 10224 9480 10224 9480 4 gnd
port 514 nsew
rlabel metal2 s 10224 7347 10224 7347 4 gnd
port 514 nsew
rlabel metal2 s 11472 8453 11472 8453 4 gnd
port 514 nsew
rlabel metal2 s 10224 7663 10224 7663 4 gnd
port 514 nsew
rlabel metal2 s 10992 7347 10992 7347 4 gnd
port 514 nsew
rlabel metal2 s 12240 7347 12240 7347 4 gnd
port 514 nsew
rlabel metal2 s 10992 8453 10992 8453 4 gnd
port 514 nsew
rlabel metal2 s 10992 8137 10992 8137 4 gnd
port 514 nsew
rlabel metal2 s 12240 8453 12240 8453 4 gnd
port 514 nsew
rlabel metal2 s 11472 6557 11472 6557 4 gnd
port 514 nsew
rlabel metal2 s 10992 7663 10992 7663 4 gnd
port 514 nsew
rlabel metal2 s 12240 6557 12240 6557 4 gnd
port 514 nsew
rlabel metal2 s 10224 7900 10224 7900 4 gnd
port 514 nsew
rlabel metal2 s 10992 7110 10992 7110 4 gnd
port 514 nsew
rlabel metal2 s 11472 9480 11472 9480 4 gnd
port 514 nsew
rlabel metal2 s 11472 8927 11472 8927 4 gnd
port 514 nsew
rlabel metal2 s 11472 7347 11472 7347 4 gnd
port 514 nsew
rlabel metal2 s 10224 8690 10224 8690 4 gnd
port 514 nsew
rlabel metal2 s 10224 7110 10224 7110 4 gnd
port 514 nsew
rlabel metal2 s 11472 7110 11472 7110 4 gnd
port 514 nsew
rlabel metal2 s 10992 6873 10992 6873 4 gnd
port 514 nsew
rlabel metal2 s 10224 6557 10224 6557 4 gnd
port 514 nsew
rlabel metal2 s 13968 7110 13968 7110 4 gnd
port 514 nsew
rlabel metal2 s 13968 7347 13968 7347 4 gnd
port 514 nsew
rlabel metal2 s 12720 6557 12720 6557 4 gnd
port 514 nsew
rlabel metal2 s 13488 7110 13488 7110 4 gnd
port 514 nsew
rlabel metal2 s 14736 9243 14736 9243 4 gnd
port 514 nsew
rlabel metal2 s 14736 8927 14736 8927 4 gnd
port 514 nsew
rlabel metal2 s 13488 8137 13488 8137 4 gnd
port 514 nsew
rlabel metal2 s 13968 8137 13968 8137 4 gnd
port 514 nsew
rlabel metal2 s 13968 7900 13968 7900 4 gnd
port 514 nsew
rlabel metal2 s 12720 7900 12720 7900 4 gnd
port 514 nsew
rlabel metal2 s 12720 8927 12720 8927 4 gnd
port 514 nsew
rlabel metal2 s 14736 7110 14736 7110 4 gnd
port 514 nsew
rlabel metal2 s 13968 6557 13968 6557 4 gnd
port 514 nsew
rlabel metal2 s 13488 7347 13488 7347 4 gnd
port 514 nsew
rlabel metal2 s 13968 9243 13968 9243 4 gnd
port 514 nsew
rlabel metal2 s 14736 6557 14736 6557 4 gnd
port 514 nsew
rlabel metal2 s 12720 7663 12720 7663 4 gnd
port 514 nsew
rlabel metal2 s 13968 8927 13968 8927 4 gnd
port 514 nsew
rlabel metal2 s 14736 8453 14736 8453 4 gnd
port 514 nsew
rlabel metal2 s 12720 9243 12720 9243 4 gnd
port 514 nsew
rlabel metal2 s 12720 8137 12720 8137 4 gnd
port 514 nsew
rlabel metal2 s 13488 8927 13488 8927 4 gnd
port 514 nsew
rlabel metal2 s 12720 6873 12720 6873 4 gnd
port 514 nsew
rlabel metal2 s 13968 9480 13968 9480 4 gnd
port 514 nsew
rlabel metal2 s 13968 8690 13968 8690 4 gnd
port 514 nsew
rlabel metal2 s 12720 8690 12720 8690 4 gnd
port 514 nsew
rlabel metal2 s 12720 7110 12720 7110 4 gnd
port 514 nsew
rlabel metal2 s 13488 7900 13488 7900 4 gnd
port 514 nsew
rlabel metal2 s 14736 8690 14736 8690 4 gnd
port 514 nsew
rlabel metal2 s 13488 6873 13488 6873 4 gnd
port 514 nsew
rlabel metal2 s 13968 6873 13968 6873 4 gnd
port 514 nsew
rlabel metal2 s 13968 8453 13968 8453 4 gnd
port 514 nsew
rlabel metal2 s 12720 7347 12720 7347 4 gnd
port 514 nsew
rlabel metal2 s 14736 7900 14736 7900 4 gnd
port 514 nsew
rlabel metal2 s 14736 9480 14736 9480 4 gnd
port 514 nsew
rlabel metal2 s 14736 7663 14736 7663 4 gnd
port 514 nsew
rlabel metal2 s 13968 7663 13968 7663 4 gnd
port 514 nsew
rlabel metal2 s 12720 9480 12720 9480 4 gnd
port 514 nsew
rlabel metal2 s 14736 7347 14736 7347 4 gnd
port 514 nsew
rlabel metal2 s 12720 8453 12720 8453 4 gnd
port 514 nsew
rlabel metal2 s 13488 9243 13488 9243 4 gnd
port 514 nsew
rlabel metal2 s 13488 8690 13488 8690 4 gnd
port 514 nsew
rlabel metal2 s 13488 6557 13488 6557 4 gnd
port 514 nsew
rlabel metal2 s 13488 8453 13488 8453 4 gnd
port 514 nsew
rlabel metal2 s 13488 9480 13488 9480 4 gnd
port 514 nsew
rlabel metal2 s 13488 7663 13488 7663 4 gnd
port 514 nsew
rlabel metal2 s 14736 6873 14736 6873 4 gnd
port 514 nsew
rlabel metal2 s 14736 8137 14736 8137 4 gnd
port 514 nsew
rlabel metal2 s 13488 3713 13488 3713 4 gnd
port 514 nsew
rlabel metal2 s 13488 5293 13488 5293 4 gnd
port 514 nsew
rlabel metal2 s 12720 4740 12720 4740 4 gnd
port 514 nsew
rlabel metal2 s 14736 3397 14736 3397 4 gnd
port 514 nsew
rlabel metal2 s 13968 3713 13968 3713 4 gnd
port 514 nsew
rlabel metal2 s 13968 6320 13968 6320 4 gnd
port 514 nsew
rlabel metal2 s 14736 4503 14736 4503 4 gnd
port 514 nsew
rlabel metal2 s 13488 6320 13488 6320 4 gnd
port 514 nsew
rlabel metal2 s 13488 3950 13488 3950 4 gnd
port 514 nsew
rlabel metal2 s 12720 5767 12720 5767 4 gnd
port 514 nsew
rlabel metal2 s 14736 4977 14736 4977 4 gnd
port 514 nsew
rlabel metal2 s 13968 4503 13968 4503 4 gnd
port 514 nsew
rlabel metal2 s 13968 3397 13968 3397 4 gnd
port 514 nsew
rlabel metal2 s 13968 5293 13968 5293 4 gnd
port 514 nsew
rlabel metal2 s 14736 4740 14736 4740 4 gnd
port 514 nsew
rlabel metal2 s 13968 4977 13968 4977 4 gnd
port 514 nsew
rlabel metal2 s 13968 3950 13968 3950 4 gnd
port 514 nsew
rlabel metal2 s 14736 5530 14736 5530 4 gnd
port 514 nsew
rlabel metal2 s 13488 3397 13488 3397 4 gnd
port 514 nsew
rlabel metal2 s 12720 5530 12720 5530 4 gnd
port 514 nsew
rlabel metal2 s 13488 6083 13488 6083 4 gnd
port 514 nsew
rlabel metal2 s 13968 6083 13968 6083 4 gnd
port 514 nsew
rlabel metal2 s 12720 3950 12720 3950 4 gnd
port 514 nsew
rlabel metal2 s 13488 4977 13488 4977 4 gnd
port 514 nsew
rlabel metal2 s 13488 4740 13488 4740 4 gnd
port 514 nsew
rlabel metal2 s 14736 4187 14736 4187 4 gnd
port 514 nsew
rlabel metal2 s 14736 3713 14736 3713 4 gnd
port 514 nsew
rlabel metal2 s 13968 4740 13968 4740 4 gnd
port 514 nsew
rlabel metal2 s 13968 5530 13968 5530 4 gnd
port 514 nsew
rlabel metal2 s 13968 5767 13968 5767 4 gnd
port 514 nsew
rlabel metal2 s 14736 5767 14736 5767 4 gnd
port 514 nsew
rlabel metal2 s 14736 6083 14736 6083 4 gnd
port 514 nsew
rlabel metal2 s 12720 6320 12720 6320 4 gnd
port 514 nsew
rlabel metal2 s 12720 5293 12720 5293 4 gnd
port 514 nsew
rlabel metal2 s 14736 3950 14736 3950 4 gnd
port 514 nsew
rlabel metal2 s 14736 6320 14736 6320 4 gnd
port 514 nsew
rlabel metal2 s 13488 5767 13488 5767 4 gnd
port 514 nsew
rlabel metal2 s 13968 4187 13968 4187 4 gnd
port 514 nsew
rlabel metal2 s 14736 5293 14736 5293 4 gnd
port 514 nsew
rlabel metal2 s 13488 4503 13488 4503 4 gnd
port 514 nsew
rlabel metal2 s 12720 3713 12720 3713 4 gnd
port 514 nsew
rlabel metal2 s 12720 4187 12720 4187 4 gnd
port 514 nsew
rlabel metal2 s 12720 6083 12720 6083 4 gnd
port 514 nsew
rlabel metal2 s 13488 5530 13488 5530 4 gnd
port 514 nsew
rlabel metal2 s 12720 4503 12720 4503 4 gnd
port 514 nsew
rlabel metal2 s 12720 4977 12720 4977 4 gnd
port 514 nsew
rlabel metal2 s 12720 3397 12720 3397 4 gnd
port 514 nsew
rlabel metal2 s 13488 4187 13488 4187 4 gnd
port 514 nsew
rlabel metal2 s 12240 5530 12240 5530 4 gnd
port 514 nsew
rlabel metal2 s 10992 3950 10992 3950 4 gnd
port 514 nsew
rlabel metal2 s 10992 6083 10992 6083 4 gnd
port 514 nsew
rlabel metal2 s 12240 3397 12240 3397 4 gnd
port 514 nsew
rlabel metal2 s 10224 4977 10224 4977 4 gnd
port 514 nsew
rlabel metal2 s 10224 3713 10224 3713 4 gnd
port 514 nsew
rlabel metal2 s 12240 4187 12240 4187 4 gnd
port 514 nsew
rlabel metal2 s 11472 3950 11472 3950 4 gnd
port 514 nsew
rlabel metal2 s 10992 4503 10992 4503 4 gnd
port 514 nsew
rlabel metal2 s 11472 6320 11472 6320 4 gnd
port 514 nsew
rlabel metal2 s 10992 6320 10992 6320 4 gnd
port 514 nsew
rlabel metal2 s 10992 3397 10992 3397 4 gnd
port 514 nsew
rlabel metal2 s 10224 6083 10224 6083 4 gnd
port 514 nsew
rlabel metal2 s 11472 6083 11472 6083 4 gnd
port 514 nsew
rlabel metal2 s 11472 4977 11472 4977 4 gnd
port 514 nsew
rlabel metal2 s 10224 5530 10224 5530 4 gnd
port 514 nsew
rlabel metal2 s 12240 6320 12240 6320 4 gnd
port 514 nsew
rlabel metal2 s 12240 4740 12240 4740 4 gnd
port 514 nsew
rlabel metal2 s 11472 5530 11472 5530 4 gnd
port 514 nsew
rlabel metal2 s 12240 5767 12240 5767 4 gnd
port 514 nsew
rlabel metal2 s 12240 5293 12240 5293 4 gnd
port 514 nsew
rlabel metal2 s 10992 4187 10992 4187 4 gnd
port 514 nsew
rlabel metal2 s 10992 5293 10992 5293 4 gnd
port 514 nsew
rlabel metal2 s 10992 5767 10992 5767 4 gnd
port 514 nsew
rlabel metal2 s 11472 4187 11472 4187 4 gnd
port 514 nsew
rlabel metal2 s 10224 4503 10224 4503 4 gnd
port 514 nsew
rlabel metal2 s 11472 3713 11472 3713 4 gnd
port 514 nsew
rlabel metal2 s 10224 4740 10224 4740 4 gnd
port 514 nsew
rlabel metal2 s 10224 3950 10224 3950 4 gnd
port 514 nsew
rlabel metal2 s 10992 5530 10992 5530 4 gnd
port 514 nsew
rlabel metal2 s 11472 4740 11472 4740 4 gnd
port 514 nsew
rlabel metal2 s 11472 4503 11472 4503 4 gnd
port 514 nsew
rlabel metal2 s 10224 5293 10224 5293 4 gnd
port 514 nsew
rlabel metal2 s 12240 4977 12240 4977 4 gnd
port 514 nsew
rlabel metal2 s 12240 3950 12240 3950 4 gnd
port 514 nsew
rlabel metal2 s 12240 4503 12240 4503 4 gnd
port 514 nsew
rlabel metal2 s 10224 3397 10224 3397 4 gnd
port 514 nsew
rlabel metal2 s 11472 3397 11472 3397 4 gnd
port 514 nsew
rlabel metal2 s 11472 5767 11472 5767 4 gnd
port 514 nsew
rlabel metal2 s 10992 3713 10992 3713 4 gnd
port 514 nsew
rlabel metal2 s 10992 4977 10992 4977 4 gnd
port 514 nsew
rlabel metal2 s 10992 4740 10992 4740 4 gnd
port 514 nsew
rlabel metal2 s 10224 6320 10224 6320 4 gnd
port 514 nsew
rlabel metal2 s 10224 5767 10224 5767 4 gnd
port 514 nsew
rlabel metal2 s 12240 6083 12240 6083 4 gnd
port 514 nsew
rlabel metal2 s 10224 4187 10224 4187 4 gnd
port 514 nsew
rlabel metal2 s 12240 3713 12240 3713 4 gnd
port 514 nsew
rlabel metal2 s 11472 5293 11472 5293 4 gnd
port 514 nsew
rlabel metal2 s 11472 2133 11472 2133 4 gnd
port 514 nsew
rlabel metal2 s 10992 1027 10992 1027 4 gnd
port 514 nsew
rlabel metal2 s 10992 1580 10992 1580 4 gnd
port 514 nsew
rlabel metal2 s 10224 0 10224 0 4 gnd
port 514 nsew
rlabel metal2 s 10224 1817 10224 1817 4 gnd
port 514 nsew
rlabel metal2 s 11472 237 11472 237 4 gnd
port 514 nsew
rlabel metal2 s 11472 1027 11472 1027 4 gnd
port 514 nsew
rlabel metal2 s 10224 1580 10224 1580 4 gnd
port 514 nsew
rlabel metal2 s 10224 790 10224 790 4 gnd
port 514 nsew
rlabel metal2 s 10992 3160 10992 3160 4 gnd
port 514 nsew
rlabel metal2 s 10992 0 10992 0 4 gnd
port 514 nsew
rlabel metal2 s 10224 2133 10224 2133 4 gnd
port 514 nsew
rlabel metal2 s 11472 790 11472 790 4 gnd
port 514 nsew
rlabel metal2 s 12240 1027 12240 1027 4 gnd
port 514 nsew
rlabel metal2 s 10992 2370 10992 2370 4 gnd
port 514 nsew
rlabel metal2 s 12240 2370 12240 2370 4 gnd
port 514 nsew
rlabel metal2 s 10992 1343 10992 1343 4 gnd
port 514 nsew
rlabel metal2 s 11472 2923 11472 2923 4 gnd
port 514 nsew
rlabel metal2 s 12240 237 12240 237 4 gnd
port 514 nsew
rlabel metal2 s 10992 1817 10992 1817 4 gnd
port 514 nsew
rlabel metal2 s 10224 2923 10224 2923 4 gnd
port 514 nsew
rlabel metal2 s 10224 2370 10224 2370 4 gnd
port 514 nsew
rlabel metal2 s 12240 1580 12240 1580 4 gnd
port 514 nsew
rlabel metal2 s 12240 0 12240 0 4 gnd
port 514 nsew
rlabel metal2 s 10224 1343 10224 1343 4 gnd
port 514 nsew
rlabel metal2 s 11472 2607 11472 2607 4 gnd
port 514 nsew
rlabel metal2 s 12240 1343 12240 1343 4 gnd
port 514 nsew
rlabel metal2 s 11472 1817 11472 1817 4 gnd
port 514 nsew
rlabel metal2 s 12240 553 12240 553 4 gnd
port 514 nsew
rlabel metal2 s 11472 0 11472 0 4 gnd
port 514 nsew
rlabel metal2 s 12240 2607 12240 2607 4 gnd
port 514 nsew
rlabel metal2 s 10992 237 10992 237 4 gnd
port 514 nsew
rlabel metal2 s 10992 553 10992 553 4 gnd
port 514 nsew
rlabel metal2 s 12240 1817 12240 1817 4 gnd
port 514 nsew
rlabel metal2 s 11472 3160 11472 3160 4 gnd
port 514 nsew
rlabel metal2 s 12240 2923 12240 2923 4 gnd
port 514 nsew
rlabel metal2 s 10224 3160 10224 3160 4 gnd
port 514 nsew
rlabel metal2 s 11472 553 11472 553 4 gnd
port 514 nsew
rlabel metal2 s 10224 553 10224 553 4 gnd
port 514 nsew
rlabel metal2 s 10992 2923 10992 2923 4 gnd
port 514 nsew
rlabel metal2 s 11472 1580 11472 1580 4 gnd
port 514 nsew
rlabel metal2 s 10992 2607 10992 2607 4 gnd
port 514 nsew
rlabel metal2 s 10224 2607 10224 2607 4 gnd
port 514 nsew
rlabel metal2 s 10224 237 10224 237 4 gnd
port 514 nsew
rlabel metal2 s 10992 790 10992 790 4 gnd
port 514 nsew
rlabel metal2 s 11472 2370 11472 2370 4 gnd
port 514 nsew
rlabel metal2 s 12240 3160 12240 3160 4 gnd
port 514 nsew
rlabel metal2 s 12240 790 12240 790 4 gnd
port 514 nsew
rlabel metal2 s 11472 1343 11472 1343 4 gnd
port 514 nsew
rlabel metal2 s 10992 2133 10992 2133 4 gnd
port 514 nsew
rlabel metal2 s 12240 2133 12240 2133 4 gnd
port 514 nsew
rlabel metal2 s 10224 1027 10224 1027 4 gnd
port 514 nsew
rlabel metal2 s 14736 2923 14736 2923 4 gnd
port 514 nsew
rlabel metal2 s 12720 3160 12720 3160 4 gnd
port 514 nsew
rlabel metal2 s 13488 2370 13488 2370 4 gnd
port 514 nsew
rlabel metal2 s 13968 2607 13968 2607 4 gnd
port 514 nsew
rlabel metal2 s 12720 237 12720 237 4 gnd
port 514 nsew
rlabel metal2 s 13968 237 13968 237 4 gnd
port 514 nsew
rlabel metal2 s 14736 2607 14736 2607 4 gnd
port 514 nsew
rlabel metal2 s 13968 2133 13968 2133 4 gnd
port 514 nsew
rlabel metal2 s 13488 2133 13488 2133 4 gnd
port 514 nsew
rlabel metal2 s 13968 3160 13968 3160 4 gnd
port 514 nsew
rlabel metal2 s 14736 1343 14736 1343 4 gnd
port 514 nsew
rlabel metal2 s 13968 1027 13968 1027 4 gnd
port 514 nsew
rlabel metal2 s 13488 1580 13488 1580 4 gnd
port 514 nsew
rlabel metal2 s 13968 2370 13968 2370 4 gnd
port 514 nsew
rlabel metal2 s 14736 0 14736 0 4 gnd
port 514 nsew
rlabel metal2 s 13968 1343 13968 1343 4 gnd
port 514 nsew
rlabel metal2 s 12720 1817 12720 1817 4 gnd
port 514 nsew
rlabel metal2 s 12720 0 12720 0 4 gnd
port 514 nsew
rlabel metal2 s 13488 1343 13488 1343 4 gnd
port 514 nsew
rlabel metal2 s 14736 1580 14736 1580 4 gnd
port 514 nsew
rlabel metal2 s 12720 2133 12720 2133 4 gnd
port 514 nsew
rlabel metal2 s 13488 0 13488 0 4 gnd
port 514 nsew
rlabel metal2 s 13968 553 13968 553 4 gnd
port 514 nsew
rlabel metal2 s 14736 2133 14736 2133 4 gnd
port 514 nsew
rlabel metal2 s 13488 790 13488 790 4 gnd
port 514 nsew
rlabel metal2 s 13968 2923 13968 2923 4 gnd
port 514 nsew
rlabel metal2 s 14736 1817 14736 1817 4 gnd
port 514 nsew
rlabel metal2 s 13488 3160 13488 3160 4 gnd
port 514 nsew
rlabel metal2 s 12720 1343 12720 1343 4 gnd
port 514 nsew
rlabel metal2 s 12720 1027 12720 1027 4 gnd
port 514 nsew
rlabel metal2 s 13968 1817 13968 1817 4 gnd
port 514 nsew
rlabel metal2 s 13488 553 13488 553 4 gnd
port 514 nsew
rlabel metal2 s 13488 1817 13488 1817 4 gnd
port 514 nsew
rlabel metal2 s 13488 2607 13488 2607 4 gnd
port 514 nsew
rlabel metal2 s 12720 790 12720 790 4 gnd
port 514 nsew
rlabel metal2 s 13488 2923 13488 2923 4 gnd
port 514 nsew
rlabel metal2 s 12720 2370 12720 2370 4 gnd
port 514 nsew
rlabel metal2 s 13968 790 13968 790 4 gnd
port 514 nsew
rlabel metal2 s 14736 2370 14736 2370 4 gnd
port 514 nsew
rlabel metal2 s 14736 1027 14736 1027 4 gnd
port 514 nsew
rlabel metal2 s 14736 790 14736 790 4 gnd
port 514 nsew
rlabel metal2 s 12720 553 12720 553 4 gnd
port 514 nsew
rlabel metal2 s 13968 0 13968 0 4 gnd
port 514 nsew
rlabel metal2 s 14736 553 14736 553 4 gnd
port 514 nsew
rlabel metal2 s 12720 1580 12720 1580 4 gnd
port 514 nsew
rlabel metal2 s 13488 237 13488 237 4 gnd
port 514 nsew
rlabel metal2 s 13488 1027 13488 1027 4 gnd
port 514 nsew
rlabel metal2 s 14736 237 14736 237 4 gnd
port 514 nsew
rlabel metal2 s 14736 3160 14736 3160 4 gnd
port 514 nsew
rlabel metal2 s 12720 2923 12720 2923 4 gnd
port 514 nsew
rlabel metal2 s 12720 2607 12720 2607 4 gnd
port 514 nsew
rlabel metal2 s 13968 1580 13968 1580 4 gnd
port 514 nsew
rlabel metal2 s 19728 5530 19728 5530 4 gnd
port 514 nsew
rlabel metal2 s 17712 5530 17712 5530 4 gnd
port 514 nsew
rlabel metal2 s 18960 5293 18960 5293 4 gnd
port 514 nsew
rlabel metal2 s 17712 4740 17712 4740 4 gnd
port 514 nsew
rlabel metal2 s 18960 4977 18960 4977 4 gnd
port 514 nsew
rlabel metal2 s 19968 3287 19968 3287 4 wl1_8
port 274 nsew
rlabel metal2 s 19728 4187 19728 4187 4 gnd
port 514 nsew
rlabel metal2 s 18480 5530 18480 5530 4 gnd
port 514 nsew
rlabel metal2 s 18960 5530 18960 5530 4 gnd
port 514 nsew
rlabel metal2 s 19968 5657 19968 5657 4 wl1_14
port 286 nsew
rlabel metal2 s 18480 5767 18480 5767 4 gnd
port 514 nsew
rlabel metal2 s 19968 3603 19968 3603 4 wl0_9
port 275 nsew
rlabel metal2 s 18960 4503 18960 4503 4 gnd
port 514 nsew
rlabel metal2 s 17712 5767 17712 5767 4 gnd
port 514 nsew
rlabel metal2 s 19968 5403 19968 5403 4 wl1_13
port 284 nsew
rlabel metal2 s 19968 5183 19968 5183 4 wl0_13
port 283 nsew
rlabel metal2 s 17712 6083 17712 6083 4 gnd
port 514 nsew
rlabel metal2 s 18960 4187 18960 4187 4 gnd
port 514 nsew
rlabel metal2 s 17712 3950 17712 3950 4 gnd
port 514 nsew
rlabel metal2 s 18480 6083 18480 6083 4 gnd
port 514 nsew
rlabel metal2 s 18960 3397 18960 3397 4 gnd
port 514 nsew
rlabel metal2 s 18960 6083 18960 6083 4 gnd
port 514 nsew
rlabel metal2 s 18480 4740 18480 4740 4 gnd
port 514 nsew
rlabel metal2 s 18480 4977 18480 4977 4 gnd
port 514 nsew
rlabel metal2 s 19728 4977 19728 4977 4 gnd
port 514 nsew
rlabel metal2 s 18480 6320 18480 6320 4 gnd
port 514 nsew
rlabel metal2 s 17712 6320 17712 6320 4 gnd
port 514 nsew
rlabel metal2 s 19728 4740 19728 4740 4 gnd
port 514 nsew
rlabel metal2 s 18960 5767 18960 5767 4 gnd
port 514 nsew
rlabel metal2 s 18960 4740 18960 4740 4 gnd
port 514 nsew
rlabel metal2 s 19968 3507 19968 3507 4 wl0_8
port 273 nsew
rlabel metal2 s 19968 4297 19968 4297 4 wl0_10
port 277 nsew
rlabel metal2 s 19728 5293 19728 5293 4 gnd
port 514 nsew
rlabel metal2 s 18480 5293 18480 5293 4 gnd
port 514 nsew
rlabel metal2 s 17712 4977 17712 4977 4 gnd
port 514 nsew
rlabel metal2 s 18480 3950 18480 3950 4 gnd
port 514 nsew
rlabel metal2 s 19968 5087 19968 5087 4 wl0_12
port 281 nsew
rlabel metal2 s 19968 4077 19968 4077 4 wl1_10
port 278 nsew
rlabel metal2 s 18960 6320 18960 6320 4 gnd
port 514 nsew
rlabel metal2 s 19968 4393 19968 4393 4 wl0_11
port 279 nsew
rlabel metal2 s 17712 3397 17712 3397 4 gnd
port 514 nsew
rlabel metal2 s 19728 4503 19728 4503 4 gnd
port 514 nsew
rlabel metal2 s 19728 3397 19728 3397 4 gnd
port 514 nsew
rlabel metal2 s 19728 6083 19728 6083 4 gnd
port 514 nsew
rlabel metal2 s 18480 4187 18480 4187 4 gnd
port 514 nsew
rlabel metal2 s 17712 4503 17712 4503 4 gnd
port 514 nsew
rlabel metal2 s 19728 6320 19728 6320 4 gnd
port 514 nsew
rlabel metal2 s 19728 5767 19728 5767 4 gnd
port 514 nsew
rlabel metal2 s 19728 3713 19728 3713 4 gnd
port 514 nsew
rlabel metal2 s 19968 4613 19968 4613 4 wl1_11
port 280 nsew
rlabel metal2 s 17712 5293 17712 5293 4 gnd
port 514 nsew
rlabel metal2 s 18480 3713 18480 3713 4 gnd
port 514 nsew
rlabel metal2 s 18480 4503 18480 4503 4 gnd
port 514 nsew
rlabel metal2 s 18960 3713 18960 3713 4 gnd
port 514 nsew
rlabel metal2 s 17712 3713 17712 3713 4 gnd
port 514 nsew
rlabel metal2 s 18480 3397 18480 3397 4 gnd
port 514 nsew
rlabel metal2 s 19968 6193 19968 6193 4 wl1_15
port 288 nsew
rlabel metal2 s 19968 5877 19968 5877 4 wl0_14
port 285 nsew
rlabel metal2 s 17712 4187 17712 4187 4 gnd
port 514 nsew
rlabel metal2 s 18960 3950 18960 3950 4 gnd
port 514 nsew
rlabel metal2 s 19968 4867 19968 4867 4 wl1_12
port 282 nsew
rlabel metal2 s 19968 3823 19968 3823 4 wl1_9
port 276 nsew
rlabel metal2 s 19968 5973 19968 5973 4 wl0_15
port 287 nsew
rlabel metal2 s 19728 3950 19728 3950 4 gnd
port 514 nsew
rlabel metal2 s 16464 6083 16464 6083 4 gnd
port 514 nsew
rlabel metal2 s 15984 3397 15984 3397 4 gnd
port 514 nsew
rlabel metal2 s 15984 5293 15984 5293 4 gnd
port 514 nsew
rlabel metal2 s 15216 3397 15216 3397 4 gnd
port 514 nsew
rlabel metal2 s 17232 4740 17232 4740 4 gnd
port 514 nsew
rlabel metal2 s 15216 3950 15216 3950 4 gnd
port 514 nsew
rlabel metal2 s 16464 4740 16464 4740 4 gnd
port 514 nsew
rlabel metal2 s 17232 5767 17232 5767 4 gnd
port 514 nsew
rlabel metal2 s 17232 4977 17232 4977 4 gnd
port 514 nsew
rlabel metal2 s 16464 5767 16464 5767 4 gnd
port 514 nsew
rlabel metal2 s 16464 5293 16464 5293 4 gnd
port 514 nsew
rlabel metal2 s 15216 6083 15216 6083 4 gnd
port 514 nsew
rlabel metal2 s 15984 4977 15984 4977 4 gnd
port 514 nsew
rlabel metal2 s 16464 3713 16464 3713 4 gnd
port 514 nsew
rlabel metal2 s 15216 5767 15216 5767 4 gnd
port 514 nsew
rlabel metal2 s 15216 4187 15216 4187 4 gnd
port 514 nsew
rlabel metal2 s 15984 5530 15984 5530 4 gnd
port 514 nsew
rlabel metal2 s 17232 6083 17232 6083 4 gnd
port 514 nsew
rlabel metal2 s 16464 4503 16464 4503 4 gnd
port 514 nsew
rlabel metal2 s 17232 4503 17232 4503 4 gnd
port 514 nsew
rlabel metal2 s 15216 4503 15216 4503 4 gnd
port 514 nsew
rlabel metal2 s 17232 6320 17232 6320 4 gnd
port 514 nsew
rlabel metal2 s 16464 3950 16464 3950 4 gnd
port 514 nsew
rlabel metal2 s 15216 3713 15216 3713 4 gnd
port 514 nsew
rlabel metal2 s 15216 6320 15216 6320 4 gnd
port 514 nsew
rlabel metal2 s 15216 4740 15216 4740 4 gnd
port 514 nsew
rlabel metal2 s 16464 6320 16464 6320 4 gnd
port 514 nsew
rlabel metal2 s 15984 4503 15984 4503 4 gnd
port 514 nsew
rlabel metal2 s 16464 5530 16464 5530 4 gnd
port 514 nsew
rlabel metal2 s 16464 3397 16464 3397 4 gnd
port 514 nsew
rlabel metal2 s 15216 4977 15216 4977 4 gnd
port 514 nsew
rlabel metal2 s 15984 4740 15984 4740 4 gnd
port 514 nsew
rlabel metal2 s 15984 3713 15984 3713 4 gnd
port 514 nsew
rlabel metal2 s 17232 3950 17232 3950 4 gnd
port 514 nsew
rlabel metal2 s 17232 5530 17232 5530 4 gnd
port 514 nsew
rlabel metal2 s 16464 4977 16464 4977 4 gnd
port 514 nsew
rlabel metal2 s 15984 6083 15984 6083 4 gnd
port 514 nsew
rlabel metal2 s 15984 5767 15984 5767 4 gnd
port 514 nsew
rlabel metal2 s 17232 4187 17232 4187 4 gnd
port 514 nsew
rlabel metal2 s 15984 4187 15984 4187 4 gnd
port 514 nsew
rlabel metal2 s 15216 5293 15216 5293 4 gnd
port 514 nsew
rlabel metal2 s 15984 6320 15984 6320 4 gnd
port 514 nsew
rlabel metal2 s 17232 3397 17232 3397 4 gnd
port 514 nsew
rlabel metal2 s 16464 4187 16464 4187 4 gnd
port 514 nsew
rlabel metal2 s 17232 3713 17232 3713 4 gnd
port 514 nsew
rlabel metal2 s 17232 5293 17232 5293 4 gnd
port 514 nsew
rlabel metal2 s 15216 5530 15216 5530 4 gnd
port 514 nsew
rlabel metal2 s 15984 3950 15984 3950 4 gnd
port 514 nsew
rlabel metal2 s 16464 2607 16464 2607 4 gnd
port 514 nsew
rlabel metal2 s 16464 1817 16464 1817 4 gnd
port 514 nsew
rlabel metal2 s 15984 2607 15984 2607 4 gnd
port 514 nsew
rlabel metal2 s 16464 553 16464 553 4 gnd
port 514 nsew
rlabel metal2 s 15984 790 15984 790 4 gnd
port 514 nsew
rlabel metal2 s 15216 790 15216 790 4 gnd
port 514 nsew
rlabel metal2 s 17232 1343 17232 1343 4 gnd
port 514 nsew
rlabel metal2 s 16464 2133 16464 2133 4 gnd
port 514 nsew
rlabel metal2 s 17232 1027 17232 1027 4 gnd
port 514 nsew
rlabel metal2 s 15984 1027 15984 1027 4 gnd
port 514 nsew
rlabel metal2 s 15984 237 15984 237 4 gnd
port 514 nsew
rlabel metal2 s 17232 1580 17232 1580 4 gnd
port 514 nsew
rlabel metal2 s 16464 1580 16464 1580 4 gnd
port 514 nsew
rlabel metal2 s 15216 2607 15216 2607 4 gnd
port 514 nsew
rlabel metal2 s 15984 1817 15984 1817 4 gnd
port 514 nsew
rlabel metal2 s 16464 237 16464 237 4 gnd
port 514 nsew
rlabel metal2 s 17232 2370 17232 2370 4 gnd
port 514 nsew
rlabel metal2 s 15216 553 15216 553 4 gnd
port 514 nsew
rlabel metal2 s 15984 2370 15984 2370 4 gnd
port 514 nsew
rlabel metal2 s 15216 3160 15216 3160 4 gnd
port 514 nsew
rlabel metal2 s 15984 553 15984 553 4 gnd
port 514 nsew
rlabel metal2 s 17232 790 17232 790 4 gnd
port 514 nsew
rlabel metal2 s 15216 237 15216 237 4 gnd
port 514 nsew
rlabel metal2 s 17232 553 17232 553 4 gnd
port 514 nsew
rlabel metal2 s 16464 2923 16464 2923 4 gnd
port 514 nsew
rlabel metal2 s 17232 0 17232 0 4 gnd
port 514 nsew
rlabel metal2 s 15216 2923 15216 2923 4 gnd
port 514 nsew
rlabel metal2 s 15216 2370 15216 2370 4 gnd
port 514 nsew
rlabel metal2 s 17232 237 17232 237 4 gnd
port 514 nsew
rlabel metal2 s 16464 2370 16464 2370 4 gnd
port 514 nsew
rlabel metal2 s 17232 2607 17232 2607 4 gnd
port 514 nsew
rlabel metal2 s 15984 1343 15984 1343 4 gnd
port 514 nsew
rlabel metal2 s 15984 0 15984 0 4 gnd
port 514 nsew
rlabel metal2 s 16464 1343 16464 1343 4 gnd
port 514 nsew
rlabel metal2 s 16464 1027 16464 1027 4 gnd
port 514 nsew
rlabel metal2 s 16464 3160 16464 3160 4 gnd
port 514 nsew
rlabel metal2 s 15216 1027 15216 1027 4 gnd
port 514 nsew
rlabel metal2 s 15984 2923 15984 2923 4 gnd
port 514 nsew
rlabel metal2 s 15984 3160 15984 3160 4 gnd
port 514 nsew
rlabel metal2 s 17232 2923 17232 2923 4 gnd
port 514 nsew
rlabel metal2 s 17232 2133 17232 2133 4 gnd
port 514 nsew
rlabel metal2 s 15216 2133 15216 2133 4 gnd
port 514 nsew
rlabel metal2 s 15216 1343 15216 1343 4 gnd
port 514 nsew
rlabel metal2 s 15216 1580 15216 1580 4 gnd
port 514 nsew
rlabel metal2 s 15984 2133 15984 2133 4 gnd
port 514 nsew
rlabel metal2 s 16464 790 16464 790 4 gnd
port 514 nsew
rlabel metal2 s 17232 3160 17232 3160 4 gnd
port 514 nsew
rlabel metal2 s 17232 1817 17232 1817 4 gnd
port 514 nsew
rlabel metal2 s 15984 1580 15984 1580 4 gnd
port 514 nsew
rlabel metal2 s 15216 0 15216 0 4 gnd
port 514 nsew
rlabel metal2 s 16464 0 16464 0 4 gnd
port 514 nsew
rlabel metal2 s 15216 1817 15216 1817 4 gnd
port 514 nsew
rlabel metal2 s 19728 2923 19728 2923 4 gnd
port 514 nsew
rlabel metal2 s 18480 790 18480 790 4 gnd
port 514 nsew
rlabel metal2 s 18960 553 18960 553 4 gnd
port 514 nsew
rlabel metal2 s 18480 3160 18480 3160 4 gnd
port 514 nsew
rlabel metal2 s 18960 790 18960 790 4 gnd
port 514 nsew
rlabel metal2 s 18480 0 18480 0 4 gnd
port 514 nsew
rlabel metal2 s 19968 2813 19968 2813 4 wl0_7
port 271 nsew
rlabel metal2 s 18480 1580 18480 1580 4 gnd
port 514 nsew
rlabel metal2 s 17712 1580 17712 1580 4 gnd
port 514 nsew
rlabel metal2 s 17712 1343 17712 1343 4 gnd
port 514 nsew
rlabel metal2 s 17712 2923 17712 2923 4 gnd
port 514 nsew
rlabel metal2 s 18960 2370 18960 2370 4 gnd
port 514 nsew
rlabel metal2 s 19968 127 19968 127 4 wl1_0
port 258 nsew
rlabel metal2 s 18480 553 18480 553 4 gnd
port 514 nsew
rlabel metal2 s 17712 2370 17712 2370 4 gnd
port 514 nsew
rlabel metal2 s 18960 2607 18960 2607 4 gnd
port 514 nsew
rlabel metal2 s 19968 1927 19968 1927 4 wl0_4
port 265 nsew
rlabel metal2 s 18480 2133 18480 2133 4 gnd
port 514 nsew
rlabel metal2 s 18960 3160 18960 3160 4 gnd
port 514 nsew
rlabel metal2 s 18960 2133 18960 2133 4 gnd
port 514 nsew
rlabel metal2 s 17712 553 17712 553 4 gnd
port 514 nsew
rlabel metal2 s 17712 2133 17712 2133 4 gnd
port 514 nsew
rlabel metal2 s 19728 1580 19728 1580 4 gnd
port 514 nsew
rlabel metal2 s 18960 237 18960 237 4 gnd
port 514 nsew
rlabel metal2 s 18480 237 18480 237 4 gnd
port 514 nsew
rlabel metal2 s 17712 1817 17712 1817 4 gnd
port 514 nsew
rlabel metal2 s 19968 663 19968 663 4 wl1_1
port 260 nsew
rlabel metal2 s 19728 237 19728 237 4 gnd
port 514 nsew
rlabel metal2 s 19968 347 19968 347 4 wl0_0
port 257 nsew
rlabel metal2 s 19968 1137 19968 1137 4 wl0_2
port 261 nsew
rlabel metal2 s 19968 2243 19968 2243 4 wl1_5
port 268 nsew
rlabel metal2 s 18960 2923 18960 2923 4 gnd
port 514 nsew
rlabel metal2 s 19728 1343 19728 1343 4 gnd
port 514 nsew
rlabel metal2 s 18480 1817 18480 1817 4 gnd
port 514 nsew
rlabel metal2 s 19728 553 19728 553 4 gnd
port 514 nsew
rlabel metal2 s 18960 1817 18960 1817 4 gnd
port 514 nsew
rlabel metal2 s 19968 917 19968 917 4 wl1_2
port 262 nsew
rlabel metal2 s 19968 1707 19968 1707 4 wl1_4
port 266 nsew
rlabel metal2 s 17712 790 17712 790 4 gnd
port 514 nsew
rlabel metal2 s 19728 1817 19728 1817 4 gnd
port 514 nsew
rlabel metal2 s 17712 0 17712 0 4 gnd
port 514 nsew
rlabel metal2 s 17712 1027 17712 1027 4 gnd
port 514 nsew
rlabel metal2 s 18480 2923 18480 2923 4 gnd
port 514 nsew
rlabel metal2 s 18480 1343 18480 1343 4 gnd
port 514 nsew
rlabel metal2 s 19728 790 19728 790 4 gnd
port 514 nsew
rlabel metal2 s 19728 2370 19728 2370 4 gnd
port 514 nsew
rlabel metal2 s 19968 2497 19968 2497 4 wl1_6
port 270 nsew
rlabel metal2 s 19728 3160 19728 3160 4 gnd
port 514 nsew
rlabel metal2 s 19968 1453 19968 1453 4 wl1_3
port 264 nsew
rlabel metal2 s 18960 1580 18960 1580 4 gnd
port 514 nsew
rlabel metal2 s 18480 2607 18480 2607 4 gnd
port 514 nsew
rlabel metal2 s 19968 1233 19968 1233 4 wl0_3
port 263 nsew
rlabel metal2 s 19728 0 19728 0 4 gnd
port 514 nsew
rlabel metal2 s 17712 237 17712 237 4 gnd
port 514 nsew
rlabel metal2 s 19968 3033 19968 3033 4 wl1_7
port 272 nsew
rlabel metal2 s 19968 2023 19968 2023 4 wl0_5
port 267 nsew
rlabel metal2 s 19968 2717 19968 2717 4 wl0_6
port 269 nsew
rlabel metal2 s 19728 2607 19728 2607 4 gnd
port 514 nsew
rlabel metal2 s 17712 3160 17712 3160 4 gnd
port 514 nsew
rlabel metal2 s 19728 2133 19728 2133 4 gnd
port 514 nsew
rlabel metal2 s 19728 1027 19728 1027 4 gnd
port 514 nsew
rlabel metal2 s 18480 1027 18480 1027 4 gnd
port 514 nsew
rlabel metal2 s 18960 1027 18960 1027 4 gnd
port 514 nsew
rlabel metal2 s 17712 2607 17712 2607 4 gnd
port 514 nsew
rlabel metal2 s 18480 2370 18480 2370 4 gnd
port 514 nsew
rlabel metal2 s 18960 0 18960 0 4 gnd
port 514 nsew
rlabel metal2 s 19968 443 19968 443 4 wl0_1
port 259 nsew
rlabel metal2 s 18960 1343 18960 1343 4 gnd
port 514 nsew
rlabel metal2 s 38928 22910 38928 22910 4 gnd
port 514 nsew
rlabel metal2 s 38448 24253 38448 24253 4 gnd
port 514 nsew
rlabel metal2 s 37680 23147 37680 23147 4 gnd
port 514 nsew
rlabel metal2 s 37680 25043 37680 25043 4 gnd
port 514 nsew
rlabel metal2 s 38928 25043 38928 25043 4 gnd
port 514 nsew
rlabel metal2 s 38448 23147 38448 23147 4 gnd
port 514 nsew
rlabel metal2 s 38448 25043 38448 25043 4 gnd
port 514 nsew
rlabel metal2 s 37680 22673 37680 22673 4 gnd
port 514 nsew
rlabel metal2 s 37680 25280 37680 25280 4 gnd
port 514 nsew
rlabel metal2 s 39696 25280 39696 25280 4 gnd
port 514 nsew
rlabel metal2 s 38928 24727 38928 24727 4 gnd
port 514 nsew
rlabel metal2 s 37680 24253 37680 24253 4 gnd
port 514 nsew
rlabel metal2 s 38448 24727 38448 24727 4 gnd
port 514 nsew
rlabel metal2 s 39696 23700 39696 23700 4 gnd
port 514 nsew
rlabel metal2 s 39696 23147 39696 23147 4 gnd
port 514 nsew
rlabel metal2 s 37680 24727 37680 24727 4 gnd
port 514 nsew
rlabel metal2 s 38448 22910 38448 22910 4 gnd
port 514 nsew
rlabel metal2 s 37680 22357 37680 22357 4 gnd
port 514 nsew
rlabel metal2 s 38928 22357 38928 22357 4 gnd
port 514 nsew
rlabel metal2 s 39696 24490 39696 24490 4 gnd
port 514 nsew
rlabel metal2 s 39696 23937 39696 23937 4 gnd
port 514 nsew
rlabel metal2 s 38928 23937 38928 23937 4 gnd
port 514 nsew
rlabel metal2 s 38928 23700 38928 23700 4 gnd
port 514 nsew
rlabel metal2 s 39696 22357 39696 22357 4 gnd
port 514 nsew
rlabel metal2 s 38448 25280 38448 25280 4 gnd
port 514 nsew
rlabel metal2 s 38928 24490 38928 24490 4 gnd
port 514 nsew
rlabel metal2 s 39696 24253 39696 24253 4 gnd
port 514 nsew
rlabel metal2 s 39696 23463 39696 23463 4 gnd
port 514 nsew
rlabel metal2 s 39696 24727 39696 24727 4 gnd
port 514 nsew
rlabel metal2 s 38928 23463 38928 23463 4 gnd
port 514 nsew
rlabel metal2 s 37680 22910 37680 22910 4 gnd
port 514 nsew
rlabel metal2 s 37680 23463 37680 23463 4 gnd
port 514 nsew
rlabel metal2 s 37680 24490 37680 24490 4 gnd
port 514 nsew
rlabel metal2 s 38448 23937 38448 23937 4 gnd
port 514 nsew
rlabel metal2 s 38448 23700 38448 23700 4 gnd
port 514 nsew
rlabel metal2 s 38448 22673 38448 22673 4 gnd
port 514 nsew
rlabel metal2 s 38448 22357 38448 22357 4 gnd
port 514 nsew
rlabel metal2 s 38928 25280 38928 25280 4 gnd
port 514 nsew
rlabel metal2 s 38448 23463 38448 23463 4 gnd
port 514 nsew
rlabel metal2 s 38928 22673 38928 22673 4 gnd
port 514 nsew
rlabel metal2 s 39696 25043 39696 25043 4 gnd
port 514 nsew
rlabel metal2 s 38928 24253 38928 24253 4 gnd
port 514 nsew
rlabel metal2 s 37680 23700 37680 23700 4 gnd
port 514 nsew
rlabel metal2 s 39696 22910 39696 22910 4 gnd
port 514 nsew
rlabel metal2 s 38448 24490 38448 24490 4 gnd
port 514 nsew
rlabel metal2 s 37680 23937 37680 23937 4 gnd
port 514 nsew
rlabel metal2 s 39696 22673 39696 22673 4 gnd
port 514 nsew
rlabel metal2 s 38928 23147 38928 23147 4 gnd
port 514 nsew
rlabel metal2 s 37200 24253 37200 24253 4 gnd
port 514 nsew
rlabel metal2 s 36432 22357 36432 22357 4 gnd
port 514 nsew
rlabel metal2 s 35184 25043 35184 25043 4 gnd
port 514 nsew
rlabel metal2 s 35952 25280 35952 25280 4 gnd
port 514 nsew
rlabel metal2 s 35952 24253 35952 24253 4 gnd
port 514 nsew
rlabel metal2 s 37200 22673 37200 22673 4 gnd
port 514 nsew
rlabel metal2 s 35184 23937 35184 23937 4 gnd
port 514 nsew
rlabel metal2 s 35952 23147 35952 23147 4 gnd
port 514 nsew
rlabel metal2 s 35952 22357 35952 22357 4 gnd
port 514 nsew
rlabel metal2 s 37200 23463 37200 23463 4 gnd
port 514 nsew
rlabel metal2 s 35952 25043 35952 25043 4 gnd
port 514 nsew
rlabel metal2 s 36432 25043 36432 25043 4 gnd
port 514 nsew
rlabel metal2 s 36432 23147 36432 23147 4 gnd
port 514 nsew
rlabel metal2 s 36432 24490 36432 24490 4 gnd
port 514 nsew
rlabel metal2 s 35184 23700 35184 23700 4 gnd
port 514 nsew
rlabel metal2 s 35184 22910 35184 22910 4 gnd
port 514 nsew
rlabel metal2 s 35952 24727 35952 24727 4 gnd
port 514 nsew
rlabel metal2 s 37200 24727 37200 24727 4 gnd
port 514 nsew
rlabel metal2 s 35184 24727 35184 24727 4 gnd
port 514 nsew
rlabel metal2 s 37200 25280 37200 25280 4 gnd
port 514 nsew
rlabel metal2 s 36432 24727 36432 24727 4 gnd
port 514 nsew
rlabel metal2 s 36432 25280 36432 25280 4 gnd
port 514 nsew
rlabel metal2 s 37200 23937 37200 23937 4 gnd
port 514 nsew
rlabel metal2 s 36432 23937 36432 23937 4 gnd
port 514 nsew
rlabel metal2 s 35184 25280 35184 25280 4 gnd
port 514 nsew
rlabel metal2 s 35952 22673 35952 22673 4 gnd
port 514 nsew
rlabel metal2 s 37200 22357 37200 22357 4 gnd
port 514 nsew
rlabel metal2 s 35184 24490 35184 24490 4 gnd
port 514 nsew
rlabel metal2 s 35184 23463 35184 23463 4 gnd
port 514 nsew
rlabel metal2 s 35952 23700 35952 23700 4 gnd
port 514 nsew
rlabel metal2 s 37200 23147 37200 23147 4 gnd
port 514 nsew
rlabel metal2 s 36432 24253 36432 24253 4 gnd
port 514 nsew
rlabel metal2 s 35952 24490 35952 24490 4 gnd
port 514 nsew
rlabel metal2 s 35952 23463 35952 23463 4 gnd
port 514 nsew
rlabel metal2 s 35184 23147 35184 23147 4 gnd
port 514 nsew
rlabel metal2 s 35184 22357 35184 22357 4 gnd
port 514 nsew
rlabel metal2 s 37200 22910 37200 22910 4 gnd
port 514 nsew
rlabel metal2 s 35952 22910 35952 22910 4 gnd
port 514 nsew
rlabel metal2 s 35952 23937 35952 23937 4 gnd
port 514 nsew
rlabel metal2 s 36432 23463 36432 23463 4 gnd
port 514 nsew
rlabel metal2 s 36432 22673 36432 22673 4 gnd
port 514 nsew
rlabel metal2 s 35184 24253 35184 24253 4 gnd
port 514 nsew
rlabel metal2 s 36432 23700 36432 23700 4 gnd
port 514 nsew
rlabel metal2 s 37200 23700 37200 23700 4 gnd
port 514 nsew
rlabel metal2 s 37200 24490 37200 24490 4 gnd
port 514 nsew
rlabel metal2 s 35184 22673 35184 22673 4 gnd
port 514 nsew
rlabel metal2 s 37200 25043 37200 25043 4 gnd
port 514 nsew
rlabel metal2 s 36432 22910 36432 22910 4 gnd
port 514 nsew
rlabel metal2 s 35184 20540 35184 20540 4 gnd
port 514 nsew
rlabel metal2 s 37200 21330 37200 21330 4 gnd
port 514 nsew
rlabel metal2 s 35184 19513 35184 19513 4 gnd
port 514 nsew
rlabel metal2 s 37200 21093 37200 21093 4 gnd
port 514 nsew
rlabel metal2 s 35184 20777 35184 20777 4 gnd
port 514 nsew
rlabel metal2 s 36432 20303 36432 20303 4 gnd
port 514 nsew
rlabel metal2 s 37200 19513 37200 19513 4 gnd
port 514 nsew
rlabel metal2 s 35184 19197 35184 19197 4 gnd
port 514 nsew
rlabel metal2 s 35184 21883 35184 21883 4 gnd
port 514 nsew
rlabel metal2 s 37200 21567 37200 21567 4 gnd
port 514 nsew
rlabel metal2 s 36432 21330 36432 21330 4 gnd
port 514 nsew
rlabel metal2 s 35952 21883 35952 21883 4 gnd
port 514 nsew
rlabel metal2 s 36432 19197 36432 19197 4 gnd
port 514 nsew
rlabel metal2 s 36432 21567 36432 21567 4 gnd
port 514 nsew
rlabel metal2 s 35184 21567 35184 21567 4 gnd
port 514 nsew
rlabel metal2 s 35184 19750 35184 19750 4 gnd
port 514 nsew
rlabel metal2 s 37200 22120 37200 22120 4 gnd
port 514 nsew
rlabel metal2 s 37200 20777 37200 20777 4 gnd
port 514 nsew
rlabel metal2 s 37200 19750 37200 19750 4 gnd
port 514 nsew
rlabel metal2 s 36432 19987 36432 19987 4 gnd
port 514 nsew
rlabel metal2 s 35952 20540 35952 20540 4 gnd
port 514 nsew
rlabel metal2 s 36432 20540 36432 20540 4 gnd
port 514 nsew
rlabel metal2 s 37200 21883 37200 21883 4 gnd
port 514 nsew
rlabel metal2 s 35952 20303 35952 20303 4 gnd
port 514 nsew
rlabel metal2 s 37200 19987 37200 19987 4 gnd
port 514 nsew
rlabel metal2 s 35952 21567 35952 21567 4 gnd
port 514 nsew
rlabel metal2 s 35184 20303 35184 20303 4 gnd
port 514 nsew
rlabel metal2 s 35184 22120 35184 22120 4 gnd
port 514 nsew
rlabel metal2 s 35952 19987 35952 19987 4 gnd
port 514 nsew
rlabel metal2 s 35952 20777 35952 20777 4 gnd
port 514 nsew
rlabel metal2 s 36432 19513 36432 19513 4 gnd
port 514 nsew
rlabel metal2 s 35952 19750 35952 19750 4 gnd
port 514 nsew
rlabel metal2 s 35952 19197 35952 19197 4 gnd
port 514 nsew
rlabel metal2 s 37200 19197 37200 19197 4 gnd
port 514 nsew
rlabel metal2 s 35952 19513 35952 19513 4 gnd
port 514 nsew
rlabel metal2 s 36432 20777 36432 20777 4 gnd
port 514 nsew
rlabel metal2 s 36432 21093 36432 21093 4 gnd
port 514 nsew
rlabel metal2 s 37200 20303 37200 20303 4 gnd
port 514 nsew
rlabel metal2 s 36432 22120 36432 22120 4 gnd
port 514 nsew
rlabel metal2 s 35952 21093 35952 21093 4 gnd
port 514 nsew
rlabel metal2 s 35184 21330 35184 21330 4 gnd
port 514 nsew
rlabel metal2 s 35952 21330 35952 21330 4 gnd
port 514 nsew
rlabel metal2 s 35184 19987 35184 19987 4 gnd
port 514 nsew
rlabel metal2 s 36432 21883 36432 21883 4 gnd
port 514 nsew
rlabel metal2 s 35952 22120 35952 22120 4 gnd
port 514 nsew
rlabel metal2 s 35184 21093 35184 21093 4 gnd
port 514 nsew
rlabel metal2 s 36432 19750 36432 19750 4 gnd
port 514 nsew
rlabel metal2 s 37200 20540 37200 20540 4 gnd
port 514 nsew
rlabel metal2 s 38928 19197 38928 19197 4 gnd
port 514 nsew
rlabel metal2 s 39696 21883 39696 21883 4 gnd
port 514 nsew
rlabel metal2 s 38928 20777 38928 20777 4 gnd
port 514 nsew
rlabel metal2 s 38928 21093 38928 21093 4 gnd
port 514 nsew
rlabel metal2 s 38448 20303 38448 20303 4 gnd
port 514 nsew
rlabel metal2 s 37680 21567 37680 21567 4 gnd
port 514 nsew
rlabel metal2 s 39696 20540 39696 20540 4 gnd
port 514 nsew
rlabel metal2 s 39696 20777 39696 20777 4 gnd
port 514 nsew
rlabel metal2 s 38928 21330 38928 21330 4 gnd
port 514 nsew
rlabel metal2 s 39696 20303 39696 20303 4 gnd
port 514 nsew
rlabel metal2 s 38448 20777 38448 20777 4 gnd
port 514 nsew
rlabel metal2 s 39696 19750 39696 19750 4 gnd
port 514 nsew
rlabel metal2 s 37680 21330 37680 21330 4 gnd
port 514 nsew
rlabel metal2 s 38448 21093 38448 21093 4 gnd
port 514 nsew
rlabel metal2 s 38448 20540 38448 20540 4 gnd
port 514 nsew
rlabel metal2 s 39696 19197 39696 19197 4 gnd
port 514 nsew
rlabel metal2 s 37680 19987 37680 19987 4 gnd
port 514 nsew
rlabel metal2 s 38928 20303 38928 20303 4 gnd
port 514 nsew
rlabel metal2 s 37680 22120 37680 22120 4 gnd
port 514 nsew
rlabel metal2 s 38448 19987 38448 19987 4 gnd
port 514 nsew
rlabel metal2 s 38448 21330 38448 21330 4 gnd
port 514 nsew
rlabel metal2 s 37680 21093 37680 21093 4 gnd
port 514 nsew
rlabel metal2 s 37680 19197 37680 19197 4 gnd
port 514 nsew
rlabel metal2 s 38928 22120 38928 22120 4 gnd
port 514 nsew
rlabel metal2 s 38448 19513 38448 19513 4 gnd
port 514 nsew
rlabel metal2 s 39696 22120 39696 22120 4 gnd
port 514 nsew
rlabel metal2 s 38928 20540 38928 20540 4 gnd
port 514 nsew
rlabel metal2 s 38928 21567 38928 21567 4 gnd
port 514 nsew
rlabel metal2 s 37680 20777 37680 20777 4 gnd
port 514 nsew
rlabel metal2 s 39696 19987 39696 19987 4 gnd
port 514 nsew
rlabel metal2 s 38448 19750 38448 19750 4 gnd
port 514 nsew
rlabel metal2 s 39696 21093 39696 21093 4 gnd
port 514 nsew
rlabel metal2 s 37680 19513 37680 19513 4 gnd
port 514 nsew
rlabel metal2 s 37680 21883 37680 21883 4 gnd
port 514 nsew
rlabel metal2 s 38448 21883 38448 21883 4 gnd
port 514 nsew
rlabel metal2 s 38448 22120 38448 22120 4 gnd
port 514 nsew
rlabel metal2 s 38448 19197 38448 19197 4 gnd
port 514 nsew
rlabel metal2 s 37680 19750 37680 19750 4 gnd
port 514 nsew
rlabel metal2 s 37680 20540 37680 20540 4 gnd
port 514 nsew
rlabel metal2 s 38928 19513 38928 19513 4 gnd
port 514 nsew
rlabel metal2 s 38448 21567 38448 21567 4 gnd
port 514 nsew
rlabel metal2 s 38928 21883 38928 21883 4 gnd
port 514 nsew
rlabel metal2 s 37680 20303 37680 20303 4 gnd
port 514 nsew
rlabel metal2 s 39696 21567 39696 21567 4 gnd
port 514 nsew
rlabel metal2 s 39696 19513 39696 19513 4 gnd
port 514 nsew
rlabel metal2 s 39696 21330 39696 21330 4 gnd
port 514 nsew
rlabel metal2 s 38928 19750 38928 19750 4 gnd
port 514 nsew
rlabel metal2 s 38928 19987 38928 19987 4 gnd
port 514 nsew
rlabel metal2 s 34704 23147 34704 23147 4 gnd
port 514 nsew
rlabel metal2 s 33936 23147 33936 23147 4 gnd
port 514 nsew
rlabel metal2 s 32688 22357 32688 22357 4 gnd
port 514 nsew
rlabel metal2 s 32688 24727 32688 24727 4 gnd
port 514 nsew
rlabel metal2 s 33936 25280 33936 25280 4 gnd
port 514 nsew
rlabel metal2 s 33936 24253 33936 24253 4 gnd
port 514 nsew
rlabel metal2 s 34704 25280 34704 25280 4 gnd
port 514 nsew
rlabel metal2 s 32688 24490 32688 24490 4 gnd
port 514 nsew
rlabel metal2 s 33936 23937 33936 23937 4 gnd
port 514 nsew
rlabel metal2 s 33936 24727 33936 24727 4 gnd
port 514 nsew
rlabel metal2 s 33456 23463 33456 23463 4 gnd
port 514 nsew
rlabel metal2 s 32688 23147 32688 23147 4 gnd
port 514 nsew
rlabel metal2 s 34704 24253 34704 24253 4 gnd
port 514 nsew
rlabel metal2 s 33936 23700 33936 23700 4 gnd
port 514 nsew
rlabel metal2 s 32688 23937 32688 23937 4 gnd
port 514 nsew
rlabel metal2 s 34704 23463 34704 23463 4 gnd
port 514 nsew
rlabel metal2 s 34704 23937 34704 23937 4 gnd
port 514 nsew
rlabel metal2 s 34704 24727 34704 24727 4 gnd
port 514 nsew
rlabel metal2 s 33936 22673 33936 22673 4 gnd
port 514 nsew
rlabel metal2 s 32688 23700 32688 23700 4 gnd
port 514 nsew
rlabel metal2 s 33456 23937 33456 23937 4 gnd
port 514 nsew
rlabel metal2 s 33456 24727 33456 24727 4 gnd
port 514 nsew
rlabel metal2 s 34704 22910 34704 22910 4 gnd
port 514 nsew
rlabel metal2 s 33456 23147 33456 23147 4 gnd
port 514 nsew
rlabel metal2 s 33456 23700 33456 23700 4 gnd
port 514 nsew
rlabel metal2 s 32688 24253 32688 24253 4 gnd
port 514 nsew
rlabel metal2 s 34704 24490 34704 24490 4 gnd
port 514 nsew
rlabel metal2 s 33456 25043 33456 25043 4 gnd
port 514 nsew
rlabel metal2 s 34704 25043 34704 25043 4 gnd
port 514 nsew
rlabel metal2 s 34704 22357 34704 22357 4 gnd
port 514 nsew
rlabel metal2 s 32688 22910 32688 22910 4 gnd
port 514 nsew
rlabel metal2 s 33456 25280 33456 25280 4 gnd
port 514 nsew
rlabel metal2 s 33936 23463 33936 23463 4 gnd
port 514 nsew
rlabel metal2 s 32688 23463 32688 23463 4 gnd
port 514 nsew
rlabel metal2 s 33456 22357 33456 22357 4 gnd
port 514 nsew
rlabel metal2 s 33456 22673 33456 22673 4 gnd
port 514 nsew
rlabel metal2 s 34704 23700 34704 23700 4 gnd
port 514 nsew
rlabel metal2 s 33936 22910 33936 22910 4 gnd
port 514 nsew
rlabel metal2 s 33936 22357 33936 22357 4 gnd
port 514 nsew
rlabel metal2 s 32688 22673 32688 22673 4 gnd
port 514 nsew
rlabel metal2 s 32688 25280 32688 25280 4 gnd
port 514 nsew
rlabel metal2 s 33456 22910 33456 22910 4 gnd
port 514 nsew
rlabel metal2 s 33936 24490 33936 24490 4 gnd
port 514 nsew
rlabel metal2 s 34704 22673 34704 22673 4 gnd
port 514 nsew
rlabel metal2 s 32688 25043 32688 25043 4 gnd
port 514 nsew
rlabel metal2 s 33936 25043 33936 25043 4 gnd
port 514 nsew
rlabel metal2 s 33456 24253 33456 24253 4 gnd
port 514 nsew
rlabel metal2 s 33456 24490 33456 24490 4 gnd
port 514 nsew
rlabel metal2 s 32208 23463 32208 23463 4 gnd
port 514 nsew
rlabel metal2 s 30192 22910 30192 22910 4 gnd
port 514 nsew
rlabel metal2 s 30960 22357 30960 22357 4 gnd
port 514 nsew
rlabel metal2 s 30192 23937 30192 23937 4 gnd
port 514 nsew
rlabel metal2 s 31440 24253 31440 24253 4 gnd
port 514 nsew
rlabel metal2 s 32208 24253 32208 24253 4 gnd
port 514 nsew
rlabel metal2 s 31440 24490 31440 24490 4 gnd
port 514 nsew
rlabel metal2 s 30960 23700 30960 23700 4 gnd
port 514 nsew
rlabel metal2 s 30192 24490 30192 24490 4 gnd
port 514 nsew
rlabel metal2 s 30960 25043 30960 25043 4 gnd
port 514 nsew
rlabel metal2 s 32208 22673 32208 22673 4 gnd
port 514 nsew
rlabel metal2 s 32208 23937 32208 23937 4 gnd
port 514 nsew
rlabel metal2 s 32208 23700 32208 23700 4 gnd
port 514 nsew
rlabel metal2 s 30960 24253 30960 24253 4 gnd
port 514 nsew
rlabel metal2 s 32208 25043 32208 25043 4 gnd
port 514 nsew
rlabel metal2 s 32208 22910 32208 22910 4 gnd
port 514 nsew
rlabel metal2 s 31440 25280 31440 25280 4 gnd
port 514 nsew
rlabel metal2 s 31440 23700 31440 23700 4 gnd
port 514 nsew
rlabel metal2 s 30960 25280 30960 25280 4 gnd
port 514 nsew
rlabel metal2 s 30960 24490 30960 24490 4 gnd
port 514 nsew
rlabel metal2 s 30960 22673 30960 22673 4 gnd
port 514 nsew
rlabel metal2 s 32208 24490 32208 24490 4 gnd
port 514 nsew
rlabel metal2 s 32208 22357 32208 22357 4 gnd
port 514 nsew
rlabel metal2 s 30192 22357 30192 22357 4 gnd
port 514 nsew
rlabel metal2 s 30192 25280 30192 25280 4 gnd
port 514 nsew
rlabel metal2 s 31440 22673 31440 22673 4 gnd
port 514 nsew
rlabel metal2 s 30192 25043 30192 25043 4 gnd
port 514 nsew
rlabel metal2 s 30192 22673 30192 22673 4 gnd
port 514 nsew
rlabel metal2 s 30192 23700 30192 23700 4 gnd
port 514 nsew
rlabel metal2 s 31440 24727 31440 24727 4 gnd
port 514 nsew
rlabel metal2 s 31440 25043 31440 25043 4 gnd
port 514 nsew
rlabel metal2 s 31440 23937 31440 23937 4 gnd
port 514 nsew
rlabel metal2 s 30960 23147 30960 23147 4 gnd
port 514 nsew
rlabel metal2 s 31440 22357 31440 22357 4 gnd
port 514 nsew
rlabel metal2 s 32208 25280 32208 25280 4 gnd
port 514 nsew
rlabel metal2 s 32208 24727 32208 24727 4 gnd
port 514 nsew
rlabel metal2 s 30192 23147 30192 23147 4 gnd
port 514 nsew
rlabel metal2 s 31440 22910 31440 22910 4 gnd
port 514 nsew
rlabel metal2 s 30960 23463 30960 23463 4 gnd
port 514 nsew
rlabel metal2 s 30960 23937 30960 23937 4 gnd
port 514 nsew
rlabel metal2 s 32208 23147 32208 23147 4 gnd
port 514 nsew
rlabel metal2 s 30192 24253 30192 24253 4 gnd
port 514 nsew
rlabel metal2 s 31440 23147 31440 23147 4 gnd
port 514 nsew
rlabel metal2 s 30960 22910 30960 22910 4 gnd
port 514 nsew
rlabel metal2 s 30960 24727 30960 24727 4 gnd
port 514 nsew
rlabel metal2 s 31440 23463 31440 23463 4 gnd
port 514 nsew
rlabel metal2 s 30192 24727 30192 24727 4 gnd
port 514 nsew
rlabel metal2 s 30192 23463 30192 23463 4 gnd
port 514 nsew
rlabel metal2 s 30192 21883 30192 21883 4 gnd
port 514 nsew
rlabel metal2 s 30960 20777 30960 20777 4 gnd
port 514 nsew
rlabel metal2 s 30192 19197 30192 19197 4 gnd
port 514 nsew
rlabel metal2 s 30960 21883 30960 21883 4 gnd
port 514 nsew
rlabel metal2 s 30960 21330 30960 21330 4 gnd
port 514 nsew
rlabel metal2 s 30192 22120 30192 22120 4 gnd
port 514 nsew
rlabel metal2 s 31440 21883 31440 21883 4 gnd
port 514 nsew
rlabel metal2 s 30192 20777 30192 20777 4 gnd
port 514 nsew
rlabel metal2 s 32208 19197 32208 19197 4 gnd
port 514 nsew
rlabel metal2 s 30960 21093 30960 21093 4 gnd
port 514 nsew
rlabel metal2 s 32208 19750 32208 19750 4 gnd
port 514 nsew
rlabel metal2 s 31440 19197 31440 19197 4 gnd
port 514 nsew
rlabel metal2 s 31440 21330 31440 21330 4 gnd
port 514 nsew
rlabel metal2 s 31440 19750 31440 19750 4 gnd
port 514 nsew
rlabel metal2 s 30192 20303 30192 20303 4 gnd
port 514 nsew
rlabel metal2 s 30192 19513 30192 19513 4 gnd
port 514 nsew
rlabel metal2 s 30960 19513 30960 19513 4 gnd
port 514 nsew
rlabel metal2 s 32208 21883 32208 21883 4 gnd
port 514 nsew
rlabel metal2 s 30960 20540 30960 20540 4 gnd
port 514 nsew
rlabel metal2 s 32208 20303 32208 20303 4 gnd
port 514 nsew
rlabel metal2 s 30192 21093 30192 21093 4 gnd
port 514 nsew
rlabel metal2 s 32208 19513 32208 19513 4 gnd
port 514 nsew
rlabel metal2 s 31440 21093 31440 21093 4 gnd
port 514 nsew
rlabel metal2 s 30192 19750 30192 19750 4 gnd
port 514 nsew
rlabel metal2 s 30960 19197 30960 19197 4 gnd
port 514 nsew
rlabel metal2 s 30960 19750 30960 19750 4 gnd
port 514 nsew
rlabel metal2 s 32208 21093 32208 21093 4 gnd
port 514 nsew
rlabel metal2 s 31440 19987 31440 19987 4 gnd
port 514 nsew
rlabel metal2 s 32208 20777 32208 20777 4 gnd
port 514 nsew
rlabel metal2 s 30960 19987 30960 19987 4 gnd
port 514 nsew
rlabel metal2 s 30960 20303 30960 20303 4 gnd
port 514 nsew
rlabel metal2 s 30192 19987 30192 19987 4 gnd
port 514 nsew
rlabel metal2 s 31440 21567 31440 21567 4 gnd
port 514 nsew
rlabel metal2 s 31440 20777 31440 20777 4 gnd
port 514 nsew
rlabel metal2 s 31440 22120 31440 22120 4 gnd
port 514 nsew
rlabel metal2 s 30192 21330 30192 21330 4 gnd
port 514 nsew
rlabel metal2 s 31440 20303 31440 20303 4 gnd
port 514 nsew
rlabel metal2 s 32208 21330 32208 21330 4 gnd
port 514 nsew
rlabel metal2 s 31440 19513 31440 19513 4 gnd
port 514 nsew
rlabel metal2 s 30960 22120 30960 22120 4 gnd
port 514 nsew
rlabel metal2 s 32208 20540 32208 20540 4 gnd
port 514 nsew
rlabel metal2 s 30960 21567 30960 21567 4 gnd
port 514 nsew
rlabel metal2 s 32208 21567 32208 21567 4 gnd
port 514 nsew
rlabel metal2 s 30192 20540 30192 20540 4 gnd
port 514 nsew
rlabel metal2 s 30192 21567 30192 21567 4 gnd
port 514 nsew
rlabel metal2 s 32208 22120 32208 22120 4 gnd
port 514 nsew
rlabel metal2 s 32208 19987 32208 19987 4 gnd
port 514 nsew
rlabel metal2 s 31440 20540 31440 20540 4 gnd
port 514 nsew
rlabel metal2 s 33456 21093 33456 21093 4 gnd
port 514 nsew
rlabel metal2 s 34704 21330 34704 21330 4 gnd
port 514 nsew
rlabel metal2 s 32688 21330 32688 21330 4 gnd
port 514 nsew
rlabel metal2 s 34704 22120 34704 22120 4 gnd
port 514 nsew
rlabel metal2 s 32688 21883 32688 21883 4 gnd
port 514 nsew
rlabel metal2 s 33456 21567 33456 21567 4 gnd
port 514 nsew
rlabel metal2 s 33936 19750 33936 19750 4 gnd
port 514 nsew
rlabel metal2 s 34704 21883 34704 21883 4 gnd
port 514 nsew
rlabel metal2 s 33456 21883 33456 21883 4 gnd
port 514 nsew
rlabel metal2 s 33456 19750 33456 19750 4 gnd
port 514 nsew
rlabel metal2 s 33936 21567 33936 21567 4 gnd
port 514 nsew
rlabel metal2 s 33936 21093 33936 21093 4 gnd
port 514 nsew
rlabel metal2 s 32688 20303 32688 20303 4 gnd
port 514 nsew
rlabel metal2 s 33936 19987 33936 19987 4 gnd
port 514 nsew
rlabel metal2 s 33456 19987 33456 19987 4 gnd
port 514 nsew
rlabel metal2 s 34704 21567 34704 21567 4 gnd
port 514 nsew
rlabel metal2 s 33456 22120 33456 22120 4 gnd
port 514 nsew
rlabel metal2 s 33936 22120 33936 22120 4 gnd
port 514 nsew
rlabel metal2 s 33456 21330 33456 21330 4 gnd
port 514 nsew
rlabel metal2 s 33456 19197 33456 19197 4 gnd
port 514 nsew
rlabel metal2 s 34704 19197 34704 19197 4 gnd
port 514 nsew
rlabel metal2 s 32688 19197 32688 19197 4 gnd
port 514 nsew
rlabel metal2 s 33456 19513 33456 19513 4 gnd
port 514 nsew
rlabel metal2 s 32688 22120 32688 22120 4 gnd
port 514 nsew
rlabel metal2 s 33456 20540 33456 20540 4 gnd
port 514 nsew
rlabel metal2 s 34704 21093 34704 21093 4 gnd
port 514 nsew
rlabel metal2 s 33936 20540 33936 20540 4 gnd
port 514 nsew
rlabel metal2 s 33936 20303 33936 20303 4 gnd
port 514 nsew
rlabel metal2 s 32688 20540 32688 20540 4 gnd
port 514 nsew
rlabel metal2 s 33936 20777 33936 20777 4 gnd
port 514 nsew
rlabel metal2 s 34704 20777 34704 20777 4 gnd
port 514 nsew
rlabel metal2 s 32688 19750 32688 19750 4 gnd
port 514 nsew
rlabel metal2 s 32688 20777 32688 20777 4 gnd
port 514 nsew
rlabel metal2 s 32688 21567 32688 21567 4 gnd
port 514 nsew
rlabel metal2 s 33936 21883 33936 21883 4 gnd
port 514 nsew
rlabel metal2 s 32688 19513 32688 19513 4 gnd
port 514 nsew
rlabel metal2 s 33456 20303 33456 20303 4 gnd
port 514 nsew
rlabel metal2 s 34704 20540 34704 20540 4 gnd
port 514 nsew
rlabel metal2 s 34704 19987 34704 19987 4 gnd
port 514 nsew
rlabel metal2 s 34704 19513 34704 19513 4 gnd
port 514 nsew
rlabel metal2 s 33936 19513 33936 19513 4 gnd
port 514 nsew
rlabel metal2 s 32688 19987 32688 19987 4 gnd
port 514 nsew
rlabel metal2 s 34704 19750 34704 19750 4 gnd
port 514 nsew
rlabel metal2 s 33936 19197 33936 19197 4 gnd
port 514 nsew
rlabel metal2 s 33936 21330 33936 21330 4 gnd
port 514 nsew
rlabel metal2 s 33456 20777 33456 20777 4 gnd
port 514 nsew
rlabel metal2 s 32688 21093 32688 21093 4 gnd
port 514 nsew
rlabel metal2 s 34704 20303 34704 20303 4 gnd
port 514 nsew
rlabel metal2 s 33936 16037 33936 16037 4 gnd
port 514 nsew
rlabel metal2 s 32688 18723 32688 18723 4 gnd
port 514 nsew
rlabel metal2 s 33456 16037 33456 16037 4 gnd
port 514 nsew
rlabel metal2 s 32688 16827 32688 16827 4 gnd
port 514 nsew
rlabel metal2 s 33456 17143 33456 17143 4 gnd
port 514 nsew
rlabel metal2 s 33936 18407 33936 18407 4 gnd
port 514 nsew
rlabel metal2 s 33456 17380 33456 17380 4 gnd
port 514 nsew
rlabel metal2 s 33456 17617 33456 17617 4 gnd
port 514 nsew
rlabel metal2 s 33456 18723 33456 18723 4 gnd
port 514 nsew
rlabel metal2 s 34704 18960 34704 18960 4 gnd
port 514 nsew
rlabel metal2 s 33936 17380 33936 17380 4 gnd
port 514 nsew
rlabel metal2 s 33456 18170 33456 18170 4 gnd
port 514 nsew
rlabel metal2 s 32688 16590 32688 16590 4 gnd
port 514 nsew
rlabel metal2 s 34704 17617 34704 17617 4 gnd
port 514 nsew
rlabel metal2 s 34704 18723 34704 18723 4 gnd
port 514 nsew
rlabel metal2 s 32688 18960 32688 18960 4 gnd
port 514 nsew
rlabel metal2 s 32688 17933 32688 17933 4 gnd
port 514 nsew
rlabel metal2 s 33936 16590 33936 16590 4 gnd
port 514 nsew
rlabel metal2 s 34704 18407 34704 18407 4 gnd
port 514 nsew
rlabel metal2 s 32688 18407 32688 18407 4 gnd
port 514 nsew
rlabel metal2 s 33936 16827 33936 16827 4 gnd
port 514 nsew
rlabel metal2 s 34704 16590 34704 16590 4 gnd
port 514 nsew
rlabel metal2 s 33456 17933 33456 17933 4 gnd
port 514 nsew
rlabel metal2 s 33456 16590 33456 16590 4 gnd
port 514 nsew
rlabel metal2 s 33936 17143 33936 17143 4 gnd
port 514 nsew
rlabel metal2 s 34704 18170 34704 18170 4 gnd
port 514 nsew
rlabel metal2 s 34704 17380 34704 17380 4 gnd
port 514 nsew
rlabel metal2 s 33936 18170 33936 18170 4 gnd
port 514 nsew
rlabel metal2 s 32688 17617 32688 17617 4 gnd
port 514 nsew
rlabel metal2 s 32688 16037 32688 16037 4 gnd
port 514 nsew
rlabel metal2 s 32688 18170 32688 18170 4 gnd
port 514 nsew
rlabel metal2 s 33456 16353 33456 16353 4 gnd
port 514 nsew
rlabel metal2 s 33936 18960 33936 18960 4 gnd
port 514 nsew
rlabel metal2 s 34704 16353 34704 16353 4 gnd
port 514 nsew
rlabel metal2 s 32688 17143 32688 17143 4 gnd
port 514 nsew
rlabel metal2 s 33936 16353 33936 16353 4 gnd
port 514 nsew
rlabel metal2 s 34704 17933 34704 17933 4 gnd
port 514 nsew
rlabel metal2 s 32688 16353 32688 16353 4 gnd
port 514 nsew
rlabel metal2 s 33936 17933 33936 17933 4 gnd
port 514 nsew
rlabel metal2 s 34704 17143 34704 17143 4 gnd
port 514 nsew
rlabel metal2 s 33456 16827 33456 16827 4 gnd
port 514 nsew
rlabel metal2 s 34704 16037 34704 16037 4 gnd
port 514 nsew
rlabel metal2 s 33936 17617 33936 17617 4 gnd
port 514 nsew
rlabel metal2 s 33456 18407 33456 18407 4 gnd
port 514 nsew
rlabel metal2 s 34704 16827 34704 16827 4 gnd
port 514 nsew
rlabel metal2 s 33456 18960 33456 18960 4 gnd
port 514 nsew
rlabel metal2 s 32688 17380 32688 17380 4 gnd
port 514 nsew
rlabel metal2 s 33936 18723 33936 18723 4 gnd
port 514 nsew
rlabel metal2 s 31440 17380 31440 17380 4 gnd
port 514 nsew
rlabel metal2 s 30192 16353 30192 16353 4 gnd
port 514 nsew
rlabel metal2 s 32208 16037 32208 16037 4 gnd
port 514 nsew
rlabel metal2 s 31440 16590 31440 16590 4 gnd
port 514 nsew
rlabel metal2 s 30960 16590 30960 16590 4 gnd
port 514 nsew
rlabel metal2 s 30192 17143 30192 17143 4 gnd
port 514 nsew
rlabel metal2 s 30192 18407 30192 18407 4 gnd
port 514 nsew
rlabel metal2 s 30192 16827 30192 16827 4 gnd
port 514 nsew
rlabel metal2 s 30192 18723 30192 18723 4 gnd
port 514 nsew
rlabel metal2 s 30960 17933 30960 17933 4 gnd
port 514 nsew
rlabel metal2 s 30192 18960 30192 18960 4 gnd
port 514 nsew
rlabel metal2 s 30960 16037 30960 16037 4 gnd
port 514 nsew
rlabel metal2 s 31440 17143 31440 17143 4 gnd
port 514 nsew
rlabel metal2 s 32208 17933 32208 17933 4 gnd
port 514 nsew
rlabel metal2 s 30960 18723 30960 18723 4 gnd
port 514 nsew
rlabel metal2 s 30192 17933 30192 17933 4 gnd
port 514 nsew
rlabel metal2 s 31440 18960 31440 18960 4 gnd
port 514 nsew
rlabel metal2 s 32208 18723 32208 18723 4 gnd
port 514 nsew
rlabel metal2 s 30192 16037 30192 16037 4 gnd
port 514 nsew
rlabel metal2 s 30960 18170 30960 18170 4 gnd
port 514 nsew
rlabel metal2 s 31440 17617 31440 17617 4 gnd
port 514 nsew
rlabel metal2 s 32208 18960 32208 18960 4 gnd
port 514 nsew
rlabel metal2 s 32208 18407 32208 18407 4 gnd
port 514 nsew
rlabel metal2 s 30960 16353 30960 16353 4 gnd
port 514 nsew
rlabel metal2 s 31440 16353 31440 16353 4 gnd
port 514 nsew
rlabel metal2 s 30192 18170 30192 18170 4 gnd
port 514 nsew
rlabel metal2 s 30960 17617 30960 17617 4 gnd
port 514 nsew
rlabel metal2 s 31440 18170 31440 18170 4 gnd
port 514 nsew
rlabel metal2 s 30960 17143 30960 17143 4 gnd
port 514 nsew
rlabel metal2 s 31440 16037 31440 16037 4 gnd
port 514 nsew
rlabel metal2 s 32208 17143 32208 17143 4 gnd
port 514 nsew
rlabel metal2 s 30960 16827 30960 16827 4 gnd
port 514 nsew
rlabel metal2 s 30960 18960 30960 18960 4 gnd
port 514 nsew
rlabel metal2 s 30192 17617 30192 17617 4 gnd
port 514 nsew
rlabel metal2 s 31440 16827 31440 16827 4 gnd
port 514 nsew
rlabel metal2 s 30960 18407 30960 18407 4 gnd
port 514 nsew
rlabel metal2 s 32208 16353 32208 16353 4 gnd
port 514 nsew
rlabel metal2 s 32208 16827 32208 16827 4 gnd
port 514 nsew
rlabel metal2 s 32208 17617 32208 17617 4 gnd
port 514 nsew
rlabel metal2 s 31440 18407 31440 18407 4 gnd
port 514 nsew
rlabel metal2 s 31440 17933 31440 17933 4 gnd
port 514 nsew
rlabel metal2 s 32208 18170 32208 18170 4 gnd
port 514 nsew
rlabel metal2 s 31440 18723 31440 18723 4 gnd
port 514 nsew
rlabel metal2 s 30192 16590 30192 16590 4 gnd
port 514 nsew
rlabel metal2 s 32208 16590 32208 16590 4 gnd
port 514 nsew
rlabel metal2 s 32208 17380 32208 17380 4 gnd
port 514 nsew
rlabel metal2 s 30192 17380 30192 17380 4 gnd
port 514 nsew
rlabel metal2 s 30960 17380 30960 17380 4 gnd
port 514 nsew
rlabel metal2 s 30192 14457 30192 14457 4 gnd
port 514 nsew
rlabel metal2 s 30960 14220 30960 14220 4 gnd
port 514 nsew
rlabel metal2 s 32208 13667 32208 13667 4 gnd
port 514 nsew
rlabel metal2 s 32208 15247 32208 15247 4 gnd
port 514 nsew
rlabel metal2 s 31440 14457 31440 14457 4 gnd
port 514 nsew
rlabel metal2 s 32208 14220 32208 14220 4 gnd
port 514 nsew
rlabel metal2 s 30192 15563 30192 15563 4 gnd
port 514 nsew
rlabel metal2 s 32208 12877 32208 12877 4 gnd
port 514 nsew
rlabel metal2 s 31440 13430 31440 13430 4 gnd
port 514 nsew
rlabel metal2 s 30192 13983 30192 13983 4 gnd
port 514 nsew
rlabel metal2 s 32208 15010 32208 15010 4 gnd
port 514 nsew
rlabel metal2 s 30960 15800 30960 15800 4 gnd
port 514 nsew
rlabel metal2 s 31440 15563 31440 15563 4 gnd
port 514 nsew
rlabel metal2 s 30960 15247 30960 15247 4 gnd
port 514 nsew
rlabel metal2 s 31440 13193 31440 13193 4 gnd
port 514 nsew
rlabel metal2 s 30192 14220 30192 14220 4 gnd
port 514 nsew
rlabel metal2 s 30960 13430 30960 13430 4 gnd
port 514 nsew
rlabel metal2 s 30192 13430 30192 13430 4 gnd
port 514 nsew
rlabel metal2 s 30192 15010 30192 15010 4 gnd
port 514 nsew
rlabel metal2 s 32208 13983 32208 13983 4 gnd
port 514 nsew
rlabel metal2 s 31440 13667 31440 13667 4 gnd
port 514 nsew
rlabel metal2 s 32208 14773 32208 14773 4 gnd
port 514 nsew
rlabel metal2 s 31440 15010 31440 15010 4 gnd
port 514 nsew
rlabel metal2 s 30960 13667 30960 13667 4 gnd
port 514 nsew
rlabel metal2 s 32208 13430 32208 13430 4 gnd
port 514 nsew
rlabel metal2 s 30192 13667 30192 13667 4 gnd
port 514 nsew
rlabel metal2 s 30192 12877 30192 12877 4 gnd
port 514 nsew
rlabel metal2 s 32208 15800 32208 15800 4 gnd
port 514 nsew
rlabel metal2 s 32208 14457 32208 14457 4 gnd
port 514 nsew
rlabel metal2 s 31440 13983 31440 13983 4 gnd
port 514 nsew
rlabel metal2 s 30960 15010 30960 15010 4 gnd
port 514 nsew
rlabel metal2 s 31440 15800 31440 15800 4 gnd
port 514 nsew
rlabel metal2 s 30192 15800 30192 15800 4 gnd
port 514 nsew
rlabel metal2 s 30192 15247 30192 15247 4 gnd
port 514 nsew
rlabel metal2 s 30192 13193 30192 13193 4 gnd
port 514 nsew
rlabel metal2 s 30960 13193 30960 13193 4 gnd
port 514 nsew
rlabel metal2 s 32208 15563 32208 15563 4 gnd
port 514 nsew
rlabel metal2 s 30960 14773 30960 14773 4 gnd
port 514 nsew
rlabel metal2 s 32208 13193 32208 13193 4 gnd
port 514 nsew
rlabel metal2 s 30192 14773 30192 14773 4 gnd
port 514 nsew
rlabel metal2 s 31440 15247 31440 15247 4 gnd
port 514 nsew
rlabel metal2 s 30960 13983 30960 13983 4 gnd
port 514 nsew
rlabel metal2 s 30960 15563 30960 15563 4 gnd
port 514 nsew
rlabel metal2 s 31440 12877 31440 12877 4 gnd
port 514 nsew
rlabel metal2 s 30960 14457 30960 14457 4 gnd
port 514 nsew
rlabel metal2 s 31440 14773 31440 14773 4 gnd
port 514 nsew
rlabel metal2 s 31440 14220 31440 14220 4 gnd
port 514 nsew
rlabel metal2 s 30960 12877 30960 12877 4 gnd
port 514 nsew
rlabel metal2 s 33456 14773 33456 14773 4 gnd
port 514 nsew
rlabel metal2 s 34704 12877 34704 12877 4 gnd
port 514 nsew
rlabel metal2 s 34704 14457 34704 14457 4 gnd
port 514 nsew
rlabel metal2 s 34704 13667 34704 13667 4 gnd
port 514 nsew
rlabel metal2 s 32688 13430 32688 13430 4 gnd
port 514 nsew
rlabel metal2 s 33456 14220 33456 14220 4 gnd
port 514 nsew
rlabel metal2 s 32688 14773 32688 14773 4 gnd
port 514 nsew
rlabel metal2 s 33936 15247 33936 15247 4 gnd
port 514 nsew
rlabel metal2 s 34704 15800 34704 15800 4 gnd
port 514 nsew
rlabel metal2 s 34704 15563 34704 15563 4 gnd
port 514 nsew
rlabel metal2 s 32688 12877 32688 12877 4 gnd
port 514 nsew
rlabel metal2 s 33936 14773 33936 14773 4 gnd
port 514 nsew
rlabel metal2 s 32688 13667 32688 13667 4 gnd
port 514 nsew
rlabel metal2 s 32688 14457 32688 14457 4 gnd
port 514 nsew
rlabel metal2 s 33936 13983 33936 13983 4 gnd
port 514 nsew
rlabel metal2 s 33456 13983 33456 13983 4 gnd
port 514 nsew
rlabel metal2 s 33456 15247 33456 15247 4 gnd
port 514 nsew
rlabel metal2 s 34704 15247 34704 15247 4 gnd
port 514 nsew
rlabel metal2 s 34704 14220 34704 14220 4 gnd
port 514 nsew
rlabel metal2 s 33936 12877 33936 12877 4 gnd
port 514 nsew
rlabel metal2 s 34704 14773 34704 14773 4 gnd
port 514 nsew
rlabel metal2 s 33456 13430 33456 13430 4 gnd
port 514 nsew
rlabel metal2 s 33456 15800 33456 15800 4 gnd
port 514 nsew
rlabel metal2 s 34704 13193 34704 13193 4 gnd
port 514 nsew
rlabel metal2 s 33456 15563 33456 15563 4 gnd
port 514 nsew
rlabel metal2 s 32688 15247 32688 15247 4 gnd
port 514 nsew
rlabel metal2 s 32688 15800 32688 15800 4 gnd
port 514 nsew
rlabel metal2 s 34704 15010 34704 15010 4 gnd
port 514 nsew
rlabel metal2 s 33456 13667 33456 13667 4 gnd
port 514 nsew
rlabel metal2 s 34704 13983 34704 13983 4 gnd
port 514 nsew
rlabel metal2 s 32688 14220 32688 14220 4 gnd
port 514 nsew
rlabel metal2 s 32688 13193 32688 13193 4 gnd
port 514 nsew
rlabel metal2 s 33936 13430 33936 13430 4 gnd
port 514 nsew
rlabel metal2 s 33936 14457 33936 14457 4 gnd
port 514 nsew
rlabel metal2 s 33456 12877 33456 12877 4 gnd
port 514 nsew
rlabel metal2 s 33936 13193 33936 13193 4 gnd
port 514 nsew
rlabel metal2 s 33936 13667 33936 13667 4 gnd
port 514 nsew
rlabel metal2 s 33456 13193 33456 13193 4 gnd
port 514 nsew
rlabel metal2 s 33456 15010 33456 15010 4 gnd
port 514 nsew
rlabel metal2 s 32688 15010 32688 15010 4 gnd
port 514 nsew
rlabel metal2 s 33936 15563 33936 15563 4 gnd
port 514 nsew
rlabel metal2 s 33456 14457 33456 14457 4 gnd
port 514 nsew
rlabel metal2 s 33936 15800 33936 15800 4 gnd
port 514 nsew
rlabel metal2 s 33936 14220 33936 14220 4 gnd
port 514 nsew
rlabel metal2 s 32688 13983 32688 13983 4 gnd
port 514 nsew
rlabel metal2 s 33936 15010 33936 15010 4 gnd
port 514 nsew
rlabel metal2 s 34704 13430 34704 13430 4 gnd
port 514 nsew
rlabel metal2 s 32688 15563 32688 15563 4 gnd
port 514 nsew
rlabel metal2 s 38448 17933 38448 17933 4 gnd
port 514 nsew
rlabel metal2 s 38928 16037 38928 16037 4 gnd
port 514 nsew
rlabel metal2 s 37680 17143 37680 17143 4 gnd
port 514 nsew
rlabel metal2 s 38448 17380 38448 17380 4 gnd
port 514 nsew
rlabel metal2 s 39696 17617 39696 17617 4 gnd
port 514 nsew
rlabel metal2 s 38928 17933 38928 17933 4 gnd
port 514 nsew
rlabel metal2 s 37680 18723 37680 18723 4 gnd
port 514 nsew
rlabel metal2 s 38448 18960 38448 18960 4 gnd
port 514 nsew
rlabel metal2 s 39696 16590 39696 16590 4 gnd
port 514 nsew
rlabel metal2 s 38928 17617 38928 17617 4 gnd
port 514 nsew
rlabel metal2 s 37680 18960 37680 18960 4 gnd
port 514 nsew
rlabel metal2 s 38928 16590 38928 16590 4 gnd
port 514 nsew
rlabel metal2 s 38448 16590 38448 16590 4 gnd
port 514 nsew
rlabel metal2 s 38448 16037 38448 16037 4 gnd
port 514 nsew
rlabel metal2 s 39696 17143 39696 17143 4 gnd
port 514 nsew
rlabel metal2 s 38448 17143 38448 17143 4 gnd
port 514 nsew
rlabel metal2 s 39696 18170 39696 18170 4 gnd
port 514 nsew
rlabel metal2 s 38928 18407 38928 18407 4 gnd
port 514 nsew
rlabel metal2 s 38928 18170 38928 18170 4 gnd
port 514 nsew
rlabel metal2 s 38448 16827 38448 16827 4 gnd
port 514 nsew
rlabel metal2 s 39696 18407 39696 18407 4 gnd
port 514 nsew
rlabel metal2 s 38928 18723 38928 18723 4 gnd
port 514 nsew
rlabel metal2 s 39696 18723 39696 18723 4 gnd
port 514 nsew
rlabel metal2 s 37680 18170 37680 18170 4 gnd
port 514 nsew
rlabel metal2 s 38448 18170 38448 18170 4 gnd
port 514 nsew
rlabel metal2 s 37680 17380 37680 17380 4 gnd
port 514 nsew
rlabel metal2 s 38448 17617 38448 17617 4 gnd
port 514 nsew
rlabel metal2 s 37680 17933 37680 17933 4 gnd
port 514 nsew
rlabel metal2 s 37680 16037 37680 16037 4 gnd
port 514 nsew
rlabel metal2 s 39696 18960 39696 18960 4 gnd
port 514 nsew
rlabel metal2 s 37680 16827 37680 16827 4 gnd
port 514 nsew
rlabel metal2 s 38928 18960 38928 18960 4 gnd
port 514 nsew
rlabel metal2 s 38448 18407 38448 18407 4 gnd
port 514 nsew
rlabel metal2 s 39696 16037 39696 16037 4 gnd
port 514 nsew
rlabel metal2 s 38928 17380 38928 17380 4 gnd
port 514 nsew
rlabel metal2 s 38928 16353 38928 16353 4 gnd
port 514 nsew
rlabel metal2 s 38928 17143 38928 17143 4 gnd
port 514 nsew
rlabel metal2 s 39696 17380 39696 17380 4 gnd
port 514 nsew
rlabel metal2 s 38448 18723 38448 18723 4 gnd
port 514 nsew
rlabel metal2 s 39696 16827 39696 16827 4 gnd
port 514 nsew
rlabel metal2 s 37680 18407 37680 18407 4 gnd
port 514 nsew
rlabel metal2 s 37680 16353 37680 16353 4 gnd
port 514 nsew
rlabel metal2 s 39696 16353 39696 16353 4 gnd
port 514 nsew
rlabel metal2 s 37680 17617 37680 17617 4 gnd
port 514 nsew
rlabel metal2 s 38448 16353 38448 16353 4 gnd
port 514 nsew
rlabel metal2 s 37680 16590 37680 16590 4 gnd
port 514 nsew
rlabel metal2 s 39696 17933 39696 17933 4 gnd
port 514 nsew
rlabel metal2 s 38928 16827 38928 16827 4 gnd
port 514 nsew
rlabel metal2 s 35952 18170 35952 18170 4 gnd
port 514 nsew
rlabel metal2 s 35184 18407 35184 18407 4 gnd
port 514 nsew
rlabel metal2 s 35952 17933 35952 17933 4 gnd
port 514 nsew
rlabel metal2 s 37200 18407 37200 18407 4 gnd
port 514 nsew
rlabel metal2 s 35952 16590 35952 16590 4 gnd
port 514 nsew
rlabel metal2 s 35184 16827 35184 16827 4 gnd
port 514 nsew
rlabel metal2 s 36432 17617 36432 17617 4 gnd
port 514 nsew
rlabel metal2 s 35952 18407 35952 18407 4 gnd
port 514 nsew
rlabel metal2 s 37200 16827 37200 16827 4 gnd
port 514 nsew
rlabel metal2 s 36432 16353 36432 16353 4 gnd
port 514 nsew
rlabel metal2 s 35952 17617 35952 17617 4 gnd
port 514 nsew
rlabel metal2 s 37200 16037 37200 16037 4 gnd
port 514 nsew
rlabel metal2 s 35952 18960 35952 18960 4 gnd
port 514 nsew
rlabel metal2 s 35184 16037 35184 16037 4 gnd
port 514 nsew
rlabel metal2 s 35952 16037 35952 16037 4 gnd
port 514 nsew
rlabel metal2 s 35184 18170 35184 18170 4 gnd
port 514 nsew
rlabel metal2 s 36432 16827 36432 16827 4 gnd
port 514 nsew
rlabel metal2 s 37200 18960 37200 18960 4 gnd
port 514 nsew
rlabel metal2 s 36432 17933 36432 17933 4 gnd
port 514 nsew
rlabel metal2 s 36432 16037 36432 16037 4 gnd
port 514 nsew
rlabel metal2 s 35952 17143 35952 17143 4 gnd
port 514 nsew
rlabel metal2 s 37200 17617 37200 17617 4 gnd
port 514 nsew
rlabel metal2 s 36432 18170 36432 18170 4 gnd
port 514 nsew
rlabel metal2 s 37200 18723 37200 18723 4 gnd
port 514 nsew
rlabel metal2 s 36432 18723 36432 18723 4 gnd
port 514 nsew
rlabel metal2 s 37200 17143 37200 17143 4 gnd
port 514 nsew
rlabel metal2 s 35184 18723 35184 18723 4 gnd
port 514 nsew
rlabel metal2 s 35184 17933 35184 17933 4 gnd
port 514 nsew
rlabel metal2 s 37200 16590 37200 16590 4 gnd
port 514 nsew
rlabel metal2 s 35184 17380 35184 17380 4 gnd
port 514 nsew
rlabel metal2 s 35952 17380 35952 17380 4 gnd
port 514 nsew
rlabel metal2 s 37200 17933 37200 17933 4 gnd
port 514 nsew
rlabel metal2 s 35184 16353 35184 16353 4 gnd
port 514 nsew
rlabel metal2 s 36432 17143 36432 17143 4 gnd
port 514 nsew
rlabel metal2 s 37200 18170 37200 18170 4 gnd
port 514 nsew
rlabel metal2 s 35952 18723 35952 18723 4 gnd
port 514 nsew
rlabel metal2 s 35952 16353 35952 16353 4 gnd
port 514 nsew
rlabel metal2 s 35184 16590 35184 16590 4 gnd
port 514 nsew
rlabel metal2 s 35184 17617 35184 17617 4 gnd
port 514 nsew
rlabel metal2 s 36432 17380 36432 17380 4 gnd
port 514 nsew
rlabel metal2 s 35184 17143 35184 17143 4 gnd
port 514 nsew
rlabel metal2 s 35184 18960 35184 18960 4 gnd
port 514 nsew
rlabel metal2 s 37200 17380 37200 17380 4 gnd
port 514 nsew
rlabel metal2 s 35952 16827 35952 16827 4 gnd
port 514 nsew
rlabel metal2 s 36432 16590 36432 16590 4 gnd
port 514 nsew
rlabel metal2 s 36432 18960 36432 18960 4 gnd
port 514 nsew
rlabel metal2 s 36432 18407 36432 18407 4 gnd
port 514 nsew
rlabel metal2 s 37200 16353 37200 16353 4 gnd
port 514 nsew
rlabel metal2 s 35952 13430 35952 13430 4 gnd
port 514 nsew
rlabel metal2 s 37200 15010 37200 15010 4 gnd
port 514 nsew
rlabel metal2 s 37200 13430 37200 13430 4 gnd
port 514 nsew
rlabel metal2 s 35952 12877 35952 12877 4 gnd
port 514 nsew
rlabel metal2 s 35184 14457 35184 14457 4 gnd
port 514 nsew
rlabel metal2 s 35184 13430 35184 13430 4 gnd
port 514 nsew
rlabel metal2 s 35184 15010 35184 15010 4 gnd
port 514 nsew
rlabel metal2 s 36432 14457 36432 14457 4 gnd
port 514 nsew
rlabel metal2 s 37200 15247 37200 15247 4 gnd
port 514 nsew
rlabel metal2 s 35184 15247 35184 15247 4 gnd
port 514 nsew
rlabel metal2 s 37200 14773 37200 14773 4 gnd
port 514 nsew
rlabel metal2 s 36432 14220 36432 14220 4 gnd
port 514 nsew
rlabel metal2 s 36432 13667 36432 13667 4 gnd
port 514 nsew
rlabel metal2 s 36432 13983 36432 13983 4 gnd
port 514 nsew
rlabel metal2 s 37200 13983 37200 13983 4 gnd
port 514 nsew
rlabel metal2 s 37200 15800 37200 15800 4 gnd
port 514 nsew
rlabel metal2 s 36432 15247 36432 15247 4 gnd
port 514 nsew
rlabel metal2 s 35952 15800 35952 15800 4 gnd
port 514 nsew
rlabel metal2 s 35184 13667 35184 13667 4 gnd
port 514 nsew
rlabel metal2 s 35952 14457 35952 14457 4 gnd
port 514 nsew
rlabel metal2 s 37200 14220 37200 14220 4 gnd
port 514 nsew
rlabel metal2 s 35184 15563 35184 15563 4 gnd
port 514 nsew
rlabel metal2 s 36432 15010 36432 15010 4 gnd
port 514 nsew
rlabel metal2 s 35952 13193 35952 13193 4 gnd
port 514 nsew
rlabel metal2 s 37200 12877 37200 12877 4 gnd
port 514 nsew
rlabel metal2 s 36432 12877 36432 12877 4 gnd
port 514 nsew
rlabel metal2 s 35952 15247 35952 15247 4 gnd
port 514 nsew
rlabel metal2 s 35184 12877 35184 12877 4 gnd
port 514 nsew
rlabel metal2 s 35184 13193 35184 13193 4 gnd
port 514 nsew
rlabel metal2 s 35184 15800 35184 15800 4 gnd
port 514 nsew
rlabel metal2 s 36432 13430 36432 13430 4 gnd
port 514 nsew
rlabel metal2 s 36432 15800 36432 15800 4 gnd
port 514 nsew
rlabel metal2 s 37200 15563 37200 15563 4 gnd
port 514 nsew
rlabel metal2 s 35952 13983 35952 13983 4 gnd
port 514 nsew
rlabel metal2 s 35184 13983 35184 13983 4 gnd
port 514 nsew
rlabel metal2 s 35952 15563 35952 15563 4 gnd
port 514 nsew
rlabel metal2 s 35952 13667 35952 13667 4 gnd
port 514 nsew
rlabel metal2 s 35952 14220 35952 14220 4 gnd
port 514 nsew
rlabel metal2 s 35952 14773 35952 14773 4 gnd
port 514 nsew
rlabel metal2 s 37200 13193 37200 13193 4 gnd
port 514 nsew
rlabel metal2 s 35184 14220 35184 14220 4 gnd
port 514 nsew
rlabel metal2 s 35184 14773 35184 14773 4 gnd
port 514 nsew
rlabel metal2 s 37200 14457 37200 14457 4 gnd
port 514 nsew
rlabel metal2 s 36432 15563 36432 15563 4 gnd
port 514 nsew
rlabel metal2 s 36432 14773 36432 14773 4 gnd
port 514 nsew
rlabel metal2 s 36432 13193 36432 13193 4 gnd
port 514 nsew
rlabel metal2 s 37200 13667 37200 13667 4 gnd
port 514 nsew
rlabel metal2 s 35952 15010 35952 15010 4 gnd
port 514 nsew
rlabel metal2 s 38928 15800 38928 15800 4 gnd
port 514 nsew
rlabel metal2 s 38928 14773 38928 14773 4 gnd
port 514 nsew
rlabel metal2 s 38448 13983 38448 13983 4 gnd
port 514 nsew
rlabel metal2 s 38448 14457 38448 14457 4 gnd
port 514 nsew
rlabel metal2 s 38448 13193 38448 13193 4 gnd
port 514 nsew
rlabel metal2 s 39696 15010 39696 15010 4 gnd
port 514 nsew
rlabel metal2 s 37680 15800 37680 15800 4 gnd
port 514 nsew
rlabel metal2 s 39696 14220 39696 14220 4 gnd
port 514 nsew
rlabel metal2 s 37680 13430 37680 13430 4 gnd
port 514 nsew
rlabel metal2 s 39696 15563 39696 15563 4 gnd
port 514 nsew
rlabel metal2 s 39696 14773 39696 14773 4 gnd
port 514 nsew
rlabel metal2 s 39696 12877 39696 12877 4 gnd
port 514 nsew
rlabel metal2 s 38928 14220 38928 14220 4 gnd
port 514 nsew
rlabel metal2 s 38448 12877 38448 12877 4 gnd
port 514 nsew
rlabel metal2 s 37680 13193 37680 13193 4 gnd
port 514 nsew
rlabel metal2 s 39696 14457 39696 14457 4 gnd
port 514 nsew
rlabel metal2 s 38448 13430 38448 13430 4 gnd
port 514 nsew
rlabel metal2 s 39696 15247 39696 15247 4 gnd
port 514 nsew
rlabel metal2 s 39696 13667 39696 13667 4 gnd
port 514 nsew
rlabel metal2 s 38928 15247 38928 15247 4 gnd
port 514 nsew
rlabel metal2 s 37680 15563 37680 15563 4 gnd
port 514 nsew
rlabel metal2 s 37680 14220 37680 14220 4 gnd
port 514 nsew
rlabel metal2 s 37680 12877 37680 12877 4 gnd
port 514 nsew
rlabel metal2 s 37680 14457 37680 14457 4 gnd
port 514 nsew
rlabel metal2 s 38928 13193 38928 13193 4 gnd
port 514 nsew
rlabel metal2 s 38448 15247 38448 15247 4 gnd
port 514 nsew
rlabel metal2 s 38928 13983 38928 13983 4 gnd
port 514 nsew
rlabel metal2 s 38448 15800 38448 15800 4 gnd
port 514 nsew
rlabel metal2 s 37680 15010 37680 15010 4 gnd
port 514 nsew
rlabel metal2 s 38928 15010 38928 15010 4 gnd
port 514 nsew
rlabel metal2 s 37680 13667 37680 13667 4 gnd
port 514 nsew
rlabel metal2 s 38448 15010 38448 15010 4 gnd
port 514 nsew
rlabel metal2 s 38928 13430 38928 13430 4 gnd
port 514 nsew
rlabel metal2 s 39696 13983 39696 13983 4 gnd
port 514 nsew
rlabel metal2 s 38928 13667 38928 13667 4 gnd
port 514 nsew
rlabel metal2 s 37680 15247 37680 15247 4 gnd
port 514 nsew
rlabel metal2 s 38448 14220 38448 14220 4 gnd
port 514 nsew
rlabel metal2 s 39696 13430 39696 13430 4 gnd
port 514 nsew
rlabel metal2 s 39696 15800 39696 15800 4 gnd
port 514 nsew
rlabel metal2 s 38448 15563 38448 15563 4 gnd
port 514 nsew
rlabel metal2 s 38928 14457 38928 14457 4 gnd
port 514 nsew
rlabel metal2 s 37680 14773 37680 14773 4 gnd
port 514 nsew
rlabel metal2 s 37680 13983 37680 13983 4 gnd
port 514 nsew
rlabel metal2 s 38448 14773 38448 14773 4 gnd
port 514 nsew
rlabel metal2 s 38448 13667 38448 13667 4 gnd
port 514 nsew
rlabel metal2 s 39696 13193 39696 13193 4 gnd
port 514 nsew
rlabel metal2 s 38928 12877 38928 12877 4 gnd
port 514 nsew
rlabel metal2 s 38928 15563 38928 15563 4 gnd
port 514 nsew
rlabel metal2 s 28944 23147 28944 23147 4 gnd
port 514 nsew
rlabel metal2 s 29712 23147 29712 23147 4 gnd
port 514 nsew
rlabel metal2 s 27696 24490 27696 24490 4 gnd
port 514 nsew
rlabel metal2 s 28944 24727 28944 24727 4 gnd
port 514 nsew
rlabel metal2 s 29712 24727 29712 24727 4 gnd
port 514 nsew
rlabel metal2 s 28464 25043 28464 25043 4 gnd
port 514 nsew
rlabel metal2 s 28944 25280 28944 25280 4 gnd
port 514 nsew
rlabel metal2 s 28464 22357 28464 22357 4 gnd
port 514 nsew
rlabel metal2 s 29712 25043 29712 25043 4 gnd
port 514 nsew
rlabel metal2 s 27696 23937 27696 23937 4 gnd
port 514 nsew
rlabel metal2 s 29712 22357 29712 22357 4 gnd
port 514 nsew
rlabel metal2 s 27696 22357 27696 22357 4 gnd
port 514 nsew
rlabel metal2 s 29712 23463 29712 23463 4 gnd
port 514 nsew
rlabel metal2 s 28464 23147 28464 23147 4 gnd
port 514 nsew
rlabel metal2 s 27696 25043 27696 25043 4 gnd
port 514 nsew
rlabel metal2 s 27696 24253 27696 24253 4 gnd
port 514 nsew
rlabel metal2 s 28944 22357 28944 22357 4 gnd
port 514 nsew
rlabel metal2 s 29712 23937 29712 23937 4 gnd
port 514 nsew
rlabel metal2 s 28464 22910 28464 22910 4 gnd
port 514 nsew
rlabel metal2 s 28464 24490 28464 24490 4 gnd
port 514 nsew
rlabel metal2 s 28464 23937 28464 23937 4 gnd
port 514 nsew
rlabel metal2 s 28944 25043 28944 25043 4 gnd
port 514 nsew
rlabel metal2 s 27696 22673 27696 22673 4 gnd
port 514 nsew
rlabel metal2 s 28944 24253 28944 24253 4 gnd
port 514 nsew
rlabel metal2 s 28464 23700 28464 23700 4 gnd
port 514 nsew
rlabel metal2 s 27696 23463 27696 23463 4 gnd
port 514 nsew
rlabel metal2 s 28944 22673 28944 22673 4 gnd
port 514 nsew
rlabel metal2 s 29712 24253 29712 24253 4 gnd
port 514 nsew
rlabel metal2 s 29712 22910 29712 22910 4 gnd
port 514 nsew
rlabel metal2 s 28944 23700 28944 23700 4 gnd
port 514 nsew
rlabel metal2 s 29712 25280 29712 25280 4 gnd
port 514 nsew
rlabel metal2 s 28464 23463 28464 23463 4 gnd
port 514 nsew
rlabel metal2 s 28464 25280 28464 25280 4 gnd
port 514 nsew
rlabel metal2 s 28944 23463 28944 23463 4 gnd
port 514 nsew
rlabel metal2 s 29712 24490 29712 24490 4 gnd
port 514 nsew
rlabel metal2 s 27696 25280 27696 25280 4 gnd
port 514 nsew
rlabel metal2 s 27696 23700 27696 23700 4 gnd
port 514 nsew
rlabel metal2 s 27696 23147 27696 23147 4 gnd
port 514 nsew
rlabel metal2 s 27696 24727 27696 24727 4 gnd
port 514 nsew
rlabel metal2 s 28464 24253 28464 24253 4 gnd
port 514 nsew
rlabel metal2 s 28944 23937 28944 23937 4 gnd
port 514 nsew
rlabel metal2 s 27696 22910 27696 22910 4 gnd
port 514 nsew
rlabel metal2 s 29712 23700 29712 23700 4 gnd
port 514 nsew
rlabel metal2 s 28944 24490 28944 24490 4 gnd
port 514 nsew
rlabel metal2 s 28944 22910 28944 22910 4 gnd
port 514 nsew
rlabel metal2 s 28464 24727 28464 24727 4 gnd
port 514 nsew
rlabel metal2 s 28464 22673 28464 22673 4 gnd
port 514 nsew
rlabel metal2 s 29712 22673 29712 22673 4 gnd
port 514 nsew
rlabel metal2 s 25968 22357 25968 22357 4 gnd
port 514 nsew
rlabel metal2 s 27216 22357 27216 22357 4 gnd
port 514 nsew
rlabel metal2 s 27216 24490 27216 24490 4 gnd
port 514 nsew
rlabel metal2 s 27216 23937 27216 23937 4 gnd
port 514 nsew
rlabel metal2 s 25200 24490 25200 24490 4 gnd
port 514 nsew
rlabel metal2 s 26448 25280 26448 25280 4 gnd
port 514 nsew
rlabel metal2 s 26448 23700 26448 23700 4 gnd
port 514 nsew
rlabel metal2 s 25200 24727 25200 24727 4 gnd
port 514 nsew
rlabel metal2 s 25968 23147 25968 23147 4 gnd
port 514 nsew
rlabel metal2 s 25200 23147 25200 23147 4 gnd
port 514 nsew
rlabel metal2 s 25200 22910 25200 22910 4 gnd
port 514 nsew
rlabel metal2 s 26448 23463 26448 23463 4 gnd
port 514 nsew
rlabel metal2 s 25200 22357 25200 22357 4 gnd
port 514 nsew
rlabel metal2 s 25200 24253 25200 24253 4 gnd
port 514 nsew
rlabel metal2 s 27216 24727 27216 24727 4 gnd
port 514 nsew
rlabel metal2 s 25968 23700 25968 23700 4 gnd
port 514 nsew
rlabel metal2 s 25968 24727 25968 24727 4 gnd
port 514 nsew
rlabel metal2 s 25968 25043 25968 25043 4 gnd
port 514 nsew
rlabel metal2 s 25968 24253 25968 24253 4 gnd
port 514 nsew
rlabel metal2 s 27216 22910 27216 22910 4 gnd
port 514 nsew
rlabel metal2 s 27216 22673 27216 22673 4 gnd
port 514 nsew
rlabel metal2 s 26448 24490 26448 24490 4 gnd
port 514 nsew
rlabel metal2 s 26448 23937 26448 23937 4 gnd
port 514 nsew
rlabel metal2 s 26448 22357 26448 22357 4 gnd
port 514 nsew
rlabel metal2 s 25200 23463 25200 23463 4 gnd
port 514 nsew
rlabel metal2 s 27216 25280 27216 25280 4 gnd
port 514 nsew
rlabel metal2 s 26448 25043 26448 25043 4 gnd
port 514 nsew
rlabel metal2 s 27216 24253 27216 24253 4 gnd
port 514 nsew
rlabel metal2 s 27216 23463 27216 23463 4 gnd
port 514 nsew
rlabel metal2 s 25200 25280 25200 25280 4 gnd
port 514 nsew
rlabel metal2 s 25968 22910 25968 22910 4 gnd
port 514 nsew
rlabel metal2 s 27216 25043 27216 25043 4 gnd
port 514 nsew
rlabel metal2 s 25200 22673 25200 22673 4 gnd
port 514 nsew
rlabel metal2 s 26448 23147 26448 23147 4 gnd
port 514 nsew
rlabel metal2 s 25200 25043 25200 25043 4 gnd
port 514 nsew
rlabel metal2 s 26448 22910 26448 22910 4 gnd
port 514 nsew
rlabel metal2 s 25200 23700 25200 23700 4 gnd
port 514 nsew
rlabel metal2 s 25968 22673 25968 22673 4 gnd
port 514 nsew
rlabel metal2 s 27216 23700 27216 23700 4 gnd
port 514 nsew
rlabel metal2 s 25968 24490 25968 24490 4 gnd
port 514 nsew
rlabel metal2 s 26448 24253 26448 24253 4 gnd
port 514 nsew
rlabel metal2 s 27216 23147 27216 23147 4 gnd
port 514 nsew
rlabel metal2 s 25200 23937 25200 23937 4 gnd
port 514 nsew
rlabel metal2 s 26448 22673 26448 22673 4 gnd
port 514 nsew
rlabel metal2 s 25968 23937 25968 23937 4 gnd
port 514 nsew
rlabel metal2 s 25968 23463 25968 23463 4 gnd
port 514 nsew
rlabel metal2 s 25968 25280 25968 25280 4 gnd
port 514 nsew
rlabel metal2 s 26448 24727 26448 24727 4 gnd
port 514 nsew
rlabel metal2 s 27216 21567 27216 21567 4 gnd
port 514 nsew
rlabel metal2 s 25200 21883 25200 21883 4 gnd
port 514 nsew
rlabel metal2 s 25200 19197 25200 19197 4 gnd
port 514 nsew
rlabel metal2 s 25200 22120 25200 22120 4 gnd
port 514 nsew
rlabel metal2 s 26448 21883 26448 21883 4 gnd
port 514 nsew
rlabel metal2 s 27216 21093 27216 21093 4 gnd
port 514 nsew
rlabel metal2 s 26448 21330 26448 21330 4 gnd
port 514 nsew
rlabel metal2 s 25968 20303 25968 20303 4 gnd
port 514 nsew
rlabel metal2 s 27216 20303 27216 20303 4 gnd
port 514 nsew
rlabel metal2 s 26448 19197 26448 19197 4 gnd
port 514 nsew
rlabel metal2 s 27216 19987 27216 19987 4 gnd
port 514 nsew
rlabel metal2 s 25200 20777 25200 20777 4 gnd
port 514 nsew
rlabel metal2 s 25200 19750 25200 19750 4 gnd
port 514 nsew
rlabel metal2 s 27216 19513 27216 19513 4 gnd
port 514 nsew
rlabel metal2 s 25968 20540 25968 20540 4 gnd
port 514 nsew
rlabel metal2 s 25968 20777 25968 20777 4 gnd
port 514 nsew
rlabel metal2 s 25968 22120 25968 22120 4 gnd
port 514 nsew
rlabel metal2 s 26448 19513 26448 19513 4 gnd
port 514 nsew
rlabel metal2 s 25968 21567 25968 21567 4 gnd
port 514 nsew
rlabel metal2 s 26448 20777 26448 20777 4 gnd
port 514 nsew
rlabel metal2 s 25968 19513 25968 19513 4 gnd
port 514 nsew
rlabel metal2 s 26448 19750 26448 19750 4 gnd
port 514 nsew
rlabel metal2 s 25200 20540 25200 20540 4 gnd
port 514 nsew
rlabel metal2 s 27216 21330 27216 21330 4 gnd
port 514 nsew
rlabel metal2 s 25968 21093 25968 21093 4 gnd
port 514 nsew
rlabel metal2 s 26448 22120 26448 22120 4 gnd
port 514 nsew
rlabel metal2 s 25200 19513 25200 19513 4 gnd
port 514 nsew
rlabel metal2 s 25200 20303 25200 20303 4 gnd
port 514 nsew
rlabel metal2 s 25968 19750 25968 19750 4 gnd
port 514 nsew
rlabel metal2 s 25200 21567 25200 21567 4 gnd
port 514 nsew
rlabel metal2 s 25968 21883 25968 21883 4 gnd
port 514 nsew
rlabel metal2 s 26448 21567 26448 21567 4 gnd
port 514 nsew
rlabel metal2 s 25968 19197 25968 19197 4 gnd
port 514 nsew
rlabel metal2 s 25200 21330 25200 21330 4 gnd
port 514 nsew
rlabel metal2 s 25968 19987 25968 19987 4 gnd
port 514 nsew
rlabel metal2 s 25200 19987 25200 19987 4 gnd
port 514 nsew
rlabel metal2 s 27216 19197 27216 19197 4 gnd
port 514 nsew
rlabel metal2 s 27216 20777 27216 20777 4 gnd
port 514 nsew
rlabel metal2 s 27216 19750 27216 19750 4 gnd
port 514 nsew
rlabel metal2 s 27216 22120 27216 22120 4 gnd
port 514 nsew
rlabel metal2 s 26448 20303 26448 20303 4 gnd
port 514 nsew
rlabel metal2 s 25968 21330 25968 21330 4 gnd
port 514 nsew
rlabel metal2 s 25200 21093 25200 21093 4 gnd
port 514 nsew
rlabel metal2 s 27216 20540 27216 20540 4 gnd
port 514 nsew
rlabel metal2 s 27216 21883 27216 21883 4 gnd
port 514 nsew
rlabel metal2 s 26448 21093 26448 21093 4 gnd
port 514 nsew
rlabel metal2 s 26448 19987 26448 19987 4 gnd
port 514 nsew
rlabel metal2 s 26448 20540 26448 20540 4 gnd
port 514 nsew
rlabel metal2 s 28464 20540 28464 20540 4 gnd
port 514 nsew
rlabel metal2 s 28464 19513 28464 19513 4 gnd
port 514 nsew
rlabel metal2 s 29712 19513 29712 19513 4 gnd
port 514 nsew
rlabel metal2 s 27696 21093 27696 21093 4 gnd
port 514 nsew
rlabel metal2 s 28464 22120 28464 22120 4 gnd
port 514 nsew
rlabel metal2 s 27696 21567 27696 21567 4 gnd
port 514 nsew
rlabel metal2 s 29712 20303 29712 20303 4 gnd
port 514 nsew
rlabel metal2 s 28944 19513 28944 19513 4 gnd
port 514 nsew
rlabel metal2 s 27696 21330 27696 21330 4 gnd
port 514 nsew
rlabel metal2 s 28464 20303 28464 20303 4 gnd
port 514 nsew
rlabel metal2 s 29712 20540 29712 20540 4 gnd
port 514 nsew
rlabel metal2 s 28464 21883 28464 21883 4 gnd
port 514 nsew
rlabel metal2 s 28944 21883 28944 21883 4 gnd
port 514 nsew
rlabel metal2 s 28944 22120 28944 22120 4 gnd
port 514 nsew
rlabel metal2 s 29712 19197 29712 19197 4 gnd
port 514 nsew
rlabel metal2 s 27696 20303 27696 20303 4 gnd
port 514 nsew
rlabel metal2 s 28464 20777 28464 20777 4 gnd
port 514 nsew
rlabel metal2 s 29712 21093 29712 21093 4 gnd
port 514 nsew
rlabel metal2 s 29712 19987 29712 19987 4 gnd
port 514 nsew
rlabel metal2 s 28464 19750 28464 19750 4 gnd
port 514 nsew
rlabel metal2 s 29712 21330 29712 21330 4 gnd
port 514 nsew
rlabel metal2 s 29712 20777 29712 20777 4 gnd
port 514 nsew
rlabel metal2 s 29712 22120 29712 22120 4 gnd
port 514 nsew
rlabel metal2 s 28944 21330 28944 21330 4 gnd
port 514 nsew
rlabel metal2 s 27696 20777 27696 20777 4 gnd
port 514 nsew
rlabel metal2 s 27696 19513 27696 19513 4 gnd
port 514 nsew
rlabel metal2 s 27696 22120 27696 22120 4 gnd
port 514 nsew
rlabel metal2 s 27696 19987 27696 19987 4 gnd
port 514 nsew
rlabel metal2 s 29712 21883 29712 21883 4 gnd
port 514 nsew
rlabel metal2 s 28944 19987 28944 19987 4 gnd
port 514 nsew
rlabel metal2 s 28944 20777 28944 20777 4 gnd
port 514 nsew
rlabel metal2 s 28944 19750 28944 19750 4 gnd
port 514 nsew
rlabel metal2 s 28944 21567 28944 21567 4 gnd
port 514 nsew
rlabel metal2 s 28464 21567 28464 21567 4 gnd
port 514 nsew
rlabel metal2 s 27696 20540 27696 20540 4 gnd
port 514 nsew
rlabel metal2 s 28464 19987 28464 19987 4 gnd
port 514 nsew
rlabel metal2 s 28944 19197 28944 19197 4 gnd
port 514 nsew
rlabel metal2 s 27696 21883 27696 21883 4 gnd
port 514 nsew
rlabel metal2 s 28944 21093 28944 21093 4 gnd
port 514 nsew
rlabel metal2 s 29712 19750 29712 19750 4 gnd
port 514 nsew
rlabel metal2 s 28944 20540 28944 20540 4 gnd
port 514 nsew
rlabel metal2 s 27696 19750 27696 19750 4 gnd
port 514 nsew
rlabel metal2 s 28464 21330 28464 21330 4 gnd
port 514 nsew
rlabel metal2 s 28464 21093 28464 21093 4 gnd
port 514 nsew
rlabel metal2 s 27696 19197 27696 19197 4 gnd
port 514 nsew
rlabel metal2 s 29712 21567 29712 21567 4 gnd
port 514 nsew
rlabel metal2 s 28944 20303 28944 20303 4 gnd
port 514 nsew
rlabel metal2 s 28464 19197 28464 19197 4 gnd
port 514 nsew
rlabel metal2 s 23472 23147 23472 23147 4 gnd
port 514 nsew
rlabel metal2 s 23472 24490 23472 24490 4 gnd
port 514 nsew
rlabel metal2 s 23952 23937 23952 23937 4 gnd
port 514 nsew
rlabel metal2 s 23472 22673 23472 22673 4 gnd
port 514 nsew
rlabel metal2 s 23472 24253 23472 24253 4 gnd
port 514 nsew
rlabel metal2 s 22704 23700 22704 23700 4 gnd
port 514 nsew
rlabel metal2 s 22704 22357 22704 22357 4 gnd
port 514 nsew
rlabel metal2 s 23952 23463 23952 23463 4 gnd
port 514 nsew
rlabel metal2 s 22704 24727 22704 24727 4 gnd
port 514 nsew
rlabel metal2 s 23472 22357 23472 22357 4 gnd
port 514 nsew
rlabel metal2 s 23952 25043 23952 25043 4 gnd
port 514 nsew
rlabel metal2 s 22704 23463 22704 23463 4 gnd
port 514 nsew
rlabel metal2 s 22704 22673 22704 22673 4 gnd
port 514 nsew
rlabel metal2 s 23472 24727 23472 24727 4 gnd
port 514 nsew
rlabel metal2 s 23952 23700 23952 23700 4 gnd
port 514 nsew
rlabel metal2 s 23472 23463 23472 23463 4 gnd
port 514 nsew
rlabel metal2 s 24720 23937 24720 23937 4 gnd
port 514 nsew
rlabel metal2 s 23472 25043 23472 25043 4 gnd
port 514 nsew
rlabel metal2 s 24720 24727 24720 24727 4 gnd
port 514 nsew
rlabel metal2 s 23952 22357 23952 22357 4 gnd
port 514 nsew
rlabel metal2 s 24720 24490 24720 24490 4 gnd
port 514 nsew
rlabel metal2 s 23472 23700 23472 23700 4 gnd
port 514 nsew
rlabel metal2 s 23952 25280 23952 25280 4 gnd
port 514 nsew
rlabel metal2 s 24720 25280 24720 25280 4 gnd
port 514 nsew
rlabel metal2 s 22704 25280 22704 25280 4 gnd
port 514 nsew
rlabel metal2 s 24720 23147 24720 23147 4 gnd
port 514 nsew
rlabel metal2 s 24720 22673 24720 22673 4 gnd
port 514 nsew
rlabel metal2 s 23952 24253 23952 24253 4 gnd
port 514 nsew
rlabel metal2 s 24720 22910 24720 22910 4 gnd
port 514 nsew
rlabel metal2 s 22704 22910 22704 22910 4 gnd
port 514 nsew
rlabel metal2 s 24720 23700 24720 23700 4 gnd
port 514 nsew
rlabel metal2 s 24720 24253 24720 24253 4 gnd
port 514 nsew
rlabel metal2 s 22704 23937 22704 23937 4 gnd
port 514 nsew
rlabel metal2 s 22704 23147 22704 23147 4 gnd
port 514 nsew
rlabel metal2 s 22704 25043 22704 25043 4 gnd
port 514 nsew
rlabel metal2 s 23952 22673 23952 22673 4 gnd
port 514 nsew
rlabel metal2 s 23952 23147 23952 23147 4 gnd
port 514 nsew
rlabel metal2 s 23472 23937 23472 23937 4 gnd
port 514 nsew
rlabel metal2 s 24720 23463 24720 23463 4 gnd
port 514 nsew
rlabel metal2 s 22704 24253 22704 24253 4 gnd
port 514 nsew
rlabel metal2 s 24720 25043 24720 25043 4 gnd
port 514 nsew
rlabel metal2 s 22704 24490 22704 24490 4 gnd
port 514 nsew
rlabel metal2 s 23472 25280 23472 25280 4 gnd
port 514 nsew
rlabel metal2 s 23952 24490 23952 24490 4 gnd
port 514 nsew
rlabel metal2 s 23952 22910 23952 22910 4 gnd
port 514 nsew
rlabel metal2 s 23952 24727 23952 24727 4 gnd
port 514 nsew
rlabel metal2 s 24720 22357 24720 22357 4 gnd
port 514 nsew
rlabel metal2 s 23472 22910 23472 22910 4 gnd
port 514 nsew
rlabel metal2 s 20976 24490 20976 24490 4 gnd
port 514 nsew
rlabel metal2 s 22224 24727 22224 24727 4 gnd
port 514 nsew
rlabel metal2 s 21456 22910 21456 22910 4 gnd
port 514 nsew
rlabel metal2 s 22224 23463 22224 23463 4 gnd
port 514 nsew
rlabel metal2 s 21456 23147 21456 23147 4 gnd
port 514 nsew
rlabel metal2 s 20976 25043 20976 25043 4 gnd
port 514 nsew
rlabel metal2 s 20976 24253 20976 24253 4 gnd
port 514 nsew
rlabel metal2 s 21456 24253 21456 24253 4 gnd
port 514 nsew
rlabel metal2 s 20208 22357 20208 22357 4 gnd
port 514 nsew
rlabel metal2 s 20976 23937 20976 23937 4 gnd
port 514 nsew
rlabel metal2 s 20208 23937 20208 23937 4 gnd
port 514 nsew
rlabel metal2 s 20208 25280 20208 25280 4 gnd
port 514 nsew
rlabel metal2 s 20208 23463 20208 23463 4 gnd
port 514 nsew
rlabel metal2 s 20976 24727 20976 24727 4 gnd
port 514 nsew
rlabel metal2 s 21456 23937 21456 23937 4 gnd
port 514 nsew
rlabel metal2 s 22224 23937 22224 23937 4 gnd
port 514 nsew
rlabel metal2 s 20976 22673 20976 22673 4 gnd
port 514 nsew
rlabel metal2 s 21456 24490 21456 24490 4 gnd
port 514 nsew
rlabel metal2 s 20976 23147 20976 23147 4 gnd
port 514 nsew
rlabel metal2 s 20208 22910 20208 22910 4 gnd
port 514 nsew
rlabel metal2 s 20976 23700 20976 23700 4 gnd
port 514 nsew
rlabel metal2 s 22224 24253 22224 24253 4 gnd
port 514 nsew
rlabel metal2 s 21456 22357 21456 22357 4 gnd
port 514 nsew
rlabel metal2 s 20208 23147 20208 23147 4 gnd
port 514 nsew
rlabel metal2 s 20208 24253 20208 24253 4 gnd
port 514 nsew
rlabel metal2 s 20208 24727 20208 24727 4 gnd
port 514 nsew
rlabel metal2 s 22224 24490 22224 24490 4 gnd
port 514 nsew
rlabel metal2 s 22224 25043 22224 25043 4 gnd
port 514 nsew
rlabel metal2 s 20208 25043 20208 25043 4 gnd
port 514 nsew
rlabel metal2 s 21456 22673 21456 22673 4 gnd
port 514 nsew
rlabel metal2 s 21456 25043 21456 25043 4 gnd
port 514 nsew
rlabel metal2 s 20208 23700 20208 23700 4 gnd
port 514 nsew
rlabel metal2 s 22224 22357 22224 22357 4 gnd
port 514 nsew
rlabel metal2 s 22224 23700 22224 23700 4 gnd
port 514 nsew
rlabel metal2 s 21456 24727 21456 24727 4 gnd
port 514 nsew
rlabel metal2 s 20208 24490 20208 24490 4 gnd
port 514 nsew
rlabel metal2 s 22224 22673 22224 22673 4 gnd
port 514 nsew
rlabel metal2 s 21456 23463 21456 23463 4 gnd
port 514 nsew
rlabel metal2 s 22224 23147 22224 23147 4 gnd
port 514 nsew
rlabel metal2 s 20976 22910 20976 22910 4 gnd
port 514 nsew
rlabel metal2 s 21456 25280 21456 25280 4 gnd
port 514 nsew
rlabel metal2 s 20208 22673 20208 22673 4 gnd
port 514 nsew
rlabel metal2 s 20976 22357 20976 22357 4 gnd
port 514 nsew
rlabel metal2 s 20976 25280 20976 25280 4 gnd
port 514 nsew
rlabel metal2 s 22224 25280 22224 25280 4 gnd
port 514 nsew
rlabel metal2 s 21456 23700 21456 23700 4 gnd
port 514 nsew
rlabel metal2 s 22224 22910 22224 22910 4 gnd
port 514 nsew
rlabel metal2 s 20976 23463 20976 23463 4 gnd
port 514 nsew
rlabel metal2 s 21456 22120 21456 22120 4 gnd
port 514 nsew
rlabel metal2 s 20208 19750 20208 19750 4 gnd
port 514 nsew
rlabel metal2 s 21456 21330 21456 21330 4 gnd
port 514 nsew
rlabel metal2 s 21456 19987 21456 19987 4 gnd
port 514 nsew
rlabel metal2 s 22224 21330 22224 21330 4 gnd
port 514 nsew
rlabel metal2 s 20976 21330 20976 21330 4 gnd
port 514 nsew
rlabel metal2 s 21456 19197 21456 19197 4 gnd
port 514 nsew
rlabel metal2 s 20976 19987 20976 19987 4 gnd
port 514 nsew
rlabel metal2 s 20208 20540 20208 20540 4 gnd
port 514 nsew
rlabel metal2 s 21456 21567 21456 21567 4 gnd
port 514 nsew
rlabel metal2 s 20208 21883 20208 21883 4 gnd
port 514 nsew
rlabel metal2 s 20208 21330 20208 21330 4 gnd
port 514 nsew
rlabel metal2 s 21456 21883 21456 21883 4 gnd
port 514 nsew
rlabel metal2 s 20208 19197 20208 19197 4 gnd
port 514 nsew
rlabel metal2 s 21456 20540 21456 20540 4 gnd
port 514 nsew
rlabel metal2 s 20208 20777 20208 20777 4 gnd
port 514 nsew
rlabel metal2 s 20976 21567 20976 21567 4 gnd
port 514 nsew
rlabel metal2 s 20976 20540 20976 20540 4 gnd
port 514 nsew
rlabel metal2 s 20976 19750 20976 19750 4 gnd
port 514 nsew
rlabel metal2 s 20208 19513 20208 19513 4 gnd
port 514 nsew
rlabel metal2 s 21456 19750 21456 19750 4 gnd
port 514 nsew
rlabel metal2 s 22224 21883 22224 21883 4 gnd
port 514 nsew
rlabel metal2 s 20976 21093 20976 21093 4 gnd
port 514 nsew
rlabel metal2 s 22224 20540 22224 20540 4 gnd
port 514 nsew
rlabel metal2 s 22224 21093 22224 21093 4 gnd
port 514 nsew
rlabel metal2 s 21456 20777 21456 20777 4 gnd
port 514 nsew
rlabel metal2 s 22224 21567 22224 21567 4 gnd
port 514 nsew
rlabel metal2 s 20976 20777 20976 20777 4 gnd
port 514 nsew
rlabel metal2 s 22224 20777 22224 20777 4 gnd
port 514 nsew
rlabel metal2 s 20208 22120 20208 22120 4 gnd
port 514 nsew
rlabel metal2 s 20208 21567 20208 21567 4 gnd
port 514 nsew
rlabel metal2 s 22224 19513 22224 19513 4 gnd
port 514 nsew
rlabel metal2 s 20976 19197 20976 19197 4 gnd
port 514 nsew
rlabel metal2 s 20208 20303 20208 20303 4 gnd
port 514 nsew
rlabel metal2 s 21456 20303 21456 20303 4 gnd
port 514 nsew
rlabel metal2 s 20976 19513 20976 19513 4 gnd
port 514 nsew
rlabel metal2 s 21456 21093 21456 21093 4 gnd
port 514 nsew
rlabel metal2 s 22224 19750 22224 19750 4 gnd
port 514 nsew
rlabel metal2 s 22224 22120 22224 22120 4 gnd
port 514 nsew
rlabel metal2 s 20208 19987 20208 19987 4 gnd
port 514 nsew
rlabel metal2 s 21456 19513 21456 19513 4 gnd
port 514 nsew
rlabel metal2 s 22224 20303 22224 20303 4 gnd
port 514 nsew
rlabel metal2 s 20208 21093 20208 21093 4 gnd
port 514 nsew
rlabel metal2 s 20976 22120 20976 22120 4 gnd
port 514 nsew
rlabel metal2 s 22224 19197 22224 19197 4 gnd
port 514 nsew
rlabel metal2 s 22224 19987 22224 19987 4 gnd
port 514 nsew
rlabel metal2 s 20976 20303 20976 20303 4 gnd
port 514 nsew
rlabel metal2 s 20976 21883 20976 21883 4 gnd
port 514 nsew
rlabel metal2 s 23952 21567 23952 21567 4 gnd
port 514 nsew
rlabel metal2 s 23472 20540 23472 20540 4 gnd
port 514 nsew
rlabel metal2 s 22704 21567 22704 21567 4 gnd
port 514 nsew
rlabel metal2 s 24720 21883 24720 21883 4 gnd
port 514 nsew
rlabel metal2 s 24720 19197 24720 19197 4 gnd
port 514 nsew
rlabel metal2 s 23952 21330 23952 21330 4 gnd
port 514 nsew
rlabel metal2 s 22704 19197 22704 19197 4 gnd
port 514 nsew
rlabel metal2 s 23472 21093 23472 21093 4 gnd
port 514 nsew
rlabel metal2 s 24720 21093 24720 21093 4 gnd
port 514 nsew
rlabel metal2 s 23952 22120 23952 22120 4 gnd
port 514 nsew
rlabel metal2 s 23472 20777 23472 20777 4 gnd
port 514 nsew
rlabel metal2 s 22704 19987 22704 19987 4 gnd
port 514 nsew
rlabel metal2 s 22704 20303 22704 20303 4 gnd
port 514 nsew
rlabel metal2 s 23952 19197 23952 19197 4 gnd
port 514 nsew
rlabel metal2 s 24720 20777 24720 20777 4 gnd
port 514 nsew
rlabel metal2 s 24720 21330 24720 21330 4 gnd
port 514 nsew
rlabel metal2 s 22704 19750 22704 19750 4 gnd
port 514 nsew
rlabel metal2 s 23952 19750 23952 19750 4 gnd
port 514 nsew
rlabel metal2 s 23952 20540 23952 20540 4 gnd
port 514 nsew
rlabel metal2 s 23472 22120 23472 22120 4 gnd
port 514 nsew
rlabel metal2 s 24720 21567 24720 21567 4 gnd
port 514 nsew
rlabel metal2 s 23472 20303 23472 20303 4 gnd
port 514 nsew
rlabel metal2 s 23472 21883 23472 21883 4 gnd
port 514 nsew
rlabel metal2 s 23952 21093 23952 21093 4 gnd
port 514 nsew
rlabel metal2 s 24720 22120 24720 22120 4 gnd
port 514 nsew
rlabel metal2 s 24720 20540 24720 20540 4 gnd
port 514 nsew
rlabel metal2 s 24720 19750 24720 19750 4 gnd
port 514 nsew
rlabel metal2 s 23952 19513 23952 19513 4 gnd
port 514 nsew
rlabel metal2 s 23952 20777 23952 20777 4 gnd
port 514 nsew
rlabel metal2 s 22704 21093 22704 21093 4 gnd
port 514 nsew
rlabel metal2 s 24720 19513 24720 19513 4 gnd
port 514 nsew
rlabel metal2 s 22704 20540 22704 20540 4 gnd
port 514 nsew
rlabel metal2 s 24720 19987 24720 19987 4 gnd
port 514 nsew
rlabel metal2 s 24720 20303 24720 20303 4 gnd
port 514 nsew
rlabel metal2 s 22704 21330 22704 21330 4 gnd
port 514 nsew
rlabel metal2 s 23472 21330 23472 21330 4 gnd
port 514 nsew
rlabel metal2 s 22704 22120 22704 22120 4 gnd
port 514 nsew
rlabel metal2 s 23472 19197 23472 19197 4 gnd
port 514 nsew
rlabel metal2 s 22704 19513 22704 19513 4 gnd
port 514 nsew
rlabel metal2 s 22704 20777 22704 20777 4 gnd
port 514 nsew
rlabel metal2 s 23472 19513 23472 19513 4 gnd
port 514 nsew
rlabel metal2 s 23472 19987 23472 19987 4 gnd
port 514 nsew
rlabel metal2 s 23952 21883 23952 21883 4 gnd
port 514 nsew
rlabel metal2 s 22704 21883 22704 21883 4 gnd
port 514 nsew
rlabel metal2 s 23472 19750 23472 19750 4 gnd
port 514 nsew
rlabel metal2 s 23472 21567 23472 21567 4 gnd
port 514 nsew
rlabel metal2 s 23952 20303 23952 20303 4 gnd
port 514 nsew
rlabel metal2 s 23952 19987 23952 19987 4 gnd
port 514 nsew
rlabel metal2 s 23952 17933 23952 17933 4 gnd
port 514 nsew
rlabel metal2 s 24720 18960 24720 18960 4 gnd
port 514 nsew
rlabel metal2 s 22704 18723 22704 18723 4 gnd
port 514 nsew
rlabel metal2 s 23472 18407 23472 18407 4 gnd
port 514 nsew
rlabel metal2 s 22704 17143 22704 17143 4 gnd
port 514 nsew
rlabel metal2 s 23472 16827 23472 16827 4 gnd
port 514 nsew
rlabel metal2 s 24720 17617 24720 17617 4 gnd
port 514 nsew
rlabel metal2 s 23472 16037 23472 16037 4 gnd
port 514 nsew
rlabel metal2 s 22704 16590 22704 16590 4 gnd
port 514 nsew
rlabel metal2 s 23952 18170 23952 18170 4 gnd
port 514 nsew
rlabel metal2 s 23472 16590 23472 16590 4 gnd
port 514 nsew
rlabel metal2 s 23952 17143 23952 17143 4 gnd
port 514 nsew
rlabel metal2 s 23952 18723 23952 18723 4 gnd
port 514 nsew
rlabel metal2 s 24720 18170 24720 18170 4 gnd
port 514 nsew
rlabel metal2 s 23952 16590 23952 16590 4 gnd
port 514 nsew
rlabel metal2 s 23472 17617 23472 17617 4 gnd
port 514 nsew
rlabel metal2 s 24720 18407 24720 18407 4 gnd
port 514 nsew
rlabel metal2 s 22704 16353 22704 16353 4 gnd
port 514 nsew
rlabel metal2 s 23952 18407 23952 18407 4 gnd
port 514 nsew
rlabel metal2 s 23472 17143 23472 17143 4 gnd
port 514 nsew
rlabel metal2 s 22704 16827 22704 16827 4 gnd
port 514 nsew
rlabel metal2 s 22704 17617 22704 17617 4 gnd
port 514 nsew
rlabel metal2 s 23952 16827 23952 16827 4 gnd
port 514 nsew
rlabel metal2 s 23952 16037 23952 16037 4 gnd
port 514 nsew
rlabel metal2 s 23952 17380 23952 17380 4 gnd
port 514 nsew
rlabel metal2 s 22704 17933 22704 17933 4 gnd
port 514 nsew
rlabel metal2 s 24720 17933 24720 17933 4 gnd
port 514 nsew
rlabel metal2 s 23952 17617 23952 17617 4 gnd
port 514 nsew
rlabel metal2 s 23952 18960 23952 18960 4 gnd
port 514 nsew
rlabel metal2 s 24720 17380 24720 17380 4 gnd
port 514 nsew
rlabel metal2 s 23472 17380 23472 17380 4 gnd
port 514 nsew
rlabel metal2 s 23472 18170 23472 18170 4 gnd
port 514 nsew
rlabel metal2 s 22704 17380 22704 17380 4 gnd
port 514 nsew
rlabel metal2 s 22704 16037 22704 16037 4 gnd
port 514 nsew
rlabel metal2 s 23472 18723 23472 18723 4 gnd
port 514 nsew
rlabel metal2 s 22704 18407 22704 18407 4 gnd
port 514 nsew
rlabel metal2 s 24720 18723 24720 18723 4 gnd
port 514 nsew
rlabel metal2 s 22704 18960 22704 18960 4 gnd
port 514 nsew
rlabel metal2 s 22704 18170 22704 18170 4 gnd
port 514 nsew
rlabel metal2 s 24720 16590 24720 16590 4 gnd
port 514 nsew
rlabel metal2 s 24720 16827 24720 16827 4 gnd
port 514 nsew
rlabel metal2 s 24720 17143 24720 17143 4 gnd
port 514 nsew
rlabel metal2 s 24720 16353 24720 16353 4 gnd
port 514 nsew
rlabel metal2 s 23472 18960 23472 18960 4 gnd
port 514 nsew
rlabel metal2 s 23472 16353 23472 16353 4 gnd
port 514 nsew
rlabel metal2 s 24720 16037 24720 16037 4 gnd
port 514 nsew
rlabel metal2 s 23472 17933 23472 17933 4 gnd
port 514 nsew
rlabel metal2 s 23952 16353 23952 16353 4 gnd
port 514 nsew
rlabel metal2 s 21456 17143 21456 17143 4 gnd
port 514 nsew
rlabel metal2 s 20976 17933 20976 17933 4 gnd
port 514 nsew
rlabel metal2 s 21456 16037 21456 16037 4 gnd
port 514 nsew
rlabel metal2 s 22224 18723 22224 18723 4 gnd
port 514 nsew
rlabel metal2 s 21456 16353 21456 16353 4 gnd
port 514 nsew
rlabel metal2 s 20208 18407 20208 18407 4 gnd
port 514 nsew
rlabel metal2 s 21456 18407 21456 18407 4 gnd
port 514 nsew
rlabel metal2 s 20976 16353 20976 16353 4 gnd
port 514 nsew
rlabel metal2 s 21456 18723 21456 18723 4 gnd
port 514 nsew
rlabel metal2 s 20208 17143 20208 17143 4 gnd
port 514 nsew
rlabel metal2 s 20208 18723 20208 18723 4 gnd
port 514 nsew
rlabel metal2 s 20208 16037 20208 16037 4 gnd
port 514 nsew
rlabel metal2 s 22224 18407 22224 18407 4 gnd
port 514 nsew
rlabel metal2 s 20976 18960 20976 18960 4 gnd
port 514 nsew
rlabel metal2 s 20976 17143 20976 17143 4 gnd
port 514 nsew
rlabel metal2 s 22224 16590 22224 16590 4 gnd
port 514 nsew
rlabel metal2 s 22224 16827 22224 16827 4 gnd
port 514 nsew
rlabel metal2 s 22224 17933 22224 17933 4 gnd
port 514 nsew
rlabel metal2 s 22224 17617 22224 17617 4 gnd
port 514 nsew
rlabel metal2 s 20976 17380 20976 17380 4 gnd
port 514 nsew
rlabel metal2 s 20208 18170 20208 18170 4 gnd
port 514 nsew
rlabel metal2 s 20208 17617 20208 17617 4 gnd
port 514 nsew
rlabel metal2 s 20976 18407 20976 18407 4 gnd
port 514 nsew
rlabel metal2 s 20208 17380 20208 17380 4 gnd
port 514 nsew
rlabel metal2 s 20208 17933 20208 17933 4 gnd
port 514 nsew
rlabel metal2 s 20208 16353 20208 16353 4 gnd
port 514 nsew
rlabel metal2 s 21456 17933 21456 17933 4 gnd
port 514 nsew
rlabel metal2 s 22224 17380 22224 17380 4 gnd
port 514 nsew
rlabel metal2 s 21456 16827 21456 16827 4 gnd
port 514 nsew
rlabel metal2 s 22224 18170 22224 18170 4 gnd
port 514 nsew
rlabel metal2 s 20208 16827 20208 16827 4 gnd
port 514 nsew
rlabel metal2 s 21456 18170 21456 18170 4 gnd
port 514 nsew
rlabel metal2 s 20976 17617 20976 17617 4 gnd
port 514 nsew
rlabel metal2 s 20208 16590 20208 16590 4 gnd
port 514 nsew
rlabel metal2 s 21456 17380 21456 17380 4 gnd
port 514 nsew
rlabel metal2 s 20976 18170 20976 18170 4 gnd
port 514 nsew
rlabel metal2 s 21456 16590 21456 16590 4 gnd
port 514 nsew
rlabel metal2 s 21456 18960 21456 18960 4 gnd
port 514 nsew
rlabel metal2 s 22224 16037 22224 16037 4 gnd
port 514 nsew
rlabel metal2 s 22224 18960 22224 18960 4 gnd
port 514 nsew
rlabel metal2 s 22224 16353 22224 16353 4 gnd
port 514 nsew
rlabel metal2 s 20208 18960 20208 18960 4 gnd
port 514 nsew
rlabel metal2 s 20976 18723 20976 18723 4 gnd
port 514 nsew
rlabel metal2 s 20976 16827 20976 16827 4 gnd
port 514 nsew
rlabel metal2 s 21456 17617 21456 17617 4 gnd
port 514 nsew
rlabel metal2 s 20976 16037 20976 16037 4 gnd
port 514 nsew
rlabel metal2 s 22224 17143 22224 17143 4 gnd
port 514 nsew
rlabel metal2 s 20976 16590 20976 16590 4 gnd
port 514 nsew
rlabel metal2 s 22224 12877 22224 12877 4 gnd
port 514 nsew
rlabel metal2 s 21456 15563 21456 15563 4 gnd
port 514 nsew
rlabel metal2 s 21456 14773 21456 14773 4 gnd
port 514 nsew
rlabel metal2 s 21456 15010 21456 15010 4 gnd
port 514 nsew
rlabel metal2 s 20976 14773 20976 14773 4 gnd
port 514 nsew
rlabel metal2 s 21456 13667 21456 13667 4 gnd
port 514 nsew
rlabel metal2 s 20976 13193 20976 13193 4 gnd
port 514 nsew
rlabel metal2 s 21456 14220 21456 14220 4 gnd
port 514 nsew
rlabel metal2 s 22224 13667 22224 13667 4 gnd
port 514 nsew
rlabel metal2 s 22224 15010 22224 15010 4 gnd
port 514 nsew
rlabel metal2 s 20976 13667 20976 13667 4 gnd
port 514 nsew
rlabel metal2 s 22224 14457 22224 14457 4 gnd
port 514 nsew
rlabel metal2 s 20976 13430 20976 13430 4 gnd
port 514 nsew
rlabel metal2 s 21456 13983 21456 13983 4 gnd
port 514 nsew
rlabel metal2 s 22224 15800 22224 15800 4 gnd
port 514 nsew
rlabel metal2 s 21456 13430 21456 13430 4 gnd
port 514 nsew
rlabel metal2 s 21456 12877 21456 12877 4 gnd
port 514 nsew
rlabel metal2 s 21456 15247 21456 15247 4 gnd
port 514 nsew
rlabel metal2 s 20208 14220 20208 14220 4 gnd
port 514 nsew
rlabel metal2 s 22224 15247 22224 15247 4 gnd
port 514 nsew
rlabel metal2 s 22224 13983 22224 13983 4 gnd
port 514 nsew
rlabel metal2 s 22224 14220 22224 14220 4 gnd
port 514 nsew
rlabel metal2 s 21456 13193 21456 13193 4 gnd
port 514 nsew
rlabel metal2 s 20976 14220 20976 14220 4 gnd
port 514 nsew
rlabel metal2 s 20208 15010 20208 15010 4 gnd
port 514 nsew
rlabel metal2 s 20208 15800 20208 15800 4 gnd
port 514 nsew
rlabel metal2 s 20208 15563 20208 15563 4 gnd
port 514 nsew
rlabel metal2 s 20976 15800 20976 15800 4 gnd
port 514 nsew
rlabel metal2 s 22224 13193 22224 13193 4 gnd
port 514 nsew
rlabel metal2 s 20208 14457 20208 14457 4 gnd
port 514 nsew
rlabel metal2 s 20208 13667 20208 13667 4 gnd
port 514 nsew
rlabel metal2 s 20208 13193 20208 13193 4 gnd
port 514 nsew
rlabel metal2 s 20976 15563 20976 15563 4 gnd
port 514 nsew
rlabel metal2 s 20208 12877 20208 12877 4 gnd
port 514 nsew
rlabel metal2 s 20208 15247 20208 15247 4 gnd
port 514 nsew
rlabel metal2 s 21456 14457 21456 14457 4 gnd
port 514 nsew
rlabel metal2 s 20208 13983 20208 13983 4 gnd
port 514 nsew
rlabel metal2 s 22224 14773 22224 14773 4 gnd
port 514 nsew
rlabel metal2 s 20976 15010 20976 15010 4 gnd
port 514 nsew
rlabel metal2 s 20976 13983 20976 13983 4 gnd
port 514 nsew
rlabel metal2 s 20976 15247 20976 15247 4 gnd
port 514 nsew
rlabel metal2 s 20208 14773 20208 14773 4 gnd
port 514 nsew
rlabel metal2 s 20976 12877 20976 12877 4 gnd
port 514 nsew
rlabel metal2 s 20976 14457 20976 14457 4 gnd
port 514 nsew
rlabel metal2 s 22224 13430 22224 13430 4 gnd
port 514 nsew
rlabel metal2 s 20208 13430 20208 13430 4 gnd
port 514 nsew
rlabel metal2 s 22224 15563 22224 15563 4 gnd
port 514 nsew
rlabel metal2 s 21456 15800 21456 15800 4 gnd
port 514 nsew
rlabel metal2 s 24720 12877 24720 12877 4 gnd
port 514 nsew
rlabel metal2 s 22704 14457 22704 14457 4 gnd
port 514 nsew
rlabel metal2 s 24720 15010 24720 15010 4 gnd
port 514 nsew
rlabel metal2 s 22704 13430 22704 13430 4 gnd
port 514 nsew
rlabel metal2 s 23952 14220 23952 14220 4 gnd
port 514 nsew
rlabel metal2 s 22704 13193 22704 13193 4 gnd
port 514 nsew
rlabel metal2 s 23952 12877 23952 12877 4 gnd
port 514 nsew
rlabel metal2 s 24720 13430 24720 13430 4 gnd
port 514 nsew
rlabel metal2 s 22704 15563 22704 15563 4 gnd
port 514 nsew
rlabel metal2 s 23952 15800 23952 15800 4 gnd
port 514 nsew
rlabel metal2 s 23952 15010 23952 15010 4 gnd
port 514 nsew
rlabel metal2 s 23472 12877 23472 12877 4 gnd
port 514 nsew
rlabel metal2 s 23472 15563 23472 15563 4 gnd
port 514 nsew
rlabel metal2 s 24720 14773 24720 14773 4 gnd
port 514 nsew
rlabel metal2 s 24720 15247 24720 15247 4 gnd
port 514 nsew
rlabel metal2 s 22704 13983 22704 13983 4 gnd
port 514 nsew
rlabel metal2 s 22704 13667 22704 13667 4 gnd
port 514 nsew
rlabel metal2 s 22704 14773 22704 14773 4 gnd
port 514 nsew
rlabel metal2 s 23952 14457 23952 14457 4 gnd
port 514 nsew
rlabel metal2 s 24720 13193 24720 13193 4 gnd
port 514 nsew
rlabel metal2 s 22704 15800 22704 15800 4 gnd
port 514 nsew
rlabel metal2 s 23952 13430 23952 13430 4 gnd
port 514 nsew
rlabel metal2 s 22704 15247 22704 15247 4 gnd
port 514 nsew
rlabel metal2 s 22704 15010 22704 15010 4 gnd
port 514 nsew
rlabel metal2 s 23472 13667 23472 13667 4 gnd
port 514 nsew
rlabel metal2 s 23472 13430 23472 13430 4 gnd
port 514 nsew
rlabel metal2 s 23472 15247 23472 15247 4 gnd
port 514 nsew
rlabel metal2 s 24720 15563 24720 15563 4 gnd
port 514 nsew
rlabel metal2 s 23952 13193 23952 13193 4 gnd
port 514 nsew
rlabel metal2 s 24720 15800 24720 15800 4 gnd
port 514 nsew
rlabel metal2 s 23952 14773 23952 14773 4 gnd
port 514 nsew
rlabel metal2 s 23952 15247 23952 15247 4 gnd
port 514 nsew
rlabel metal2 s 23952 13983 23952 13983 4 gnd
port 514 nsew
rlabel metal2 s 22704 14220 22704 14220 4 gnd
port 514 nsew
rlabel metal2 s 24720 14457 24720 14457 4 gnd
port 514 nsew
rlabel metal2 s 24720 14220 24720 14220 4 gnd
port 514 nsew
rlabel metal2 s 23472 15010 23472 15010 4 gnd
port 514 nsew
rlabel metal2 s 23952 13667 23952 13667 4 gnd
port 514 nsew
rlabel metal2 s 23472 15800 23472 15800 4 gnd
port 514 nsew
rlabel metal2 s 23952 15563 23952 15563 4 gnd
port 514 nsew
rlabel metal2 s 24720 13667 24720 13667 4 gnd
port 514 nsew
rlabel metal2 s 23472 14220 23472 14220 4 gnd
port 514 nsew
rlabel metal2 s 23472 13983 23472 13983 4 gnd
port 514 nsew
rlabel metal2 s 23472 14457 23472 14457 4 gnd
port 514 nsew
rlabel metal2 s 22704 12877 22704 12877 4 gnd
port 514 nsew
rlabel metal2 s 23472 14773 23472 14773 4 gnd
port 514 nsew
rlabel metal2 s 23472 13193 23472 13193 4 gnd
port 514 nsew
rlabel metal2 s 24720 13983 24720 13983 4 gnd
port 514 nsew
rlabel metal2 s 28464 18407 28464 18407 4 gnd
port 514 nsew
rlabel metal2 s 27696 17933 27696 17933 4 gnd
port 514 nsew
rlabel metal2 s 28944 18170 28944 18170 4 gnd
port 514 nsew
rlabel metal2 s 27696 16827 27696 16827 4 gnd
port 514 nsew
rlabel metal2 s 29712 17143 29712 17143 4 gnd
port 514 nsew
rlabel metal2 s 29712 18723 29712 18723 4 gnd
port 514 nsew
rlabel metal2 s 28464 18723 28464 18723 4 gnd
port 514 nsew
rlabel metal2 s 28464 17143 28464 17143 4 gnd
port 514 nsew
rlabel metal2 s 27696 18170 27696 18170 4 gnd
port 514 nsew
rlabel metal2 s 28944 18407 28944 18407 4 gnd
port 514 nsew
rlabel metal2 s 28944 17380 28944 17380 4 gnd
port 514 nsew
rlabel metal2 s 28464 16037 28464 16037 4 gnd
port 514 nsew
rlabel metal2 s 28464 17617 28464 17617 4 gnd
port 514 nsew
rlabel metal2 s 27696 16590 27696 16590 4 gnd
port 514 nsew
rlabel metal2 s 29712 18170 29712 18170 4 gnd
port 514 nsew
rlabel metal2 s 27696 18960 27696 18960 4 gnd
port 514 nsew
rlabel metal2 s 29712 16353 29712 16353 4 gnd
port 514 nsew
rlabel metal2 s 29712 16037 29712 16037 4 gnd
port 514 nsew
rlabel metal2 s 28464 18170 28464 18170 4 gnd
port 514 nsew
rlabel metal2 s 28464 17380 28464 17380 4 gnd
port 514 nsew
rlabel metal2 s 28944 16590 28944 16590 4 gnd
port 514 nsew
rlabel metal2 s 29712 16827 29712 16827 4 gnd
port 514 nsew
rlabel metal2 s 27696 17617 27696 17617 4 gnd
port 514 nsew
rlabel metal2 s 28944 18960 28944 18960 4 gnd
port 514 nsew
rlabel metal2 s 28944 17143 28944 17143 4 gnd
port 514 nsew
rlabel metal2 s 29712 18960 29712 18960 4 gnd
port 514 nsew
rlabel metal2 s 27696 18723 27696 18723 4 gnd
port 514 nsew
rlabel metal2 s 28944 17933 28944 17933 4 gnd
port 514 nsew
rlabel metal2 s 29712 17380 29712 17380 4 gnd
port 514 nsew
rlabel metal2 s 28944 16037 28944 16037 4 gnd
port 514 nsew
rlabel metal2 s 27696 17380 27696 17380 4 gnd
port 514 nsew
rlabel metal2 s 27696 16353 27696 16353 4 gnd
port 514 nsew
rlabel metal2 s 28464 16827 28464 16827 4 gnd
port 514 nsew
rlabel metal2 s 29712 18407 29712 18407 4 gnd
port 514 nsew
rlabel metal2 s 28944 18723 28944 18723 4 gnd
port 514 nsew
rlabel metal2 s 29712 17617 29712 17617 4 gnd
port 514 nsew
rlabel metal2 s 28944 16353 28944 16353 4 gnd
port 514 nsew
rlabel metal2 s 29712 16590 29712 16590 4 gnd
port 514 nsew
rlabel metal2 s 27696 18407 27696 18407 4 gnd
port 514 nsew
rlabel metal2 s 28464 16353 28464 16353 4 gnd
port 514 nsew
rlabel metal2 s 29712 17933 29712 17933 4 gnd
port 514 nsew
rlabel metal2 s 28464 18960 28464 18960 4 gnd
port 514 nsew
rlabel metal2 s 27696 17143 27696 17143 4 gnd
port 514 nsew
rlabel metal2 s 27696 16037 27696 16037 4 gnd
port 514 nsew
rlabel metal2 s 28464 16590 28464 16590 4 gnd
port 514 nsew
rlabel metal2 s 28944 17617 28944 17617 4 gnd
port 514 nsew
rlabel metal2 s 28464 17933 28464 17933 4 gnd
port 514 nsew
rlabel metal2 s 28944 16827 28944 16827 4 gnd
port 514 nsew
rlabel metal2 s 26448 18723 26448 18723 4 gnd
port 514 nsew
rlabel metal2 s 26448 16353 26448 16353 4 gnd
port 514 nsew
rlabel metal2 s 25200 16353 25200 16353 4 gnd
port 514 nsew
rlabel metal2 s 27216 18170 27216 18170 4 gnd
port 514 nsew
rlabel metal2 s 25968 16037 25968 16037 4 gnd
port 514 nsew
rlabel metal2 s 26448 17617 26448 17617 4 gnd
port 514 nsew
rlabel metal2 s 25968 17143 25968 17143 4 gnd
port 514 nsew
rlabel metal2 s 26448 18960 26448 18960 4 gnd
port 514 nsew
rlabel metal2 s 25968 16827 25968 16827 4 gnd
port 514 nsew
rlabel metal2 s 27216 17143 27216 17143 4 gnd
port 514 nsew
rlabel metal2 s 25968 18407 25968 18407 4 gnd
port 514 nsew
rlabel metal2 s 27216 17380 27216 17380 4 gnd
port 514 nsew
rlabel metal2 s 25968 18170 25968 18170 4 gnd
port 514 nsew
rlabel metal2 s 25968 18960 25968 18960 4 gnd
port 514 nsew
rlabel metal2 s 27216 18960 27216 18960 4 gnd
port 514 nsew
rlabel metal2 s 26448 18170 26448 18170 4 gnd
port 514 nsew
rlabel metal2 s 25968 18723 25968 18723 4 gnd
port 514 nsew
rlabel metal2 s 25200 16590 25200 16590 4 gnd
port 514 nsew
rlabel metal2 s 25200 17143 25200 17143 4 gnd
port 514 nsew
rlabel metal2 s 26448 16590 26448 16590 4 gnd
port 514 nsew
rlabel metal2 s 27216 16353 27216 16353 4 gnd
port 514 nsew
rlabel metal2 s 25968 16590 25968 16590 4 gnd
port 514 nsew
rlabel metal2 s 25968 17933 25968 17933 4 gnd
port 514 nsew
rlabel metal2 s 27216 16827 27216 16827 4 gnd
port 514 nsew
rlabel metal2 s 25200 16037 25200 16037 4 gnd
port 514 nsew
rlabel metal2 s 26448 16037 26448 16037 4 gnd
port 514 nsew
rlabel metal2 s 25968 17617 25968 17617 4 gnd
port 514 nsew
rlabel metal2 s 25200 18960 25200 18960 4 gnd
port 514 nsew
rlabel metal2 s 25200 18407 25200 18407 4 gnd
port 514 nsew
rlabel metal2 s 27216 18723 27216 18723 4 gnd
port 514 nsew
rlabel metal2 s 25968 17380 25968 17380 4 gnd
port 514 nsew
rlabel metal2 s 27216 16037 27216 16037 4 gnd
port 514 nsew
rlabel metal2 s 25200 17933 25200 17933 4 gnd
port 514 nsew
rlabel metal2 s 26448 17933 26448 17933 4 gnd
port 514 nsew
rlabel metal2 s 25200 18723 25200 18723 4 gnd
port 514 nsew
rlabel metal2 s 26448 17380 26448 17380 4 gnd
port 514 nsew
rlabel metal2 s 25200 18170 25200 18170 4 gnd
port 514 nsew
rlabel metal2 s 27216 17933 27216 17933 4 gnd
port 514 nsew
rlabel metal2 s 26448 17143 26448 17143 4 gnd
port 514 nsew
rlabel metal2 s 25200 17617 25200 17617 4 gnd
port 514 nsew
rlabel metal2 s 27216 17617 27216 17617 4 gnd
port 514 nsew
rlabel metal2 s 27216 18407 27216 18407 4 gnd
port 514 nsew
rlabel metal2 s 26448 18407 26448 18407 4 gnd
port 514 nsew
rlabel metal2 s 26448 16827 26448 16827 4 gnd
port 514 nsew
rlabel metal2 s 27216 16590 27216 16590 4 gnd
port 514 nsew
rlabel metal2 s 25200 16827 25200 16827 4 gnd
port 514 nsew
rlabel metal2 s 25200 17380 25200 17380 4 gnd
port 514 nsew
rlabel metal2 s 25968 16353 25968 16353 4 gnd
port 514 nsew
rlabel metal2 s 25200 15247 25200 15247 4 gnd
port 514 nsew
rlabel metal2 s 27216 15010 27216 15010 4 gnd
port 514 nsew
rlabel metal2 s 26448 14457 26448 14457 4 gnd
port 514 nsew
rlabel metal2 s 26448 15563 26448 15563 4 gnd
port 514 nsew
rlabel metal2 s 25200 13193 25200 13193 4 gnd
port 514 nsew
rlabel metal2 s 25968 12877 25968 12877 4 gnd
port 514 nsew
rlabel metal2 s 27216 13193 27216 13193 4 gnd
port 514 nsew
rlabel metal2 s 25968 13667 25968 13667 4 gnd
port 514 nsew
rlabel metal2 s 27216 13430 27216 13430 4 gnd
port 514 nsew
rlabel metal2 s 26448 15800 26448 15800 4 gnd
port 514 nsew
rlabel metal2 s 27216 12877 27216 12877 4 gnd
port 514 nsew
rlabel metal2 s 25968 14457 25968 14457 4 gnd
port 514 nsew
rlabel metal2 s 27216 15563 27216 15563 4 gnd
port 514 nsew
rlabel metal2 s 25968 15010 25968 15010 4 gnd
port 514 nsew
rlabel metal2 s 26448 14773 26448 14773 4 gnd
port 514 nsew
rlabel metal2 s 27216 14220 27216 14220 4 gnd
port 514 nsew
rlabel metal2 s 26448 13193 26448 13193 4 gnd
port 514 nsew
rlabel metal2 s 26448 13667 26448 13667 4 gnd
port 514 nsew
rlabel metal2 s 26448 15247 26448 15247 4 gnd
port 514 nsew
rlabel metal2 s 26448 12877 26448 12877 4 gnd
port 514 nsew
rlabel metal2 s 26448 14220 26448 14220 4 gnd
port 514 nsew
rlabel metal2 s 26448 15010 26448 15010 4 gnd
port 514 nsew
rlabel metal2 s 25968 13193 25968 13193 4 gnd
port 514 nsew
rlabel metal2 s 25200 12877 25200 12877 4 gnd
port 514 nsew
rlabel metal2 s 25968 13983 25968 13983 4 gnd
port 514 nsew
rlabel metal2 s 27216 15800 27216 15800 4 gnd
port 514 nsew
rlabel metal2 s 25968 14220 25968 14220 4 gnd
port 514 nsew
rlabel metal2 s 27216 13667 27216 13667 4 gnd
port 514 nsew
rlabel metal2 s 26448 13983 26448 13983 4 gnd
port 514 nsew
rlabel metal2 s 25968 15563 25968 15563 4 gnd
port 514 nsew
rlabel metal2 s 25200 15800 25200 15800 4 gnd
port 514 nsew
rlabel metal2 s 25200 13430 25200 13430 4 gnd
port 514 nsew
rlabel metal2 s 27216 14457 27216 14457 4 gnd
port 514 nsew
rlabel metal2 s 27216 15247 27216 15247 4 gnd
port 514 nsew
rlabel metal2 s 25200 15563 25200 15563 4 gnd
port 514 nsew
rlabel metal2 s 25200 13983 25200 13983 4 gnd
port 514 nsew
rlabel metal2 s 25968 14773 25968 14773 4 gnd
port 514 nsew
rlabel metal2 s 25200 14220 25200 14220 4 gnd
port 514 nsew
rlabel metal2 s 27216 14773 27216 14773 4 gnd
port 514 nsew
rlabel metal2 s 27216 13983 27216 13983 4 gnd
port 514 nsew
rlabel metal2 s 25968 15800 25968 15800 4 gnd
port 514 nsew
rlabel metal2 s 25968 15247 25968 15247 4 gnd
port 514 nsew
rlabel metal2 s 25200 14773 25200 14773 4 gnd
port 514 nsew
rlabel metal2 s 25968 13430 25968 13430 4 gnd
port 514 nsew
rlabel metal2 s 25200 14457 25200 14457 4 gnd
port 514 nsew
rlabel metal2 s 25200 13667 25200 13667 4 gnd
port 514 nsew
rlabel metal2 s 25200 15010 25200 15010 4 gnd
port 514 nsew
rlabel metal2 s 26448 13430 26448 13430 4 gnd
port 514 nsew
rlabel metal2 s 29712 14773 29712 14773 4 gnd
port 514 nsew
rlabel metal2 s 28464 14220 28464 14220 4 gnd
port 514 nsew
rlabel metal2 s 28464 13667 28464 13667 4 gnd
port 514 nsew
rlabel metal2 s 28944 12877 28944 12877 4 gnd
port 514 nsew
rlabel metal2 s 29712 14457 29712 14457 4 gnd
port 514 nsew
rlabel metal2 s 28464 13430 28464 13430 4 gnd
port 514 nsew
rlabel metal2 s 27696 13667 27696 13667 4 gnd
port 514 nsew
rlabel metal2 s 27696 13430 27696 13430 4 gnd
port 514 nsew
rlabel metal2 s 28944 14773 28944 14773 4 gnd
port 514 nsew
rlabel metal2 s 29712 15010 29712 15010 4 gnd
port 514 nsew
rlabel metal2 s 28944 15010 28944 15010 4 gnd
port 514 nsew
rlabel metal2 s 29712 15800 29712 15800 4 gnd
port 514 nsew
rlabel metal2 s 28944 13667 28944 13667 4 gnd
port 514 nsew
rlabel metal2 s 29712 15247 29712 15247 4 gnd
port 514 nsew
rlabel metal2 s 27696 13983 27696 13983 4 gnd
port 514 nsew
rlabel metal2 s 29712 13193 29712 13193 4 gnd
port 514 nsew
rlabel metal2 s 29712 15563 29712 15563 4 gnd
port 514 nsew
rlabel metal2 s 27696 14773 27696 14773 4 gnd
port 514 nsew
rlabel metal2 s 28464 13193 28464 13193 4 gnd
port 514 nsew
rlabel metal2 s 28944 15247 28944 15247 4 gnd
port 514 nsew
rlabel metal2 s 27696 13193 27696 13193 4 gnd
port 514 nsew
rlabel metal2 s 28944 13430 28944 13430 4 gnd
port 514 nsew
rlabel metal2 s 28464 15563 28464 15563 4 gnd
port 514 nsew
rlabel metal2 s 28944 13193 28944 13193 4 gnd
port 514 nsew
rlabel metal2 s 28464 14773 28464 14773 4 gnd
port 514 nsew
rlabel metal2 s 27696 14457 27696 14457 4 gnd
port 514 nsew
rlabel metal2 s 28464 13983 28464 13983 4 gnd
port 514 nsew
rlabel metal2 s 29712 13430 29712 13430 4 gnd
port 514 nsew
rlabel metal2 s 27696 15563 27696 15563 4 gnd
port 514 nsew
rlabel metal2 s 29712 12877 29712 12877 4 gnd
port 514 nsew
rlabel metal2 s 29712 13983 29712 13983 4 gnd
port 514 nsew
rlabel metal2 s 29712 13667 29712 13667 4 gnd
port 514 nsew
rlabel metal2 s 28944 15800 28944 15800 4 gnd
port 514 nsew
rlabel metal2 s 28464 14457 28464 14457 4 gnd
port 514 nsew
rlabel metal2 s 27696 12877 27696 12877 4 gnd
port 514 nsew
rlabel metal2 s 28464 15010 28464 15010 4 gnd
port 514 nsew
rlabel metal2 s 27696 14220 27696 14220 4 gnd
port 514 nsew
rlabel metal2 s 27696 15010 27696 15010 4 gnd
port 514 nsew
rlabel metal2 s 28944 15563 28944 15563 4 gnd
port 514 nsew
rlabel metal2 s 29712 14220 29712 14220 4 gnd
port 514 nsew
rlabel metal2 s 28464 12877 28464 12877 4 gnd
port 514 nsew
rlabel metal2 s 27696 15800 27696 15800 4 gnd
port 514 nsew
rlabel metal2 s 28944 14220 28944 14220 4 gnd
port 514 nsew
rlabel metal2 s 27696 15247 27696 15247 4 gnd
port 514 nsew
rlabel metal2 s 28464 15800 28464 15800 4 gnd
port 514 nsew
rlabel metal2 s 28944 13983 28944 13983 4 gnd
port 514 nsew
rlabel metal2 s 28944 14457 28944 14457 4 gnd
port 514 nsew
rlabel metal2 s 28464 15247 28464 15247 4 gnd
port 514 nsew
rlabel metal2 s 27696 10270 27696 10270 4 gnd
port 514 nsew
rlabel metal2 s 28944 11060 28944 11060 4 gnd
port 514 nsew
rlabel metal2 s 28944 11850 28944 11850 4 gnd
port 514 nsew
rlabel metal2 s 27696 10823 27696 10823 4 gnd
port 514 nsew
rlabel metal2 s 28464 12640 28464 12640 4 gnd
port 514 nsew
rlabel metal2 s 27696 10507 27696 10507 4 gnd
port 514 nsew
rlabel metal2 s 28944 12403 28944 12403 4 gnd
port 514 nsew
rlabel metal2 s 28944 9717 28944 9717 4 gnd
port 514 nsew
rlabel metal2 s 28464 12087 28464 12087 4 gnd
port 514 nsew
rlabel metal2 s 29712 10507 29712 10507 4 gnd
port 514 nsew
rlabel metal2 s 28464 11613 28464 11613 4 gnd
port 514 nsew
rlabel metal2 s 27696 11850 27696 11850 4 gnd
port 514 nsew
rlabel metal2 s 28944 11613 28944 11613 4 gnd
port 514 nsew
rlabel metal2 s 27696 12087 27696 12087 4 gnd
port 514 nsew
rlabel metal2 s 28464 12403 28464 12403 4 gnd
port 514 nsew
rlabel metal2 s 29712 12640 29712 12640 4 gnd
port 514 nsew
rlabel metal2 s 28944 11297 28944 11297 4 gnd
port 514 nsew
rlabel metal2 s 29712 10270 29712 10270 4 gnd
port 514 nsew
rlabel metal2 s 29712 11297 29712 11297 4 gnd
port 514 nsew
rlabel metal2 s 28464 11850 28464 11850 4 gnd
port 514 nsew
rlabel metal2 s 28944 10270 28944 10270 4 gnd
port 514 nsew
rlabel metal2 s 29712 10823 29712 10823 4 gnd
port 514 nsew
rlabel metal2 s 27696 11297 27696 11297 4 gnd
port 514 nsew
rlabel metal2 s 27696 11613 27696 11613 4 gnd
port 514 nsew
rlabel metal2 s 28464 10033 28464 10033 4 gnd
port 514 nsew
rlabel metal2 s 28944 12087 28944 12087 4 gnd
port 514 nsew
rlabel metal2 s 28944 12640 28944 12640 4 gnd
port 514 nsew
rlabel metal2 s 28464 11297 28464 11297 4 gnd
port 514 nsew
rlabel metal2 s 27696 12640 27696 12640 4 gnd
port 514 nsew
rlabel metal2 s 27696 10033 27696 10033 4 gnd
port 514 nsew
rlabel metal2 s 27696 11060 27696 11060 4 gnd
port 514 nsew
rlabel metal2 s 29712 9717 29712 9717 4 gnd
port 514 nsew
rlabel metal2 s 29712 11060 29712 11060 4 gnd
port 514 nsew
rlabel metal2 s 29712 12403 29712 12403 4 gnd
port 514 nsew
rlabel metal2 s 29712 11613 29712 11613 4 gnd
port 514 nsew
rlabel metal2 s 28464 11060 28464 11060 4 gnd
port 514 nsew
rlabel metal2 s 28944 10033 28944 10033 4 gnd
port 514 nsew
rlabel metal2 s 28464 10823 28464 10823 4 gnd
port 514 nsew
rlabel metal2 s 29712 11850 29712 11850 4 gnd
port 514 nsew
rlabel metal2 s 28464 9717 28464 9717 4 gnd
port 514 nsew
rlabel metal2 s 27696 12403 27696 12403 4 gnd
port 514 nsew
rlabel metal2 s 28464 10507 28464 10507 4 gnd
port 514 nsew
rlabel metal2 s 29712 12087 29712 12087 4 gnd
port 514 nsew
rlabel metal2 s 27696 9717 27696 9717 4 gnd
port 514 nsew
rlabel metal2 s 28944 10507 28944 10507 4 gnd
port 514 nsew
rlabel metal2 s 29712 10033 29712 10033 4 gnd
port 514 nsew
rlabel metal2 s 28944 10823 28944 10823 4 gnd
port 514 nsew
rlabel metal2 s 28464 10270 28464 10270 4 gnd
port 514 nsew
rlabel metal2 s 25200 12640 25200 12640 4 gnd
port 514 nsew
rlabel metal2 s 25968 12640 25968 12640 4 gnd
port 514 nsew
rlabel metal2 s 27216 11297 27216 11297 4 gnd
port 514 nsew
rlabel metal2 s 25968 10823 25968 10823 4 gnd
port 514 nsew
rlabel metal2 s 27216 11613 27216 11613 4 gnd
port 514 nsew
rlabel metal2 s 27216 12403 27216 12403 4 gnd
port 514 nsew
rlabel metal2 s 26448 10507 26448 10507 4 gnd
port 514 nsew
rlabel metal2 s 25200 11060 25200 11060 4 gnd
port 514 nsew
rlabel metal2 s 27216 11850 27216 11850 4 gnd
port 514 nsew
rlabel metal2 s 25200 11613 25200 11613 4 gnd
port 514 nsew
rlabel metal2 s 26448 11613 26448 11613 4 gnd
port 514 nsew
rlabel metal2 s 26448 12640 26448 12640 4 gnd
port 514 nsew
rlabel metal2 s 27216 11060 27216 11060 4 gnd
port 514 nsew
rlabel metal2 s 25200 9717 25200 9717 4 gnd
port 514 nsew
rlabel metal2 s 27216 9717 27216 9717 4 gnd
port 514 nsew
rlabel metal2 s 26448 10270 26448 10270 4 gnd
port 514 nsew
rlabel metal2 s 26448 11297 26448 11297 4 gnd
port 514 nsew
rlabel metal2 s 25200 12403 25200 12403 4 gnd
port 514 nsew
rlabel metal2 s 27216 10270 27216 10270 4 gnd
port 514 nsew
rlabel metal2 s 27216 10823 27216 10823 4 gnd
port 514 nsew
rlabel metal2 s 25200 10507 25200 10507 4 gnd
port 514 nsew
rlabel metal2 s 26448 12403 26448 12403 4 gnd
port 514 nsew
rlabel metal2 s 26448 12087 26448 12087 4 gnd
port 514 nsew
rlabel metal2 s 25968 12087 25968 12087 4 gnd
port 514 nsew
rlabel metal2 s 26448 11060 26448 11060 4 gnd
port 514 nsew
rlabel metal2 s 27216 10507 27216 10507 4 gnd
port 514 nsew
rlabel metal2 s 26448 10823 26448 10823 4 gnd
port 514 nsew
rlabel metal2 s 25200 12087 25200 12087 4 gnd
port 514 nsew
rlabel metal2 s 25968 11297 25968 11297 4 gnd
port 514 nsew
rlabel metal2 s 25968 12403 25968 12403 4 gnd
port 514 nsew
rlabel metal2 s 25968 10270 25968 10270 4 gnd
port 514 nsew
rlabel metal2 s 25200 10823 25200 10823 4 gnd
port 514 nsew
rlabel metal2 s 25968 11850 25968 11850 4 gnd
port 514 nsew
rlabel metal2 s 25200 11850 25200 11850 4 gnd
port 514 nsew
rlabel metal2 s 26448 9717 26448 9717 4 gnd
port 514 nsew
rlabel metal2 s 25968 9717 25968 9717 4 gnd
port 514 nsew
rlabel metal2 s 26448 11850 26448 11850 4 gnd
port 514 nsew
rlabel metal2 s 25200 10270 25200 10270 4 gnd
port 514 nsew
rlabel metal2 s 26448 10033 26448 10033 4 gnd
port 514 nsew
rlabel metal2 s 25968 11613 25968 11613 4 gnd
port 514 nsew
rlabel metal2 s 27216 12087 27216 12087 4 gnd
port 514 nsew
rlabel metal2 s 25968 10033 25968 10033 4 gnd
port 514 nsew
rlabel metal2 s 25968 11060 25968 11060 4 gnd
port 514 nsew
rlabel metal2 s 27216 12640 27216 12640 4 gnd
port 514 nsew
rlabel metal2 s 25200 11297 25200 11297 4 gnd
port 514 nsew
rlabel metal2 s 25200 10033 25200 10033 4 gnd
port 514 nsew
rlabel metal2 s 25968 10507 25968 10507 4 gnd
port 514 nsew
rlabel metal2 s 27216 10033 27216 10033 4 gnd
port 514 nsew
rlabel metal2 s 26448 8137 26448 8137 4 gnd
port 514 nsew
rlabel metal2 s 27216 9243 27216 9243 4 gnd
port 514 nsew
rlabel metal2 s 25200 8927 25200 8927 4 gnd
port 514 nsew
rlabel metal2 s 25968 8137 25968 8137 4 gnd
port 514 nsew
rlabel metal2 s 27216 8690 27216 8690 4 gnd
port 514 nsew
rlabel metal2 s 25200 8453 25200 8453 4 gnd
port 514 nsew
rlabel metal2 s 26448 6873 26448 6873 4 gnd
port 514 nsew
rlabel metal2 s 25200 9243 25200 9243 4 gnd
port 514 nsew
rlabel metal2 s 25968 6557 25968 6557 4 gnd
port 514 nsew
rlabel metal2 s 25200 7663 25200 7663 4 gnd
port 514 nsew
rlabel metal2 s 25968 7900 25968 7900 4 gnd
port 514 nsew
rlabel metal2 s 27216 7347 27216 7347 4 gnd
port 514 nsew
rlabel metal2 s 27216 7110 27216 7110 4 gnd
port 514 nsew
rlabel metal2 s 25968 7663 25968 7663 4 gnd
port 514 nsew
rlabel metal2 s 27216 8453 27216 8453 4 gnd
port 514 nsew
rlabel metal2 s 27216 8927 27216 8927 4 gnd
port 514 nsew
rlabel metal2 s 25200 6873 25200 6873 4 gnd
port 514 nsew
rlabel metal2 s 26448 8453 26448 8453 4 gnd
port 514 nsew
rlabel metal2 s 26448 7110 26448 7110 4 gnd
port 514 nsew
rlabel metal2 s 25968 7347 25968 7347 4 gnd
port 514 nsew
rlabel metal2 s 26448 8690 26448 8690 4 gnd
port 514 nsew
rlabel metal2 s 27216 8137 27216 8137 4 gnd
port 514 nsew
rlabel metal2 s 25200 6557 25200 6557 4 gnd
port 514 nsew
rlabel metal2 s 25968 9243 25968 9243 4 gnd
port 514 nsew
rlabel metal2 s 25200 8137 25200 8137 4 gnd
port 514 nsew
rlabel metal2 s 27216 6873 27216 6873 4 gnd
port 514 nsew
rlabel metal2 s 27216 7900 27216 7900 4 gnd
port 514 nsew
rlabel metal2 s 26448 7663 26448 7663 4 gnd
port 514 nsew
rlabel metal2 s 25968 8453 25968 8453 4 gnd
port 514 nsew
rlabel metal2 s 26448 6557 26448 6557 4 gnd
port 514 nsew
rlabel metal2 s 25200 7347 25200 7347 4 gnd
port 514 nsew
rlabel metal2 s 25968 8927 25968 8927 4 gnd
port 514 nsew
rlabel metal2 s 27216 9480 27216 9480 4 gnd
port 514 nsew
rlabel metal2 s 27216 7663 27216 7663 4 gnd
port 514 nsew
rlabel metal2 s 26448 7347 26448 7347 4 gnd
port 514 nsew
rlabel metal2 s 25968 8690 25968 8690 4 gnd
port 514 nsew
rlabel metal2 s 26448 7900 26448 7900 4 gnd
port 514 nsew
rlabel metal2 s 26448 9243 26448 9243 4 gnd
port 514 nsew
rlabel metal2 s 25200 7900 25200 7900 4 gnd
port 514 nsew
rlabel metal2 s 25968 7110 25968 7110 4 gnd
port 514 nsew
rlabel metal2 s 25968 6873 25968 6873 4 gnd
port 514 nsew
rlabel metal2 s 27216 6557 27216 6557 4 gnd
port 514 nsew
rlabel metal2 s 25200 9480 25200 9480 4 gnd
port 514 nsew
rlabel metal2 s 26448 8927 26448 8927 4 gnd
port 514 nsew
rlabel metal2 s 26448 9480 26448 9480 4 gnd
port 514 nsew
rlabel metal2 s 25968 9480 25968 9480 4 gnd
port 514 nsew
rlabel metal2 s 25200 8690 25200 8690 4 gnd
port 514 nsew
rlabel metal2 s 25200 7110 25200 7110 4 gnd
port 514 nsew
rlabel metal2 s 28944 7663 28944 7663 4 gnd
port 514 nsew
rlabel metal2 s 28464 8137 28464 8137 4 gnd
port 514 nsew
rlabel metal2 s 29712 7110 29712 7110 4 gnd
port 514 nsew
rlabel metal2 s 29712 7900 29712 7900 4 gnd
port 514 nsew
rlabel metal2 s 27696 8137 27696 8137 4 gnd
port 514 nsew
rlabel metal2 s 29712 8927 29712 8927 4 gnd
port 514 nsew
rlabel metal2 s 28944 8137 28944 8137 4 gnd
port 514 nsew
rlabel metal2 s 28464 7663 28464 7663 4 gnd
port 514 nsew
rlabel metal2 s 28464 6873 28464 6873 4 gnd
port 514 nsew
rlabel metal2 s 27696 7900 27696 7900 4 gnd
port 514 nsew
rlabel metal2 s 29712 8453 29712 8453 4 gnd
port 514 nsew
rlabel metal2 s 28944 9480 28944 9480 4 gnd
port 514 nsew
rlabel metal2 s 28944 7347 28944 7347 4 gnd
port 514 nsew
rlabel metal2 s 28464 7110 28464 7110 4 gnd
port 514 nsew
rlabel metal2 s 28464 6557 28464 6557 4 gnd
port 514 nsew
rlabel metal2 s 28464 8927 28464 8927 4 gnd
port 514 nsew
rlabel metal2 s 29712 8137 29712 8137 4 gnd
port 514 nsew
rlabel metal2 s 28944 8453 28944 8453 4 gnd
port 514 nsew
rlabel metal2 s 28944 6557 28944 6557 4 gnd
port 514 nsew
rlabel metal2 s 28464 7900 28464 7900 4 gnd
port 514 nsew
rlabel metal2 s 29712 7347 29712 7347 4 gnd
port 514 nsew
rlabel metal2 s 28944 7900 28944 7900 4 gnd
port 514 nsew
rlabel metal2 s 27696 7110 27696 7110 4 gnd
port 514 nsew
rlabel metal2 s 29712 6873 29712 6873 4 gnd
port 514 nsew
rlabel metal2 s 29712 6557 29712 6557 4 gnd
port 514 nsew
rlabel metal2 s 27696 7347 27696 7347 4 gnd
port 514 nsew
rlabel metal2 s 28464 9480 28464 9480 4 gnd
port 514 nsew
rlabel metal2 s 28464 9243 28464 9243 4 gnd
port 514 nsew
rlabel metal2 s 28944 9243 28944 9243 4 gnd
port 514 nsew
rlabel metal2 s 27696 9480 27696 9480 4 gnd
port 514 nsew
rlabel metal2 s 27696 6873 27696 6873 4 gnd
port 514 nsew
rlabel metal2 s 29712 8690 29712 8690 4 gnd
port 514 nsew
rlabel metal2 s 28464 8453 28464 8453 4 gnd
port 514 nsew
rlabel metal2 s 27696 6557 27696 6557 4 gnd
port 514 nsew
rlabel metal2 s 28944 6873 28944 6873 4 gnd
port 514 nsew
rlabel metal2 s 27696 8453 27696 8453 4 gnd
port 514 nsew
rlabel metal2 s 29712 9480 29712 9480 4 gnd
port 514 nsew
rlabel metal2 s 29712 9243 29712 9243 4 gnd
port 514 nsew
rlabel metal2 s 28464 8690 28464 8690 4 gnd
port 514 nsew
rlabel metal2 s 28944 8927 28944 8927 4 gnd
port 514 nsew
rlabel metal2 s 28464 7347 28464 7347 4 gnd
port 514 nsew
rlabel metal2 s 27696 8690 27696 8690 4 gnd
port 514 nsew
rlabel metal2 s 28944 7110 28944 7110 4 gnd
port 514 nsew
rlabel metal2 s 27696 8927 27696 8927 4 gnd
port 514 nsew
rlabel metal2 s 29712 7663 29712 7663 4 gnd
port 514 nsew
rlabel metal2 s 27696 9243 27696 9243 4 gnd
port 514 nsew
rlabel metal2 s 27696 7663 27696 7663 4 gnd
port 514 nsew
rlabel metal2 s 28944 8690 28944 8690 4 gnd
port 514 nsew
rlabel metal2 s 24720 9717 24720 9717 4 gnd
port 514 nsew
rlabel metal2 s 23472 10507 23472 10507 4 gnd
port 514 nsew
rlabel metal2 s 24720 10270 24720 10270 4 gnd
port 514 nsew
rlabel metal2 s 23472 10033 23472 10033 4 gnd
port 514 nsew
rlabel metal2 s 24720 11850 24720 11850 4 gnd
port 514 nsew
rlabel metal2 s 23472 12087 23472 12087 4 gnd
port 514 nsew
rlabel metal2 s 23472 11613 23472 11613 4 gnd
port 514 nsew
rlabel metal2 s 23952 10823 23952 10823 4 gnd
port 514 nsew
rlabel metal2 s 23952 10033 23952 10033 4 gnd
port 514 nsew
rlabel metal2 s 24720 12403 24720 12403 4 gnd
port 514 nsew
rlabel metal2 s 22704 11060 22704 11060 4 gnd
port 514 nsew
rlabel metal2 s 23472 10270 23472 10270 4 gnd
port 514 nsew
rlabel metal2 s 23952 11060 23952 11060 4 gnd
port 514 nsew
rlabel metal2 s 22704 12087 22704 12087 4 gnd
port 514 nsew
rlabel metal2 s 23952 11613 23952 11613 4 gnd
port 514 nsew
rlabel metal2 s 22704 11613 22704 11613 4 gnd
port 514 nsew
rlabel metal2 s 23952 9717 23952 9717 4 gnd
port 514 nsew
rlabel metal2 s 22704 10507 22704 10507 4 gnd
port 514 nsew
rlabel metal2 s 23472 12640 23472 12640 4 gnd
port 514 nsew
rlabel metal2 s 23952 12087 23952 12087 4 gnd
port 514 nsew
rlabel metal2 s 22704 11297 22704 11297 4 gnd
port 514 nsew
rlabel metal2 s 22704 10033 22704 10033 4 gnd
port 514 nsew
rlabel metal2 s 24720 11297 24720 11297 4 gnd
port 514 nsew
rlabel metal2 s 22704 10823 22704 10823 4 gnd
port 514 nsew
rlabel metal2 s 23472 11297 23472 11297 4 gnd
port 514 nsew
rlabel metal2 s 23472 11060 23472 11060 4 gnd
port 514 nsew
rlabel metal2 s 22704 12640 22704 12640 4 gnd
port 514 nsew
rlabel metal2 s 22704 12403 22704 12403 4 gnd
port 514 nsew
rlabel metal2 s 23952 12640 23952 12640 4 gnd
port 514 nsew
rlabel metal2 s 23952 11850 23952 11850 4 gnd
port 514 nsew
rlabel metal2 s 23952 11297 23952 11297 4 gnd
port 514 nsew
rlabel metal2 s 24720 12640 24720 12640 4 gnd
port 514 nsew
rlabel metal2 s 23952 10507 23952 10507 4 gnd
port 514 nsew
rlabel metal2 s 22704 11850 22704 11850 4 gnd
port 514 nsew
rlabel metal2 s 24720 12087 24720 12087 4 gnd
port 514 nsew
rlabel metal2 s 22704 9717 22704 9717 4 gnd
port 514 nsew
rlabel metal2 s 23472 12403 23472 12403 4 gnd
port 514 nsew
rlabel metal2 s 23952 10270 23952 10270 4 gnd
port 514 nsew
rlabel metal2 s 24720 10823 24720 10823 4 gnd
port 514 nsew
rlabel metal2 s 23952 12403 23952 12403 4 gnd
port 514 nsew
rlabel metal2 s 24720 10507 24720 10507 4 gnd
port 514 nsew
rlabel metal2 s 24720 11060 24720 11060 4 gnd
port 514 nsew
rlabel metal2 s 23472 10823 23472 10823 4 gnd
port 514 nsew
rlabel metal2 s 24720 10033 24720 10033 4 gnd
port 514 nsew
rlabel metal2 s 22704 10270 22704 10270 4 gnd
port 514 nsew
rlabel metal2 s 24720 11613 24720 11613 4 gnd
port 514 nsew
rlabel metal2 s 23472 9717 23472 9717 4 gnd
port 514 nsew
rlabel metal2 s 23472 11850 23472 11850 4 gnd
port 514 nsew
rlabel metal2 s 20208 12087 20208 12087 4 gnd
port 514 nsew
rlabel metal2 s 21456 11297 21456 11297 4 gnd
port 514 nsew
rlabel metal2 s 22224 11297 22224 11297 4 gnd
port 514 nsew
rlabel metal2 s 21456 11850 21456 11850 4 gnd
port 514 nsew
rlabel metal2 s 21456 11613 21456 11613 4 gnd
port 514 nsew
rlabel metal2 s 20208 10823 20208 10823 4 gnd
port 514 nsew
rlabel metal2 s 20976 10507 20976 10507 4 gnd
port 514 nsew
rlabel metal2 s 22224 11850 22224 11850 4 gnd
port 514 nsew
rlabel metal2 s 22224 12087 22224 12087 4 gnd
port 514 nsew
rlabel metal2 s 21456 11060 21456 11060 4 gnd
port 514 nsew
rlabel metal2 s 22224 10033 22224 10033 4 gnd
port 514 nsew
rlabel metal2 s 20976 11297 20976 11297 4 gnd
port 514 nsew
rlabel metal2 s 20208 11850 20208 11850 4 gnd
port 514 nsew
rlabel metal2 s 21456 9717 21456 9717 4 gnd
port 514 nsew
rlabel metal2 s 20976 10270 20976 10270 4 gnd
port 514 nsew
rlabel metal2 s 20208 10033 20208 10033 4 gnd
port 514 nsew
rlabel metal2 s 20208 11297 20208 11297 4 gnd
port 514 nsew
rlabel metal2 s 21456 10507 21456 10507 4 gnd
port 514 nsew
rlabel metal2 s 22224 10270 22224 10270 4 gnd
port 514 nsew
rlabel metal2 s 22224 11060 22224 11060 4 gnd
port 514 nsew
rlabel metal2 s 22224 12640 22224 12640 4 gnd
port 514 nsew
rlabel metal2 s 20976 12403 20976 12403 4 gnd
port 514 nsew
rlabel metal2 s 20976 12087 20976 12087 4 gnd
port 514 nsew
rlabel metal2 s 20976 9717 20976 9717 4 gnd
port 514 nsew
rlabel metal2 s 21456 12640 21456 12640 4 gnd
port 514 nsew
rlabel metal2 s 21456 12403 21456 12403 4 gnd
port 514 nsew
rlabel metal2 s 22224 9717 22224 9717 4 gnd
port 514 nsew
rlabel metal2 s 21456 12087 21456 12087 4 gnd
port 514 nsew
rlabel metal2 s 22224 11613 22224 11613 4 gnd
port 514 nsew
rlabel metal2 s 20976 10823 20976 10823 4 gnd
port 514 nsew
rlabel metal2 s 20208 9717 20208 9717 4 gnd
port 514 nsew
rlabel metal2 s 20208 10270 20208 10270 4 gnd
port 514 nsew
rlabel metal2 s 20976 10033 20976 10033 4 gnd
port 514 nsew
rlabel metal2 s 22224 12403 22224 12403 4 gnd
port 514 nsew
rlabel metal2 s 20208 10507 20208 10507 4 gnd
port 514 nsew
rlabel metal2 s 20208 12640 20208 12640 4 gnd
port 514 nsew
rlabel metal2 s 22224 10823 22224 10823 4 gnd
port 514 nsew
rlabel metal2 s 20976 11850 20976 11850 4 gnd
port 514 nsew
rlabel metal2 s 20976 11613 20976 11613 4 gnd
port 514 nsew
rlabel metal2 s 21456 10823 21456 10823 4 gnd
port 514 nsew
rlabel metal2 s 21456 10270 21456 10270 4 gnd
port 514 nsew
rlabel metal2 s 20976 11060 20976 11060 4 gnd
port 514 nsew
rlabel metal2 s 20208 11613 20208 11613 4 gnd
port 514 nsew
rlabel metal2 s 20208 11060 20208 11060 4 gnd
port 514 nsew
rlabel metal2 s 20208 12403 20208 12403 4 gnd
port 514 nsew
rlabel metal2 s 21456 10033 21456 10033 4 gnd
port 514 nsew
rlabel metal2 s 20976 12640 20976 12640 4 gnd
port 514 nsew
rlabel metal2 s 22224 10507 22224 10507 4 gnd
port 514 nsew
rlabel metal2 s 22224 8690 22224 8690 4 gnd
port 514 nsew
rlabel metal2 s 20976 9480 20976 9480 4 gnd
port 514 nsew
rlabel metal2 s 21456 6557 21456 6557 4 gnd
port 514 nsew
rlabel metal2 s 20208 8927 20208 8927 4 gnd
port 514 nsew
rlabel metal2 s 22224 7110 22224 7110 4 gnd
port 514 nsew
rlabel metal2 s 21456 9480 21456 9480 4 gnd
port 514 nsew
rlabel metal2 s 22224 8137 22224 8137 4 gnd
port 514 nsew
rlabel metal2 s 20208 7900 20208 7900 4 gnd
port 514 nsew
rlabel metal2 s 20208 7663 20208 7663 4 gnd
port 514 nsew
rlabel metal2 s 20976 8453 20976 8453 4 gnd
port 514 nsew
rlabel metal2 s 21456 7900 21456 7900 4 gnd
port 514 nsew
rlabel metal2 s 21456 9243 21456 9243 4 gnd
port 514 nsew
rlabel metal2 s 20976 7900 20976 7900 4 gnd
port 514 nsew
rlabel metal2 s 21456 6873 21456 6873 4 gnd
port 514 nsew
rlabel metal2 s 21456 8137 21456 8137 4 gnd
port 514 nsew
rlabel metal2 s 22224 7663 22224 7663 4 gnd
port 514 nsew
rlabel metal2 s 21456 8690 21456 8690 4 gnd
port 514 nsew
rlabel metal2 s 20208 8137 20208 8137 4 gnd
port 514 nsew
rlabel metal2 s 22224 7900 22224 7900 4 gnd
port 514 nsew
rlabel metal2 s 20976 7110 20976 7110 4 gnd
port 514 nsew
rlabel metal2 s 20208 9243 20208 9243 4 gnd
port 514 nsew
rlabel metal2 s 20208 6873 20208 6873 4 gnd
port 514 nsew
rlabel metal2 s 20976 8927 20976 8927 4 gnd
port 514 nsew
rlabel metal2 s 22224 9480 22224 9480 4 gnd
port 514 nsew
rlabel metal2 s 22224 8453 22224 8453 4 gnd
port 514 nsew
rlabel metal2 s 21456 8927 21456 8927 4 gnd
port 514 nsew
rlabel metal2 s 22224 6557 22224 6557 4 gnd
port 514 nsew
rlabel metal2 s 22224 9243 22224 9243 4 gnd
port 514 nsew
rlabel metal2 s 20208 7347 20208 7347 4 gnd
port 514 nsew
rlabel metal2 s 20208 9480 20208 9480 4 gnd
port 514 nsew
rlabel metal2 s 20208 8453 20208 8453 4 gnd
port 514 nsew
rlabel metal2 s 20976 6557 20976 6557 4 gnd
port 514 nsew
rlabel metal2 s 21456 7663 21456 7663 4 gnd
port 514 nsew
rlabel metal2 s 22224 6873 22224 6873 4 gnd
port 514 nsew
rlabel metal2 s 21456 7347 21456 7347 4 gnd
port 514 nsew
rlabel metal2 s 21456 8453 21456 8453 4 gnd
port 514 nsew
rlabel metal2 s 22224 7347 22224 7347 4 gnd
port 514 nsew
rlabel metal2 s 21456 7110 21456 7110 4 gnd
port 514 nsew
rlabel metal2 s 20976 8137 20976 8137 4 gnd
port 514 nsew
rlabel metal2 s 20976 7663 20976 7663 4 gnd
port 514 nsew
rlabel metal2 s 20976 7347 20976 7347 4 gnd
port 514 nsew
rlabel metal2 s 20208 7110 20208 7110 4 gnd
port 514 nsew
rlabel metal2 s 22224 8927 22224 8927 4 gnd
port 514 nsew
rlabel metal2 s 20208 8690 20208 8690 4 gnd
port 514 nsew
rlabel metal2 s 20976 8690 20976 8690 4 gnd
port 514 nsew
rlabel metal2 s 20976 9243 20976 9243 4 gnd
port 514 nsew
rlabel metal2 s 20976 6873 20976 6873 4 gnd
port 514 nsew
rlabel metal2 s 20208 6557 20208 6557 4 gnd
port 514 nsew
rlabel metal2 s 24720 8690 24720 8690 4 gnd
port 514 nsew
rlabel metal2 s 22704 8690 22704 8690 4 gnd
port 514 nsew
rlabel metal2 s 23472 8690 23472 8690 4 gnd
port 514 nsew
rlabel metal2 s 23952 7110 23952 7110 4 gnd
port 514 nsew
rlabel metal2 s 22704 7663 22704 7663 4 gnd
port 514 nsew
rlabel metal2 s 23472 7900 23472 7900 4 gnd
port 514 nsew
rlabel metal2 s 23472 8453 23472 8453 4 gnd
port 514 nsew
rlabel metal2 s 24720 7900 24720 7900 4 gnd
port 514 nsew
rlabel metal2 s 22704 9243 22704 9243 4 gnd
port 514 nsew
rlabel metal2 s 24720 8453 24720 8453 4 gnd
port 514 nsew
rlabel metal2 s 24720 6557 24720 6557 4 gnd
port 514 nsew
rlabel metal2 s 23472 6557 23472 6557 4 gnd
port 514 nsew
rlabel metal2 s 22704 7110 22704 7110 4 gnd
port 514 nsew
rlabel metal2 s 23952 7663 23952 7663 4 gnd
port 514 nsew
rlabel metal2 s 23472 9243 23472 9243 4 gnd
port 514 nsew
rlabel metal2 s 23952 8137 23952 8137 4 gnd
port 514 nsew
rlabel metal2 s 23472 6873 23472 6873 4 gnd
port 514 nsew
rlabel metal2 s 24720 6873 24720 6873 4 gnd
port 514 nsew
rlabel metal2 s 22704 8453 22704 8453 4 gnd
port 514 nsew
rlabel metal2 s 22704 8927 22704 8927 4 gnd
port 514 nsew
rlabel metal2 s 23472 7110 23472 7110 4 gnd
port 514 nsew
rlabel metal2 s 24720 7663 24720 7663 4 gnd
port 514 nsew
rlabel metal2 s 23472 7347 23472 7347 4 gnd
port 514 nsew
rlabel metal2 s 23472 9480 23472 9480 4 gnd
port 514 nsew
rlabel metal2 s 22704 6557 22704 6557 4 gnd
port 514 nsew
rlabel metal2 s 22704 6873 22704 6873 4 gnd
port 514 nsew
rlabel metal2 s 22704 7900 22704 7900 4 gnd
port 514 nsew
rlabel metal2 s 23952 8453 23952 8453 4 gnd
port 514 nsew
rlabel metal2 s 22704 8137 22704 8137 4 gnd
port 514 nsew
rlabel metal2 s 24720 9243 24720 9243 4 gnd
port 514 nsew
rlabel metal2 s 22704 7347 22704 7347 4 gnd
port 514 nsew
rlabel metal2 s 23952 6873 23952 6873 4 gnd
port 514 nsew
rlabel metal2 s 24720 8137 24720 8137 4 gnd
port 514 nsew
rlabel metal2 s 23952 7900 23952 7900 4 gnd
port 514 nsew
rlabel metal2 s 23952 8927 23952 8927 4 gnd
port 514 nsew
rlabel metal2 s 23952 6557 23952 6557 4 gnd
port 514 nsew
rlabel metal2 s 23952 9243 23952 9243 4 gnd
port 514 nsew
rlabel metal2 s 23472 7663 23472 7663 4 gnd
port 514 nsew
rlabel metal2 s 23952 8690 23952 8690 4 gnd
port 514 nsew
rlabel metal2 s 24720 7347 24720 7347 4 gnd
port 514 nsew
rlabel metal2 s 24720 8927 24720 8927 4 gnd
port 514 nsew
rlabel metal2 s 23952 7347 23952 7347 4 gnd
port 514 nsew
rlabel metal2 s 22704 9480 22704 9480 4 gnd
port 514 nsew
rlabel metal2 s 24720 9480 24720 9480 4 gnd
port 514 nsew
rlabel metal2 s 23472 8927 23472 8927 4 gnd
port 514 nsew
rlabel metal2 s 23952 9480 23952 9480 4 gnd
port 514 nsew
rlabel metal2 s 24720 7110 24720 7110 4 gnd
port 514 nsew
rlabel metal2 s 23472 8137 23472 8137 4 gnd
port 514 nsew
rlabel metal2 s 23472 4503 23472 4503 4 gnd
port 514 nsew
rlabel metal2 s 23472 4187 23472 4187 4 gnd
port 514 nsew
rlabel metal2 s 23952 6320 23952 6320 4 gnd
port 514 nsew
rlabel metal2 s 24720 4187 24720 4187 4 gnd
port 514 nsew
rlabel metal2 s 22704 4740 22704 4740 4 gnd
port 514 nsew
rlabel metal2 s 24720 3950 24720 3950 4 gnd
port 514 nsew
rlabel metal2 s 23472 5767 23472 5767 4 gnd
port 514 nsew
rlabel metal2 s 24720 4977 24720 4977 4 gnd
port 514 nsew
rlabel metal2 s 23952 3397 23952 3397 4 gnd
port 514 nsew
rlabel metal2 s 23952 5767 23952 5767 4 gnd
port 514 nsew
rlabel metal2 s 22704 4977 22704 4977 4 gnd
port 514 nsew
rlabel metal2 s 24720 4740 24720 4740 4 gnd
port 514 nsew
rlabel metal2 s 23952 4977 23952 4977 4 gnd
port 514 nsew
rlabel metal2 s 24720 3397 24720 3397 4 gnd
port 514 nsew
rlabel metal2 s 22704 5530 22704 5530 4 gnd
port 514 nsew
rlabel metal2 s 23472 6083 23472 6083 4 gnd
port 514 nsew
rlabel metal2 s 22704 5293 22704 5293 4 gnd
port 514 nsew
rlabel metal2 s 23952 6083 23952 6083 4 gnd
port 514 nsew
rlabel metal2 s 23472 3950 23472 3950 4 gnd
port 514 nsew
rlabel metal2 s 23472 5530 23472 5530 4 gnd
port 514 nsew
rlabel metal2 s 22704 3397 22704 3397 4 gnd
port 514 nsew
rlabel metal2 s 22704 3950 22704 3950 4 gnd
port 514 nsew
rlabel metal2 s 23952 5530 23952 5530 4 gnd
port 514 nsew
rlabel metal2 s 22704 6083 22704 6083 4 gnd
port 514 nsew
rlabel metal2 s 24720 6083 24720 6083 4 gnd
port 514 nsew
rlabel metal2 s 23472 6320 23472 6320 4 gnd
port 514 nsew
rlabel metal2 s 23952 3950 23952 3950 4 gnd
port 514 nsew
rlabel metal2 s 23952 4503 23952 4503 4 gnd
port 514 nsew
rlabel metal2 s 23952 4740 23952 4740 4 gnd
port 514 nsew
rlabel metal2 s 23472 5293 23472 5293 4 gnd
port 514 nsew
rlabel metal2 s 24720 4503 24720 4503 4 gnd
port 514 nsew
rlabel metal2 s 22704 3713 22704 3713 4 gnd
port 514 nsew
rlabel metal2 s 24720 6320 24720 6320 4 gnd
port 514 nsew
rlabel metal2 s 23472 3397 23472 3397 4 gnd
port 514 nsew
rlabel metal2 s 22704 5767 22704 5767 4 gnd
port 514 nsew
rlabel metal2 s 24720 5767 24720 5767 4 gnd
port 514 nsew
rlabel metal2 s 22704 4503 22704 4503 4 gnd
port 514 nsew
rlabel metal2 s 23472 4977 23472 4977 4 gnd
port 514 nsew
rlabel metal2 s 24720 5293 24720 5293 4 gnd
port 514 nsew
rlabel metal2 s 22704 6320 22704 6320 4 gnd
port 514 nsew
rlabel metal2 s 22704 4187 22704 4187 4 gnd
port 514 nsew
rlabel metal2 s 23952 4187 23952 4187 4 gnd
port 514 nsew
rlabel metal2 s 23952 3713 23952 3713 4 gnd
port 514 nsew
rlabel metal2 s 23472 4740 23472 4740 4 gnd
port 514 nsew
rlabel metal2 s 23952 5293 23952 5293 4 gnd
port 514 nsew
rlabel metal2 s 24720 5530 24720 5530 4 gnd
port 514 nsew
rlabel metal2 s 23472 3713 23472 3713 4 gnd
port 514 nsew
rlabel metal2 s 24720 3713 24720 3713 4 gnd
port 514 nsew
rlabel metal2 s 21456 3397 21456 3397 4 gnd
port 514 nsew
rlabel metal2 s 20976 3950 20976 3950 4 gnd
port 514 nsew
rlabel metal2 s 20208 4187 20208 4187 4 gnd
port 514 nsew
rlabel metal2 s 22224 4977 22224 4977 4 gnd
port 514 nsew
rlabel metal2 s 22224 6320 22224 6320 4 gnd
port 514 nsew
rlabel metal2 s 21456 6083 21456 6083 4 gnd
port 514 nsew
rlabel metal2 s 20208 3397 20208 3397 4 gnd
port 514 nsew
rlabel metal2 s 22224 3397 22224 3397 4 gnd
port 514 nsew
rlabel metal2 s 21456 4503 21456 4503 4 gnd
port 514 nsew
rlabel metal2 s 20208 4740 20208 4740 4 gnd
port 514 nsew
rlabel metal2 s 22224 4503 22224 4503 4 gnd
port 514 nsew
rlabel metal2 s 20976 3397 20976 3397 4 gnd
port 514 nsew
rlabel metal2 s 22224 4187 22224 4187 4 gnd
port 514 nsew
rlabel metal2 s 21456 3713 21456 3713 4 gnd
port 514 nsew
rlabel metal2 s 20976 6320 20976 6320 4 gnd
port 514 nsew
rlabel metal2 s 21456 6320 21456 6320 4 gnd
port 514 nsew
rlabel metal2 s 20976 5530 20976 5530 4 gnd
port 514 nsew
rlabel metal2 s 20208 5767 20208 5767 4 gnd
port 514 nsew
rlabel metal2 s 22224 5293 22224 5293 4 gnd
port 514 nsew
rlabel metal2 s 20976 3713 20976 3713 4 gnd
port 514 nsew
rlabel metal2 s 20208 6320 20208 6320 4 gnd
port 514 nsew
rlabel metal2 s 20208 3950 20208 3950 4 gnd
port 514 nsew
rlabel metal2 s 20208 5530 20208 5530 4 gnd
port 514 nsew
rlabel metal2 s 20976 4187 20976 4187 4 gnd
port 514 nsew
rlabel metal2 s 20976 4977 20976 4977 4 gnd
port 514 nsew
rlabel metal2 s 20976 4503 20976 4503 4 gnd
port 514 nsew
rlabel metal2 s 20976 5767 20976 5767 4 gnd
port 514 nsew
rlabel metal2 s 21456 5293 21456 5293 4 gnd
port 514 nsew
rlabel metal2 s 21456 4977 21456 4977 4 gnd
port 514 nsew
rlabel metal2 s 21456 5767 21456 5767 4 gnd
port 514 nsew
rlabel metal2 s 22224 4740 22224 4740 4 gnd
port 514 nsew
rlabel metal2 s 22224 5530 22224 5530 4 gnd
port 514 nsew
rlabel metal2 s 20208 4977 20208 4977 4 gnd
port 514 nsew
rlabel metal2 s 21456 4740 21456 4740 4 gnd
port 514 nsew
rlabel metal2 s 20208 6083 20208 6083 4 gnd
port 514 nsew
rlabel metal2 s 20976 4740 20976 4740 4 gnd
port 514 nsew
rlabel metal2 s 22224 3713 22224 3713 4 gnd
port 514 nsew
rlabel metal2 s 22224 6083 22224 6083 4 gnd
port 514 nsew
rlabel metal2 s 20208 4503 20208 4503 4 gnd
port 514 nsew
rlabel metal2 s 20976 5293 20976 5293 4 gnd
port 514 nsew
rlabel metal2 s 20976 6083 20976 6083 4 gnd
port 514 nsew
rlabel metal2 s 21456 4187 21456 4187 4 gnd
port 514 nsew
rlabel metal2 s 21456 5530 21456 5530 4 gnd
port 514 nsew
rlabel metal2 s 22224 5767 22224 5767 4 gnd
port 514 nsew
rlabel metal2 s 20208 5293 20208 5293 4 gnd
port 514 nsew
rlabel metal2 s 22224 3950 22224 3950 4 gnd
port 514 nsew
rlabel metal2 s 21456 3950 21456 3950 4 gnd
port 514 nsew
rlabel metal2 s 20208 3713 20208 3713 4 gnd
port 514 nsew
rlabel metal2 s 20976 553 20976 553 4 gnd
port 514 nsew
rlabel metal2 s 22224 237 22224 237 4 gnd
port 514 nsew
rlabel metal2 s 20208 553 20208 553 4 gnd
port 514 nsew
rlabel metal2 s 21456 1580 21456 1580 4 gnd
port 514 nsew
rlabel metal2 s 20208 1580 20208 1580 4 gnd
port 514 nsew
rlabel metal2 s 22224 2923 22224 2923 4 gnd
port 514 nsew
rlabel metal2 s 20208 2923 20208 2923 4 gnd
port 514 nsew
rlabel metal2 s 20976 0 20976 0 4 gnd
port 514 nsew
rlabel metal2 s 20976 2607 20976 2607 4 gnd
port 514 nsew
rlabel metal2 s 20208 790 20208 790 4 gnd
port 514 nsew
rlabel metal2 s 22224 1580 22224 1580 4 gnd
port 514 nsew
rlabel metal2 s 20208 2370 20208 2370 4 gnd
port 514 nsew
rlabel metal2 s 21456 1343 21456 1343 4 gnd
port 514 nsew
rlabel metal2 s 21456 2607 21456 2607 4 gnd
port 514 nsew
rlabel metal2 s 22224 2370 22224 2370 4 gnd
port 514 nsew
rlabel metal2 s 21456 0 21456 0 4 gnd
port 514 nsew
rlabel metal2 s 20208 2607 20208 2607 4 gnd
port 514 nsew
rlabel metal2 s 21456 553 21456 553 4 gnd
port 514 nsew
rlabel metal2 s 20976 2133 20976 2133 4 gnd
port 514 nsew
rlabel metal2 s 22224 1027 22224 1027 4 gnd
port 514 nsew
rlabel metal2 s 22224 0 22224 0 4 gnd
port 514 nsew
rlabel metal2 s 20208 237 20208 237 4 gnd
port 514 nsew
rlabel metal2 s 22224 2607 22224 2607 4 gnd
port 514 nsew
rlabel metal2 s 21456 790 21456 790 4 gnd
port 514 nsew
rlabel metal2 s 20208 2133 20208 2133 4 gnd
port 514 nsew
rlabel metal2 s 21456 237 21456 237 4 gnd
port 514 nsew
rlabel metal2 s 20976 1027 20976 1027 4 gnd
port 514 nsew
rlabel metal2 s 20208 1343 20208 1343 4 gnd
port 514 nsew
rlabel metal2 s 21456 1817 21456 1817 4 gnd
port 514 nsew
rlabel metal2 s 21456 2370 21456 2370 4 gnd
port 514 nsew
rlabel metal2 s 20208 3160 20208 3160 4 gnd
port 514 nsew
rlabel metal2 s 22224 3160 22224 3160 4 gnd
port 514 nsew
rlabel metal2 s 20208 1027 20208 1027 4 gnd
port 514 nsew
rlabel metal2 s 20208 1817 20208 1817 4 gnd
port 514 nsew
rlabel metal2 s 20976 1817 20976 1817 4 gnd
port 514 nsew
rlabel metal2 s 22224 1343 22224 1343 4 gnd
port 514 nsew
rlabel metal2 s 22224 553 22224 553 4 gnd
port 514 nsew
rlabel metal2 s 20976 790 20976 790 4 gnd
port 514 nsew
rlabel metal2 s 20976 1343 20976 1343 4 gnd
port 514 nsew
rlabel metal2 s 21456 2923 21456 2923 4 gnd
port 514 nsew
rlabel metal2 s 20976 1580 20976 1580 4 gnd
port 514 nsew
rlabel metal2 s 21456 1027 21456 1027 4 gnd
port 514 nsew
rlabel metal2 s 20976 2923 20976 2923 4 gnd
port 514 nsew
rlabel metal2 s 22224 1817 22224 1817 4 gnd
port 514 nsew
rlabel metal2 s 22224 790 22224 790 4 gnd
port 514 nsew
rlabel metal2 s 20976 3160 20976 3160 4 gnd
port 514 nsew
rlabel metal2 s 22224 2133 22224 2133 4 gnd
port 514 nsew
rlabel metal2 s 21456 2133 21456 2133 4 gnd
port 514 nsew
rlabel metal2 s 20976 2370 20976 2370 4 gnd
port 514 nsew
rlabel metal2 s 20208 0 20208 0 4 gnd
port 514 nsew
rlabel metal2 s 21456 3160 21456 3160 4 gnd
port 514 nsew
rlabel metal2 s 20976 237 20976 237 4 gnd
port 514 nsew
rlabel metal2 s 24720 1580 24720 1580 4 gnd
port 514 nsew
rlabel metal2 s 23952 1027 23952 1027 4 gnd
port 514 nsew
rlabel metal2 s 23952 237 23952 237 4 gnd
port 514 nsew
rlabel metal2 s 24720 3160 24720 3160 4 gnd
port 514 nsew
rlabel metal2 s 24720 237 24720 237 4 gnd
port 514 nsew
rlabel metal2 s 23952 790 23952 790 4 gnd
port 514 nsew
rlabel metal2 s 23472 3160 23472 3160 4 gnd
port 514 nsew
rlabel metal2 s 22704 237 22704 237 4 gnd
port 514 nsew
rlabel metal2 s 23472 1580 23472 1580 4 gnd
port 514 nsew
rlabel metal2 s 23952 0 23952 0 4 gnd
port 514 nsew
rlabel metal2 s 23952 1580 23952 1580 4 gnd
port 514 nsew
rlabel metal2 s 23472 237 23472 237 4 gnd
port 514 nsew
rlabel metal2 s 22704 1580 22704 1580 4 gnd
port 514 nsew
rlabel metal2 s 22704 2607 22704 2607 4 gnd
port 514 nsew
rlabel metal2 s 22704 790 22704 790 4 gnd
port 514 nsew
rlabel metal2 s 22704 2133 22704 2133 4 gnd
port 514 nsew
rlabel metal2 s 24720 1817 24720 1817 4 gnd
port 514 nsew
rlabel metal2 s 23952 3160 23952 3160 4 gnd
port 514 nsew
rlabel metal2 s 23952 1817 23952 1817 4 gnd
port 514 nsew
rlabel metal2 s 23472 1027 23472 1027 4 gnd
port 514 nsew
rlabel metal2 s 23472 1817 23472 1817 4 gnd
port 514 nsew
rlabel metal2 s 23952 1343 23952 1343 4 gnd
port 514 nsew
rlabel metal2 s 24720 0 24720 0 4 gnd
port 514 nsew
rlabel metal2 s 23952 2370 23952 2370 4 gnd
port 514 nsew
rlabel metal2 s 22704 3160 22704 3160 4 gnd
port 514 nsew
rlabel metal2 s 23472 1343 23472 1343 4 gnd
port 514 nsew
rlabel metal2 s 23472 2133 23472 2133 4 gnd
port 514 nsew
rlabel metal2 s 23472 2370 23472 2370 4 gnd
port 514 nsew
rlabel metal2 s 24720 790 24720 790 4 gnd
port 514 nsew
rlabel metal2 s 22704 1027 22704 1027 4 gnd
port 514 nsew
rlabel metal2 s 22704 1343 22704 1343 4 gnd
port 514 nsew
rlabel metal2 s 23952 2133 23952 2133 4 gnd
port 514 nsew
rlabel metal2 s 24720 553 24720 553 4 gnd
port 514 nsew
rlabel metal2 s 24720 2133 24720 2133 4 gnd
port 514 nsew
rlabel metal2 s 24720 2923 24720 2923 4 gnd
port 514 nsew
rlabel metal2 s 22704 2370 22704 2370 4 gnd
port 514 nsew
rlabel metal2 s 24720 1027 24720 1027 4 gnd
port 514 nsew
rlabel metal2 s 24720 1343 24720 1343 4 gnd
port 514 nsew
rlabel metal2 s 23472 0 23472 0 4 gnd
port 514 nsew
rlabel metal2 s 23952 2923 23952 2923 4 gnd
port 514 nsew
rlabel metal2 s 23472 2923 23472 2923 4 gnd
port 514 nsew
rlabel metal2 s 22704 2923 22704 2923 4 gnd
port 514 nsew
rlabel metal2 s 24720 2370 24720 2370 4 gnd
port 514 nsew
rlabel metal2 s 24720 2607 24720 2607 4 gnd
port 514 nsew
rlabel metal2 s 22704 0 22704 0 4 gnd
port 514 nsew
rlabel metal2 s 22704 553 22704 553 4 gnd
port 514 nsew
rlabel metal2 s 23952 553 23952 553 4 gnd
port 514 nsew
rlabel metal2 s 23472 2607 23472 2607 4 gnd
port 514 nsew
rlabel metal2 s 22704 1817 22704 1817 4 gnd
port 514 nsew
rlabel metal2 s 23472 553 23472 553 4 gnd
port 514 nsew
rlabel metal2 s 23952 2607 23952 2607 4 gnd
port 514 nsew
rlabel metal2 s 23472 790 23472 790 4 gnd
port 514 nsew
rlabel metal2 s 27696 4977 27696 4977 4 gnd
port 514 nsew
rlabel metal2 s 28944 3950 28944 3950 4 gnd
port 514 nsew
rlabel metal2 s 28944 6320 28944 6320 4 gnd
port 514 nsew
rlabel metal2 s 29712 3950 29712 3950 4 gnd
port 514 nsew
rlabel metal2 s 29712 3713 29712 3713 4 gnd
port 514 nsew
rlabel metal2 s 28464 4740 28464 4740 4 gnd
port 514 nsew
rlabel metal2 s 28464 6083 28464 6083 4 gnd
port 514 nsew
rlabel metal2 s 28944 4503 28944 4503 4 gnd
port 514 nsew
rlabel metal2 s 28944 4740 28944 4740 4 gnd
port 514 nsew
rlabel metal2 s 27696 4503 27696 4503 4 gnd
port 514 nsew
rlabel metal2 s 27696 3397 27696 3397 4 gnd
port 514 nsew
rlabel metal2 s 27696 5530 27696 5530 4 gnd
port 514 nsew
rlabel metal2 s 27696 4740 27696 4740 4 gnd
port 514 nsew
rlabel metal2 s 27696 3950 27696 3950 4 gnd
port 514 nsew
rlabel metal2 s 29712 4187 29712 4187 4 gnd
port 514 nsew
rlabel metal2 s 28464 3950 28464 3950 4 gnd
port 514 nsew
rlabel metal2 s 29712 3397 29712 3397 4 gnd
port 514 nsew
rlabel metal2 s 27696 5293 27696 5293 4 gnd
port 514 nsew
rlabel metal2 s 29712 6083 29712 6083 4 gnd
port 514 nsew
rlabel metal2 s 29712 5767 29712 5767 4 gnd
port 514 nsew
rlabel metal2 s 27696 3713 27696 3713 4 gnd
port 514 nsew
rlabel metal2 s 27696 5767 27696 5767 4 gnd
port 514 nsew
rlabel metal2 s 28464 4187 28464 4187 4 gnd
port 514 nsew
rlabel metal2 s 28944 4977 28944 4977 4 gnd
port 514 nsew
rlabel metal2 s 28944 5767 28944 5767 4 gnd
port 514 nsew
rlabel metal2 s 28464 3397 28464 3397 4 gnd
port 514 nsew
rlabel metal2 s 28944 3713 28944 3713 4 gnd
port 514 nsew
rlabel metal2 s 29712 5530 29712 5530 4 gnd
port 514 nsew
rlabel metal2 s 28464 3713 28464 3713 4 gnd
port 514 nsew
rlabel metal2 s 28464 5530 28464 5530 4 gnd
port 514 nsew
rlabel metal2 s 29712 4977 29712 4977 4 gnd
port 514 nsew
rlabel metal2 s 27696 6320 27696 6320 4 gnd
port 514 nsew
rlabel metal2 s 28464 6320 28464 6320 4 gnd
port 514 nsew
rlabel metal2 s 27696 6083 27696 6083 4 gnd
port 514 nsew
rlabel metal2 s 29712 4740 29712 4740 4 gnd
port 514 nsew
rlabel metal2 s 28944 4187 28944 4187 4 gnd
port 514 nsew
rlabel metal2 s 28464 4503 28464 4503 4 gnd
port 514 nsew
rlabel metal2 s 28944 3397 28944 3397 4 gnd
port 514 nsew
rlabel metal2 s 27696 4187 27696 4187 4 gnd
port 514 nsew
rlabel metal2 s 28464 5767 28464 5767 4 gnd
port 514 nsew
rlabel metal2 s 28944 5530 28944 5530 4 gnd
port 514 nsew
rlabel metal2 s 29712 6320 29712 6320 4 gnd
port 514 nsew
rlabel metal2 s 28464 4977 28464 4977 4 gnd
port 514 nsew
rlabel metal2 s 28464 5293 28464 5293 4 gnd
port 514 nsew
rlabel metal2 s 29712 4503 29712 4503 4 gnd
port 514 nsew
rlabel metal2 s 28944 5293 28944 5293 4 gnd
port 514 nsew
rlabel metal2 s 28944 6083 28944 6083 4 gnd
port 514 nsew
rlabel metal2 s 29712 5293 29712 5293 4 gnd
port 514 nsew
rlabel metal2 s 26448 4503 26448 4503 4 gnd
port 514 nsew
rlabel metal2 s 25200 3950 25200 3950 4 gnd
port 514 nsew
rlabel metal2 s 25968 3713 25968 3713 4 gnd
port 514 nsew
rlabel metal2 s 25200 3397 25200 3397 4 gnd
port 514 nsew
rlabel metal2 s 27216 3950 27216 3950 4 gnd
port 514 nsew
rlabel metal2 s 26448 5293 26448 5293 4 gnd
port 514 nsew
rlabel metal2 s 25968 4187 25968 4187 4 gnd
port 514 nsew
rlabel metal2 s 25968 5767 25968 5767 4 gnd
port 514 nsew
rlabel metal2 s 26448 4740 26448 4740 4 gnd
port 514 nsew
rlabel metal2 s 25968 6083 25968 6083 4 gnd
port 514 nsew
rlabel metal2 s 27216 4187 27216 4187 4 gnd
port 514 nsew
rlabel metal2 s 26448 6320 26448 6320 4 gnd
port 514 nsew
rlabel metal2 s 25968 6320 25968 6320 4 gnd
port 514 nsew
rlabel metal2 s 27216 3713 27216 3713 4 gnd
port 514 nsew
rlabel metal2 s 27216 4977 27216 4977 4 gnd
port 514 nsew
rlabel metal2 s 26448 3950 26448 3950 4 gnd
port 514 nsew
rlabel metal2 s 25200 4187 25200 4187 4 gnd
port 514 nsew
rlabel metal2 s 25200 4503 25200 4503 4 gnd
port 514 nsew
rlabel metal2 s 26448 4187 26448 4187 4 gnd
port 514 nsew
rlabel metal2 s 26448 4977 26448 4977 4 gnd
port 514 nsew
rlabel metal2 s 25200 4740 25200 4740 4 gnd
port 514 nsew
rlabel metal2 s 25968 5530 25968 5530 4 gnd
port 514 nsew
rlabel metal2 s 25200 5293 25200 5293 4 gnd
port 514 nsew
rlabel metal2 s 25200 3713 25200 3713 4 gnd
port 514 nsew
rlabel metal2 s 25200 6320 25200 6320 4 gnd
port 514 nsew
rlabel metal2 s 25968 5293 25968 5293 4 gnd
port 514 nsew
rlabel metal2 s 25200 5767 25200 5767 4 gnd
port 514 nsew
rlabel metal2 s 25968 3397 25968 3397 4 gnd
port 514 nsew
rlabel metal2 s 27216 3397 27216 3397 4 gnd
port 514 nsew
rlabel metal2 s 27216 5767 27216 5767 4 gnd
port 514 nsew
rlabel metal2 s 26448 5530 26448 5530 4 gnd
port 514 nsew
rlabel metal2 s 27216 6083 27216 6083 4 gnd
port 514 nsew
rlabel metal2 s 27216 5530 27216 5530 4 gnd
port 514 nsew
rlabel metal2 s 25968 4503 25968 4503 4 gnd
port 514 nsew
rlabel metal2 s 25968 4977 25968 4977 4 gnd
port 514 nsew
rlabel metal2 s 25200 6083 25200 6083 4 gnd
port 514 nsew
rlabel metal2 s 27216 6320 27216 6320 4 gnd
port 514 nsew
rlabel metal2 s 25968 4740 25968 4740 4 gnd
port 514 nsew
rlabel metal2 s 25200 5530 25200 5530 4 gnd
port 514 nsew
rlabel metal2 s 26448 5767 26448 5767 4 gnd
port 514 nsew
rlabel metal2 s 26448 3713 26448 3713 4 gnd
port 514 nsew
rlabel metal2 s 27216 4503 27216 4503 4 gnd
port 514 nsew
rlabel metal2 s 26448 6083 26448 6083 4 gnd
port 514 nsew
rlabel metal2 s 25968 3950 25968 3950 4 gnd
port 514 nsew
rlabel metal2 s 25200 4977 25200 4977 4 gnd
port 514 nsew
rlabel metal2 s 27216 5293 27216 5293 4 gnd
port 514 nsew
rlabel metal2 s 27216 4740 27216 4740 4 gnd
port 514 nsew
rlabel metal2 s 26448 3397 26448 3397 4 gnd
port 514 nsew
rlabel metal2 s 26448 1027 26448 1027 4 gnd
port 514 nsew
rlabel metal2 s 27216 1343 27216 1343 4 gnd
port 514 nsew
rlabel metal2 s 26448 1580 26448 1580 4 gnd
port 514 nsew
rlabel metal2 s 27216 2370 27216 2370 4 gnd
port 514 nsew
rlabel metal2 s 27216 1027 27216 1027 4 gnd
port 514 nsew
rlabel metal2 s 27216 237 27216 237 4 gnd
port 514 nsew
rlabel metal2 s 25968 0 25968 0 4 gnd
port 514 nsew
rlabel metal2 s 25968 1817 25968 1817 4 gnd
port 514 nsew
rlabel metal2 s 27216 790 27216 790 4 gnd
port 514 nsew
rlabel metal2 s 25200 1027 25200 1027 4 gnd
port 514 nsew
rlabel metal2 s 25968 2370 25968 2370 4 gnd
port 514 nsew
rlabel metal2 s 25968 1027 25968 1027 4 gnd
port 514 nsew
rlabel metal2 s 25968 237 25968 237 4 gnd
port 514 nsew
rlabel metal2 s 26448 553 26448 553 4 gnd
port 514 nsew
rlabel metal2 s 25968 1343 25968 1343 4 gnd
port 514 nsew
rlabel metal2 s 27216 1817 27216 1817 4 gnd
port 514 nsew
rlabel metal2 s 27216 2133 27216 2133 4 gnd
port 514 nsew
rlabel metal2 s 25968 2607 25968 2607 4 gnd
port 514 nsew
rlabel metal2 s 25968 790 25968 790 4 gnd
port 514 nsew
rlabel metal2 s 25200 2370 25200 2370 4 gnd
port 514 nsew
rlabel metal2 s 25200 3160 25200 3160 4 gnd
port 514 nsew
rlabel metal2 s 25968 1580 25968 1580 4 gnd
port 514 nsew
rlabel metal2 s 25968 2923 25968 2923 4 gnd
port 514 nsew
rlabel metal2 s 25200 237 25200 237 4 gnd
port 514 nsew
rlabel metal2 s 25200 1817 25200 1817 4 gnd
port 514 nsew
rlabel metal2 s 25200 2133 25200 2133 4 gnd
port 514 nsew
rlabel metal2 s 26448 3160 26448 3160 4 gnd
port 514 nsew
rlabel metal2 s 27216 2923 27216 2923 4 gnd
port 514 nsew
rlabel metal2 s 25968 3160 25968 3160 4 gnd
port 514 nsew
rlabel metal2 s 26448 2370 26448 2370 4 gnd
port 514 nsew
rlabel metal2 s 25200 2923 25200 2923 4 gnd
port 514 nsew
rlabel metal2 s 26448 2607 26448 2607 4 gnd
port 514 nsew
rlabel metal2 s 26448 1817 26448 1817 4 gnd
port 514 nsew
rlabel metal2 s 25200 1580 25200 1580 4 gnd
port 514 nsew
rlabel metal2 s 27216 1580 27216 1580 4 gnd
port 514 nsew
rlabel metal2 s 25200 1343 25200 1343 4 gnd
port 514 nsew
rlabel metal2 s 25968 553 25968 553 4 gnd
port 514 nsew
rlabel metal2 s 26448 790 26448 790 4 gnd
port 514 nsew
rlabel metal2 s 26448 2923 26448 2923 4 gnd
port 514 nsew
rlabel metal2 s 26448 237 26448 237 4 gnd
port 514 nsew
rlabel metal2 s 25200 2607 25200 2607 4 gnd
port 514 nsew
rlabel metal2 s 27216 2607 27216 2607 4 gnd
port 514 nsew
rlabel metal2 s 25200 553 25200 553 4 gnd
port 514 nsew
rlabel metal2 s 25200 790 25200 790 4 gnd
port 514 nsew
rlabel metal2 s 27216 553 27216 553 4 gnd
port 514 nsew
rlabel metal2 s 26448 1343 26448 1343 4 gnd
port 514 nsew
rlabel metal2 s 26448 2133 26448 2133 4 gnd
port 514 nsew
rlabel metal2 s 27216 0 27216 0 4 gnd
port 514 nsew
rlabel metal2 s 26448 0 26448 0 4 gnd
port 514 nsew
rlabel metal2 s 25968 2133 25968 2133 4 gnd
port 514 nsew
rlabel metal2 s 25200 0 25200 0 4 gnd
port 514 nsew
rlabel metal2 s 27216 3160 27216 3160 4 gnd
port 514 nsew
rlabel metal2 s 28464 0 28464 0 4 gnd
port 514 nsew
rlabel metal2 s 27696 1027 27696 1027 4 gnd
port 514 nsew
rlabel metal2 s 27696 2370 27696 2370 4 gnd
port 514 nsew
rlabel metal2 s 28464 790 28464 790 4 gnd
port 514 nsew
rlabel metal2 s 28464 2370 28464 2370 4 gnd
port 514 nsew
rlabel metal2 s 28944 0 28944 0 4 gnd
port 514 nsew
rlabel metal2 s 28944 790 28944 790 4 gnd
port 514 nsew
rlabel metal2 s 28944 2923 28944 2923 4 gnd
port 514 nsew
rlabel metal2 s 28944 1580 28944 1580 4 gnd
port 514 nsew
rlabel metal2 s 29712 1817 29712 1817 4 gnd
port 514 nsew
rlabel metal2 s 27696 3160 27696 3160 4 gnd
port 514 nsew
rlabel metal2 s 29712 2607 29712 2607 4 gnd
port 514 nsew
rlabel metal2 s 28464 237 28464 237 4 gnd
port 514 nsew
rlabel metal2 s 29712 3160 29712 3160 4 gnd
port 514 nsew
rlabel metal2 s 28944 1343 28944 1343 4 gnd
port 514 nsew
rlabel metal2 s 28464 1817 28464 1817 4 gnd
port 514 nsew
rlabel metal2 s 27696 2607 27696 2607 4 gnd
port 514 nsew
rlabel metal2 s 29712 1027 29712 1027 4 gnd
port 514 nsew
rlabel metal2 s 28944 1027 28944 1027 4 gnd
port 514 nsew
rlabel metal2 s 28944 3160 28944 3160 4 gnd
port 514 nsew
rlabel metal2 s 29712 0 29712 0 4 gnd
port 514 nsew
rlabel metal2 s 28464 553 28464 553 4 gnd
port 514 nsew
rlabel metal2 s 28944 2607 28944 2607 4 gnd
port 514 nsew
rlabel metal2 s 29712 2370 29712 2370 4 gnd
port 514 nsew
rlabel metal2 s 28944 237 28944 237 4 gnd
port 514 nsew
rlabel metal2 s 28464 2133 28464 2133 4 gnd
port 514 nsew
rlabel metal2 s 27696 1580 27696 1580 4 gnd
port 514 nsew
rlabel metal2 s 29712 237 29712 237 4 gnd
port 514 nsew
rlabel metal2 s 28464 2923 28464 2923 4 gnd
port 514 nsew
rlabel metal2 s 29712 1580 29712 1580 4 gnd
port 514 nsew
rlabel metal2 s 28464 1343 28464 1343 4 gnd
port 514 nsew
rlabel metal2 s 28464 3160 28464 3160 4 gnd
port 514 nsew
rlabel metal2 s 28944 2133 28944 2133 4 gnd
port 514 nsew
rlabel metal2 s 29712 2133 29712 2133 4 gnd
port 514 nsew
rlabel metal2 s 27696 237 27696 237 4 gnd
port 514 nsew
rlabel metal2 s 27696 0 27696 0 4 gnd
port 514 nsew
rlabel metal2 s 27696 2133 27696 2133 4 gnd
port 514 nsew
rlabel metal2 s 29712 790 29712 790 4 gnd
port 514 nsew
rlabel metal2 s 27696 553 27696 553 4 gnd
port 514 nsew
rlabel metal2 s 28944 1817 28944 1817 4 gnd
port 514 nsew
rlabel metal2 s 28944 2370 28944 2370 4 gnd
port 514 nsew
rlabel metal2 s 28464 1580 28464 1580 4 gnd
port 514 nsew
rlabel metal2 s 29712 1343 29712 1343 4 gnd
port 514 nsew
rlabel metal2 s 27696 1343 27696 1343 4 gnd
port 514 nsew
rlabel metal2 s 29712 553 29712 553 4 gnd
port 514 nsew
rlabel metal2 s 28464 1027 28464 1027 4 gnd
port 514 nsew
rlabel metal2 s 28464 2607 28464 2607 4 gnd
port 514 nsew
rlabel metal2 s 27696 1817 27696 1817 4 gnd
port 514 nsew
rlabel metal2 s 27696 790 27696 790 4 gnd
port 514 nsew
rlabel metal2 s 28944 553 28944 553 4 gnd
port 514 nsew
rlabel metal2 s 29712 2923 29712 2923 4 gnd
port 514 nsew
rlabel metal2 s 27696 2923 27696 2923 4 gnd
port 514 nsew
rlabel metal2 s 38448 12640 38448 12640 4 gnd
port 514 nsew
rlabel metal2 s 37680 10507 37680 10507 4 gnd
port 514 nsew
rlabel metal2 s 39696 11613 39696 11613 4 gnd
port 514 nsew
rlabel metal2 s 39696 11297 39696 11297 4 gnd
port 514 nsew
rlabel metal2 s 37680 10823 37680 10823 4 gnd
port 514 nsew
rlabel metal2 s 38928 11613 38928 11613 4 gnd
port 514 nsew
rlabel metal2 s 39696 12640 39696 12640 4 gnd
port 514 nsew
rlabel metal2 s 38448 12403 38448 12403 4 gnd
port 514 nsew
rlabel metal2 s 38928 10270 38928 10270 4 gnd
port 514 nsew
rlabel metal2 s 37680 12087 37680 12087 4 gnd
port 514 nsew
rlabel metal2 s 37680 11060 37680 11060 4 gnd
port 514 nsew
rlabel metal2 s 37680 11850 37680 11850 4 gnd
port 514 nsew
rlabel metal2 s 38928 11297 38928 11297 4 gnd
port 514 nsew
rlabel metal2 s 39696 12403 39696 12403 4 gnd
port 514 nsew
rlabel metal2 s 38448 11850 38448 11850 4 gnd
port 514 nsew
rlabel metal2 s 38928 10033 38928 10033 4 gnd
port 514 nsew
rlabel metal2 s 37680 10270 37680 10270 4 gnd
port 514 nsew
rlabel metal2 s 37680 12403 37680 12403 4 gnd
port 514 nsew
rlabel metal2 s 38928 11850 38928 11850 4 gnd
port 514 nsew
rlabel metal2 s 38448 10270 38448 10270 4 gnd
port 514 nsew
rlabel metal2 s 38928 11060 38928 11060 4 gnd
port 514 nsew
rlabel metal2 s 38928 12403 38928 12403 4 gnd
port 514 nsew
rlabel metal2 s 38928 12640 38928 12640 4 gnd
port 514 nsew
rlabel metal2 s 39696 9717 39696 9717 4 gnd
port 514 nsew
rlabel metal2 s 38448 9717 38448 9717 4 gnd
port 514 nsew
rlabel metal2 s 39696 10823 39696 10823 4 gnd
port 514 nsew
rlabel metal2 s 38448 12087 38448 12087 4 gnd
port 514 nsew
rlabel metal2 s 39696 10033 39696 10033 4 gnd
port 514 nsew
rlabel metal2 s 38448 10507 38448 10507 4 gnd
port 514 nsew
rlabel metal2 s 39696 10507 39696 10507 4 gnd
port 514 nsew
rlabel metal2 s 38928 12087 38928 12087 4 gnd
port 514 nsew
rlabel metal2 s 38928 10507 38928 10507 4 gnd
port 514 nsew
rlabel metal2 s 39696 10270 39696 10270 4 gnd
port 514 nsew
rlabel metal2 s 37680 9717 37680 9717 4 gnd
port 514 nsew
rlabel metal2 s 39696 11060 39696 11060 4 gnd
port 514 nsew
rlabel metal2 s 39696 12087 39696 12087 4 gnd
port 514 nsew
rlabel metal2 s 38928 10823 38928 10823 4 gnd
port 514 nsew
rlabel metal2 s 37680 11613 37680 11613 4 gnd
port 514 nsew
rlabel metal2 s 38448 11060 38448 11060 4 gnd
port 514 nsew
rlabel metal2 s 39696 11850 39696 11850 4 gnd
port 514 nsew
rlabel metal2 s 37680 12640 37680 12640 4 gnd
port 514 nsew
rlabel metal2 s 37680 11297 37680 11297 4 gnd
port 514 nsew
rlabel metal2 s 37680 10033 37680 10033 4 gnd
port 514 nsew
rlabel metal2 s 38448 11613 38448 11613 4 gnd
port 514 nsew
rlabel metal2 s 38448 10823 38448 10823 4 gnd
port 514 nsew
rlabel metal2 s 38448 10033 38448 10033 4 gnd
port 514 nsew
rlabel metal2 s 38928 9717 38928 9717 4 gnd
port 514 nsew
rlabel metal2 s 38448 11297 38448 11297 4 gnd
port 514 nsew
rlabel metal2 s 36432 10507 36432 10507 4 gnd
port 514 nsew
rlabel metal2 s 35952 11613 35952 11613 4 gnd
port 514 nsew
rlabel metal2 s 36432 10823 36432 10823 4 gnd
port 514 nsew
rlabel metal2 s 36432 9717 36432 9717 4 gnd
port 514 nsew
rlabel metal2 s 35184 9717 35184 9717 4 gnd
port 514 nsew
rlabel metal2 s 35184 12403 35184 12403 4 gnd
port 514 nsew
rlabel metal2 s 35184 10507 35184 10507 4 gnd
port 514 nsew
rlabel metal2 s 36432 12640 36432 12640 4 gnd
port 514 nsew
rlabel metal2 s 35952 12640 35952 12640 4 gnd
port 514 nsew
rlabel metal2 s 35952 10270 35952 10270 4 gnd
port 514 nsew
rlabel metal2 s 35952 9717 35952 9717 4 gnd
port 514 nsew
rlabel metal2 s 37200 12087 37200 12087 4 gnd
port 514 nsew
rlabel metal2 s 35952 12403 35952 12403 4 gnd
port 514 nsew
rlabel metal2 s 35952 11060 35952 11060 4 gnd
port 514 nsew
rlabel metal2 s 35184 12087 35184 12087 4 gnd
port 514 nsew
rlabel metal2 s 36432 11297 36432 11297 4 gnd
port 514 nsew
rlabel metal2 s 35184 11060 35184 11060 4 gnd
port 514 nsew
rlabel metal2 s 35184 10033 35184 10033 4 gnd
port 514 nsew
rlabel metal2 s 35952 10823 35952 10823 4 gnd
port 514 nsew
rlabel metal2 s 35184 11613 35184 11613 4 gnd
port 514 nsew
rlabel metal2 s 36432 11060 36432 11060 4 gnd
port 514 nsew
rlabel metal2 s 37200 10823 37200 10823 4 gnd
port 514 nsew
rlabel metal2 s 37200 10507 37200 10507 4 gnd
port 514 nsew
rlabel metal2 s 35184 10823 35184 10823 4 gnd
port 514 nsew
rlabel metal2 s 36432 11850 36432 11850 4 gnd
port 514 nsew
rlabel metal2 s 37200 10033 37200 10033 4 gnd
port 514 nsew
rlabel metal2 s 37200 12403 37200 12403 4 gnd
port 514 nsew
rlabel metal2 s 35184 11850 35184 11850 4 gnd
port 514 nsew
rlabel metal2 s 35952 11297 35952 11297 4 gnd
port 514 nsew
rlabel metal2 s 37200 12640 37200 12640 4 gnd
port 514 nsew
rlabel metal2 s 37200 9717 37200 9717 4 gnd
port 514 nsew
rlabel metal2 s 35952 12087 35952 12087 4 gnd
port 514 nsew
rlabel metal2 s 37200 11850 37200 11850 4 gnd
port 514 nsew
rlabel metal2 s 36432 12087 36432 12087 4 gnd
port 514 nsew
rlabel metal2 s 35952 10507 35952 10507 4 gnd
port 514 nsew
rlabel metal2 s 36432 11613 36432 11613 4 gnd
port 514 nsew
rlabel metal2 s 35184 11297 35184 11297 4 gnd
port 514 nsew
rlabel metal2 s 36432 10033 36432 10033 4 gnd
port 514 nsew
rlabel metal2 s 35184 12640 35184 12640 4 gnd
port 514 nsew
rlabel metal2 s 35184 10270 35184 10270 4 gnd
port 514 nsew
rlabel metal2 s 37200 11060 37200 11060 4 gnd
port 514 nsew
rlabel metal2 s 36432 10270 36432 10270 4 gnd
port 514 nsew
rlabel metal2 s 35952 11850 35952 11850 4 gnd
port 514 nsew
rlabel metal2 s 35952 10033 35952 10033 4 gnd
port 514 nsew
rlabel metal2 s 37200 11297 37200 11297 4 gnd
port 514 nsew
rlabel metal2 s 37200 10270 37200 10270 4 gnd
port 514 nsew
rlabel metal2 s 37200 11613 37200 11613 4 gnd
port 514 nsew
rlabel metal2 s 36432 12403 36432 12403 4 gnd
port 514 nsew
rlabel metal2 s 36432 8927 36432 8927 4 gnd
port 514 nsew
rlabel metal2 s 35952 7110 35952 7110 4 gnd
port 514 nsew
rlabel metal2 s 35952 9243 35952 9243 4 gnd
port 514 nsew
rlabel metal2 s 37200 7900 37200 7900 4 gnd
port 514 nsew
rlabel metal2 s 35952 8927 35952 8927 4 gnd
port 514 nsew
rlabel metal2 s 37200 9243 37200 9243 4 gnd
port 514 nsew
rlabel metal2 s 36432 9243 36432 9243 4 gnd
port 514 nsew
rlabel metal2 s 35952 9480 35952 9480 4 gnd
port 514 nsew
rlabel metal2 s 35952 7663 35952 7663 4 gnd
port 514 nsew
rlabel metal2 s 35184 6873 35184 6873 4 gnd
port 514 nsew
rlabel metal2 s 35952 8690 35952 8690 4 gnd
port 514 nsew
rlabel metal2 s 35184 7347 35184 7347 4 gnd
port 514 nsew
rlabel metal2 s 37200 9480 37200 9480 4 gnd
port 514 nsew
rlabel metal2 s 37200 8690 37200 8690 4 gnd
port 514 nsew
rlabel metal2 s 37200 8453 37200 8453 4 gnd
port 514 nsew
rlabel metal2 s 36432 8453 36432 8453 4 gnd
port 514 nsew
rlabel metal2 s 35184 9243 35184 9243 4 gnd
port 514 nsew
rlabel metal2 s 36432 7663 36432 7663 4 gnd
port 514 nsew
rlabel metal2 s 36432 6873 36432 6873 4 gnd
port 514 nsew
rlabel metal2 s 37200 7347 37200 7347 4 gnd
port 514 nsew
rlabel metal2 s 35184 7110 35184 7110 4 gnd
port 514 nsew
rlabel metal2 s 36432 8137 36432 8137 4 gnd
port 514 nsew
rlabel metal2 s 36432 7900 36432 7900 4 gnd
port 514 nsew
rlabel metal2 s 36432 7110 36432 7110 4 gnd
port 514 nsew
rlabel metal2 s 35952 7347 35952 7347 4 gnd
port 514 nsew
rlabel metal2 s 35952 8137 35952 8137 4 gnd
port 514 nsew
rlabel metal2 s 35184 7900 35184 7900 4 gnd
port 514 nsew
rlabel metal2 s 36432 8690 36432 8690 4 gnd
port 514 nsew
rlabel metal2 s 37200 8137 37200 8137 4 gnd
port 514 nsew
rlabel metal2 s 35952 7900 35952 7900 4 gnd
port 514 nsew
rlabel metal2 s 36432 6557 36432 6557 4 gnd
port 514 nsew
rlabel metal2 s 35184 9480 35184 9480 4 gnd
port 514 nsew
rlabel metal2 s 37200 6873 37200 6873 4 gnd
port 514 nsew
rlabel metal2 s 37200 7663 37200 7663 4 gnd
port 514 nsew
rlabel metal2 s 37200 6557 37200 6557 4 gnd
port 514 nsew
rlabel metal2 s 35184 8927 35184 8927 4 gnd
port 514 nsew
rlabel metal2 s 36432 7347 36432 7347 4 gnd
port 514 nsew
rlabel metal2 s 35952 6557 35952 6557 4 gnd
port 514 nsew
rlabel metal2 s 35184 6557 35184 6557 4 gnd
port 514 nsew
rlabel metal2 s 37200 7110 37200 7110 4 gnd
port 514 nsew
rlabel metal2 s 35952 6873 35952 6873 4 gnd
port 514 nsew
rlabel metal2 s 35184 8690 35184 8690 4 gnd
port 514 nsew
rlabel metal2 s 36432 9480 36432 9480 4 gnd
port 514 nsew
rlabel metal2 s 35952 8453 35952 8453 4 gnd
port 514 nsew
rlabel metal2 s 35184 8453 35184 8453 4 gnd
port 514 nsew
rlabel metal2 s 35184 8137 35184 8137 4 gnd
port 514 nsew
rlabel metal2 s 37200 8927 37200 8927 4 gnd
port 514 nsew
rlabel metal2 s 35184 7663 35184 7663 4 gnd
port 514 nsew
rlabel metal2 s 38928 9480 38928 9480 4 gnd
port 514 nsew
rlabel metal2 s 38448 7900 38448 7900 4 gnd
port 514 nsew
rlabel metal2 s 37680 9243 37680 9243 4 gnd
port 514 nsew
rlabel metal2 s 39696 6873 39696 6873 4 gnd
port 514 nsew
rlabel metal2 s 37680 8137 37680 8137 4 gnd
port 514 nsew
rlabel metal2 s 37680 9480 37680 9480 4 gnd
port 514 nsew
rlabel metal2 s 37680 8453 37680 8453 4 gnd
port 514 nsew
rlabel metal2 s 38448 8137 38448 8137 4 gnd
port 514 nsew
rlabel metal2 s 38448 6557 38448 6557 4 gnd
port 514 nsew
rlabel metal2 s 39696 7900 39696 7900 4 gnd
port 514 nsew
rlabel metal2 s 38448 8927 38448 8927 4 gnd
port 514 nsew
rlabel metal2 s 38928 7663 38928 7663 4 gnd
port 514 nsew
rlabel metal2 s 37680 7110 37680 7110 4 gnd
port 514 nsew
rlabel metal2 s 38448 6873 38448 6873 4 gnd
port 514 nsew
rlabel metal2 s 37680 6557 37680 6557 4 gnd
port 514 nsew
rlabel metal2 s 38928 7347 38928 7347 4 gnd
port 514 nsew
rlabel metal2 s 38928 9243 38928 9243 4 gnd
port 514 nsew
rlabel metal2 s 37680 6873 37680 6873 4 gnd
port 514 nsew
rlabel metal2 s 39696 7663 39696 7663 4 gnd
port 514 nsew
rlabel metal2 s 39696 8690 39696 8690 4 gnd
port 514 nsew
rlabel metal2 s 39696 9243 39696 9243 4 gnd
port 514 nsew
rlabel metal2 s 38448 7110 38448 7110 4 gnd
port 514 nsew
rlabel metal2 s 38928 6557 38928 6557 4 gnd
port 514 nsew
rlabel metal2 s 38448 8690 38448 8690 4 gnd
port 514 nsew
rlabel metal2 s 37680 7347 37680 7347 4 gnd
port 514 nsew
rlabel metal2 s 38928 6873 38928 6873 4 gnd
port 514 nsew
rlabel metal2 s 37680 8927 37680 8927 4 gnd
port 514 nsew
rlabel metal2 s 38448 9480 38448 9480 4 gnd
port 514 nsew
rlabel metal2 s 37680 7663 37680 7663 4 gnd
port 514 nsew
rlabel metal2 s 39696 6557 39696 6557 4 gnd
port 514 nsew
rlabel metal2 s 38928 8927 38928 8927 4 gnd
port 514 nsew
rlabel metal2 s 38928 8690 38928 8690 4 gnd
port 514 nsew
rlabel metal2 s 38928 8137 38928 8137 4 gnd
port 514 nsew
rlabel metal2 s 38928 7900 38928 7900 4 gnd
port 514 nsew
rlabel metal2 s 38928 7110 38928 7110 4 gnd
port 514 nsew
rlabel metal2 s 39696 7110 39696 7110 4 gnd
port 514 nsew
rlabel metal2 s 38448 7663 38448 7663 4 gnd
port 514 nsew
rlabel metal2 s 38928 8453 38928 8453 4 gnd
port 514 nsew
rlabel metal2 s 38448 7347 38448 7347 4 gnd
port 514 nsew
rlabel metal2 s 39696 8137 39696 8137 4 gnd
port 514 nsew
rlabel metal2 s 38448 9243 38448 9243 4 gnd
port 514 nsew
rlabel metal2 s 39696 8927 39696 8927 4 gnd
port 514 nsew
rlabel metal2 s 38448 8453 38448 8453 4 gnd
port 514 nsew
rlabel metal2 s 37680 8690 37680 8690 4 gnd
port 514 nsew
rlabel metal2 s 39696 9480 39696 9480 4 gnd
port 514 nsew
rlabel metal2 s 37680 7900 37680 7900 4 gnd
port 514 nsew
rlabel metal2 s 39696 8453 39696 8453 4 gnd
port 514 nsew
rlabel metal2 s 39696 7347 39696 7347 4 gnd
port 514 nsew
rlabel metal2 s 32688 10033 32688 10033 4 gnd
port 514 nsew
rlabel metal2 s 33456 11850 33456 11850 4 gnd
port 514 nsew
rlabel metal2 s 33936 11613 33936 11613 4 gnd
port 514 nsew
rlabel metal2 s 32688 10270 32688 10270 4 gnd
port 514 nsew
rlabel metal2 s 34704 11060 34704 11060 4 gnd
port 514 nsew
rlabel metal2 s 33936 10823 33936 10823 4 gnd
port 514 nsew
rlabel metal2 s 34704 11850 34704 11850 4 gnd
port 514 nsew
rlabel metal2 s 33936 9717 33936 9717 4 gnd
port 514 nsew
rlabel metal2 s 34704 12087 34704 12087 4 gnd
port 514 nsew
rlabel metal2 s 32688 10823 32688 10823 4 gnd
port 514 nsew
rlabel metal2 s 33456 9717 33456 9717 4 gnd
port 514 nsew
rlabel metal2 s 32688 12403 32688 12403 4 gnd
port 514 nsew
rlabel metal2 s 32688 12640 32688 12640 4 gnd
port 514 nsew
rlabel metal2 s 33936 11297 33936 11297 4 gnd
port 514 nsew
rlabel metal2 s 33456 12640 33456 12640 4 gnd
port 514 nsew
rlabel metal2 s 34704 12640 34704 12640 4 gnd
port 514 nsew
rlabel metal2 s 34704 10033 34704 10033 4 gnd
port 514 nsew
rlabel metal2 s 33936 10507 33936 10507 4 gnd
port 514 nsew
rlabel metal2 s 34704 10823 34704 10823 4 gnd
port 514 nsew
rlabel metal2 s 32688 11613 32688 11613 4 gnd
port 514 nsew
rlabel metal2 s 33456 10270 33456 10270 4 gnd
port 514 nsew
rlabel metal2 s 34704 10507 34704 10507 4 gnd
port 514 nsew
rlabel metal2 s 32688 12087 32688 12087 4 gnd
port 514 nsew
rlabel metal2 s 33456 11297 33456 11297 4 gnd
port 514 nsew
rlabel metal2 s 33456 11060 33456 11060 4 gnd
port 514 nsew
rlabel metal2 s 33456 12403 33456 12403 4 gnd
port 514 nsew
rlabel metal2 s 32688 10507 32688 10507 4 gnd
port 514 nsew
rlabel metal2 s 34704 12403 34704 12403 4 gnd
port 514 nsew
rlabel metal2 s 33456 12087 33456 12087 4 gnd
port 514 nsew
rlabel metal2 s 34704 9717 34704 9717 4 gnd
port 514 nsew
rlabel metal2 s 33936 10033 33936 10033 4 gnd
port 514 nsew
rlabel metal2 s 33456 10823 33456 10823 4 gnd
port 514 nsew
rlabel metal2 s 32688 11850 32688 11850 4 gnd
port 514 nsew
rlabel metal2 s 32688 11297 32688 11297 4 gnd
port 514 nsew
rlabel metal2 s 33936 12640 33936 12640 4 gnd
port 514 nsew
rlabel metal2 s 33456 10033 33456 10033 4 gnd
port 514 nsew
rlabel metal2 s 34704 11613 34704 11613 4 gnd
port 514 nsew
rlabel metal2 s 34704 11297 34704 11297 4 gnd
port 514 nsew
rlabel metal2 s 33936 12403 33936 12403 4 gnd
port 514 nsew
rlabel metal2 s 33456 10507 33456 10507 4 gnd
port 514 nsew
rlabel metal2 s 33936 12087 33936 12087 4 gnd
port 514 nsew
rlabel metal2 s 33936 11060 33936 11060 4 gnd
port 514 nsew
rlabel metal2 s 32688 9717 32688 9717 4 gnd
port 514 nsew
rlabel metal2 s 34704 10270 34704 10270 4 gnd
port 514 nsew
rlabel metal2 s 33936 10270 33936 10270 4 gnd
port 514 nsew
rlabel metal2 s 33936 11850 33936 11850 4 gnd
port 514 nsew
rlabel metal2 s 33456 11613 33456 11613 4 gnd
port 514 nsew
rlabel metal2 s 32688 11060 32688 11060 4 gnd
port 514 nsew
rlabel metal2 s 30192 9717 30192 9717 4 gnd
port 514 nsew
rlabel metal2 s 30192 11060 30192 11060 4 gnd
port 514 nsew
rlabel metal2 s 31440 11850 31440 11850 4 gnd
port 514 nsew
rlabel metal2 s 31440 12640 31440 12640 4 gnd
port 514 nsew
rlabel metal2 s 30960 11060 30960 11060 4 gnd
port 514 nsew
rlabel metal2 s 31440 12403 31440 12403 4 gnd
port 514 nsew
rlabel metal2 s 30960 10507 30960 10507 4 gnd
port 514 nsew
rlabel metal2 s 30192 12403 30192 12403 4 gnd
port 514 nsew
rlabel metal2 s 32208 10507 32208 10507 4 gnd
port 514 nsew
rlabel metal2 s 32208 10823 32208 10823 4 gnd
port 514 nsew
rlabel metal2 s 32208 11297 32208 11297 4 gnd
port 514 nsew
rlabel metal2 s 31440 11060 31440 11060 4 gnd
port 514 nsew
rlabel metal2 s 30192 12087 30192 12087 4 gnd
port 514 nsew
rlabel metal2 s 32208 10270 32208 10270 4 gnd
port 514 nsew
rlabel metal2 s 31440 10823 31440 10823 4 gnd
port 514 nsew
rlabel metal2 s 30960 11613 30960 11613 4 gnd
port 514 nsew
rlabel metal2 s 30192 10033 30192 10033 4 gnd
port 514 nsew
rlabel metal2 s 30960 9717 30960 9717 4 gnd
port 514 nsew
rlabel metal2 s 30960 10270 30960 10270 4 gnd
port 514 nsew
rlabel metal2 s 32208 12640 32208 12640 4 gnd
port 514 nsew
rlabel metal2 s 30192 10823 30192 10823 4 gnd
port 514 nsew
rlabel metal2 s 32208 11613 32208 11613 4 gnd
port 514 nsew
rlabel metal2 s 32208 9717 32208 9717 4 gnd
port 514 nsew
rlabel metal2 s 32208 12087 32208 12087 4 gnd
port 514 nsew
rlabel metal2 s 32208 11060 32208 11060 4 gnd
port 514 nsew
rlabel metal2 s 30192 11297 30192 11297 4 gnd
port 514 nsew
rlabel metal2 s 30960 10823 30960 10823 4 gnd
port 514 nsew
rlabel metal2 s 31440 10507 31440 10507 4 gnd
port 514 nsew
rlabel metal2 s 31440 11613 31440 11613 4 gnd
port 514 nsew
rlabel metal2 s 32208 10033 32208 10033 4 gnd
port 514 nsew
rlabel metal2 s 31440 10033 31440 10033 4 gnd
port 514 nsew
rlabel metal2 s 30192 11850 30192 11850 4 gnd
port 514 nsew
rlabel metal2 s 30960 12640 30960 12640 4 gnd
port 514 nsew
rlabel metal2 s 30960 12087 30960 12087 4 gnd
port 514 nsew
rlabel metal2 s 30960 12403 30960 12403 4 gnd
port 514 nsew
rlabel metal2 s 30960 10033 30960 10033 4 gnd
port 514 nsew
rlabel metal2 s 30192 12640 30192 12640 4 gnd
port 514 nsew
rlabel metal2 s 31440 10270 31440 10270 4 gnd
port 514 nsew
rlabel metal2 s 31440 11297 31440 11297 4 gnd
port 514 nsew
rlabel metal2 s 30960 11850 30960 11850 4 gnd
port 514 nsew
rlabel metal2 s 30192 10270 30192 10270 4 gnd
port 514 nsew
rlabel metal2 s 32208 12403 32208 12403 4 gnd
port 514 nsew
rlabel metal2 s 30192 10507 30192 10507 4 gnd
port 514 nsew
rlabel metal2 s 30192 11613 30192 11613 4 gnd
port 514 nsew
rlabel metal2 s 30960 11297 30960 11297 4 gnd
port 514 nsew
rlabel metal2 s 32208 11850 32208 11850 4 gnd
port 514 nsew
rlabel metal2 s 31440 12087 31440 12087 4 gnd
port 514 nsew
rlabel metal2 s 31440 9717 31440 9717 4 gnd
port 514 nsew
rlabel metal2 s 32208 7663 32208 7663 4 gnd
port 514 nsew
rlabel metal2 s 31440 7110 31440 7110 4 gnd
port 514 nsew
rlabel metal2 s 31440 6557 31440 6557 4 gnd
port 514 nsew
rlabel metal2 s 32208 6873 32208 6873 4 gnd
port 514 nsew
rlabel metal2 s 30960 6557 30960 6557 4 gnd
port 514 nsew
rlabel metal2 s 31440 8453 31440 8453 4 gnd
port 514 nsew
rlabel metal2 s 30960 8927 30960 8927 4 gnd
port 514 nsew
rlabel metal2 s 30960 8690 30960 8690 4 gnd
port 514 nsew
rlabel metal2 s 32208 7900 32208 7900 4 gnd
port 514 nsew
rlabel metal2 s 30192 9480 30192 9480 4 gnd
port 514 nsew
rlabel metal2 s 30960 8453 30960 8453 4 gnd
port 514 nsew
rlabel metal2 s 30960 7900 30960 7900 4 gnd
port 514 nsew
rlabel metal2 s 32208 7347 32208 7347 4 gnd
port 514 nsew
rlabel metal2 s 30960 8137 30960 8137 4 gnd
port 514 nsew
rlabel metal2 s 30192 7110 30192 7110 4 gnd
port 514 nsew
rlabel metal2 s 30960 6873 30960 6873 4 gnd
port 514 nsew
rlabel metal2 s 31440 8137 31440 8137 4 gnd
port 514 nsew
rlabel metal2 s 30192 8690 30192 8690 4 gnd
port 514 nsew
rlabel metal2 s 32208 9243 32208 9243 4 gnd
port 514 nsew
rlabel metal2 s 30192 8927 30192 8927 4 gnd
port 514 nsew
rlabel metal2 s 30192 7663 30192 7663 4 gnd
port 514 nsew
rlabel metal2 s 30192 7900 30192 7900 4 gnd
port 514 nsew
rlabel metal2 s 30192 8137 30192 8137 4 gnd
port 514 nsew
rlabel metal2 s 30960 9480 30960 9480 4 gnd
port 514 nsew
rlabel metal2 s 30960 7663 30960 7663 4 gnd
port 514 nsew
rlabel metal2 s 32208 7110 32208 7110 4 gnd
port 514 nsew
rlabel metal2 s 31440 7900 31440 7900 4 gnd
port 514 nsew
rlabel metal2 s 30960 7347 30960 7347 4 gnd
port 514 nsew
rlabel metal2 s 32208 8137 32208 8137 4 gnd
port 514 nsew
rlabel metal2 s 30960 7110 30960 7110 4 gnd
port 514 nsew
rlabel metal2 s 32208 8453 32208 8453 4 gnd
port 514 nsew
rlabel metal2 s 32208 8927 32208 8927 4 gnd
port 514 nsew
rlabel metal2 s 31440 8927 31440 8927 4 gnd
port 514 nsew
rlabel metal2 s 31440 9243 31440 9243 4 gnd
port 514 nsew
rlabel metal2 s 30192 7347 30192 7347 4 gnd
port 514 nsew
rlabel metal2 s 30192 9243 30192 9243 4 gnd
port 514 nsew
rlabel metal2 s 32208 8690 32208 8690 4 gnd
port 514 nsew
rlabel metal2 s 32208 9480 32208 9480 4 gnd
port 514 nsew
rlabel metal2 s 31440 7663 31440 7663 4 gnd
port 514 nsew
rlabel metal2 s 32208 6557 32208 6557 4 gnd
port 514 nsew
rlabel metal2 s 30192 8453 30192 8453 4 gnd
port 514 nsew
rlabel metal2 s 30192 6557 30192 6557 4 gnd
port 514 nsew
rlabel metal2 s 31440 9480 31440 9480 4 gnd
port 514 nsew
rlabel metal2 s 30192 6873 30192 6873 4 gnd
port 514 nsew
rlabel metal2 s 30960 9243 30960 9243 4 gnd
port 514 nsew
rlabel metal2 s 31440 8690 31440 8690 4 gnd
port 514 nsew
rlabel metal2 s 31440 6873 31440 6873 4 gnd
port 514 nsew
rlabel metal2 s 31440 7347 31440 7347 4 gnd
port 514 nsew
rlabel metal2 s 33936 6873 33936 6873 4 gnd
port 514 nsew
rlabel metal2 s 32688 6557 32688 6557 4 gnd
port 514 nsew
rlabel metal2 s 32688 9243 32688 9243 4 gnd
port 514 nsew
rlabel metal2 s 33456 7110 33456 7110 4 gnd
port 514 nsew
rlabel metal2 s 34704 7110 34704 7110 4 gnd
port 514 nsew
rlabel metal2 s 33456 7900 33456 7900 4 gnd
port 514 nsew
rlabel metal2 s 32688 9480 32688 9480 4 gnd
port 514 nsew
rlabel metal2 s 33456 6873 33456 6873 4 gnd
port 514 nsew
rlabel metal2 s 32688 7663 32688 7663 4 gnd
port 514 nsew
rlabel metal2 s 33456 9243 33456 9243 4 gnd
port 514 nsew
rlabel metal2 s 33456 8137 33456 8137 4 gnd
port 514 nsew
rlabel metal2 s 33936 9243 33936 9243 4 gnd
port 514 nsew
rlabel metal2 s 33456 7663 33456 7663 4 gnd
port 514 nsew
rlabel metal2 s 33936 9480 33936 9480 4 gnd
port 514 nsew
rlabel metal2 s 32688 8690 32688 8690 4 gnd
port 514 nsew
rlabel metal2 s 33936 7347 33936 7347 4 gnd
port 514 nsew
rlabel metal2 s 32688 7110 32688 7110 4 gnd
port 514 nsew
rlabel metal2 s 32688 7347 32688 7347 4 gnd
port 514 nsew
rlabel metal2 s 32688 7900 32688 7900 4 gnd
port 514 nsew
rlabel metal2 s 34704 7347 34704 7347 4 gnd
port 514 nsew
rlabel metal2 s 34704 8927 34704 8927 4 gnd
port 514 nsew
rlabel metal2 s 34704 9480 34704 9480 4 gnd
port 514 nsew
rlabel metal2 s 34704 8453 34704 8453 4 gnd
port 514 nsew
rlabel metal2 s 34704 6557 34704 6557 4 gnd
port 514 nsew
rlabel metal2 s 34704 7663 34704 7663 4 gnd
port 514 nsew
rlabel metal2 s 33936 7900 33936 7900 4 gnd
port 514 nsew
rlabel metal2 s 32688 6873 32688 6873 4 gnd
port 514 nsew
rlabel metal2 s 33936 8690 33936 8690 4 gnd
port 514 nsew
rlabel metal2 s 33456 8690 33456 8690 4 gnd
port 514 nsew
rlabel metal2 s 32688 8137 32688 8137 4 gnd
port 514 nsew
rlabel metal2 s 33456 8927 33456 8927 4 gnd
port 514 nsew
rlabel metal2 s 33936 7110 33936 7110 4 gnd
port 514 nsew
rlabel metal2 s 33936 8927 33936 8927 4 gnd
port 514 nsew
rlabel metal2 s 34704 8137 34704 8137 4 gnd
port 514 nsew
rlabel metal2 s 33936 6557 33936 6557 4 gnd
port 514 nsew
rlabel metal2 s 34704 6873 34704 6873 4 gnd
port 514 nsew
rlabel metal2 s 33936 8137 33936 8137 4 gnd
port 514 nsew
rlabel metal2 s 33936 7663 33936 7663 4 gnd
port 514 nsew
rlabel metal2 s 34704 7900 34704 7900 4 gnd
port 514 nsew
rlabel metal2 s 33456 7347 33456 7347 4 gnd
port 514 nsew
rlabel metal2 s 33456 8453 33456 8453 4 gnd
port 514 nsew
rlabel metal2 s 33936 8453 33936 8453 4 gnd
port 514 nsew
rlabel metal2 s 32688 8453 32688 8453 4 gnd
port 514 nsew
rlabel metal2 s 32688 8927 32688 8927 4 gnd
port 514 nsew
rlabel metal2 s 33456 9480 33456 9480 4 gnd
port 514 nsew
rlabel metal2 s 34704 8690 34704 8690 4 gnd
port 514 nsew
rlabel metal2 s 33456 6557 33456 6557 4 gnd
port 514 nsew
rlabel metal2 s 34704 9243 34704 9243 4 gnd
port 514 nsew
rlabel metal2 s 32688 4503 32688 4503 4 gnd
port 514 nsew
rlabel metal2 s 34704 5293 34704 5293 4 gnd
port 514 nsew
rlabel metal2 s 32688 3713 32688 3713 4 gnd
port 514 nsew
rlabel metal2 s 33456 4503 33456 4503 4 gnd
port 514 nsew
rlabel metal2 s 33456 3397 33456 3397 4 gnd
port 514 nsew
rlabel metal2 s 33936 4977 33936 4977 4 gnd
port 514 nsew
rlabel metal2 s 32688 3397 32688 3397 4 gnd
port 514 nsew
rlabel metal2 s 34704 3950 34704 3950 4 gnd
port 514 nsew
rlabel metal2 s 33936 5530 33936 5530 4 gnd
port 514 nsew
rlabel metal2 s 32688 6083 32688 6083 4 gnd
port 514 nsew
rlabel metal2 s 34704 3713 34704 3713 4 gnd
port 514 nsew
rlabel metal2 s 32688 3950 32688 3950 4 gnd
port 514 nsew
rlabel metal2 s 33936 5293 33936 5293 4 gnd
port 514 nsew
rlabel metal2 s 33936 4740 33936 4740 4 gnd
port 514 nsew
rlabel metal2 s 32688 5530 32688 5530 4 gnd
port 514 nsew
rlabel metal2 s 33456 3713 33456 3713 4 gnd
port 514 nsew
rlabel metal2 s 32688 6320 32688 6320 4 gnd
port 514 nsew
rlabel metal2 s 34704 4740 34704 4740 4 gnd
port 514 nsew
rlabel metal2 s 33456 5530 33456 5530 4 gnd
port 514 nsew
rlabel metal2 s 33456 6083 33456 6083 4 gnd
port 514 nsew
rlabel metal2 s 33936 5767 33936 5767 4 gnd
port 514 nsew
rlabel metal2 s 34704 4187 34704 4187 4 gnd
port 514 nsew
rlabel metal2 s 33936 6320 33936 6320 4 gnd
port 514 nsew
rlabel metal2 s 32688 4187 32688 4187 4 gnd
port 514 nsew
rlabel metal2 s 32688 5767 32688 5767 4 gnd
port 514 nsew
rlabel metal2 s 34704 4977 34704 4977 4 gnd
port 514 nsew
rlabel metal2 s 34704 5767 34704 5767 4 gnd
port 514 nsew
rlabel metal2 s 34704 6320 34704 6320 4 gnd
port 514 nsew
rlabel metal2 s 33456 4187 33456 4187 4 gnd
port 514 nsew
rlabel metal2 s 34704 6083 34704 6083 4 gnd
port 514 nsew
rlabel metal2 s 33936 3713 33936 3713 4 gnd
port 514 nsew
rlabel metal2 s 33936 6083 33936 6083 4 gnd
port 514 nsew
rlabel metal2 s 33456 4740 33456 4740 4 gnd
port 514 nsew
rlabel metal2 s 33936 3950 33936 3950 4 gnd
port 514 nsew
rlabel metal2 s 32688 4977 32688 4977 4 gnd
port 514 nsew
rlabel metal2 s 33456 5293 33456 5293 4 gnd
port 514 nsew
rlabel metal2 s 33456 6320 33456 6320 4 gnd
port 514 nsew
rlabel metal2 s 33936 4187 33936 4187 4 gnd
port 514 nsew
rlabel metal2 s 33936 4503 33936 4503 4 gnd
port 514 nsew
rlabel metal2 s 34704 3397 34704 3397 4 gnd
port 514 nsew
rlabel metal2 s 34704 5530 34704 5530 4 gnd
port 514 nsew
rlabel metal2 s 33456 5767 33456 5767 4 gnd
port 514 nsew
rlabel metal2 s 33456 3950 33456 3950 4 gnd
port 514 nsew
rlabel metal2 s 33456 4977 33456 4977 4 gnd
port 514 nsew
rlabel metal2 s 32688 4740 32688 4740 4 gnd
port 514 nsew
rlabel metal2 s 32688 5293 32688 5293 4 gnd
port 514 nsew
rlabel metal2 s 34704 4503 34704 4503 4 gnd
port 514 nsew
rlabel metal2 s 33936 3397 33936 3397 4 gnd
port 514 nsew
rlabel metal2 s 30192 4740 30192 4740 4 gnd
port 514 nsew
rlabel metal2 s 30960 3713 30960 3713 4 gnd
port 514 nsew
rlabel metal2 s 32208 6320 32208 6320 4 gnd
port 514 nsew
rlabel metal2 s 31440 6320 31440 6320 4 gnd
port 514 nsew
rlabel metal2 s 31440 4503 31440 4503 4 gnd
port 514 nsew
rlabel metal2 s 32208 3713 32208 3713 4 gnd
port 514 nsew
rlabel metal2 s 32208 5293 32208 5293 4 gnd
port 514 nsew
rlabel metal2 s 32208 3397 32208 3397 4 gnd
port 514 nsew
rlabel metal2 s 30960 4187 30960 4187 4 gnd
port 514 nsew
rlabel metal2 s 32208 5767 32208 5767 4 gnd
port 514 nsew
rlabel metal2 s 30960 5530 30960 5530 4 gnd
port 514 nsew
rlabel metal2 s 30192 4187 30192 4187 4 gnd
port 514 nsew
rlabel metal2 s 32208 5530 32208 5530 4 gnd
port 514 nsew
rlabel metal2 s 31440 4740 31440 4740 4 gnd
port 514 nsew
rlabel metal2 s 31440 6083 31440 6083 4 gnd
port 514 nsew
rlabel metal2 s 31440 3950 31440 3950 4 gnd
port 514 nsew
rlabel metal2 s 30960 4977 30960 4977 4 gnd
port 514 nsew
rlabel metal2 s 30960 5767 30960 5767 4 gnd
port 514 nsew
rlabel metal2 s 30960 3950 30960 3950 4 gnd
port 514 nsew
rlabel metal2 s 30192 6320 30192 6320 4 gnd
port 514 nsew
rlabel metal2 s 32208 3950 32208 3950 4 gnd
port 514 nsew
rlabel metal2 s 32208 6083 32208 6083 4 gnd
port 514 nsew
rlabel metal2 s 30960 5293 30960 5293 4 gnd
port 514 nsew
rlabel metal2 s 31440 4187 31440 4187 4 gnd
port 514 nsew
rlabel metal2 s 31440 5293 31440 5293 4 gnd
port 514 nsew
rlabel metal2 s 30192 5767 30192 5767 4 gnd
port 514 nsew
rlabel metal2 s 30192 3713 30192 3713 4 gnd
port 514 nsew
rlabel metal2 s 31440 5767 31440 5767 4 gnd
port 514 nsew
rlabel metal2 s 30192 4503 30192 4503 4 gnd
port 514 nsew
rlabel metal2 s 30192 4977 30192 4977 4 gnd
port 514 nsew
rlabel metal2 s 31440 4977 31440 4977 4 gnd
port 514 nsew
rlabel metal2 s 30960 6083 30960 6083 4 gnd
port 514 nsew
rlabel metal2 s 30960 6320 30960 6320 4 gnd
port 514 nsew
rlabel metal2 s 30960 4740 30960 4740 4 gnd
port 514 nsew
rlabel metal2 s 32208 4187 32208 4187 4 gnd
port 514 nsew
rlabel metal2 s 31440 3713 31440 3713 4 gnd
port 514 nsew
rlabel metal2 s 32208 4977 32208 4977 4 gnd
port 514 nsew
rlabel metal2 s 31440 3397 31440 3397 4 gnd
port 514 nsew
rlabel metal2 s 30192 6083 30192 6083 4 gnd
port 514 nsew
rlabel metal2 s 30960 3397 30960 3397 4 gnd
port 514 nsew
rlabel metal2 s 30192 3950 30192 3950 4 gnd
port 514 nsew
rlabel metal2 s 30960 4503 30960 4503 4 gnd
port 514 nsew
rlabel metal2 s 32208 4740 32208 4740 4 gnd
port 514 nsew
rlabel metal2 s 32208 4503 32208 4503 4 gnd
port 514 nsew
rlabel metal2 s 30192 3397 30192 3397 4 gnd
port 514 nsew
rlabel metal2 s 30192 5530 30192 5530 4 gnd
port 514 nsew
rlabel metal2 s 30192 5293 30192 5293 4 gnd
port 514 nsew
rlabel metal2 s 31440 5530 31440 5530 4 gnd
port 514 nsew
rlabel metal2 s 30192 3160 30192 3160 4 gnd
port 514 nsew
rlabel metal2 s 30192 237 30192 237 4 gnd
port 514 nsew
rlabel metal2 s 31440 237 31440 237 4 gnd
port 514 nsew
rlabel metal2 s 31440 0 31440 0 4 gnd
port 514 nsew
rlabel metal2 s 30960 2607 30960 2607 4 gnd
port 514 nsew
rlabel metal2 s 32208 3160 32208 3160 4 gnd
port 514 nsew
rlabel metal2 s 32208 1027 32208 1027 4 gnd
port 514 nsew
rlabel metal2 s 30960 2923 30960 2923 4 gnd
port 514 nsew
rlabel metal2 s 30960 1343 30960 1343 4 gnd
port 514 nsew
rlabel metal2 s 31440 2607 31440 2607 4 gnd
port 514 nsew
rlabel metal2 s 30960 0 30960 0 4 gnd
port 514 nsew
rlabel metal2 s 30192 1817 30192 1817 4 gnd
port 514 nsew
rlabel metal2 s 30960 553 30960 553 4 gnd
port 514 nsew
rlabel metal2 s 30192 1027 30192 1027 4 gnd
port 514 nsew
rlabel metal2 s 32208 1817 32208 1817 4 gnd
port 514 nsew
rlabel metal2 s 32208 553 32208 553 4 gnd
port 514 nsew
rlabel metal2 s 30192 553 30192 553 4 gnd
port 514 nsew
rlabel metal2 s 30192 2370 30192 2370 4 gnd
port 514 nsew
rlabel metal2 s 32208 2607 32208 2607 4 gnd
port 514 nsew
rlabel metal2 s 30192 2607 30192 2607 4 gnd
port 514 nsew
rlabel metal2 s 32208 2133 32208 2133 4 gnd
port 514 nsew
rlabel metal2 s 30960 237 30960 237 4 gnd
port 514 nsew
rlabel metal2 s 30960 2370 30960 2370 4 gnd
port 514 nsew
rlabel metal2 s 31440 1817 31440 1817 4 gnd
port 514 nsew
rlabel metal2 s 30192 1580 30192 1580 4 gnd
port 514 nsew
rlabel metal2 s 30960 2133 30960 2133 4 gnd
port 514 nsew
rlabel metal2 s 31440 2370 31440 2370 4 gnd
port 514 nsew
rlabel metal2 s 31440 1027 31440 1027 4 gnd
port 514 nsew
rlabel metal2 s 31440 1343 31440 1343 4 gnd
port 514 nsew
rlabel metal2 s 30192 2133 30192 2133 4 gnd
port 514 nsew
rlabel metal2 s 30960 3160 30960 3160 4 gnd
port 514 nsew
rlabel metal2 s 32208 2923 32208 2923 4 gnd
port 514 nsew
rlabel metal2 s 31440 2133 31440 2133 4 gnd
port 514 nsew
rlabel metal2 s 32208 0 32208 0 4 gnd
port 514 nsew
rlabel metal2 s 30192 1343 30192 1343 4 gnd
port 514 nsew
rlabel metal2 s 32208 790 32208 790 4 gnd
port 514 nsew
rlabel metal2 s 31440 790 31440 790 4 gnd
port 514 nsew
rlabel metal2 s 30960 1817 30960 1817 4 gnd
port 514 nsew
rlabel metal2 s 32208 1580 32208 1580 4 gnd
port 514 nsew
rlabel metal2 s 32208 1343 32208 1343 4 gnd
port 514 nsew
rlabel metal2 s 30960 790 30960 790 4 gnd
port 514 nsew
rlabel metal2 s 31440 2923 31440 2923 4 gnd
port 514 nsew
rlabel metal2 s 30192 2923 30192 2923 4 gnd
port 514 nsew
rlabel metal2 s 30960 1580 30960 1580 4 gnd
port 514 nsew
rlabel metal2 s 30192 790 30192 790 4 gnd
port 514 nsew
rlabel metal2 s 32208 2370 32208 2370 4 gnd
port 514 nsew
rlabel metal2 s 32208 237 32208 237 4 gnd
port 514 nsew
rlabel metal2 s 31440 3160 31440 3160 4 gnd
port 514 nsew
rlabel metal2 s 30960 1027 30960 1027 4 gnd
port 514 nsew
rlabel metal2 s 31440 553 31440 553 4 gnd
port 514 nsew
rlabel metal2 s 30192 0 30192 0 4 gnd
port 514 nsew
rlabel metal2 s 31440 1580 31440 1580 4 gnd
port 514 nsew
rlabel metal2 s 32688 1343 32688 1343 4 gnd
port 514 nsew
rlabel metal2 s 33936 2923 33936 2923 4 gnd
port 514 nsew
rlabel metal2 s 33936 1027 33936 1027 4 gnd
port 514 nsew
rlabel metal2 s 33936 3160 33936 3160 4 gnd
port 514 nsew
rlabel metal2 s 33936 1817 33936 1817 4 gnd
port 514 nsew
rlabel metal2 s 33456 0 33456 0 4 gnd
port 514 nsew
rlabel metal2 s 33936 0 33936 0 4 gnd
port 514 nsew
rlabel metal2 s 34704 790 34704 790 4 gnd
port 514 nsew
rlabel metal2 s 33936 2133 33936 2133 4 gnd
port 514 nsew
rlabel metal2 s 33936 2370 33936 2370 4 gnd
port 514 nsew
rlabel metal2 s 32688 790 32688 790 4 gnd
port 514 nsew
rlabel metal2 s 33456 1343 33456 1343 4 gnd
port 514 nsew
rlabel metal2 s 34704 1580 34704 1580 4 gnd
port 514 nsew
rlabel metal2 s 32688 2133 32688 2133 4 gnd
port 514 nsew
rlabel metal2 s 32688 237 32688 237 4 gnd
port 514 nsew
rlabel metal2 s 32688 1027 32688 1027 4 gnd
port 514 nsew
rlabel metal2 s 33456 2923 33456 2923 4 gnd
port 514 nsew
rlabel metal2 s 32688 1580 32688 1580 4 gnd
port 514 nsew
rlabel metal2 s 34704 2607 34704 2607 4 gnd
port 514 nsew
rlabel metal2 s 33456 790 33456 790 4 gnd
port 514 nsew
rlabel metal2 s 32688 2370 32688 2370 4 gnd
port 514 nsew
rlabel metal2 s 33936 790 33936 790 4 gnd
port 514 nsew
rlabel metal2 s 32688 1817 32688 1817 4 gnd
port 514 nsew
rlabel metal2 s 33936 237 33936 237 4 gnd
port 514 nsew
rlabel metal2 s 34704 1343 34704 1343 4 gnd
port 514 nsew
rlabel metal2 s 33936 1343 33936 1343 4 gnd
port 514 nsew
rlabel metal2 s 33456 2607 33456 2607 4 gnd
port 514 nsew
rlabel metal2 s 33456 1817 33456 1817 4 gnd
port 514 nsew
rlabel metal2 s 32688 0 32688 0 4 gnd
port 514 nsew
rlabel metal2 s 33456 1027 33456 1027 4 gnd
port 514 nsew
rlabel metal2 s 33456 3160 33456 3160 4 gnd
port 514 nsew
rlabel metal2 s 34704 1027 34704 1027 4 gnd
port 514 nsew
rlabel metal2 s 33456 237 33456 237 4 gnd
port 514 nsew
rlabel metal2 s 33936 2607 33936 2607 4 gnd
port 514 nsew
rlabel metal2 s 33456 2133 33456 2133 4 gnd
port 514 nsew
rlabel metal2 s 32688 2923 32688 2923 4 gnd
port 514 nsew
rlabel metal2 s 32688 553 32688 553 4 gnd
port 514 nsew
rlabel metal2 s 34704 553 34704 553 4 gnd
port 514 nsew
rlabel metal2 s 34704 1817 34704 1817 4 gnd
port 514 nsew
rlabel metal2 s 34704 237 34704 237 4 gnd
port 514 nsew
rlabel metal2 s 34704 2133 34704 2133 4 gnd
port 514 nsew
rlabel metal2 s 34704 2923 34704 2923 4 gnd
port 514 nsew
rlabel metal2 s 33456 553 33456 553 4 gnd
port 514 nsew
rlabel metal2 s 34704 3160 34704 3160 4 gnd
port 514 nsew
rlabel metal2 s 32688 3160 32688 3160 4 gnd
port 514 nsew
rlabel metal2 s 33456 2370 33456 2370 4 gnd
port 514 nsew
rlabel metal2 s 33456 1580 33456 1580 4 gnd
port 514 nsew
rlabel metal2 s 34704 0 34704 0 4 gnd
port 514 nsew
rlabel metal2 s 33936 1580 33936 1580 4 gnd
port 514 nsew
rlabel metal2 s 33936 553 33936 553 4 gnd
port 514 nsew
rlabel metal2 s 34704 2370 34704 2370 4 gnd
port 514 nsew
rlabel metal2 s 32688 2607 32688 2607 4 gnd
port 514 nsew
rlabel metal2 s 38448 3950 38448 3950 4 gnd
port 514 nsew
rlabel metal2 s 38448 6320 38448 6320 4 gnd
port 514 nsew
rlabel metal2 s 38448 4503 38448 4503 4 gnd
port 514 nsew
rlabel metal2 s 38448 4740 38448 4740 4 gnd
port 514 nsew
rlabel metal2 s 38928 3397 38928 3397 4 gnd
port 514 nsew
rlabel metal2 s 39696 6083 39696 6083 4 gnd
port 514 nsew
rlabel metal2 s 37680 5293 37680 5293 4 gnd
port 514 nsew
rlabel metal2 s 37680 4740 37680 4740 4 gnd
port 514 nsew
rlabel metal2 s 38448 6083 38448 6083 4 gnd
port 514 nsew
rlabel metal2 s 39696 3713 39696 3713 4 gnd
port 514 nsew
rlabel metal2 s 39696 3950 39696 3950 4 gnd
port 514 nsew
rlabel metal2 s 39696 5293 39696 5293 4 gnd
port 514 nsew
rlabel metal2 s 39696 4740 39696 4740 4 gnd
port 514 nsew
rlabel metal2 s 39696 6320 39696 6320 4 gnd
port 514 nsew
rlabel metal2 s 37680 3397 37680 3397 4 gnd
port 514 nsew
rlabel metal2 s 39696 4503 39696 4503 4 gnd
port 514 nsew
rlabel metal2 s 38448 4977 38448 4977 4 gnd
port 514 nsew
rlabel metal2 s 39696 3397 39696 3397 4 gnd
port 514 nsew
rlabel metal2 s 38928 5293 38928 5293 4 gnd
port 514 nsew
rlabel metal2 s 37680 3950 37680 3950 4 gnd
port 514 nsew
rlabel metal2 s 38928 6083 38928 6083 4 gnd
port 514 nsew
rlabel metal2 s 38448 3397 38448 3397 4 gnd
port 514 nsew
rlabel metal2 s 38928 4187 38928 4187 4 gnd
port 514 nsew
rlabel metal2 s 37680 4977 37680 4977 4 gnd
port 514 nsew
rlabel metal2 s 38928 6320 38928 6320 4 gnd
port 514 nsew
rlabel metal2 s 38448 4187 38448 4187 4 gnd
port 514 nsew
rlabel metal2 s 37680 4503 37680 4503 4 gnd
port 514 nsew
rlabel metal2 s 38448 3713 38448 3713 4 gnd
port 514 nsew
rlabel metal2 s 38928 4977 38928 4977 4 gnd
port 514 nsew
rlabel metal2 s 39696 5767 39696 5767 4 gnd
port 514 nsew
rlabel metal2 s 38928 3950 38928 3950 4 gnd
port 514 nsew
rlabel metal2 s 38448 5767 38448 5767 4 gnd
port 514 nsew
rlabel metal2 s 39696 4977 39696 4977 4 gnd
port 514 nsew
rlabel metal2 s 38928 3713 38928 3713 4 gnd
port 514 nsew
rlabel metal2 s 37680 6083 37680 6083 4 gnd
port 514 nsew
rlabel metal2 s 37680 3713 37680 3713 4 gnd
port 514 nsew
rlabel metal2 s 39696 4187 39696 4187 4 gnd
port 514 nsew
rlabel metal2 s 38448 5293 38448 5293 4 gnd
port 514 nsew
rlabel metal2 s 39696 5530 39696 5530 4 gnd
port 514 nsew
rlabel metal2 s 37680 4187 37680 4187 4 gnd
port 514 nsew
rlabel metal2 s 37680 5530 37680 5530 4 gnd
port 514 nsew
rlabel metal2 s 38928 4503 38928 4503 4 gnd
port 514 nsew
rlabel metal2 s 37680 6320 37680 6320 4 gnd
port 514 nsew
rlabel metal2 s 38928 4740 38928 4740 4 gnd
port 514 nsew
rlabel metal2 s 38928 5767 38928 5767 4 gnd
port 514 nsew
rlabel metal2 s 38448 5530 38448 5530 4 gnd
port 514 nsew
rlabel metal2 s 37680 5767 37680 5767 4 gnd
port 514 nsew
rlabel metal2 s 38928 5530 38928 5530 4 gnd
port 514 nsew
rlabel metal2 s 35952 3950 35952 3950 4 gnd
port 514 nsew
rlabel metal2 s 36432 4740 36432 4740 4 gnd
port 514 nsew
rlabel metal2 s 36432 3397 36432 3397 4 gnd
port 514 nsew
rlabel metal2 s 35952 4740 35952 4740 4 gnd
port 514 nsew
rlabel metal2 s 35184 3397 35184 3397 4 gnd
port 514 nsew
rlabel metal2 s 35952 4503 35952 4503 4 gnd
port 514 nsew
rlabel metal2 s 37200 3397 37200 3397 4 gnd
port 514 nsew
rlabel metal2 s 37200 5767 37200 5767 4 gnd
port 514 nsew
rlabel metal2 s 35184 6083 35184 6083 4 gnd
port 514 nsew
rlabel metal2 s 35952 5293 35952 5293 4 gnd
port 514 nsew
rlabel metal2 s 35184 5767 35184 5767 4 gnd
port 514 nsew
rlabel metal2 s 36432 6320 36432 6320 4 gnd
port 514 nsew
rlabel metal2 s 37200 4187 37200 4187 4 gnd
port 514 nsew
rlabel metal2 s 36432 4977 36432 4977 4 gnd
port 514 nsew
rlabel metal2 s 37200 3713 37200 3713 4 gnd
port 514 nsew
rlabel metal2 s 36432 5530 36432 5530 4 gnd
port 514 nsew
rlabel metal2 s 35184 4187 35184 4187 4 gnd
port 514 nsew
rlabel metal2 s 35952 6320 35952 6320 4 gnd
port 514 nsew
rlabel metal2 s 35184 6320 35184 6320 4 gnd
port 514 nsew
rlabel metal2 s 35184 4977 35184 4977 4 gnd
port 514 nsew
rlabel metal2 s 35952 3713 35952 3713 4 gnd
port 514 nsew
rlabel metal2 s 35952 6083 35952 6083 4 gnd
port 514 nsew
rlabel metal2 s 37200 4503 37200 4503 4 gnd
port 514 nsew
rlabel metal2 s 35952 5767 35952 5767 4 gnd
port 514 nsew
rlabel metal2 s 36432 6083 36432 6083 4 gnd
port 514 nsew
rlabel metal2 s 35184 4740 35184 4740 4 gnd
port 514 nsew
rlabel metal2 s 36432 4503 36432 4503 4 gnd
port 514 nsew
rlabel metal2 s 35184 4503 35184 4503 4 gnd
port 514 nsew
rlabel metal2 s 37200 6083 37200 6083 4 gnd
port 514 nsew
rlabel metal2 s 35184 3713 35184 3713 4 gnd
port 514 nsew
rlabel metal2 s 35952 5530 35952 5530 4 gnd
port 514 nsew
rlabel metal2 s 37200 5530 37200 5530 4 gnd
port 514 nsew
rlabel metal2 s 35952 4187 35952 4187 4 gnd
port 514 nsew
rlabel metal2 s 36432 3713 36432 3713 4 gnd
port 514 nsew
rlabel metal2 s 36432 4187 36432 4187 4 gnd
port 514 nsew
rlabel metal2 s 37200 3950 37200 3950 4 gnd
port 514 nsew
rlabel metal2 s 35952 4977 35952 4977 4 gnd
port 514 nsew
rlabel metal2 s 37200 4740 37200 4740 4 gnd
port 514 nsew
rlabel metal2 s 35184 5530 35184 5530 4 gnd
port 514 nsew
rlabel metal2 s 35184 5293 35184 5293 4 gnd
port 514 nsew
rlabel metal2 s 37200 6320 37200 6320 4 gnd
port 514 nsew
rlabel metal2 s 37200 5293 37200 5293 4 gnd
port 514 nsew
rlabel metal2 s 35184 3950 35184 3950 4 gnd
port 514 nsew
rlabel metal2 s 35952 3397 35952 3397 4 gnd
port 514 nsew
rlabel metal2 s 37200 4977 37200 4977 4 gnd
port 514 nsew
rlabel metal2 s 36432 5293 36432 5293 4 gnd
port 514 nsew
rlabel metal2 s 36432 3950 36432 3950 4 gnd
port 514 nsew
rlabel metal2 s 36432 5767 36432 5767 4 gnd
port 514 nsew
rlabel metal2 s 36432 237 36432 237 4 gnd
port 514 nsew
rlabel metal2 s 35184 0 35184 0 4 gnd
port 514 nsew
rlabel metal2 s 35952 2370 35952 2370 4 gnd
port 514 nsew
rlabel metal2 s 35184 2370 35184 2370 4 gnd
port 514 nsew
rlabel metal2 s 36432 0 36432 0 4 gnd
port 514 nsew
rlabel metal2 s 35184 553 35184 553 4 gnd
port 514 nsew
rlabel metal2 s 37200 237 37200 237 4 gnd
port 514 nsew
rlabel metal2 s 37200 1817 37200 1817 4 gnd
port 514 nsew
rlabel metal2 s 35184 790 35184 790 4 gnd
port 514 nsew
rlabel metal2 s 37200 1343 37200 1343 4 gnd
port 514 nsew
rlabel metal2 s 35184 1580 35184 1580 4 gnd
port 514 nsew
rlabel metal2 s 35184 2923 35184 2923 4 gnd
port 514 nsew
rlabel metal2 s 37200 2133 37200 2133 4 gnd
port 514 nsew
rlabel metal2 s 36432 2133 36432 2133 4 gnd
port 514 nsew
rlabel metal2 s 37200 1580 37200 1580 4 gnd
port 514 nsew
rlabel metal2 s 36432 2607 36432 2607 4 gnd
port 514 nsew
rlabel metal2 s 35184 1027 35184 1027 4 gnd
port 514 nsew
rlabel metal2 s 35184 237 35184 237 4 gnd
port 514 nsew
rlabel metal2 s 36432 1027 36432 1027 4 gnd
port 514 nsew
rlabel metal2 s 35952 237 35952 237 4 gnd
port 514 nsew
rlabel metal2 s 36432 1580 36432 1580 4 gnd
port 514 nsew
rlabel metal2 s 37200 0 37200 0 4 gnd
port 514 nsew
rlabel metal2 s 37200 790 37200 790 4 gnd
port 514 nsew
rlabel metal2 s 35184 2133 35184 2133 4 gnd
port 514 nsew
rlabel metal2 s 36432 1343 36432 1343 4 gnd
port 514 nsew
rlabel metal2 s 37200 3160 37200 3160 4 gnd
port 514 nsew
rlabel metal2 s 35952 1343 35952 1343 4 gnd
port 514 nsew
rlabel metal2 s 36432 790 36432 790 4 gnd
port 514 nsew
rlabel metal2 s 35952 553 35952 553 4 gnd
port 514 nsew
rlabel metal2 s 36432 553 36432 553 4 gnd
port 514 nsew
rlabel metal2 s 35952 2607 35952 2607 4 gnd
port 514 nsew
rlabel metal2 s 36432 2923 36432 2923 4 gnd
port 514 nsew
rlabel metal2 s 37200 1027 37200 1027 4 gnd
port 514 nsew
rlabel metal2 s 37200 2370 37200 2370 4 gnd
port 514 nsew
rlabel metal2 s 36432 3160 36432 3160 4 gnd
port 514 nsew
rlabel metal2 s 36432 1817 36432 1817 4 gnd
port 514 nsew
rlabel metal2 s 35952 790 35952 790 4 gnd
port 514 nsew
rlabel metal2 s 35184 3160 35184 3160 4 gnd
port 514 nsew
rlabel metal2 s 35952 2133 35952 2133 4 gnd
port 514 nsew
rlabel metal2 s 35952 3160 35952 3160 4 gnd
port 514 nsew
rlabel metal2 s 35184 2607 35184 2607 4 gnd
port 514 nsew
rlabel metal2 s 37200 2607 37200 2607 4 gnd
port 514 nsew
rlabel metal2 s 35184 1817 35184 1817 4 gnd
port 514 nsew
rlabel metal2 s 35952 1027 35952 1027 4 gnd
port 514 nsew
rlabel metal2 s 35952 0 35952 0 4 gnd
port 514 nsew
rlabel metal2 s 37200 553 37200 553 4 gnd
port 514 nsew
rlabel metal2 s 35952 2923 35952 2923 4 gnd
port 514 nsew
rlabel metal2 s 35184 1343 35184 1343 4 gnd
port 514 nsew
rlabel metal2 s 37200 2923 37200 2923 4 gnd
port 514 nsew
rlabel metal2 s 36432 2370 36432 2370 4 gnd
port 514 nsew
rlabel metal2 s 35952 1580 35952 1580 4 gnd
port 514 nsew
rlabel metal2 s 35952 1817 35952 1817 4 gnd
port 514 nsew
rlabel metal2 s 37680 1817 37680 1817 4 gnd
port 514 nsew
rlabel metal2 s 38928 1580 38928 1580 4 gnd
port 514 nsew
rlabel metal2 s 38448 2607 38448 2607 4 gnd
port 514 nsew
rlabel metal2 s 39696 1817 39696 1817 4 gnd
port 514 nsew
rlabel metal2 s 39696 1027 39696 1027 4 gnd
port 514 nsew
rlabel metal2 s 38448 1027 38448 1027 4 gnd
port 514 nsew
rlabel metal2 s 38448 553 38448 553 4 gnd
port 514 nsew
rlabel metal2 s 39696 1580 39696 1580 4 gnd
port 514 nsew
rlabel metal2 s 38928 1027 38928 1027 4 gnd
port 514 nsew
rlabel metal2 s 38928 3160 38928 3160 4 gnd
port 514 nsew
rlabel metal2 s 38928 237 38928 237 4 gnd
port 514 nsew
rlabel metal2 s 39696 3160 39696 3160 4 gnd
port 514 nsew
rlabel metal2 s 38928 2370 38928 2370 4 gnd
port 514 nsew
rlabel metal2 s 38448 0 38448 0 4 gnd
port 514 nsew
rlabel metal2 s 39696 2607 39696 2607 4 gnd
port 514 nsew
rlabel metal2 s 38448 1580 38448 1580 4 gnd
port 514 nsew
rlabel metal2 s 37680 237 37680 237 4 gnd
port 514 nsew
rlabel metal2 s 38448 1343 38448 1343 4 gnd
port 514 nsew
rlabel metal2 s 39696 790 39696 790 4 gnd
port 514 nsew
rlabel metal2 s 38448 2923 38448 2923 4 gnd
port 514 nsew
rlabel metal2 s 38448 237 38448 237 4 gnd
port 514 nsew
rlabel metal2 s 38448 2370 38448 2370 4 gnd
port 514 nsew
rlabel metal2 s 37680 1343 37680 1343 4 gnd
port 514 nsew
rlabel metal2 s 38928 2923 38928 2923 4 gnd
port 514 nsew
rlabel metal2 s 38928 553 38928 553 4 gnd
port 514 nsew
rlabel metal2 s 39696 1343 39696 1343 4 gnd
port 514 nsew
rlabel metal2 s 38928 1343 38928 1343 4 gnd
port 514 nsew
rlabel metal2 s 39696 2370 39696 2370 4 gnd
port 514 nsew
rlabel metal2 s 37680 1580 37680 1580 4 gnd
port 514 nsew
rlabel metal2 s 38928 1817 38928 1817 4 gnd
port 514 nsew
rlabel metal2 s 37680 1027 37680 1027 4 gnd
port 514 nsew
rlabel metal2 s 38448 1817 38448 1817 4 gnd
port 514 nsew
rlabel metal2 s 38928 0 38928 0 4 gnd
port 514 nsew
rlabel metal2 s 39696 2923 39696 2923 4 gnd
port 514 nsew
rlabel metal2 s 38448 3160 38448 3160 4 gnd
port 514 nsew
rlabel metal2 s 37680 2370 37680 2370 4 gnd
port 514 nsew
rlabel metal2 s 39696 0 39696 0 4 gnd
port 514 nsew
rlabel metal2 s 38928 2133 38928 2133 4 gnd
port 514 nsew
rlabel metal2 s 39696 553 39696 553 4 gnd
port 514 nsew
rlabel metal2 s 38448 790 38448 790 4 gnd
port 514 nsew
rlabel metal2 s 37680 2133 37680 2133 4 gnd
port 514 nsew
rlabel metal2 s 38448 2133 38448 2133 4 gnd
port 514 nsew
rlabel metal2 s 39696 237 39696 237 4 gnd
port 514 nsew
rlabel metal2 s 37680 3160 37680 3160 4 gnd
port 514 nsew
rlabel metal2 s 37680 2923 37680 2923 4 gnd
port 514 nsew
rlabel metal2 s 38928 790 38928 790 4 gnd
port 514 nsew
rlabel metal2 s 37680 0 37680 0 4 gnd
port 514 nsew
rlabel metal2 s 39696 2133 39696 2133 4 gnd
port 514 nsew
rlabel metal2 s 38928 2607 38928 2607 4 gnd
port 514 nsew
rlabel metal2 s 37680 2607 37680 2607 4 gnd
port 514 nsew
rlabel metal2 s 37680 790 37680 790 4 gnd
port 514 nsew
rlabel metal2 s 37680 553 37680 553 4 gnd
port 514 nsew
<< properties >>
string FIXED_BBOX 0 0 39936 50560
string GDS_END 3370912
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 239660
<< end >>
