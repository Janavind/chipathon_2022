magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -54 252 420 390
rect -59 84 425 252
rect -54 -54 420 84
<< scpmos >>
rect 60 0 90 336
rect 168 0 198 336
rect 276 0 306 336
<< pdiff >>
rect 0 185 60 336
rect 0 151 8 185
rect 42 151 60 185
rect 0 0 60 151
rect 90 185 168 336
rect 90 151 112 185
rect 146 151 168 185
rect 90 0 168 151
rect 198 185 276 336
rect 198 151 220 185
rect 254 151 276 185
rect 198 0 276 151
rect 306 185 366 336
rect 306 151 324 185
rect 358 151 366 185
rect 306 0 366 151
<< pdiffc >>
rect 8 151 42 185
rect 112 151 146 185
rect 220 151 254 185
rect 324 151 358 185
<< poly >>
rect 60 336 90 362
rect 168 336 198 362
rect 276 336 306 362
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 60 -56 306 -26
<< locali >>
rect 8 185 42 201
rect 8 135 42 151
rect 112 185 146 201
rect 112 101 146 151
rect 220 185 254 201
rect 220 135 254 151
rect 324 185 358 201
rect 324 101 358 151
rect 112 67 358 101
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_12  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_12_0
timestamp 1666199351
transform 1 0 316 0 1 135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_12  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_12_1
timestamp 1666199351
transform 1 0 212 0 1 135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_12  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_12_2
timestamp 1666199351
transform 1 0 104 0 1 135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_12  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_12_3
timestamp 1666199351
transform 1 0 0 0 1 135
box 0 0 1 1
<< labels >>
rlabel locali s 25 168 25 168 4 S
port 1 nsew
rlabel locali s 237 168 237 168 4 S
port 1 nsew
rlabel locali s 235 84 235 84 4 D
port 2 nsew
rlabel poly s 183 -41 183 -41 4 G
port 3 nsew
<< properties >>
string FIXED_BBOX -54 -56 420 84
string GDS_END 42980
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 41608
<< end >>
