magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 98 157 940 203
rect 1 21 1195 157
rect 30 -17 64 21
<< locali >>
rect 86 153 156 327
rect 192 309 432 343
rect 192 164 248 309
rect 192 130 416 164
rect 214 51 248 130
rect 382 51 416 130
rect 536 199 616 265
rect 650 151 709 265
rect 1097 199 1169 324
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 417 69 493
rect 103 451 169 527
rect 282 451 348 527
rect 450 451 516 527
rect 666 451 732 527
rect 872 451 1074 527
rect 1127 417 1161 493
rect 17 383 898 417
rect 17 117 52 383
rect 466 309 830 343
rect 466 249 500 309
rect 864 265 898 383
rect 282 215 500 249
rect 17 51 69 117
rect 114 17 180 94
rect 282 17 348 94
rect 466 157 500 215
rect 466 123 588 157
rect 746 231 898 265
rect 990 383 1161 417
rect 746 199 780 231
rect 990 165 1024 383
rect 554 94 588 123
rect 851 94 922 162
rect 990 131 1161 165
rect 454 17 520 89
rect 554 60 922 94
rect 995 17 1061 93
rect 1127 51 1161 131
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 1097 199 1169 324 6 A_N
port 1 nsew signal input
rlabel locali s 86 153 156 327 6 B_N
port 2 nsew signal input
rlabel locali s 650 151 709 265 6 C
port 3 nsew signal input
rlabel locali s 536 199 616 265 6 D
port 4 nsew signal input
rlabel metal1 s 0 -48 1196 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 1195 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 98 157 940 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 382 51 416 130 6 X
port 9 nsew signal output
rlabel locali s 214 51 248 130 6 X
port 9 nsew signal output
rlabel locali s 192 130 416 164 6 X
port 9 nsew signal output
rlabel locali s 192 164 248 309 6 X
port 9 nsew signal output
rlabel locali s 192 309 432 343 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1196 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3106168
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3097510
<< end >>
