magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< dnwell >>
rect 214 214 1778 3178
<< nwell >>
rect 134 2898 1858 3258
rect 134 494 494 2898
rect 1498 494 1858 2898
rect 134 134 1858 494
<< pwell >>
rect 0 3258 1992 3392
rect 0 134 134 3258
rect 628 628 1364 2764
rect 1858 134 1992 3258
rect 0 0 1992 134
<< ndiff >>
rect 896 2461 1096 2496
rect 896 931 911 2461
rect 1081 931 1096 2461
rect 896 896 1096 931
<< ndiffc >>
rect 911 931 1081 2461
<< psubdiff >>
rect 26 3342 1966 3366
rect 26 3308 50 3342
rect 84 3308 129 3342
rect 163 3308 197 3342
rect 231 3308 265 3342
rect 299 3308 333 3342
rect 367 3308 401 3342
rect 435 3308 469 3342
rect 503 3308 537 3342
rect 571 3308 605 3342
rect 639 3308 673 3342
rect 707 3308 741 3342
rect 775 3308 809 3342
rect 843 3308 877 3342
rect 911 3308 945 3342
rect 979 3308 1013 3342
rect 1047 3308 1081 3342
rect 1115 3308 1149 3342
rect 1183 3308 1217 3342
rect 1251 3308 1285 3342
rect 1319 3308 1353 3342
rect 1387 3308 1421 3342
rect 1455 3308 1489 3342
rect 1523 3308 1557 3342
rect 1591 3308 1625 3342
rect 1659 3308 1693 3342
rect 1727 3308 1761 3342
rect 1795 3308 1829 3342
rect 1863 3308 1908 3342
rect 1942 3308 1966 3342
rect 26 3284 1966 3308
rect 26 3243 108 3284
rect 26 3209 50 3243
rect 84 3209 108 3243
rect 26 3175 108 3209
rect 26 3141 50 3175
rect 84 3141 108 3175
rect 26 3107 108 3141
rect 1884 3243 1966 3284
rect 1884 3209 1908 3243
rect 1942 3209 1966 3243
rect 1884 3175 1966 3209
rect 1884 3141 1908 3175
rect 1942 3141 1966 3175
rect 26 3073 50 3107
rect 84 3073 108 3107
rect 26 3039 108 3073
rect 26 3005 50 3039
rect 84 3005 108 3039
rect 26 2971 108 3005
rect 26 2937 50 2971
rect 84 2937 108 2971
rect 26 2903 108 2937
rect 26 2869 50 2903
rect 84 2869 108 2903
rect 26 2835 108 2869
rect 26 2801 50 2835
rect 84 2801 108 2835
rect 26 2767 108 2801
rect 26 2733 50 2767
rect 84 2733 108 2767
rect 26 2699 108 2733
rect 26 2665 50 2699
rect 84 2665 108 2699
rect 26 2631 108 2665
rect 26 2597 50 2631
rect 84 2597 108 2631
rect 26 2563 108 2597
rect 26 2529 50 2563
rect 84 2529 108 2563
rect 26 2495 108 2529
rect 26 2461 50 2495
rect 84 2461 108 2495
rect 26 2427 108 2461
rect 26 2393 50 2427
rect 84 2393 108 2427
rect 26 2359 108 2393
rect 26 2325 50 2359
rect 84 2325 108 2359
rect 26 2291 108 2325
rect 26 2257 50 2291
rect 84 2257 108 2291
rect 26 2223 108 2257
rect 26 2189 50 2223
rect 84 2189 108 2223
rect 26 2155 108 2189
rect 26 2121 50 2155
rect 84 2121 108 2155
rect 26 2087 108 2121
rect 26 2053 50 2087
rect 84 2053 108 2087
rect 26 2019 108 2053
rect 26 1985 50 2019
rect 84 1985 108 2019
rect 26 1951 108 1985
rect 26 1917 50 1951
rect 84 1917 108 1951
rect 26 1883 108 1917
rect 26 1849 50 1883
rect 84 1849 108 1883
rect 26 1815 108 1849
rect 26 1781 50 1815
rect 84 1781 108 1815
rect 26 1747 108 1781
rect 26 1713 50 1747
rect 84 1713 108 1747
rect 26 1679 108 1713
rect 26 1645 50 1679
rect 84 1645 108 1679
rect 26 1611 108 1645
rect 26 1577 50 1611
rect 84 1577 108 1611
rect 26 1543 108 1577
rect 26 1509 50 1543
rect 84 1509 108 1543
rect 26 1475 108 1509
rect 26 1441 50 1475
rect 84 1441 108 1475
rect 26 1407 108 1441
rect 26 1373 50 1407
rect 84 1373 108 1407
rect 26 1339 108 1373
rect 26 1305 50 1339
rect 84 1305 108 1339
rect 26 1271 108 1305
rect 26 1237 50 1271
rect 84 1237 108 1271
rect 26 1203 108 1237
rect 26 1169 50 1203
rect 84 1169 108 1203
rect 26 1135 108 1169
rect 26 1101 50 1135
rect 84 1101 108 1135
rect 26 1067 108 1101
rect 26 1033 50 1067
rect 84 1033 108 1067
rect 26 999 108 1033
rect 26 965 50 999
rect 84 965 108 999
rect 26 931 108 965
rect 26 897 50 931
rect 84 897 108 931
rect 26 863 108 897
rect 26 829 50 863
rect 84 829 108 863
rect 26 795 108 829
rect 26 761 50 795
rect 84 761 108 795
rect 26 727 108 761
rect 26 693 50 727
rect 84 693 108 727
rect 26 659 108 693
rect 26 625 50 659
rect 84 625 108 659
rect 26 591 108 625
rect 26 557 50 591
rect 84 557 108 591
rect 26 523 108 557
rect 26 489 50 523
rect 84 489 108 523
rect 26 455 108 489
rect 26 421 50 455
rect 84 421 108 455
rect 26 387 108 421
rect 26 353 50 387
rect 84 353 108 387
rect 26 319 108 353
rect 26 285 50 319
rect 84 285 108 319
rect 26 251 108 285
rect 654 2714 1338 2738
rect 654 2680 678 2714
rect 712 2680 775 2714
rect 809 2680 843 2714
rect 877 2680 911 2714
rect 945 2680 979 2714
rect 1013 2680 1047 2714
rect 1081 2680 1115 2714
rect 1149 2680 1183 2714
rect 1217 2680 1280 2714
rect 1314 2680 1338 2714
rect 654 2656 1338 2680
rect 654 2631 736 2656
rect 654 2597 678 2631
rect 712 2597 736 2631
rect 654 2563 736 2597
rect 654 2529 678 2563
rect 712 2529 736 2563
rect 654 2495 736 2529
rect 1256 2631 1338 2656
rect 1256 2597 1280 2631
rect 1314 2597 1338 2631
rect 1256 2563 1338 2597
rect 1256 2529 1280 2563
rect 1314 2529 1338 2563
rect 654 2461 678 2495
rect 712 2461 736 2495
rect 654 2427 736 2461
rect 654 2393 678 2427
rect 712 2393 736 2427
rect 654 2359 736 2393
rect 654 2325 678 2359
rect 712 2325 736 2359
rect 654 2291 736 2325
rect 654 2257 678 2291
rect 712 2257 736 2291
rect 654 2223 736 2257
rect 654 2189 678 2223
rect 712 2189 736 2223
rect 654 2155 736 2189
rect 654 2121 678 2155
rect 712 2121 736 2155
rect 654 2087 736 2121
rect 654 2053 678 2087
rect 712 2053 736 2087
rect 654 2019 736 2053
rect 654 1985 678 2019
rect 712 1985 736 2019
rect 654 1951 736 1985
rect 654 1917 678 1951
rect 712 1917 736 1951
rect 654 1883 736 1917
rect 654 1849 678 1883
rect 712 1849 736 1883
rect 654 1815 736 1849
rect 654 1781 678 1815
rect 712 1781 736 1815
rect 654 1747 736 1781
rect 654 1713 678 1747
rect 712 1713 736 1747
rect 654 1679 736 1713
rect 654 1645 678 1679
rect 712 1645 736 1679
rect 654 1611 736 1645
rect 654 1577 678 1611
rect 712 1577 736 1611
rect 654 1543 736 1577
rect 654 1509 678 1543
rect 712 1509 736 1543
rect 654 1475 736 1509
rect 654 1441 678 1475
rect 712 1441 736 1475
rect 654 1407 736 1441
rect 654 1373 678 1407
rect 712 1373 736 1407
rect 654 1339 736 1373
rect 654 1305 678 1339
rect 712 1305 736 1339
rect 654 1271 736 1305
rect 654 1237 678 1271
rect 712 1237 736 1271
rect 654 1203 736 1237
rect 654 1169 678 1203
rect 712 1169 736 1203
rect 654 1135 736 1169
rect 654 1101 678 1135
rect 712 1101 736 1135
rect 654 1067 736 1101
rect 654 1033 678 1067
rect 712 1033 736 1067
rect 654 999 736 1033
rect 654 965 678 999
rect 712 965 736 999
rect 654 931 736 965
rect 654 897 678 931
rect 712 897 736 931
rect 654 863 736 897
rect 1256 2495 1338 2529
rect 1256 2461 1280 2495
rect 1314 2461 1338 2495
rect 1256 2427 1338 2461
rect 1256 2393 1280 2427
rect 1314 2393 1338 2427
rect 1256 2359 1338 2393
rect 1256 2325 1280 2359
rect 1314 2325 1338 2359
rect 1256 2291 1338 2325
rect 1256 2257 1280 2291
rect 1314 2257 1338 2291
rect 1256 2223 1338 2257
rect 1256 2189 1280 2223
rect 1314 2189 1338 2223
rect 1256 2155 1338 2189
rect 1256 2121 1280 2155
rect 1314 2121 1338 2155
rect 1256 2087 1338 2121
rect 1256 2053 1280 2087
rect 1314 2053 1338 2087
rect 1256 2019 1338 2053
rect 1256 1985 1280 2019
rect 1314 1985 1338 2019
rect 1256 1951 1338 1985
rect 1256 1917 1280 1951
rect 1314 1917 1338 1951
rect 1256 1883 1338 1917
rect 1256 1849 1280 1883
rect 1314 1849 1338 1883
rect 1256 1815 1338 1849
rect 1256 1781 1280 1815
rect 1314 1781 1338 1815
rect 1256 1747 1338 1781
rect 1256 1713 1280 1747
rect 1314 1713 1338 1747
rect 1256 1679 1338 1713
rect 1256 1645 1280 1679
rect 1314 1645 1338 1679
rect 1256 1611 1338 1645
rect 1256 1577 1280 1611
rect 1314 1577 1338 1611
rect 1256 1543 1338 1577
rect 1256 1509 1280 1543
rect 1314 1509 1338 1543
rect 1256 1475 1338 1509
rect 1256 1441 1280 1475
rect 1314 1441 1338 1475
rect 1256 1407 1338 1441
rect 1256 1373 1280 1407
rect 1314 1373 1338 1407
rect 1256 1339 1338 1373
rect 1256 1305 1280 1339
rect 1314 1305 1338 1339
rect 1256 1271 1338 1305
rect 1256 1237 1280 1271
rect 1314 1237 1338 1271
rect 1256 1203 1338 1237
rect 1256 1169 1280 1203
rect 1314 1169 1338 1203
rect 1256 1135 1338 1169
rect 1256 1101 1280 1135
rect 1314 1101 1338 1135
rect 1256 1067 1338 1101
rect 1256 1033 1280 1067
rect 1314 1033 1338 1067
rect 1256 999 1338 1033
rect 1256 965 1280 999
rect 1314 965 1338 999
rect 1256 931 1338 965
rect 1256 897 1280 931
rect 1314 897 1338 931
rect 654 829 678 863
rect 712 829 736 863
rect 654 795 736 829
rect 654 761 678 795
rect 712 761 736 795
rect 654 736 736 761
rect 1256 863 1338 897
rect 1256 829 1280 863
rect 1314 829 1338 863
rect 1256 795 1338 829
rect 1256 761 1280 795
rect 1314 761 1338 795
rect 1256 736 1338 761
rect 654 712 1338 736
rect 654 678 678 712
rect 712 678 775 712
rect 809 678 843 712
rect 877 678 911 712
rect 945 678 979 712
rect 1013 678 1047 712
rect 1081 678 1115 712
rect 1149 678 1183 712
rect 1217 678 1280 712
rect 1314 678 1338 712
rect 654 654 1338 678
rect 1884 3107 1966 3141
rect 1884 3073 1908 3107
rect 1942 3073 1966 3107
rect 1884 3039 1966 3073
rect 1884 3005 1908 3039
rect 1942 3005 1966 3039
rect 1884 2971 1966 3005
rect 1884 2937 1908 2971
rect 1942 2937 1966 2971
rect 1884 2903 1966 2937
rect 1884 2869 1908 2903
rect 1942 2869 1966 2903
rect 1884 2835 1966 2869
rect 1884 2801 1908 2835
rect 1942 2801 1966 2835
rect 1884 2767 1966 2801
rect 1884 2733 1908 2767
rect 1942 2733 1966 2767
rect 1884 2699 1966 2733
rect 1884 2665 1908 2699
rect 1942 2665 1966 2699
rect 1884 2631 1966 2665
rect 1884 2597 1908 2631
rect 1942 2597 1966 2631
rect 1884 2563 1966 2597
rect 1884 2529 1908 2563
rect 1942 2529 1966 2563
rect 1884 2495 1966 2529
rect 1884 2461 1908 2495
rect 1942 2461 1966 2495
rect 1884 2427 1966 2461
rect 1884 2393 1908 2427
rect 1942 2393 1966 2427
rect 1884 2359 1966 2393
rect 1884 2325 1908 2359
rect 1942 2325 1966 2359
rect 1884 2291 1966 2325
rect 1884 2257 1908 2291
rect 1942 2257 1966 2291
rect 1884 2223 1966 2257
rect 1884 2189 1908 2223
rect 1942 2189 1966 2223
rect 1884 2155 1966 2189
rect 1884 2121 1908 2155
rect 1942 2121 1966 2155
rect 1884 2087 1966 2121
rect 1884 2053 1908 2087
rect 1942 2053 1966 2087
rect 1884 2019 1966 2053
rect 1884 1985 1908 2019
rect 1942 1985 1966 2019
rect 1884 1951 1966 1985
rect 1884 1917 1908 1951
rect 1942 1917 1966 1951
rect 1884 1883 1966 1917
rect 1884 1849 1908 1883
rect 1942 1849 1966 1883
rect 1884 1815 1966 1849
rect 1884 1781 1908 1815
rect 1942 1781 1966 1815
rect 1884 1747 1966 1781
rect 1884 1713 1908 1747
rect 1942 1713 1966 1747
rect 1884 1679 1966 1713
rect 1884 1645 1908 1679
rect 1942 1645 1966 1679
rect 1884 1611 1966 1645
rect 1884 1577 1908 1611
rect 1942 1577 1966 1611
rect 1884 1543 1966 1577
rect 1884 1509 1908 1543
rect 1942 1509 1966 1543
rect 1884 1475 1966 1509
rect 1884 1441 1908 1475
rect 1942 1441 1966 1475
rect 1884 1407 1966 1441
rect 1884 1373 1908 1407
rect 1942 1373 1966 1407
rect 1884 1339 1966 1373
rect 1884 1305 1908 1339
rect 1942 1305 1966 1339
rect 1884 1271 1966 1305
rect 1884 1237 1908 1271
rect 1942 1237 1966 1271
rect 1884 1203 1966 1237
rect 1884 1169 1908 1203
rect 1942 1169 1966 1203
rect 1884 1135 1966 1169
rect 1884 1101 1908 1135
rect 1942 1101 1966 1135
rect 1884 1067 1966 1101
rect 1884 1033 1908 1067
rect 1942 1033 1966 1067
rect 1884 999 1966 1033
rect 1884 965 1908 999
rect 1942 965 1966 999
rect 1884 931 1966 965
rect 1884 897 1908 931
rect 1942 897 1966 931
rect 1884 863 1966 897
rect 1884 829 1908 863
rect 1942 829 1966 863
rect 1884 795 1966 829
rect 1884 761 1908 795
rect 1942 761 1966 795
rect 1884 727 1966 761
rect 1884 693 1908 727
rect 1942 693 1966 727
rect 1884 659 1966 693
rect 1884 625 1908 659
rect 1942 625 1966 659
rect 1884 591 1966 625
rect 1884 557 1908 591
rect 1942 557 1966 591
rect 1884 523 1966 557
rect 1884 489 1908 523
rect 1942 489 1966 523
rect 1884 455 1966 489
rect 1884 421 1908 455
rect 1942 421 1966 455
rect 1884 387 1966 421
rect 1884 353 1908 387
rect 1942 353 1966 387
rect 1884 319 1966 353
rect 1884 285 1908 319
rect 1942 285 1966 319
rect 26 217 50 251
rect 84 217 108 251
rect 26 183 108 217
rect 26 149 50 183
rect 84 149 108 183
rect 26 108 108 149
rect 1884 251 1966 285
rect 1884 217 1908 251
rect 1942 217 1966 251
rect 1884 183 1966 217
rect 1884 149 1908 183
rect 1942 149 1966 183
rect 1884 108 1966 149
rect 26 84 1966 108
rect 26 50 50 84
rect 84 50 129 84
rect 163 50 197 84
rect 231 50 265 84
rect 299 50 333 84
rect 367 50 401 84
rect 435 50 469 84
rect 503 50 537 84
rect 571 50 605 84
rect 639 50 673 84
rect 707 50 741 84
rect 775 50 809 84
rect 843 50 877 84
rect 911 50 945 84
rect 979 50 1013 84
rect 1047 50 1081 84
rect 1115 50 1149 84
rect 1183 50 1217 84
rect 1251 50 1285 84
rect 1319 50 1353 84
rect 1387 50 1421 84
rect 1455 50 1489 84
rect 1523 50 1557 84
rect 1591 50 1625 84
rect 1659 50 1693 84
rect 1727 50 1761 84
rect 1795 50 1829 84
rect 1863 50 1908 84
rect 1942 50 1966 84
rect 26 26 1966 50
<< nsubdiff >>
rect 252 3116 1740 3140
rect 252 3082 276 3116
rect 310 3082 367 3116
rect 401 3082 435 3116
rect 469 3082 503 3116
rect 537 3082 571 3116
rect 605 3082 639 3116
rect 673 3082 707 3116
rect 741 3082 775 3116
rect 809 3082 843 3116
rect 877 3082 911 3116
rect 945 3082 979 3116
rect 1013 3082 1047 3116
rect 1081 3082 1115 3116
rect 1149 3082 1183 3116
rect 1217 3082 1251 3116
rect 1285 3082 1319 3116
rect 1353 3082 1387 3116
rect 1421 3082 1455 3116
rect 1489 3082 1523 3116
rect 1557 3082 1591 3116
rect 1625 3082 1682 3116
rect 1716 3082 1740 3116
rect 252 3058 1740 3082
rect 252 3039 334 3058
rect 252 3005 276 3039
rect 310 3005 334 3039
rect 252 2971 334 3005
rect 252 2937 276 2971
rect 310 2937 334 2971
rect 252 2903 334 2937
rect 252 2869 276 2903
rect 310 2869 334 2903
rect 252 2835 334 2869
rect 252 2801 276 2835
rect 310 2801 334 2835
rect 252 2767 334 2801
rect 252 2733 276 2767
rect 310 2733 334 2767
rect 1658 3039 1740 3058
rect 1658 3005 1682 3039
rect 1716 3005 1740 3039
rect 1658 2971 1740 3005
rect 1658 2937 1682 2971
rect 1716 2937 1740 2971
rect 1658 2903 1740 2937
rect 1658 2869 1682 2903
rect 1716 2869 1740 2903
rect 1658 2835 1740 2869
rect 1658 2801 1682 2835
rect 1716 2801 1740 2835
rect 1658 2767 1740 2801
rect 252 2699 334 2733
rect 252 2665 276 2699
rect 310 2665 334 2699
rect 252 2631 334 2665
rect 252 2597 276 2631
rect 310 2597 334 2631
rect 252 2563 334 2597
rect 252 2529 276 2563
rect 310 2529 334 2563
rect 252 2495 334 2529
rect 252 2461 276 2495
rect 310 2461 334 2495
rect 252 2427 334 2461
rect 252 2393 276 2427
rect 310 2393 334 2427
rect 252 2359 334 2393
rect 252 2325 276 2359
rect 310 2325 334 2359
rect 252 2291 334 2325
rect 252 2257 276 2291
rect 310 2257 334 2291
rect 252 2223 334 2257
rect 252 2189 276 2223
rect 310 2189 334 2223
rect 252 2155 334 2189
rect 252 2121 276 2155
rect 310 2121 334 2155
rect 252 2087 334 2121
rect 252 2053 276 2087
rect 310 2053 334 2087
rect 252 2019 334 2053
rect 252 1985 276 2019
rect 310 1985 334 2019
rect 252 1951 334 1985
rect 252 1917 276 1951
rect 310 1917 334 1951
rect 252 1883 334 1917
rect 252 1849 276 1883
rect 310 1849 334 1883
rect 252 1815 334 1849
rect 252 1781 276 1815
rect 310 1781 334 1815
rect 252 1747 334 1781
rect 252 1713 276 1747
rect 310 1713 334 1747
rect 252 1679 334 1713
rect 252 1645 276 1679
rect 310 1645 334 1679
rect 252 1611 334 1645
rect 252 1577 276 1611
rect 310 1577 334 1611
rect 252 1543 334 1577
rect 252 1509 276 1543
rect 310 1509 334 1543
rect 252 1475 334 1509
rect 252 1441 276 1475
rect 310 1441 334 1475
rect 252 1407 334 1441
rect 252 1373 276 1407
rect 310 1373 334 1407
rect 252 1339 334 1373
rect 252 1305 276 1339
rect 310 1305 334 1339
rect 252 1271 334 1305
rect 252 1237 276 1271
rect 310 1237 334 1271
rect 252 1203 334 1237
rect 252 1169 276 1203
rect 310 1169 334 1203
rect 252 1135 334 1169
rect 252 1101 276 1135
rect 310 1101 334 1135
rect 252 1067 334 1101
rect 252 1033 276 1067
rect 310 1033 334 1067
rect 252 999 334 1033
rect 252 965 276 999
rect 310 965 334 999
rect 252 931 334 965
rect 252 897 276 931
rect 310 897 334 931
rect 252 863 334 897
rect 252 829 276 863
rect 310 829 334 863
rect 252 795 334 829
rect 252 761 276 795
rect 310 761 334 795
rect 252 727 334 761
rect 252 693 276 727
rect 310 693 334 727
rect 252 659 334 693
rect 252 625 276 659
rect 310 625 334 659
rect 1658 2733 1682 2767
rect 1716 2733 1740 2767
rect 1658 2699 1740 2733
rect 1658 2665 1682 2699
rect 1716 2665 1740 2699
rect 1658 2631 1740 2665
rect 1658 2597 1682 2631
rect 1716 2597 1740 2631
rect 1658 2563 1740 2597
rect 1658 2529 1682 2563
rect 1716 2529 1740 2563
rect 1658 2495 1740 2529
rect 1658 2461 1682 2495
rect 1716 2461 1740 2495
rect 1658 2427 1740 2461
rect 1658 2393 1682 2427
rect 1716 2393 1740 2427
rect 1658 2359 1740 2393
rect 1658 2325 1682 2359
rect 1716 2325 1740 2359
rect 1658 2291 1740 2325
rect 1658 2257 1682 2291
rect 1716 2257 1740 2291
rect 1658 2223 1740 2257
rect 1658 2189 1682 2223
rect 1716 2189 1740 2223
rect 1658 2155 1740 2189
rect 1658 2121 1682 2155
rect 1716 2121 1740 2155
rect 1658 2087 1740 2121
rect 1658 2053 1682 2087
rect 1716 2053 1740 2087
rect 1658 2019 1740 2053
rect 1658 1985 1682 2019
rect 1716 1985 1740 2019
rect 1658 1951 1740 1985
rect 1658 1917 1682 1951
rect 1716 1917 1740 1951
rect 1658 1883 1740 1917
rect 1658 1849 1682 1883
rect 1716 1849 1740 1883
rect 1658 1815 1740 1849
rect 1658 1781 1682 1815
rect 1716 1781 1740 1815
rect 1658 1747 1740 1781
rect 1658 1713 1682 1747
rect 1716 1713 1740 1747
rect 1658 1679 1740 1713
rect 1658 1645 1682 1679
rect 1716 1645 1740 1679
rect 1658 1611 1740 1645
rect 1658 1577 1682 1611
rect 1716 1577 1740 1611
rect 1658 1543 1740 1577
rect 1658 1509 1682 1543
rect 1716 1509 1740 1543
rect 1658 1475 1740 1509
rect 1658 1441 1682 1475
rect 1716 1441 1740 1475
rect 1658 1407 1740 1441
rect 1658 1373 1682 1407
rect 1716 1373 1740 1407
rect 1658 1339 1740 1373
rect 1658 1305 1682 1339
rect 1716 1305 1740 1339
rect 1658 1271 1740 1305
rect 1658 1237 1682 1271
rect 1716 1237 1740 1271
rect 1658 1203 1740 1237
rect 1658 1169 1682 1203
rect 1716 1169 1740 1203
rect 1658 1135 1740 1169
rect 1658 1101 1682 1135
rect 1716 1101 1740 1135
rect 1658 1067 1740 1101
rect 1658 1033 1682 1067
rect 1716 1033 1740 1067
rect 1658 999 1740 1033
rect 1658 965 1682 999
rect 1716 965 1740 999
rect 1658 931 1740 965
rect 1658 897 1682 931
rect 1716 897 1740 931
rect 1658 863 1740 897
rect 1658 829 1682 863
rect 1716 829 1740 863
rect 1658 795 1740 829
rect 1658 761 1682 795
rect 1716 761 1740 795
rect 1658 727 1740 761
rect 1658 693 1682 727
rect 1716 693 1740 727
rect 1658 659 1740 693
rect 252 591 334 625
rect 252 557 276 591
rect 310 557 334 591
rect 252 523 334 557
rect 252 489 276 523
rect 310 489 334 523
rect 252 455 334 489
rect 252 421 276 455
rect 310 421 334 455
rect 252 387 334 421
rect 252 353 276 387
rect 310 353 334 387
rect 252 334 334 353
rect 1658 625 1682 659
rect 1716 625 1740 659
rect 1658 591 1740 625
rect 1658 557 1682 591
rect 1716 557 1740 591
rect 1658 523 1740 557
rect 1658 489 1682 523
rect 1716 489 1740 523
rect 1658 455 1740 489
rect 1658 421 1682 455
rect 1716 421 1740 455
rect 1658 387 1740 421
rect 1658 353 1682 387
rect 1716 353 1740 387
rect 1658 334 1740 353
rect 252 310 1740 334
rect 252 276 276 310
rect 310 276 367 310
rect 401 276 435 310
rect 469 276 503 310
rect 537 276 571 310
rect 605 276 639 310
rect 673 276 707 310
rect 741 276 775 310
rect 809 276 843 310
rect 877 276 911 310
rect 945 276 979 310
rect 1013 276 1047 310
rect 1081 276 1115 310
rect 1149 276 1183 310
rect 1217 276 1251 310
rect 1285 276 1319 310
rect 1353 276 1387 310
rect 1421 276 1455 310
rect 1489 276 1523 310
rect 1557 276 1591 310
rect 1625 276 1682 310
rect 1716 276 1740 310
rect 252 252 1740 276
<< psubdiffcont >>
rect 50 3308 84 3342
rect 129 3308 163 3342
rect 197 3308 231 3342
rect 265 3308 299 3342
rect 333 3308 367 3342
rect 401 3308 435 3342
rect 469 3308 503 3342
rect 537 3308 571 3342
rect 605 3308 639 3342
rect 673 3308 707 3342
rect 741 3308 775 3342
rect 809 3308 843 3342
rect 877 3308 911 3342
rect 945 3308 979 3342
rect 1013 3308 1047 3342
rect 1081 3308 1115 3342
rect 1149 3308 1183 3342
rect 1217 3308 1251 3342
rect 1285 3308 1319 3342
rect 1353 3308 1387 3342
rect 1421 3308 1455 3342
rect 1489 3308 1523 3342
rect 1557 3308 1591 3342
rect 1625 3308 1659 3342
rect 1693 3308 1727 3342
rect 1761 3308 1795 3342
rect 1829 3308 1863 3342
rect 1908 3308 1942 3342
rect 50 3209 84 3243
rect 50 3141 84 3175
rect 1908 3209 1942 3243
rect 1908 3141 1942 3175
rect 50 3073 84 3107
rect 50 3005 84 3039
rect 50 2937 84 2971
rect 50 2869 84 2903
rect 50 2801 84 2835
rect 50 2733 84 2767
rect 50 2665 84 2699
rect 50 2597 84 2631
rect 50 2529 84 2563
rect 50 2461 84 2495
rect 50 2393 84 2427
rect 50 2325 84 2359
rect 50 2257 84 2291
rect 50 2189 84 2223
rect 50 2121 84 2155
rect 50 2053 84 2087
rect 50 1985 84 2019
rect 50 1917 84 1951
rect 50 1849 84 1883
rect 50 1781 84 1815
rect 50 1713 84 1747
rect 50 1645 84 1679
rect 50 1577 84 1611
rect 50 1509 84 1543
rect 50 1441 84 1475
rect 50 1373 84 1407
rect 50 1305 84 1339
rect 50 1237 84 1271
rect 50 1169 84 1203
rect 50 1101 84 1135
rect 50 1033 84 1067
rect 50 965 84 999
rect 50 897 84 931
rect 50 829 84 863
rect 50 761 84 795
rect 50 693 84 727
rect 50 625 84 659
rect 50 557 84 591
rect 50 489 84 523
rect 50 421 84 455
rect 50 353 84 387
rect 50 285 84 319
rect 678 2680 712 2714
rect 775 2680 809 2714
rect 843 2680 877 2714
rect 911 2680 945 2714
rect 979 2680 1013 2714
rect 1047 2680 1081 2714
rect 1115 2680 1149 2714
rect 1183 2680 1217 2714
rect 1280 2680 1314 2714
rect 678 2597 712 2631
rect 678 2529 712 2563
rect 1280 2597 1314 2631
rect 1280 2529 1314 2563
rect 678 2461 712 2495
rect 678 2393 712 2427
rect 678 2325 712 2359
rect 678 2257 712 2291
rect 678 2189 712 2223
rect 678 2121 712 2155
rect 678 2053 712 2087
rect 678 1985 712 2019
rect 678 1917 712 1951
rect 678 1849 712 1883
rect 678 1781 712 1815
rect 678 1713 712 1747
rect 678 1645 712 1679
rect 678 1577 712 1611
rect 678 1509 712 1543
rect 678 1441 712 1475
rect 678 1373 712 1407
rect 678 1305 712 1339
rect 678 1237 712 1271
rect 678 1169 712 1203
rect 678 1101 712 1135
rect 678 1033 712 1067
rect 678 965 712 999
rect 678 897 712 931
rect 1280 2461 1314 2495
rect 1280 2393 1314 2427
rect 1280 2325 1314 2359
rect 1280 2257 1314 2291
rect 1280 2189 1314 2223
rect 1280 2121 1314 2155
rect 1280 2053 1314 2087
rect 1280 1985 1314 2019
rect 1280 1917 1314 1951
rect 1280 1849 1314 1883
rect 1280 1781 1314 1815
rect 1280 1713 1314 1747
rect 1280 1645 1314 1679
rect 1280 1577 1314 1611
rect 1280 1509 1314 1543
rect 1280 1441 1314 1475
rect 1280 1373 1314 1407
rect 1280 1305 1314 1339
rect 1280 1237 1314 1271
rect 1280 1169 1314 1203
rect 1280 1101 1314 1135
rect 1280 1033 1314 1067
rect 1280 965 1314 999
rect 1280 897 1314 931
rect 678 829 712 863
rect 678 761 712 795
rect 1280 829 1314 863
rect 1280 761 1314 795
rect 678 678 712 712
rect 775 678 809 712
rect 843 678 877 712
rect 911 678 945 712
rect 979 678 1013 712
rect 1047 678 1081 712
rect 1115 678 1149 712
rect 1183 678 1217 712
rect 1280 678 1314 712
rect 1908 3073 1942 3107
rect 1908 3005 1942 3039
rect 1908 2937 1942 2971
rect 1908 2869 1942 2903
rect 1908 2801 1942 2835
rect 1908 2733 1942 2767
rect 1908 2665 1942 2699
rect 1908 2597 1942 2631
rect 1908 2529 1942 2563
rect 1908 2461 1942 2495
rect 1908 2393 1942 2427
rect 1908 2325 1942 2359
rect 1908 2257 1942 2291
rect 1908 2189 1942 2223
rect 1908 2121 1942 2155
rect 1908 2053 1942 2087
rect 1908 1985 1942 2019
rect 1908 1917 1942 1951
rect 1908 1849 1942 1883
rect 1908 1781 1942 1815
rect 1908 1713 1942 1747
rect 1908 1645 1942 1679
rect 1908 1577 1942 1611
rect 1908 1509 1942 1543
rect 1908 1441 1942 1475
rect 1908 1373 1942 1407
rect 1908 1305 1942 1339
rect 1908 1237 1942 1271
rect 1908 1169 1942 1203
rect 1908 1101 1942 1135
rect 1908 1033 1942 1067
rect 1908 965 1942 999
rect 1908 897 1942 931
rect 1908 829 1942 863
rect 1908 761 1942 795
rect 1908 693 1942 727
rect 1908 625 1942 659
rect 1908 557 1942 591
rect 1908 489 1942 523
rect 1908 421 1942 455
rect 1908 353 1942 387
rect 1908 285 1942 319
rect 50 217 84 251
rect 50 149 84 183
rect 1908 217 1942 251
rect 1908 149 1942 183
rect 50 50 84 84
rect 129 50 163 84
rect 197 50 231 84
rect 265 50 299 84
rect 333 50 367 84
rect 401 50 435 84
rect 469 50 503 84
rect 537 50 571 84
rect 605 50 639 84
rect 673 50 707 84
rect 741 50 775 84
rect 809 50 843 84
rect 877 50 911 84
rect 945 50 979 84
rect 1013 50 1047 84
rect 1081 50 1115 84
rect 1149 50 1183 84
rect 1217 50 1251 84
rect 1285 50 1319 84
rect 1353 50 1387 84
rect 1421 50 1455 84
rect 1489 50 1523 84
rect 1557 50 1591 84
rect 1625 50 1659 84
rect 1693 50 1727 84
rect 1761 50 1795 84
rect 1829 50 1863 84
rect 1908 50 1942 84
<< nsubdiffcont >>
rect 276 3082 310 3116
rect 367 3082 401 3116
rect 435 3082 469 3116
rect 503 3082 537 3116
rect 571 3082 605 3116
rect 639 3082 673 3116
rect 707 3082 741 3116
rect 775 3082 809 3116
rect 843 3082 877 3116
rect 911 3082 945 3116
rect 979 3082 1013 3116
rect 1047 3082 1081 3116
rect 1115 3082 1149 3116
rect 1183 3082 1217 3116
rect 1251 3082 1285 3116
rect 1319 3082 1353 3116
rect 1387 3082 1421 3116
rect 1455 3082 1489 3116
rect 1523 3082 1557 3116
rect 1591 3082 1625 3116
rect 1682 3082 1716 3116
rect 276 3005 310 3039
rect 276 2937 310 2971
rect 276 2869 310 2903
rect 276 2801 310 2835
rect 276 2733 310 2767
rect 1682 3005 1716 3039
rect 1682 2937 1716 2971
rect 1682 2869 1716 2903
rect 1682 2801 1716 2835
rect 276 2665 310 2699
rect 276 2597 310 2631
rect 276 2529 310 2563
rect 276 2461 310 2495
rect 276 2393 310 2427
rect 276 2325 310 2359
rect 276 2257 310 2291
rect 276 2189 310 2223
rect 276 2121 310 2155
rect 276 2053 310 2087
rect 276 1985 310 2019
rect 276 1917 310 1951
rect 276 1849 310 1883
rect 276 1781 310 1815
rect 276 1713 310 1747
rect 276 1645 310 1679
rect 276 1577 310 1611
rect 276 1509 310 1543
rect 276 1441 310 1475
rect 276 1373 310 1407
rect 276 1305 310 1339
rect 276 1237 310 1271
rect 276 1169 310 1203
rect 276 1101 310 1135
rect 276 1033 310 1067
rect 276 965 310 999
rect 276 897 310 931
rect 276 829 310 863
rect 276 761 310 795
rect 276 693 310 727
rect 276 625 310 659
rect 1682 2733 1716 2767
rect 1682 2665 1716 2699
rect 1682 2597 1716 2631
rect 1682 2529 1716 2563
rect 1682 2461 1716 2495
rect 1682 2393 1716 2427
rect 1682 2325 1716 2359
rect 1682 2257 1716 2291
rect 1682 2189 1716 2223
rect 1682 2121 1716 2155
rect 1682 2053 1716 2087
rect 1682 1985 1716 2019
rect 1682 1917 1716 1951
rect 1682 1849 1716 1883
rect 1682 1781 1716 1815
rect 1682 1713 1716 1747
rect 1682 1645 1716 1679
rect 1682 1577 1716 1611
rect 1682 1509 1716 1543
rect 1682 1441 1716 1475
rect 1682 1373 1716 1407
rect 1682 1305 1716 1339
rect 1682 1237 1716 1271
rect 1682 1169 1716 1203
rect 1682 1101 1716 1135
rect 1682 1033 1716 1067
rect 1682 965 1716 999
rect 1682 897 1716 931
rect 1682 829 1716 863
rect 1682 761 1716 795
rect 1682 693 1716 727
rect 276 557 310 591
rect 276 489 310 523
rect 276 421 310 455
rect 276 353 310 387
rect 1682 625 1716 659
rect 1682 557 1716 591
rect 1682 489 1716 523
rect 1682 421 1716 455
rect 1682 353 1716 387
rect 276 276 310 310
rect 367 276 401 310
rect 435 276 469 310
rect 503 276 537 310
rect 571 276 605 310
rect 639 276 673 310
rect 707 276 741 310
rect 775 276 809 310
rect 843 276 877 310
rect 911 276 945 310
rect 979 276 1013 310
rect 1047 276 1081 310
rect 1115 276 1149 310
rect 1183 276 1217 310
rect 1251 276 1285 310
rect 1319 276 1353 310
rect 1387 276 1421 310
rect 1455 276 1489 310
rect 1523 276 1557 310
rect 1591 276 1625 310
rect 1682 276 1716 310
<< locali >>
rect 34 3342 1958 3358
rect 34 3308 50 3342
rect 84 3308 129 3342
rect 185 3308 197 3342
rect 257 3308 265 3342
rect 329 3308 333 3342
rect 435 3308 439 3342
rect 503 3308 511 3342
rect 571 3308 583 3342
rect 639 3308 655 3342
rect 707 3308 727 3342
rect 775 3308 799 3342
rect 843 3308 871 3342
rect 911 3308 943 3342
rect 979 3308 1013 3342
rect 1049 3308 1081 3342
rect 1121 3308 1149 3342
rect 1193 3308 1217 3342
rect 1265 3308 1285 3342
rect 1337 3308 1353 3342
rect 1409 3308 1421 3342
rect 1481 3308 1489 3342
rect 1553 3308 1557 3342
rect 1659 3308 1663 3342
rect 1727 3308 1735 3342
rect 1795 3308 1807 3342
rect 1863 3308 1908 3342
rect 1942 3308 1958 3342
rect 34 3292 1958 3308
rect 34 3261 100 3292
rect 34 3209 50 3261
rect 84 3209 100 3261
rect 34 3189 100 3209
rect 34 3141 50 3189
rect 84 3141 100 3189
rect 34 3117 100 3141
rect 1892 3261 1958 3292
rect 1892 3209 1908 3261
rect 1942 3209 1958 3261
rect 1892 3189 1958 3209
rect 1892 3141 1908 3189
rect 1942 3141 1958 3189
rect 34 3073 50 3117
rect 84 3073 100 3117
rect 34 3045 100 3073
rect 34 3005 50 3045
rect 84 3005 100 3045
rect 34 2973 100 3005
rect 34 2937 50 2973
rect 84 2937 100 2973
rect 34 2903 100 2937
rect 34 2867 50 2903
rect 84 2867 100 2903
rect 34 2835 100 2867
rect 34 2795 50 2835
rect 84 2795 100 2835
rect 34 2767 100 2795
rect 34 2723 50 2767
rect 84 2723 100 2767
rect 34 2699 100 2723
rect 34 2651 50 2699
rect 84 2651 100 2699
rect 34 2631 100 2651
rect 34 2579 50 2631
rect 84 2579 100 2631
rect 34 2563 100 2579
rect 34 2507 50 2563
rect 84 2507 100 2563
rect 34 2495 100 2507
rect 34 2435 50 2495
rect 84 2435 100 2495
rect 34 2427 100 2435
rect 34 2363 50 2427
rect 84 2363 100 2427
rect 34 2359 100 2363
rect 34 2257 50 2359
rect 84 2257 100 2359
rect 34 2253 100 2257
rect 34 2189 50 2253
rect 84 2189 100 2253
rect 34 2181 100 2189
rect 34 2121 50 2181
rect 84 2121 100 2181
rect 34 2109 100 2121
rect 34 2053 50 2109
rect 84 2053 100 2109
rect 34 2037 100 2053
rect 34 1985 50 2037
rect 84 1985 100 2037
rect 34 1965 100 1985
rect 34 1917 50 1965
rect 84 1917 100 1965
rect 34 1893 100 1917
rect 34 1849 50 1893
rect 84 1849 100 1893
rect 34 1821 100 1849
rect 34 1781 50 1821
rect 84 1781 100 1821
rect 34 1749 100 1781
rect 34 1713 50 1749
rect 84 1713 100 1749
rect 34 1679 100 1713
rect 34 1643 50 1679
rect 84 1643 100 1679
rect 34 1611 100 1643
rect 34 1571 50 1611
rect 84 1571 100 1611
rect 34 1543 100 1571
rect 34 1499 50 1543
rect 84 1499 100 1543
rect 34 1475 100 1499
rect 34 1427 50 1475
rect 84 1427 100 1475
rect 34 1407 100 1427
rect 34 1355 50 1407
rect 84 1355 100 1407
rect 34 1339 100 1355
rect 34 1283 50 1339
rect 84 1283 100 1339
rect 34 1271 100 1283
rect 34 1211 50 1271
rect 84 1211 100 1271
rect 34 1203 100 1211
rect 34 1139 50 1203
rect 84 1139 100 1203
rect 34 1135 100 1139
rect 34 1033 50 1135
rect 84 1033 100 1135
rect 34 1029 100 1033
rect 34 965 50 1029
rect 84 965 100 1029
rect 34 957 100 965
rect 34 897 50 957
rect 84 897 100 957
rect 34 885 100 897
rect 34 829 50 885
rect 84 829 100 885
rect 34 813 100 829
rect 34 761 50 813
rect 84 761 100 813
rect 34 741 100 761
rect 34 693 50 741
rect 84 693 100 741
rect 34 669 100 693
rect 34 625 50 669
rect 84 625 100 669
rect 34 597 100 625
rect 34 557 50 597
rect 84 557 100 597
rect 34 525 100 557
rect 34 489 50 525
rect 84 489 100 525
rect 34 455 100 489
rect 34 419 50 455
rect 84 419 100 455
rect 34 387 100 419
rect 34 347 50 387
rect 84 347 100 387
rect 34 319 100 347
rect 34 275 50 319
rect 84 275 100 319
rect 34 251 100 275
rect 260 3116 1732 3132
rect 260 3082 276 3116
rect 310 3082 367 3116
rect 401 3082 435 3116
rect 473 3082 503 3116
rect 545 3082 571 3116
rect 617 3082 639 3116
rect 689 3082 707 3116
rect 761 3082 775 3116
rect 833 3082 843 3116
rect 905 3082 911 3116
rect 977 3082 979 3116
rect 1013 3082 1015 3116
rect 1081 3082 1087 3116
rect 1149 3082 1159 3116
rect 1217 3082 1231 3116
rect 1285 3082 1303 3116
rect 1353 3082 1375 3116
rect 1421 3082 1447 3116
rect 1489 3082 1519 3116
rect 1557 3082 1591 3116
rect 1625 3082 1682 3116
rect 1716 3082 1732 3116
rect 260 3066 1732 3082
rect 260 3039 326 3066
rect 260 2975 276 3039
rect 310 2975 326 3039
rect 260 2971 326 2975
rect 260 2869 276 2971
rect 310 2869 326 2971
rect 260 2865 326 2869
rect 260 2801 276 2865
rect 310 2801 326 2865
rect 260 2793 326 2801
rect 260 2733 276 2793
rect 310 2733 326 2793
rect 260 2721 326 2733
rect 1666 3039 1732 3066
rect 1666 2975 1682 3039
rect 1716 2975 1732 3039
rect 1666 2971 1732 2975
rect 1666 2869 1682 2971
rect 1716 2869 1732 2971
rect 1666 2865 1732 2869
rect 1666 2801 1682 2865
rect 1716 2801 1732 2865
rect 1666 2793 1732 2801
rect 1666 2733 1682 2793
rect 1716 2733 1732 2793
rect 260 2665 276 2721
rect 310 2665 326 2721
rect 260 2649 326 2665
rect 260 2597 276 2649
rect 310 2597 326 2649
rect 260 2577 326 2597
rect 260 2529 276 2577
rect 310 2529 326 2577
rect 260 2505 326 2529
rect 260 2461 276 2505
rect 310 2461 326 2505
rect 260 2433 326 2461
rect 260 2393 276 2433
rect 310 2393 326 2433
rect 260 2361 326 2393
rect 260 2325 276 2361
rect 310 2325 326 2361
rect 260 2291 326 2325
rect 260 2255 276 2291
rect 310 2255 326 2291
rect 260 2223 326 2255
rect 260 2183 276 2223
rect 310 2183 326 2223
rect 260 2155 326 2183
rect 260 2111 276 2155
rect 310 2111 326 2155
rect 260 2087 326 2111
rect 260 2039 276 2087
rect 310 2039 326 2087
rect 260 2019 326 2039
rect 260 1967 276 2019
rect 310 1967 326 2019
rect 260 1951 326 1967
rect 260 1895 276 1951
rect 310 1895 326 1951
rect 260 1883 326 1895
rect 260 1823 276 1883
rect 310 1823 326 1883
rect 260 1815 326 1823
rect 260 1751 276 1815
rect 310 1751 326 1815
rect 260 1747 326 1751
rect 260 1645 276 1747
rect 310 1645 326 1747
rect 260 1641 326 1645
rect 260 1577 276 1641
rect 310 1577 326 1641
rect 260 1569 326 1577
rect 260 1509 276 1569
rect 310 1509 326 1569
rect 260 1497 326 1509
rect 260 1441 276 1497
rect 310 1441 326 1497
rect 260 1425 326 1441
rect 260 1373 276 1425
rect 310 1373 326 1425
rect 260 1353 326 1373
rect 260 1305 276 1353
rect 310 1305 326 1353
rect 260 1281 326 1305
rect 260 1237 276 1281
rect 310 1237 326 1281
rect 260 1209 326 1237
rect 260 1169 276 1209
rect 310 1169 326 1209
rect 260 1137 326 1169
rect 260 1101 276 1137
rect 310 1101 326 1137
rect 260 1067 326 1101
rect 260 1031 276 1067
rect 310 1031 326 1067
rect 260 999 326 1031
rect 260 959 276 999
rect 310 959 326 999
rect 260 931 326 959
rect 260 887 276 931
rect 310 887 326 931
rect 260 863 326 887
rect 260 815 276 863
rect 310 815 326 863
rect 260 795 326 815
rect 260 743 276 795
rect 310 743 326 795
rect 260 727 326 743
rect 260 671 276 727
rect 310 671 326 727
rect 260 659 326 671
rect 662 2714 1330 2730
rect 662 2680 678 2714
rect 712 2680 763 2714
rect 809 2680 835 2714
rect 877 2680 907 2714
rect 945 2680 979 2714
rect 1013 2680 1047 2714
rect 1085 2680 1115 2714
rect 1157 2680 1183 2714
rect 1229 2680 1280 2714
rect 1314 2680 1330 2714
rect 662 2664 1330 2680
rect 662 2631 728 2664
rect 662 2579 678 2631
rect 712 2579 728 2631
rect 662 2563 728 2579
rect 662 2507 678 2563
rect 712 2507 728 2563
rect 662 2495 728 2507
rect 1264 2631 1330 2664
rect 1264 2579 1280 2631
rect 1314 2579 1330 2631
rect 1264 2563 1330 2579
rect 1264 2507 1280 2563
rect 1314 2507 1330 2563
rect 662 2435 678 2495
rect 712 2435 728 2495
rect 662 2427 728 2435
rect 662 2363 678 2427
rect 712 2363 728 2427
rect 662 2359 728 2363
rect 662 2257 678 2359
rect 712 2257 728 2359
rect 662 2253 728 2257
rect 662 2189 678 2253
rect 712 2189 728 2253
rect 662 2181 728 2189
rect 662 2121 678 2181
rect 712 2121 728 2181
rect 662 2109 728 2121
rect 662 2053 678 2109
rect 712 2053 728 2109
rect 662 2037 728 2053
rect 662 1985 678 2037
rect 712 1985 728 2037
rect 662 1965 728 1985
rect 662 1917 678 1965
rect 712 1917 728 1965
rect 662 1893 728 1917
rect 662 1849 678 1893
rect 712 1849 728 1893
rect 662 1821 728 1849
rect 662 1781 678 1821
rect 712 1781 728 1821
rect 662 1749 728 1781
rect 662 1713 678 1749
rect 712 1713 728 1749
rect 662 1679 728 1713
rect 662 1643 678 1679
rect 712 1643 728 1679
rect 662 1611 728 1643
rect 662 1571 678 1611
rect 712 1571 728 1611
rect 662 1543 728 1571
rect 662 1499 678 1543
rect 712 1499 728 1543
rect 662 1475 728 1499
rect 662 1427 678 1475
rect 712 1427 728 1475
rect 662 1407 728 1427
rect 662 1355 678 1407
rect 712 1355 728 1407
rect 662 1339 728 1355
rect 662 1283 678 1339
rect 712 1283 728 1339
rect 662 1271 728 1283
rect 662 1211 678 1271
rect 712 1211 728 1271
rect 662 1203 728 1211
rect 662 1139 678 1203
rect 712 1139 728 1203
rect 662 1135 728 1139
rect 662 1033 678 1135
rect 712 1033 728 1135
rect 662 1029 728 1033
rect 662 965 678 1029
rect 712 965 728 1029
rect 662 957 728 965
rect 662 897 678 957
rect 712 897 728 957
rect 662 885 728 897
rect 895 2469 1097 2497
rect 895 923 907 2469
rect 1085 923 1097 2469
rect 895 895 1097 923
rect 1264 2495 1330 2507
rect 1264 2435 1280 2495
rect 1314 2435 1330 2495
rect 1264 2427 1330 2435
rect 1264 2363 1280 2427
rect 1314 2363 1330 2427
rect 1264 2359 1330 2363
rect 1264 2257 1280 2359
rect 1314 2257 1330 2359
rect 1264 2253 1330 2257
rect 1264 2189 1280 2253
rect 1314 2189 1330 2253
rect 1264 2181 1330 2189
rect 1264 2121 1280 2181
rect 1314 2121 1330 2181
rect 1264 2109 1330 2121
rect 1264 2053 1280 2109
rect 1314 2053 1330 2109
rect 1264 2037 1330 2053
rect 1264 1985 1280 2037
rect 1314 1985 1330 2037
rect 1264 1965 1330 1985
rect 1264 1917 1280 1965
rect 1314 1917 1330 1965
rect 1264 1893 1330 1917
rect 1264 1849 1280 1893
rect 1314 1849 1330 1893
rect 1264 1821 1330 1849
rect 1264 1781 1280 1821
rect 1314 1781 1330 1821
rect 1264 1749 1330 1781
rect 1264 1713 1280 1749
rect 1314 1713 1330 1749
rect 1264 1679 1330 1713
rect 1264 1643 1280 1679
rect 1314 1643 1330 1679
rect 1264 1611 1330 1643
rect 1264 1571 1280 1611
rect 1314 1571 1330 1611
rect 1264 1543 1330 1571
rect 1264 1499 1280 1543
rect 1314 1499 1330 1543
rect 1264 1475 1330 1499
rect 1264 1427 1280 1475
rect 1314 1427 1330 1475
rect 1264 1407 1330 1427
rect 1264 1355 1280 1407
rect 1314 1355 1330 1407
rect 1264 1339 1330 1355
rect 1264 1283 1280 1339
rect 1314 1283 1330 1339
rect 1264 1271 1330 1283
rect 1264 1211 1280 1271
rect 1314 1211 1330 1271
rect 1264 1203 1330 1211
rect 1264 1139 1280 1203
rect 1314 1139 1330 1203
rect 1264 1135 1330 1139
rect 1264 1033 1280 1135
rect 1314 1033 1330 1135
rect 1264 1029 1330 1033
rect 1264 965 1280 1029
rect 1314 965 1330 1029
rect 1264 957 1330 965
rect 1264 897 1280 957
rect 1314 897 1330 957
rect 662 829 678 885
rect 712 829 728 885
rect 662 813 728 829
rect 662 761 678 813
rect 712 761 728 813
rect 662 728 728 761
rect 1264 885 1330 897
rect 1264 829 1280 885
rect 1314 829 1330 885
rect 1264 813 1330 829
rect 1264 761 1280 813
rect 1314 761 1330 813
rect 1264 728 1330 761
rect 662 712 1330 728
rect 662 678 678 712
rect 712 678 763 712
rect 809 678 835 712
rect 877 678 907 712
rect 945 678 979 712
rect 1013 678 1047 712
rect 1085 678 1115 712
rect 1157 678 1183 712
rect 1229 678 1280 712
rect 1314 678 1330 712
rect 662 662 1330 678
rect 1666 2721 1732 2733
rect 1666 2665 1682 2721
rect 1716 2665 1732 2721
rect 1666 2649 1732 2665
rect 1666 2597 1682 2649
rect 1716 2597 1732 2649
rect 1666 2577 1732 2597
rect 1666 2529 1682 2577
rect 1716 2529 1732 2577
rect 1666 2505 1732 2529
rect 1666 2461 1682 2505
rect 1716 2461 1732 2505
rect 1666 2433 1732 2461
rect 1666 2393 1682 2433
rect 1716 2393 1732 2433
rect 1666 2361 1732 2393
rect 1666 2325 1682 2361
rect 1716 2325 1732 2361
rect 1666 2291 1732 2325
rect 1666 2255 1682 2291
rect 1716 2255 1732 2291
rect 1666 2223 1732 2255
rect 1666 2183 1682 2223
rect 1716 2183 1732 2223
rect 1666 2155 1732 2183
rect 1666 2111 1682 2155
rect 1716 2111 1732 2155
rect 1666 2087 1732 2111
rect 1666 2039 1682 2087
rect 1716 2039 1732 2087
rect 1666 2019 1732 2039
rect 1666 1967 1682 2019
rect 1716 1967 1732 2019
rect 1666 1951 1732 1967
rect 1666 1895 1682 1951
rect 1716 1895 1732 1951
rect 1666 1883 1732 1895
rect 1666 1823 1682 1883
rect 1716 1823 1732 1883
rect 1666 1815 1732 1823
rect 1666 1751 1682 1815
rect 1716 1751 1732 1815
rect 1666 1747 1732 1751
rect 1666 1645 1682 1747
rect 1716 1645 1732 1747
rect 1666 1641 1732 1645
rect 1666 1577 1682 1641
rect 1716 1577 1732 1641
rect 1666 1569 1732 1577
rect 1666 1509 1682 1569
rect 1716 1509 1732 1569
rect 1666 1497 1732 1509
rect 1666 1441 1682 1497
rect 1716 1441 1732 1497
rect 1666 1425 1732 1441
rect 1666 1373 1682 1425
rect 1716 1373 1732 1425
rect 1666 1353 1732 1373
rect 1666 1305 1682 1353
rect 1716 1305 1732 1353
rect 1666 1281 1732 1305
rect 1666 1237 1682 1281
rect 1716 1237 1732 1281
rect 1666 1209 1732 1237
rect 1666 1169 1682 1209
rect 1716 1169 1732 1209
rect 1666 1137 1732 1169
rect 1666 1101 1682 1137
rect 1716 1101 1732 1137
rect 1666 1067 1732 1101
rect 1666 1031 1682 1067
rect 1716 1031 1732 1067
rect 1666 999 1732 1031
rect 1666 959 1682 999
rect 1716 959 1732 999
rect 1666 931 1732 959
rect 1666 887 1682 931
rect 1716 887 1732 931
rect 1666 863 1732 887
rect 1666 815 1682 863
rect 1716 815 1732 863
rect 1666 795 1732 815
rect 1666 743 1682 795
rect 1716 743 1732 795
rect 1666 727 1732 743
rect 1666 671 1682 727
rect 1716 671 1732 727
rect 260 599 276 659
rect 310 599 326 659
rect 260 591 326 599
rect 260 527 276 591
rect 310 527 326 591
rect 260 523 326 527
rect 260 421 276 523
rect 310 421 326 523
rect 260 417 326 421
rect 260 353 276 417
rect 310 353 326 417
rect 260 326 326 353
rect 1666 659 1732 671
rect 1666 599 1682 659
rect 1716 599 1732 659
rect 1666 591 1732 599
rect 1666 527 1682 591
rect 1716 527 1732 591
rect 1666 523 1732 527
rect 1666 421 1682 523
rect 1716 421 1732 523
rect 1666 417 1732 421
rect 1666 353 1682 417
rect 1716 353 1732 417
rect 1666 326 1732 353
rect 260 310 1732 326
rect 260 276 276 310
rect 310 276 367 310
rect 401 276 435 310
rect 473 276 503 310
rect 545 276 571 310
rect 617 276 639 310
rect 689 276 707 310
rect 761 276 775 310
rect 833 276 843 310
rect 905 276 911 310
rect 977 276 979 310
rect 1013 276 1015 310
rect 1081 276 1087 310
rect 1149 276 1159 310
rect 1217 276 1231 310
rect 1285 276 1303 310
rect 1353 276 1375 310
rect 1421 276 1447 310
rect 1489 276 1519 310
rect 1557 276 1591 310
rect 1625 276 1682 310
rect 1716 276 1732 310
rect 260 260 1732 276
rect 1892 3117 1958 3141
rect 1892 3073 1908 3117
rect 1942 3073 1958 3117
rect 1892 3045 1958 3073
rect 1892 3005 1908 3045
rect 1942 3005 1958 3045
rect 1892 2973 1958 3005
rect 1892 2937 1908 2973
rect 1942 2937 1958 2973
rect 1892 2903 1958 2937
rect 1892 2867 1908 2903
rect 1942 2867 1958 2903
rect 1892 2835 1958 2867
rect 1892 2795 1908 2835
rect 1942 2795 1958 2835
rect 1892 2767 1958 2795
rect 1892 2723 1908 2767
rect 1942 2723 1958 2767
rect 1892 2699 1958 2723
rect 1892 2651 1908 2699
rect 1942 2651 1958 2699
rect 1892 2631 1958 2651
rect 1892 2579 1908 2631
rect 1942 2579 1958 2631
rect 1892 2563 1958 2579
rect 1892 2507 1908 2563
rect 1942 2507 1958 2563
rect 1892 2495 1958 2507
rect 1892 2435 1908 2495
rect 1942 2435 1958 2495
rect 1892 2427 1958 2435
rect 1892 2363 1908 2427
rect 1942 2363 1958 2427
rect 1892 2359 1958 2363
rect 1892 2257 1908 2359
rect 1942 2257 1958 2359
rect 1892 2253 1958 2257
rect 1892 2189 1908 2253
rect 1942 2189 1958 2253
rect 1892 2181 1958 2189
rect 1892 2121 1908 2181
rect 1942 2121 1958 2181
rect 1892 2109 1958 2121
rect 1892 2053 1908 2109
rect 1942 2053 1958 2109
rect 1892 2037 1958 2053
rect 1892 1985 1908 2037
rect 1942 1985 1958 2037
rect 1892 1965 1958 1985
rect 1892 1917 1908 1965
rect 1942 1917 1958 1965
rect 1892 1893 1958 1917
rect 1892 1849 1908 1893
rect 1942 1849 1958 1893
rect 1892 1821 1958 1849
rect 1892 1781 1908 1821
rect 1942 1781 1958 1821
rect 1892 1749 1958 1781
rect 1892 1713 1908 1749
rect 1942 1713 1958 1749
rect 1892 1679 1958 1713
rect 1892 1643 1908 1679
rect 1942 1643 1958 1679
rect 1892 1611 1958 1643
rect 1892 1571 1908 1611
rect 1942 1571 1958 1611
rect 1892 1543 1958 1571
rect 1892 1499 1908 1543
rect 1942 1499 1958 1543
rect 1892 1475 1958 1499
rect 1892 1427 1908 1475
rect 1942 1427 1958 1475
rect 1892 1407 1958 1427
rect 1892 1355 1908 1407
rect 1942 1355 1958 1407
rect 1892 1339 1958 1355
rect 1892 1283 1908 1339
rect 1942 1283 1958 1339
rect 1892 1271 1958 1283
rect 1892 1211 1908 1271
rect 1942 1211 1958 1271
rect 1892 1203 1958 1211
rect 1892 1139 1908 1203
rect 1942 1139 1958 1203
rect 1892 1135 1958 1139
rect 1892 1033 1908 1135
rect 1942 1033 1958 1135
rect 1892 1029 1958 1033
rect 1892 965 1908 1029
rect 1942 965 1958 1029
rect 1892 957 1958 965
rect 1892 897 1908 957
rect 1942 897 1958 957
rect 1892 885 1958 897
rect 1892 829 1908 885
rect 1942 829 1958 885
rect 1892 813 1958 829
rect 1892 761 1908 813
rect 1942 761 1958 813
rect 1892 741 1958 761
rect 1892 693 1908 741
rect 1942 693 1958 741
rect 1892 669 1958 693
rect 1892 625 1908 669
rect 1942 625 1958 669
rect 1892 597 1958 625
rect 1892 557 1908 597
rect 1942 557 1958 597
rect 1892 525 1958 557
rect 1892 489 1908 525
rect 1942 489 1958 525
rect 1892 455 1958 489
rect 1892 419 1908 455
rect 1942 419 1958 455
rect 1892 387 1958 419
rect 1892 347 1908 387
rect 1942 347 1958 387
rect 1892 319 1958 347
rect 1892 275 1908 319
rect 1942 275 1958 319
rect 34 203 50 251
rect 84 203 100 251
rect 34 183 100 203
rect 34 131 50 183
rect 84 131 100 183
rect 34 100 100 131
rect 1892 251 1958 275
rect 1892 203 1908 251
rect 1942 203 1958 251
rect 1892 183 1958 203
rect 1892 131 1908 183
rect 1942 131 1958 183
rect 1892 100 1958 131
rect 34 84 1958 100
rect 34 50 50 84
rect 84 50 129 84
rect 185 50 197 84
rect 257 50 265 84
rect 329 50 333 84
rect 435 50 439 84
rect 503 50 511 84
rect 571 50 583 84
rect 639 50 655 84
rect 707 50 727 84
rect 775 50 799 84
rect 843 50 871 84
rect 911 50 943 84
rect 979 50 1013 84
rect 1049 50 1081 84
rect 1121 50 1149 84
rect 1193 50 1217 84
rect 1265 50 1285 84
rect 1337 50 1353 84
rect 1409 50 1421 84
rect 1481 50 1489 84
rect 1553 50 1557 84
rect 1659 50 1663 84
rect 1727 50 1735 84
rect 1795 50 1807 84
rect 1863 50 1908 84
rect 1942 50 1958 84
rect 34 34 1958 50
<< viali >>
rect 50 3308 84 3342
rect 151 3308 163 3342
rect 163 3308 185 3342
rect 223 3308 231 3342
rect 231 3308 257 3342
rect 295 3308 299 3342
rect 299 3308 329 3342
rect 367 3308 401 3342
rect 439 3308 469 3342
rect 469 3308 473 3342
rect 511 3308 537 3342
rect 537 3308 545 3342
rect 583 3308 605 3342
rect 605 3308 617 3342
rect 655 3308 673 3342
rect 673 3308 689 3342
rect 727 3308 741 3342
rect 741 3308 761 3342
rect 799 3308 809 3342
rect 809 3308 833 3342
rect 871 3308 877 3342
rect 877 3308 905 3342
rect 943 3308 945 3342
rect 945 3308 977 3342
rect 1015 3308 1047 3342
rect 1047 3308 1049 3342
rect 1087 3308 1115 3342
rect 1115 3308 1121 3342
rect 1159 3308 1183 3342
rect 1183 3308 1193 3342
rect 1231 3308 1251 3342
rect 1251 3308 1265 3342
rect 1303 3308 1319 3342
rect 1319 3308 1337 3342
rect 1375 3308 1387 3342
rect 1387 3308 1409 3342
rect 1447 3308 1455 3342
rect 1455 3308 1481 3342
rect 1519 3308 1523 3342
rect 1523 3308 1553 3342
rect 1591 3308 1625 3342
rect 1663 3308 1693 3342
rect 1693 3308 1697 3342
rect 1735 3308 1761 3342
rect 1761 3308 1769 3342
rect 1807 3308 1829 3342
rect 1829 3308 1841 3342
rect 1908 3308 1942 3342
rect 50 3243 84 3261
rect 50 3227 84 3243
rect 50 3175 84 3189
rect 50 3155 84 3175
rect 1908 3243 1942 3261
rect 1908 3227 1942 3243
rect 1908 3175 1942 3189
rect 1908 3155 1942 3175
rect 50 3107 84 3117
rect 50 3083 84 3107
rect 50 3039 84 3045
rect 50 3011 84 3039
rect 50 2971 84 2973
rect 50 2939 84 2971
rect 50 2869 84 2901
rect 50 2867 84 2869
rect 50 2801 84 2829
rect 50 2795 84 2801
rect 50 2733 84 2757
rect 50 2723 84 2733
rect 50 2665 84 2685
rect 50 2651 84 2665
rect 50 2597 84 2613
rect 50 2579 84 2597
rect 50 2529 84 2541
rect 50 2507 84 2529
rect 50 2461 84 2469
rect 50 2435 84 2461
rect 50 2393 84 2397
rect 50 2363 84 2393
rect 50 2291 84 2325
rect 50 2223 84 2253
rect 50 2219 84 2223
rect 50 2155 84 2181
rect 50 2147 84 2155
rect 50 2087 84 2109
rect 50 2075 84 2087
rect 50 2019 84 2037
rect 50 2003 84 2019
rect 50 1951 84 1965
rect 50 1931 84 1951
rect 50 1883 84 1893
rect 50 1859 84 1883
rect 50 1815 84 1821
rect 50 1787 84 1815
rect 50 1747 84 1749
rect 50 1715 84 1747
rect 50 1645 84 1677
rect 50 1643 84 1645
rect 50 1577 84 1605
rect 50 1571 84 1577
rect 50 1509 84 1533
rect 50 1499 84 1509
rect 50 1441 84 1461
rect 50 1427 84 1441
rect 50 1373 84 1389
rect 50 1355 84 1373
rect 50 1305 84 1317
rect 50 1283 84 1305
rect 50 1237 84 1245
rect 50 1211 84 1237
rect 50 1169 84 1173
rect 50 1139 84 1169
rect 50 1067 84 1101
rect 50 999 84 1029
rect 50 995 84 999
rect 50 931 84 957
rect 50 923 84 931
rect 50 863 84 885
rect 50 851 84 863
rect 50 795 84 813
rect 50 779 84 795
rect 50 727 84 741
rect 50 707 84 727
rect 50 659 84 669
rect 50 635 84 659
rect 50 591 84 597
rect 50 563 84 591
rect 50 523 84 525
rect 50 491 84 523
rect 50 421 84 453
rect 50 419 84 421
rect 50 353 84 381
rect 50 347 84 353
rect 50 285 84 309
rect 50 275 84 285
rect 276 3082 310 3116
rect 367 3082 401 3116
rect 439 3082 469 3116
rect 469 3082 473 3116
rect 511 3082 537 3116
rect 537 3082 545 3116
rect 583 3082 605 3116
rect 605 3082 617 3116
rect 655 3082 673 3116
rect 673 3082 689 3116
rect 727 3082 741 3116
rect 741 3082 761 3116
rect 799 3082 809 3116
rect 809 3082 833 3116
rect 871 3082 877 3116
rect 877 3082 905 3116
rect 943 3082 945 3116
rect 945 3082 977 3116
rect 1015 3082 1047 3116
rect 1047 3082 1049 3116
rect 1087 3082 1115 3116
rect 1115 3082 1121 3116
rect 1159 3082 1183 3116
rect 1183 3082 1193 3116
rect 1231 3082 1251 3116
rect 1251 3082 1265 3116
rect 1303 3082 1319 3116
rect 1319 3082 1337 3116
rect 1375 3082 1387 3116
rect 1387 3082 1409 3116
rect 1447 3082 1455 3116
rect 1455 3082 1481 3116
rect 1519 3082 1523 3116
rect 1523 3082 1553 3116
rect 1591 3082 1625 3116
rect 1682 3082 1716 3116
rect 276 3005 310 3009
rect 276 2975 310 3005
rect 276 2903 310 2937
rect 276 2835 310 2865
rect 276 2831 310 2835
rect 276 2767 310 2793
rect 276 2759 310 2767
rect 1682 3005 1716 3009
rect 1682 2975 1716 3005
rect 1682 2903 1716 2937
rect 1682 2835 1716 2865
rect 1682 2831 1716 2835
rect 1682 2767 1716 2793
rect 1682 2759 1716 2767
rect 276 2699 310 2721
rect 276 2687 310 2699
rect 276 2631 310 2649
rect 276 2615 310 2631
rect 276 2563 310 2577
rect 276 2543 310 2563
rect 276 2495 310 2505
rect 276 2471 310 2495
rect 276 2427 310 2433
rect 276 2399 310 2427
rect 276 2359 310 2361
rect 276 2327 310 2359
rect 276 2257 310 2289
rect 276 2255 310 2257
rect 276 2189 310 2217
rect 276 2183 310 2189
rect 276 2121 310 2145
rect 276 2111 310 2121
rect 276 2053 310 2073
rect 276 2039 310 2053
rect 276 1985 310 2001
rect 276 1967 310 1985
rect 276 1917 310 1929
rect 276 1895 310 1917
rect 276 1849 310 1857
rect 276 1823 310 1849
rect 276 1781 310 1785
rect 276 1751 310 1781
rect 276 1679 310 1713
rect 276 1611 310 1641
rect 276 1607 310 1611
rect 276 1543 310 1569
rect 276 1535 310 1543
rect 276 1475 310 1497
rect 276 1463 310 1475
rect 276 1407 310 1425
rect 276 1391 310 1407
rect 276 1339 310 1353
rect 276 1319 310 1339
rect 276 1271 310 1281
rect 276 1247 310 1271
rect 276 1203 310 1209
rect 276 1175 310 1203
rect 276 1135 310 1137
rect 276 1103 310 1135
rect 276 1033 310 1065
rect 276 1031 310 1033
rect 276 965 310 993
rect 276 959 310 965
rect 276 897 310 921
rect 276 887 310 897
rect 276 829 310 849
rect 276 815 310 829
rect 276 761 310 777
rect 276 743 310 761
rect 276 693 310 705
rect 276 671 310 693
rect 678 2680 712 2714
rect 763 2680 775 2714
rect 775 2680 797 2714
rect 835 2680 843 2714
rect 843 2680 869 2714
rect 907 2680 911 2714
rect 911 2680 941 2714
rect 979 2680 1013 2714
rect 1051 2680 1081 2714
rect 1081 2680 1085 2714
rect 1123 2680 1149 2714
rect 1149 2680 1157 2714
rect 1195 2680 1217 2714
rect 1217 2680 1229 2714
rect 1280 2680 1314 2714
rect 678 2597 712 2613
rect 678 2579 712 2597
rect 678 2529 712 2541
rect 678 2507 712 2529
rect 1280 2597 1314 2613
rect 1280 2579 1314 2597
rect 1280 2529 1314 2541
rect 1280 2507 1314 2529
rect 678 2461 712 2469
rect 678 2435 712 2461
rect 678 2393 712 2397
rect 678 2363 712 2393
rect 678 2291 712 2325
rect 678 2223 712 2253
rect 678 2219 712 2223
rect 678 2155 712 2181
rect 678 2147 712 2155
rect 678 2087 712 2109
rect 678 2075 712 2087
rect 678 2019 712 2037
rect 678 2003 712 2019
rect 678 1951 712 1965
rect 678 1931 712 1951
rect 678 1883 712 1893
rect 678 1859 712 1883
rect 678 1815 712 1821
rect 678 1787 712 1815
rect 678 1747 712 1749
rect 678 1715 712 1747
rect 678 1645 712 1677
rect 678 1643 712 1645
rect 678 1577 712 1605
rect 678 1571 712 1577
rect 678 1509 712 1533
rect 678 1499 712 1509
rect 678 1441 712 1461
rect 678 1427 712 1441
rect 678 1373 712 1389
rect 678 1355 712 1373
rect 678 1305 712 1317
rect 678 1283 712 1305
rect 678 1237 712 1245
rect 678 1211 712 1237
rect 678 1169 712 1173
rect 678 1139 712 1169
rect 678 1067 712 1101
rect 678 999 712 1029
rect 678 995 712 999
rect 678 931 712 957
rect 678 923 712 931
rect 907 2461 1085 2469
rect 907 931 911 2461
rect 911 931 1081 2461
rect 1081 931 1085 2461
rect 907 923 1085 931
rect 1280 2461 1314 2469
rect 1280 2435 1314 2461
rect 1280 2393 1314 2397
rect 1280 2363 1314 2393
rect 1280 2291 1314 2325
rect 1280 2223 1314 2253
rect 1280 2219 1314 2223
rect 1280 2155 1314 2181
rect 1280 2147 1314 2155
rect 1280 2087 1314 2109
rect 1280 2075 1314 2087
rect 1280 2019 1314 2037
rect 1280 2003 1314 2019
rect 1280 1951 1314 1965
rect 1280 1931 1314 1951
rect 1280 1883 1314 1893
rect 1280 1859 1314 1883
rect 1280 1815 1314 1821
rect 1280 1787 1314 1815
rect 1280 1747 1314 1749
rect 1280 1715 1314 1747
rect 1280 1645 1314 1677
rect 1280 1643 1314 1645
rect 1280 1577 1314 1605
rect 1280 1571 1314 1577
rect 1280 1509 1314 1533
rect 1280 1499 1314 1509
rect 1280 1441 1314 1461
rect 1280 1427 1314 1441
rect 1280 1373 1314 1389
rect 1280 1355 1314 1373
rect 1280 1305 1314 1317
rect 1280 1283 1314 1305
rect 1280 1237 1314 1245
rect 1280 1211 1314 1237
rect 1280 1169 1314 1173
rect 1280 1139 1314 1169
rect 1280 1067 1314 1101
rect 1280 999 1314 1029
rect 1280 995 1314 999
rect 1280 931 1314 957
rect 1280 923 1314 931
rect 678 863 712 885
rect 678 851 712 863
rect 678 795 712 813
rect 678 779 712 795
rect 1280 863 1314 885
rect 1280 851 1314 863
rect 1280 795 1314 813
rect 1280 779 1314 795
rect 678 678 712 712
rect 763 678 775 712
rect 775 678 797 712
rect 835 678 843 712
rect 843 678 869 712
rect 907 678 911 712
rect 911 678 941 712
rect 979 678 1013 712
rect 1051 678 1081 712
rect 1081 678 1085 712
rect 1123 678 1149 712
rect 1149 678 1157 712
rect 1195 678 1217 712
rect 1217 678 1229 712
rect 1280 678 1314 712
rect 1682 2699 1716 2721
rect 1682 2687 1716 2699
rect 1682 2631 1716 2649
rect 1682 2615 1716 2631
rect 1682 2563 1716 2577
rect 1682 2543 1716 2563
rect 1682 2495 1716 2505
rect 1682 2471 1716 2495
rect 1682 2427 1716 2433
rect 1682 2399 1716 2427
rect 1682 2359 1716 2361
rect 1682 2327 1716 2359
rect 1682 2257 1716 2289
rect 1682 2255 1716 2257
rect 1682 2189 1716 2217
rect 1682 2183 1716 2189
rect 1682 2121 1716 2145
rect 1682 2111 1716 2121
rect 1682 2053 1716 2073
rect 1682 2039 1716 2053
rect 1682 1985 1716 2001
rect 1682 1967 1716 1985
rect 1682 1917 1716 1929
rect 1682 1895 1716 1917
rect 1682 1849 1716 1857
rect 1682 1823 1716 1849
rect 1682 1781 1716 1785
rect 1682 1751 1716 1781
rect 1682 1679 1716 1713
rect 1682 1611 1716 1641
rect 1682 1607 1716 1611
rect 1682 1543 1716 1569
rect 1682 1535 1716 1543
rect 1682 1475 1716 1497
rect 1682 1463 1716 1475
rect 1682 1407 1716 1425
rect 1682 1391 1716 1407
rect 1682 1339 1716 1353
rect 1682 1319 1716 1339
rect 1682 1271 1716 1281
rect 1682 1247 1716 1271
rect 1682 1203 1716 1209
rect 1682 1175 1716 1203
rect 1682 1135 1716 1137
rect 1682 1103 1716 1135
rect 1682 1033 1716 1065
rect 1682 1031 1716 1033
rect 1682 965 1716 993
rect 1682 959 1716 965
rect 1682 897 1716 921
rect 1682 887 1716 897
rect 1682 829 1716 849
rect 1682 815 1716 829
rect 1682 761 1716 777
rect 1682 743 1716 761
rect 1682 693 1716 705
rect 1682 671 1716 693
rect 276 625 310 633
rect 276 599 310 625
rect 276 557 310 561
rect 276 527 310 557
rect 276 455 310 489
rect 276 387 310 417
rect 276 383 310 387
rect 1682 625 1716 633
rect 1682 599 1716 625
rect 1682 557 1716 561
rect 1682 527 1716 557
rect 1682 455 1716 489
rect 1682 387 1716 417
rect 1682 383 1716 387
rect 276 276 310 310
rect 367 276 401 310
rect 439 276 469 310
rect 469 276 473 310
rect 511 276 537 310
rect 537 276 545 310
rect 583 276 605 310
rect 605 276 617 310
rect 655 276 673 310
rect 673 276 689 310
rect 727 276 741 310
rect 741 276 761 310
rect 799 276 809 310
rect 809 276 833 310
rect 871 276 877 310
rect 877 276 905 310
rect 943 276 945 310
rect 945 276 977 310
rect 1015 276 1047 310
rect 1047 276 1049 310
rect 1087 276 1115 310
rect 1115 276 1121 310
rect 1159 276 1183 310
rect 1183 276 1193 310
rect 1231 276 1251 310
rect 1251 276 1265 310
rect 1303 276 1319 310
rect 1319 276 1337 310
rect 1375 276 1387 310
rect 1387 276 1409 310
rect 1447 276 1455 310
rect 1455 276 1481 310
rect 1519 276 1523 310
rect 1523 276 1553 310
rect 1591 276 1625 310
rect 1682 276 1716 310
rect 1908 3107 1942 3117
rect 1908 3083 1942 3107
rect 1908 3039 1942 3045
rect 1908 3011 1942 3039
rect 1908 2971 1942 2973
rect 1908 2939 1942 2971
rect 1908 2869 1942 2901
rect 1908 2867 1942 2869
rect 1908 2801 1942 2829
rect 1908 2795 1942 2801
rect 1908 2733 1942 2757
rect 1908 2723 1942 2733
rect 1908 2665 1942 2685
rect 1908 2651 1942 2665
rect 1908 2597 1942 2613
rect 1908 2579 1942 2597
rect 1908 2529 1942 2541
rect 1908 2507 1942 2529
rect 1908 2461 1942 2469
rect 1908 2435 1942 2461
rect 1908 2393 1942 2397
rect 1908 2363 1942 2393
rect 1908 2291 1942 2325
rect 1908 2223 1942 2253
rect 1908 2219 1942 2223
rect 1908 2155 1942 2181
rect 1908 2147 1942 2155
rect 1908 2087 1942 2109
rect 1908 2075 1942 2087
rect 1908 2019 1942 2037
rect 1908 2003 1942 2019
rect 1908 1951 1942 1965
rect 1908 1931 1942 1951
rect 1908 1883 1942 1893
rect 1908 1859 1942 1883
rect 1908 1815 1942 1821
rect 1908 1787 1942 1815
rect 1908 1747 1942 1749
rect 1908 1715 1942 1747
rect 1908 1645 1942 1677
rect 1908 1643 1942 1645
rect 1908 1577 1942 1605
rect 1908 1571 1942 1577
rect 1908 1509 1942 1533
rect 1908 1499 1942 1509
rect 1908 1441 1942 1461
rect 1908 1427 1942 1441
rect 1908 1373 1942 1389
rect 1908 1355 1942 1373
rect 1908 1305 1942 1317
rect 1908 1283 1942 1305
rect 1908 1237 1942 1245
rect 1908 1211 1942 1237
rect 1908 1169 1942 1173
rect 1908 1139 1942 1169
rect 1908 1067 1942 1101
rect 1908 999 1942 1029
rect 1908 995 1942 999
rect 1908 931 1942 957
rect 1908 923 1942 931
rect 1908 863 1942 885
rect 1908 851 1942 863
rect 1908 795 1942 813
rect 1908 779 1942 795
rect 1908 727 1942 741
rect 1908 707 1942 727
rect 1908 659 1942 669
rect 1908 635 1942 659
rect 1908 591 1942 597
rect 1908 563 1942 591
rect 1908 523 1942 525
rect 1908 491 1942 523
rect 1908 421 1942 453
rect 1908 419 1942 421
rect 1908 353 1942 381
rect 1908 347 1942 353
rect 1908 285 1942 309
rect 1908 275 1942 285
rect 50 217 84 237
rect 50 203 84 217
rect 50 149 84 165
rect 50 131 84 149
rect 1908 217 1942 237
rect 1908 203 1942 217
rect 1908 149 1942 165
rect 1908 131 1942 149
rect 50 50 84 84
rect 151 50 163 84
rect 163 50 185 84
rect 223 50 231 84
rect 231 50 257 84
rect 295 50 299 84
rect 299 50 329 84
rect 367 50 401 84
rect 439 50 469 84
rect 469 50 473 84
rect 511 50 537 84
rect 537 50 545 84
rect 583 50 605 84
rect 605 50 617 84
rect 655 50 673 84
rect 673 50 689 84
rect 727 50 741 84
rect 741 50 761 84
rect 799 50 809 84
rect 809 50 833 84
rect 871 50 877 84
rect 877 50 905 84
rect 943 50 945 84
rect 945 50 977 84
rect 1015 50 1047 84
rect 1047 50 1049 84
rect 1087 50 1115 84
rect 1115 50 1121 84
rect 1159 50 1183 84
rect 1183 50 1193 84
rect 1231 50 1251 84
rect 1251 50 1265 84
rect 1303 50 1319 84
rect 1319 50 1337 84
rect 1375 50 1387 84
rect 1387 50 1409 84
rect 1447 50 1455 84
rect 1455 50 1481 84
rect 1519 50 1523 84
rect 1523 50 1553 84
rect 1591 50 1625 84
rect 1663 50 1693 84
rect 1693 50 1697 84
rect 1735 50 1761 84
rect 1761 50 1769 84
rect 1807 50 1829 84
rect 1829 50 1841 84
rect 1908 50 1942 84
<< metal1 >>
rect 38 3342 1954 3354
rect 38 3308 50 3342
rect 84 3308 151 3342
rect 185 3308 223 3342
rect 257 3308 295 3342
rect 329 3308 367 3342
rect 401 3308 439 3342
rect 473 3308 511 3342
rect 545 3308 583 3342
rect 617 3308 655 3342
rect 689 3308 727 3342
rect 761 3308 799 3342
rect 833 3308 871 3342
rect 905 3308 943 3342
rect 977 3308 1015 3342
rect 1049 3308 1087 3342
rect 1121 3308 1159 3342
rect 1193 3308 1231 3342
rect 1265 3308 1303 3342
rect 1337 3308 1375 3342
rect 1409 3308 1447 3342
rect 1481 3308 1519 3342
rect 1553 3308 1591 3342
rect 1625 3308 1663 3342
rect 1697 3308 1735 3342
rect 1769 3308 1807 3342
rect 1841 3308 1908 3342
rect 1942 3308 1954 3342
rect 38 3296 1954 3308
rect 38 3261 96 3296
rect 38 3227 50 3261
rect 84 3227 96 3261
rect 38 3189 96 3227
rect 38 3155 50 3189
rect 84 3155 96 3189
rect 38 3117 96 3155
rect 1896 3261 1954 3296
rect 1896 3227 1908 3261
rect 1942 3227 1954 3261
rect 1896 3189 1954 3227
rect 1896 3155 1908 3189
rect 1942 3155 1954 3189
rect 38 3083 50 3117
rect 84 3083 96 3117
rect 38 3045 96 3083
rect 38 3011 50 3045
rect 84 3011 96 3045
rect 38 2973 96 3011
rect 38 2939 50 2973
rect 84 2939 96 2973
rect 38 2901 96 2939
rect 38 2867 50 2901
rect 84 2867 96 2901
rect 38 2829 96 2867
rect 38 2795 50 2829
rect 84 2795 96 2829
rect 38 2757 96 2795
rect 38 2723 50 2757
rect 84 2723 96 2757
rect 38 2685 96 2723
rect 38 2651 50 2685
rect 84 2651 96 2685
rect 38 2613 96 2651
rect 38 2579 50 2613
rect 84 2579 96 2613
rect 38 2541 96 2579
rect 38 2507 50 2541
rect 84 2507 96 2541
rect 38 2469 96 2507
rect 38 2435 50 2469
rect 84 2435 96 2469
rect 38 2397 96 2435
rect 38 2363 50 2397
rect 84 2363 96 2397
rect 38 2325 96 2363
rect 38 2291 50 2325
rect 84 2291 96 2325
rect 38 2253 96 2291
rect 38 2219 50 2253
rect 84 2219 96 2253
rect 38 2181 96 2219
rect 38 2147 50 2181
rect 84 2147 96 2181
rect 38 2109 96 2147
rect 38 2075 50 2109
rect 84 2075 96 2109
rect 38 2037 96 2075
rect 38 2003 50 2037
rect 84 2003 96 2037
rect 38 1965 96 2003
rect 38 1931 50 1965
rect 84 1931 96 1965
rect 38 1893 96 1931
rect 38 1859 50 1893
rect 84 1859 96 1893
rect 38 1821 96 1859
rect 38 1787 50 1821
rect 84 1787 96 1821
rect 38 1749 96 1787
rect 38 1715 50 1749
rect 84 1715 96 1749
rect 38 1677 96 1715
rect 38 1643 50 1677
rect 84 1643 96 1677
rect 38 1605 96 1643
rect 38 1571 50 1605
rect 84 1571 96 1605
rect 38 1533 96 1571
rect 38 1499 50 1533
rect 84 1499 96 1533
rect 38 1461 96 1499
rect 38 1427 50 1461
rect 84 1427 96 1461
rect 38 1389 96 1427
rect 38 1355 50 1389
rect 84 1355 96 1389
rect 38 1317 96 1355
rect 38 1283 50 1317
rect 84 1283 96 1317
rect 38 1245 96 1283
rect 38 1211 50 1245
rect 84 1211 96 1245
rect 38 1173 96 1211
rect 38 1139 50 1173
rect 84 1139 96 1173
rect 38 1101 96 1139
rect 38 1067 50 1101
rect 84 1067 96 1101
rect 38 1029 96 1067
rect 38 995 50 1029
rect 84 995 96 1029
rect 38 957 96 995
rect 38 923 50 957
rect 84 923 96 957
rect 38 885 96 923
rect 38 851 50 885
rect 84 851 96 885
rect 38 813 96 851
rect 38 779 50 813
rect 84 779 96 813
rect 38 741 96 779
rect 38 707 50 741
rect 84 707 96 741
rect 38 669 96 707
rect 38 635 50 669
rect 84 635 96 669
rect 38 597 96 635
rect 38 563 50 597
rect 84 563 96 597
rect 38 525 96 563
rect 38 491 50 525
rect 84 491 96 525
rect 38 453 96 491
rect 38 419 50 453
rect 84 419 96 453
rect 38 381 96 419
rect 38 347 50 381
rect 84 347 96 381
rect 38 309 96 347
rect 38 275 50 309
rect 84 275 96 309
rect 38 237 96 275
rect 264 3116 1728 3128
rect 264 3082 276 3116
rect 310 3082 367 3116
rect 401 3082 439 3116
rect 473 3082 511 3116
rect 545 3082 583 3116
rect 617 3082 655 3116
rect 689 3082 727 3116
rect 761 3082 799 3116
rect 833 3082 871 3116
rect 905 3082 943 3116
rect 977 3082 1015 3116
rect 1049 3082 1087 3116
rect 1121 3082 1159 3116
rect 1193 3082 1231 3116
rect 1265 3082 1303 3116
rect 1337 3082 1375 3116
rect 1409 3082 1447 3116
rect 1481 3082 1519 3116
rect 1553 3082 1591 3116
rect 1625 3082 1682 3116
rect 1716 3082 1728 3116
rect 264 3070 1728 3082
rect 264 3009 322 3070
rect 264 2975 276 3009
rect 310 2975 322 3009
rect 264 2937 322 2975
rect 264 2903 276 2937
rect 310 2903 322 2937
rect 264 2865 322 2903
rect 264 2831 276 2865
rect 310 2831 322 2865
rect 264 2793 322 2831
rect 264 2759 276 2793
rect 310 2759 322 2793
rect 264 2721 322 2759
rect 1670 3009 1728 3070
rect 1670 2975 1682 3009
rect 1716 2975 1728 3009
rect 1670 2937 1728 2975
rect 1670 2903 1682 2937
rect 1716 2903 1728 2937
rect 1670 2865 1728 2903
rect 1670 2831 1682 2865
rect 1716 2831 1728 2865
rect 1670 2793 1728 2831
rect 1670 2759 1682 2793
rect 1716 2759 1728 2793
rect 264 2687 276 2721
rect 310 2687 322 2721
rect 264 2649 322 2687
rect 264 2615 276 2649
rect 310 2615 322 2649
rect 264 2577 322 2615
rect 264 2543 276 2577
rect 310 2543 322 2577
rect 264 2505 322 2543
rect 264 2471 276 2505
rect 310 2471 322 2505
rect 264 2433 322 2471
rect 264 2399 276 2433
rect 310 2399 322 2433
rect 264 2361 322 2399
rect 264 2327 276 2361
rect 310 2327 322 2361
rect 264 2289 322 2327
rect 264 2255 276 2289
rect 310 2255 322 2289
rect 264 2217 322 2255
rect 264 2183 276 2217
rect 310 2183 322 2217
rect 264 2145 322 2183
rect 264 2111 276 2145
rect 310 2111 322 2145
rect 264 2073 322 2111
rect 264 2039 276 2073
rect 310 2039 322 2073
rect 264 2001 322 2039
rect 264 1967 276 2001
rect 310 1967 322 2001
rect 264 1929 322 1967
rect 264 1895 276 1929
rect 310 1895 322 1929
rect 264 1857 322 1895
rect 264 1823 276 1857
rect 310 1823 322 1857
rect 264 1785 322 1823
rect 264 1751 276 1785
rect 310 1751 322 1785
rect 264 1713 322 1751
rect 264 1679 276 1713
rect 310 1679 322 1713
rect 264 1641 322 1679
rect 264 1607 276 1641
rect 310 1607 322 1641
rect 264 1569 322 1607
rect 264 1535 276 1569
rect 310 1535 322 1569
rect 264 1497 322 1535
rect 264 1463 276 1497
rect 310 1463 322 1497
rect 264 1425 322 1463
rect 264 1391 276 1425
rect 310 1391 322 1425
rect 264 1353 322 1391
rect 264 1319 276 1353
rect 310 1319 322 1353
rect 264 1281 322 1319
rect 264 1247 276 1281
rect 310 1247 322 1281
rect 264 1209 322 1247
rect 264 1175 276 1209
rect 310 1175 322 1209
rect 264 1137 322 1175
rect 264 1103 276 1137
rect 310 1103 322 1137
rect 264 1065 322 1103
rect 264 1031 276 1065
rect 310 1031 322 1065
rect 264 993 322 1031
rect 264 959 276 993
rect 310 959 322 993
rect 264 921 322 959
rect 264 887 276 921
rect 310 887 322 921
rect 264 849 322 887
rect 264 815 276 849
rect 310 815 322 849
rect 264 777 322 815
rect 264 743 276 777
rect 310 743 322 777
rect 264 705 322 743
rect 264 671 276 705
rect 310 671 322 705
rect 264 633 322 671
rect 666 2714 1326 2726
rect 666 2680 678 2714
rect 712 2680 763 2714
rect 797 2680 835 2714
rect 869 2680 907 2714
rect 941 2680 979 2714
rect 1013 2680 1051 2714
rect 1085 2680 1123 2714
rect 1157 2680 1195 2714
rect 1229 2680 1280 2714
rect 1314 2680 1326 2714
rect 666 2668 1326 2680
rect 666 2613 724 2668
rect 666 2579 678 2613
rect 712 2579 724 2613
rect 666 2541 724 2579
rect 666 2507 678 2541
rect 712 2507 724 2541
rect 666 2469 724 2507
rect 1268 2613 1326 2668
rect 1268 2579 1280 2613
rect 1314 2579 1326 2613
rect 1268 2541 1326 2579
rect 1268 2507 1280 2541
rect 1314 2507 1326 2541
rect 666 2435 678 2469
rect 712 2435 724 2469
rect 666 2397 724 2435
rect 666 2363 678 2397
rect 712 2363 724 2397
rect 666 2325 724 2363
rect 666 2291 678 2325
rect 712 2291 724 2325
rect 666 2253 724 2291
rect 666 2219 678 2253
rect 712 2219 724 2253
rect 666 2181 724 2219
rect 666 2147 678 2181
rect 712 2147 724 2181
rect 666 2109 724 2147
rect 666 2075 678 2109
rect 712 2075 724 2109
rect 666 2037 724 2075
rect 666 2003 678 2037
rect 712 2003 724 2037
rect 666 1965 724 2003
rect 666 1931 678 1965
rect 712 1931 724 1965
rect 666 1893 724 1931
rect 666 1859 678 1893
rect 712 1859 724 1893
rect 666 1821 724 1859
rect 666 1787 678 1821
rect 712 1787 724 1821
rect 666 1749 724 1787
rect 666 1715 678 1749
rect 712 1715 724 1749
rect 666 1677 724 1715
rect 666 1643 678 1677
rect 712 1643 724 1677
rect 666 1605 724 1643
rect 666 1571 678 1605
rect 712 1571 724 1605
rect 666 1533 724 1571
rect 666 1499 678 1533
rect 712 1499 724 1533
rect 666 1461 724 1499
rect 666 1427 678 1461
rect 712 1427 724 1461
rect 666 1389 724 1427
rect 666 1355 678 1389
rect 712 1355 724 1389
rect 666 1317 724 1355
rect 666 1283 678 1317
rect 712 1283 724 1317
rect 666 1245 724 1283
rect 666 1211 678 1245
rect 712 1211 724 1245
rect 666 1173 724 1211
rect 666 1139 678 1173
rect 712 1139 724 1173
rect 666 1101 724 1139
rect 666 1067 678 1101
rect 712 1067 724 1101
rect 666 1029 724 1067
rect 666 995 678 1029
rect 712 995 724 1029
rect 666 957 724 995
rect 666 923 678 957
rect 712 923 724 957
rect 666 885 724 923
rect 895 2469 1097 2481
rect 895 923 907 2469
rect 1085 923 1097 2469
rect 895 911 1097 923
rect 1268 2469 1326 2507
rect 1268 2435 1280 2469
rect 1314 2435 1326 2469
rect 1268 2397 1326 2435
rect 1268 2363 1280 2397
rect 1314 2363 1326 2397
rect 1268 2325 1326 2363
rect 1268 2291 1280 2325
rect 1314 2291 1326 2325
rect 1268 2253 1326 2291
rect 1268 2219 1280 2253
rect 1314 2219 1326 2253
rect 1268 2181 1326 2219
rect 1268 2147 1280 2181
rect 1314 2147 1326 2181
rect 1268 2109 1326 2147
rect 1268 2075 1280 2109
rect 1314 2075 1326 2109
rect 1268 2037 1326 2075
rect 1268 2003 1280 2037
rect 1314 2003 1326 2037
rect 1268 1965 1326 2003
rect 1268 1931 1280 1965
rect 1314 1931 1326 1965
rect 1268 1893 1326 1931
rect 1268 1859 1280 1893
rect 1314 1859 1326 1893
rect 1268 1821 1326 1859
rect 1268 1787 1280 1821
rect 1314 1787 1326 1821
rect 1268 1749 1326 1787
rect 1268 1715 1280 1749
rect 1314 1715 1326 1749
rect 1268 1677 1326 1715
rect 1268 1643 1280 1677
rect 1314 1643 1326 1677
rect 1268 1605 1326 1643
rect 1268 1571 1280 1605
rect 1314 1571 1326 1605
rect 1268 1533 1326 1571
rect 1268 1499 1280 1533
rect 1314 1499 1326 1533
rect 1268 1461 1326 1499
rect 1268 1427 1280 1461
rect 1314 1427 1326 1461
rect 1268 1389 1326 1427
rect 1268 1355 1280 1389
rect 1314 1355 1326 1389
rect 1268 1317 1326 1355
rect 1268 1283 1280 1317
rect 1314 1283 1326 1317
rect 1268 1245 1326 1283
rect 1268 1211 1280 1245
rect 1314 1211 1326 1245
rect 1268 1173 1326 1211
rect 1268 1139 1280 1173
rect 1314 1139 1326 1173
rect 1268 1101 1326 1139
rect 1268 1067 1280 1101
rect 1314 1067 1326 1101
rect 1268 1029 1326 1067
rect 1268 995 1280 1029
rect 1314 995 1326 1029
rect 1268 957 1326 995
rect 1268 923 1280 957
rect 1314 923 1326 957
rect 666 851 678 885
rect 712 851 724 885
rect 666 813 724 851
rect 666 779 678 813
rect 712 779 724 813
rect 666 724 724 779
rect 1268 885 1326 923
rect 1268 851 1280 885
rect 1314 851 1326 885
rect 1268 813 1326 851
rect 1268 779 1280 813
rect 1314 779 1326 813
rect 1268 724 1326 779
rect 666 712 1326 724
rect 666 678 678 712
rect 712 678 763 712
rect 797 678 835 712
rect 869 678 907 712
rect 941 678 979 712
rect 1013 678 1051 712
rect 1085 678 1123 712
rect 1157 678 1195 712
rect 1229 678 1280 712
rect 1314 678 1326 712
rect 666 666 1326 678
rect 1670 2721 1728 2759
rect 1670 2687 1682 2721
rect 1716 2687 1728 2721
rect 1670 2649 1728 2687
rect 1670 2615 1682 2649
rect 1716 2615 1728 2649
rect 1670 2577 1728 2615
rect 1670 2543 1682 2577
rect 1716 2543 1728 2577
rect 1670 2505 1728 2543
rect 1670 2471 1682 2505
rect 1716 2471 1728 2505
rect 1670 2433 1728 2471
rect 1670 2399 1682 2433
rect 1716 2399 1728 2433
rect 1670 2361 1728 2399
rect 1670 2327 1682 2361
rect 1716 2327 1728 2361
rect 1670 2289 1728 2327
rect 1670 2255 1682 2289
rect 1716 2255 1728 2289
rect 1670 2217 1728 2255
rect 1670 2183 1682 2217
rect 1716 2183 1728 2217
rect 1670 2145 1728 2183
rect 1670 2111 1682 2145
rect 1716 2111 1728 2145
rect 1670 2073 1728 2111
rect 1670 2039 1682 2073
rect 1716 2039 1728 2073
rect 1670 2001 1728 2039
rect 1670 1967 1682 2001
rect 1716 1967 1728 2001
rect 1670 1929 1728 1967
rect 1670 1895 1682 1929
rect 1716 1895 1728 1929
rect 1670 1857 1728 1895
rect 1670 1823 1682 1857
rect 1716 1823 1728 1857
rect 1670 1785 1728 1823
rect 1670 1751 1682 1785
rect 1716 1751 1728 1785
rect 1670 1713 1728 1751
rect 1670 1679 1682 1713
rect 1716 1679 1728 1713
rect 1670 1641 1728 1679
rect 1670 1607 1682 1641
rect 1716 1607 1728 1641
rect 1670 1569 1728 1607
rect 1670 1535 1682 1569
rect 1716 1535 1728 1569
rect 1670 1497 1728 1535
rect 1670 1463 1682 1497
rect 1716 1463 1728 1497
rect 1670 1425 1728 1463
rect 1670 1391 1682 1425
rect 1716 1391 1728 1425
rect 1670 1353 1728 1391
rect 1670 1319 1682 1353
rect 1716 1319 1728 1353
rect 1670 1281 1728 1319
rect 1670 1247 1682 1281
rect 1716 1247 1728 1281
rect 1670 1209 1728 1247
rect 1670 1175 1682 1209
rect 1716 1175 1728 1209
rect 1670 1137 1728 1175
rect 1670 1103 1682 1137
rect 1716 1103 1728 1137
rect 1670 1065 1728 1103
rect 1670 1031 1682 1065
rect 1716 1031 1728 1065
rect 1670 993 1728 1031
rect 1670 959 1682 993
rect 1716 959 1728 993
rect 1670 921 1728 959
rect 1670 887 1682 921
rect 1716 887 1728 921
rect 1670 849 1728 887
rect 1670 815 1682 849
rect 1716 815 1728 849
rect 1670 777 1728 815
rect 1670 743 1682 777
rect 1716 743 1728 777
rect 1670 705 1728 743
rect 1670 671 1682 705
rect 1716 671 1728 705
rect 264 599 276 633
rect 310 599 322 633
rect 264 561 322 599
rect 264 527 276 561
rect 310 527 322 561
rect 264 489 322 527
rect 264 455 276 489
rect 310 455 322 489
rect 264 417 322 455
rect 264 383 276 417
rect 310 383 322 417
rect 264 322 322 383
rect 1670 633 1728 671
rect 1670 599 1682 633
rect 1716 599 1728 633
rect 1670 561 1728 599
rect 1670 527 1682 561
rect 1716 527 1728 561
rect 1670 489 1728 527
rect 1670 455 1682 489
rect 1716 455 1728 489
rect 1670 417 1728 455
rect 1670 383 1682 417
rect 1716 383 1728 417
rect 1670 322 1728 383
rect 264 310 1728 322
rect 264 276 276 310
rect 310 276 367 310
rect 401 276 439 310
rect 473 276 511 310
rect 545 276 583 310
rect 617 276 655 310
rect 689 276 727 310
rect 761 276 799 310
rect 833 276 871 310
rect 905 276 943 310
rect 977 276 1015 310
rect 1049 276 1087 310
rect 1121 276 1159 310
rect 1193 276 1231 310
rect 1265 276 1303 310
rect 1337 276 1375 310
rect 1409 276 1447 310
rect 1481 276 1519 310
rect 1553 276 1591 310
rect 1625 276 1682 310
rect 1716 276 1728 310
rect 264 264 1728 276
rect 1896 3117 1954 3155
rect 1896 3083 1908 3117
rect 1942 3083 1954 3117
rect 1896 3045 1954 3083
rect 1896 3011 1908 3045
rect 1942 3011 1954 3045
rect 1896 2973 1954 3011
rect 1896 2939 1908 2973
rect 1942 2939 1954 2973
rect 1896 2901 1954 2939
rect 1896 2867 1908 2901
rect 1942 2867 1954 2901
rect 1896 2829 1954 2867
rect 1896 2795 1908 2829
rect 1942 2795 1954 2829
rect 1896 2757 1954 2795
rect 1896 2723 1908 2757
rect 1942 2723 1954 2757
rect 1896 2685 1954 2723
rect 1896 2651 1908 2685
rect 1942 2651 1954 2685
rect 1896 2613 1954 2651
rect 1896 2579 1908 2613
rect 1942 2579 1954 2613
rect 1896 2541 1954 2579
rect 1896 2507 1908 2541
rect 1942 2507 1954 2541
rect 1896 2469 1954 2507
rect 1896 2435 1908 2469
rect 1942 2435 1954 2469
rect 1896 2397 1954 2435
rect 1896 2363 1908 2397
rect 1942 2363 1954 2397
rect 1896 2325 1954 2363
rect 1896 2291 1908 2325
rect 1942 2291 1954 2325
rect 1896 2253 1954 2291
rect 1896 2219 1908 2253
rect 1942 2219 1954 2253
rect 1896 2181 1954 2219
rect 1896 2147 1908 2181
rect 1942 2147 1954 2181
rect 1896 2109 1954 2147
rect 1896 2075 1908 2109
rect 1942 2075 1954 2109
rect 1896 2037 1954 2075
rect 1896 2003 1908 2037
rect 1942 2003 1954 2037
rect 1896 1965 1954 2003
rect 1896 1931 1908 1965
rect 1942 1931 1954 1965
rect 1896 1893 1954 1931
rect 1896 1859 1908 1893
rect 1942 1859 1954 1893
rect 1896 1821 1954 1859
rect 1896 1787 1908 1821
rect 1942 1787 1954 1821
rect 1896 1749 1954 1787
rect 1896 1715 1908 1749
rect 1942 1715 1954 1749
rect 1896 1677 1954 1715
rect 1896 1643 1908 1677
rect 1942 1643 1954 1677
rect 1896 1605 1954 1643
rect 1896 1571 1908 1605
rect 1942 1571 1954 1605
rect 1896 1533 1954 1571
rect 1896 1499 1908 1533
rect 1942 1499 1954 1533
rect 1896 1461 1954 1499
rect 1896 1427 1908 1461
rect 1942 1427 1954 1461
rect 1896 1389 1954 1427
rect 1896 1355 1908 1389
rect 1942 1355 1954 1389
rect 1896 1317 1954 1355
rect 1896 1283 1908 1317
rect 1942 1283 1954 1317
rect 1896 1245 1954 1283
rect 1896 1211 1908 1245
rect 1942 1211 1954 1245
rect 1896 1173 1954 1211
rect 1896 1139 1908 1173
rect 1942 1139 1954 1173
rect 1896 1101 1954 1139
rect 1896 1067 1908 1101
rect 1942 1067 1954 1101
rect 1896 1029 1954 1067
rect 1896 995 1908 1029
rect 1942 995 1954 1029
rect 1896 957 1954 995
rect 1896 923 1908 957
rect 1942 923 1954 957
rect 1896 885 1954 923
rect 1896 851 1908 885
rect 1942 851 1954 885
rect 1896 813 1954 851
rect 1896 779 1908 813
rect 1942 779 1954 813
rect 1896 741 1954 779
rect 1896 707 1908 741
rect 1942 707 1954 741
rect 1896 669 1954 707
rect 1896 635 1908 669
rect 1942 635 1954 669
rect 1896 597 1954 635
rect 1896 563 1908 597
rect 1942 563 1954 597
rect 1896 525 1954 563
rect 1896 491 1908 525
rect 1942 491 1954 525
rect 1896 453 1954 491
rect 1896 419 1908 453
rect 1942 419 1954 453
rect 1896 381 1954 419
rect 1896 347 1908 381
rect 1942 347 1954 381
rect 1896 309 1954 347
rect 1896 275 1908 309
rect 1942 275 1954 309
rect 38 203 50 237
rect 84 203 96 237
rect 38 165 96 203
rect 38 131 50 165
rect 84 131 96 165
rect 38 96 96 131
rect 1896 237 1954 275
rect 1896 203 1908 237
rect 1942 203 1954 237
rect 1896 165 1954 203
rect 1896 131 1908 165
rect 1942 131 1954 165
rect 1896 96 1954 131
rect 38 84 1954 96
rect 38 50 50 84
rect 84 50 151 84
rect 185 50 223 84
rect 257 50 295 84
rect 329 50 367 84
rect 401 50 439 84
rect 473 50 511 84
rect 545 50 583 84
rect 617 50 655 84
rect 689 50 727 84
rect 761 50 799 84
rect 833 50 871 84
rect 905 50 943 84
rect 977 50 1015 84
rect 1049 50 1087 84
rect 1121 50 1159 84
rect 1193 50 1231 84
rect 1265 50 1303 84
rect 1337 50 1375 84
rect 1409 50 1447 84
rect 1481 50 1519 84
rect 1553 50 1591 84
rect 1625 50 1663 84
rect 1697 50 1735 84
rect 1769 50 1807 84
rect 1841 50 1908 84
rect 1942 50 1954 84
rect 38 38 1954 50
<< properties >>
string GDS_END 8872010
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8811326
string path 7.850 12.350 7.850 76.950 41.950 76.950 41.950 7.850 3.350 7.850 
<< end >>
