magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< pwell >>
rect 15 163 655 545
<< nmoslvt >>
rect 171 189 201 519
rect 257 189 307 519
rect 363 189 413 519
rect 469 189 499 519
<< ndiff >>
rect 111 507 171 519
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 507 257 519
rect 201 201 212 507
rect 246 201 257 507
rect 201 189 257 201
rect 307 507 363 519
rect 307 201 318 507
rect 352 201 363 507
rect 307 189 363 201
rect 413 507 469 519
rect 413 201 424 507
rect 458 201 469 507
rect 413 189 469 201
rect 499 507 559 519
rect 499 473 510 507
rect 544 473 559 507
rect 499 439 559 473
rect 499 405 510 439
rect 544 405 559 439
rect 499 371 559 405
rect 499 337 510 371
rect 544 337 559 371
rect 499 303 559 337
rect 499 269 510 303
rect 544 269 559 303
rect 499 235 559 269
rect 499 201 510 235
rect 544 201 559 235
rect 499 189 559 201
<< ndiffc >>
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 201 246 507
rect 318 201 352 507
rect 424 201 458 507
rect 510 473 544 507
rect 510 405 544 439
rect 510 337 544 371
rect 510 269 544 303
rect 510 201 544 235
<< psubdiff >>
rect 41 507 111 519
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 559 507 629 519
rect 559 473 578 507
rect 612 473 629 507
rect 559 439 629 473
rect 559 405 578 439
rect 612 405 629 439
rect 559 371 629 405
rect 559 337 578 371
rect 612 337 629 371
rect 559 303 629 337
rect 559 269 578 303
rect 612 269 629 303
rect 559 235 629 269
rect 559 201 578 235
rect 612 201 629 235
rect 559 189 629 201
<< psubdiffcont >>
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 578 473 612 507
rect 578 405 612 439
rect 578 337 612 371
rect 578 269 612 303
rect 578 201 612 235
<< poly >>
rect 243 619 427 635
rect 120 595 201 611
rect 120 561 136 595
rect 170 561 201 595
rect 243 585 264 619
rect 406 585 427 619
rect 243 569 427 585
rect 469 595 550 611
rect 120 545 201 561
rect 171 519 201 545
rect 257 519 307 569
rect 363 519 413 569
rect 469 561 500 595
rect 534 561 550 595
rect 469 545 550 561
rect 469 519 499 545
rect 171 163 201 189
rect 120 147 201 163
rect 120 113 136 147
rect 170 113 201 147
rect 257 139 307 189
rect 363 139 413 189
rect 469 163 499 189
rect 469 147 550 163
rect 120 97 201 113
rect 243 123 427 139
rect 243 89 264 123
rect 406 89 427 123
rect 469 113 500 147
rect 534 113 550 147
rect 469 97 550 113
rect 243 73 427 89
<< polycont >>
rect 136 561 170 595
rect 264 585 406 619
rect 500 561 534 595
rect 136 113 170 147
rect 264 89 406 123
rect 500 113 534 147
<< locali >>
rect 248 689 422 708
rect 248 655 276 689
rect 310 655 360 689
rect 394 655 422 689
rect 248 619 422 655
rect 120 595 186 611
rect 120 561 136 595
rect 170 561 186 595
rect 248 585 264 619
rect 406 585 422 619
rect 248 583 276 585
rect 310 583 360 585
rect 394 583 422 585
rect 248 569 422 583
rect 484 595 550 611
rect 120 545 186 561
rect 484 561 500 595
rect 534 561 550 595
rect 484 545 550 561
rect 120 523 160 545
rect 510 523 550 545
rect 41 507 160 523
rect 41 473 58 507
rect 92 479 126 507
rect 94 473 126 479
rect 41 445 60 473
rect 94 445 160 473
rect 41 439 160 445
rect 41 405 58 439
rect 92 407 126 439
rect 94 405 126 407
rect 41 373 60 405
rect 94 373 160 405
rect 41 371 160 373
rect 41 337 58 371
rect 92 337 126 371
rect 41 335 160 337
rect 41 303 60 335
rect 94 303 160 335
rect 41 269 58 303
rect 94 301 126 303
rect 92 269 126 301
rect 41 263 160 269
rect 41 235 60 263
rect 94 235 160 263
rect 41 201 58 235
rect 94 229 126 235
rect 92 201 126 229
rect 41 185 160 201
rect 212 507 246 523
rect 212 185 246 201
rect 318 507 352 523
rect 318 185 352 201
rect 424 507 458 523
rect 424 185 458 201
rect 510 507 629 523
rect 544 479 578 507
rect 544 473 576 479
rect 612 473 629 507
rect 510 445 576 473
rect 610 445 629 473
rect 510 439 629 445
rect 544 407 578 439
rect 544 405 576 407
rect 612 405 629 439
rect 510 373 576 405
rect 610 373 629 405
rect 510 371 629 373
rect 544 337 578 371
rect 612 337 629 371
rect 510 335 629 337
rect 510 303 576 335
rect 610 303 629 335
rect 544 301 576 303
rect 544 269 578 301
rect 612 269 629 303
rect 510 263 629 269
rect 510 235 576 263
rect 610 235 629 263
rect 544 229 576 235
rect 544 201 578 229
rect 612 201 629 235
rect 510 185 629 201
rect 120 163 160 185
rect 510 163 550 185
rect 120 147 186 163
rect 120 113 136 147
rect 170 113 186 147
rect 484 147 550 163
rect 120 97 186 113
rect 248 125 422 139
rect 248 123 276 125
rect 310 123 360 125
rect 394 123 422 125
rect 248 89 264 123
rect 406 89 422 123
rect 484 113 500 147
rect 534 113 550 147
rect 484 97 550 113
rect 248 53 422 89
rect 248 19 276 53
rect 310 19 360 53
rect 394 19 422 53
rect 248 0 422 19
<< viali >>
rect 276 655 310 689
rect 360 655 394 689
rect 276 585 310 617
rect 360 585 394 617
rect 276 583 310 585
rect 360 583 394 585
rect 60 473 92 479
rect 92 473 94 479
rect 60 445 94 473
rect 60 405 92 407
rect 92 405 94 407
rect 60 373 94 405
rect 60 303 94 335
rect 60 301 92 303
rect 92 301 94 303
rect 60 235 94 263
rect 60 229 92 235
rect 92 229 94 235
rect 212 445 246 479
rect 212 373 246 407
rect 212 301 246 335
rect 212 229 246 263
rect 318 445 352 479
rect 318 373 352 407
rect 318 301 352 335
rect 318 229 352 263
rect 424 445 458 479
rect 424 373 458 407
rect 424 301 458 335
rect 424 229 458 263
rect 576 473 578 479
rect 578 473 610 479
rect 576 445 610 473
rect 576 405 578 407
rect 578 405 610 407
rect 576 373 610 405
rect 576 303 610 335
rect 576 301 578 303
rect 578 301 610 303
rect 576 235 610 263
rect 576 229 578 235
rect 578 229 610 235
rect 276 123 310 125
rect 360 123 394 125
rect 276 91 310 123
rect 360 91 394 123
rect 276 19 310 53
rect 360 19 394 53
<< metal1 >>
rect 250 689 420 708
rect 250 655 276 689
rect 310 655 360 689
rect 394 655 420 689
rect 250 617 420 655
rect 250 583 276 617
rect 310 583 360 617
rect 394 583 420 617
rect 250 571 420 583
rect 41 479 100 507
rect 41 445 60 479
rect 94 445 100 479
rect 41 407 100 445
rect 41 373 60 407
rect 94 373 100 407
rect 41 335 100 373
rect 41 301 60 335
rect 94 301 100 335
rect 41 263 100 301
rect 41 229 60 263
rect 94 229 100 263
rect 41 201 100 229
rect 203 479 255 507
rect 203 445 212 479
rect 246 445 255 479
rect 203 407 255 445
rect 203 373 212 407
rect 246 373 255 407
rect 203 335 255 373
rect 203 323 212 335
rect 246 323 255 335
rect 203 263 255 271
rect 203 259 212 263
rect 246 259 255 263
rect 203 201 255 207
rect 309 501 361 507
rect 309 445 318 449
rect 352 445 361 449
rect 309 437 361 445
rect 309 373 318 385
rect 352 373 361 385
rect 309 335 361 373
rect 309 301 318 335
rect 352 301 361 335
rect 309 263 361 301
rect 309 229 318 263
rect 352 229 361 263
rect 309 201 361 229
rect 415 479 467 507
rect 415 445 424 479
rect 458 445 467 479
rect 415 407 467 445
rect 415 373 424 407
rect 458 373 467 407
rect 415 335 467 373
rect 415 323 424 335
rect 458 323 467 335
rect 415 263 467 271
rect 415 259 424 263
rect 458 259 467 263
rect 415 201 467 207
rect 570 479 629 507
rect 570 445 576 479
rect 610 445 629 479
rect 570 407 629 445
rect 570 373 576 407
rect 610 373 629 407
rect 570 335 629 373
rect 570 301 576 335
rect 610 301 629 335
rect 570 263 629 301
rect 570 229 576 263
rect 610 229 629 263
rect 570 201 629 229
rect 250 125 420 137
rect 250 91 276 125
rect 310 91 360 125
rect 394 91 420 125
rect 250 53 420 91
rect 250 19 276 53
rect 310 19 360 53
rect 394 19 420 53
rect 250 0 420 19
<< via1 >>
rect 203 301 212 323
rect 212 301 246 323
rect 246 301 255 323
rect 203 271 255 301
rect 203 229 212 259
rect 212 229 246 259
rect 246 229 255 259
rect 203 207 255 229
rect 309 479 361 501
rect 309 449 318 479
rect 318 449 352 479
rect 352 449 361 479
rect 309 407 361 437
rect 309 385 318 407
rect 318 385 352 407
rect 352 385 361 407
rect 415 301 424 323
rect 424 301 458 323
rect 458 301 467 323
rect 415 271 467 301
rect 415 229 424 259
rect 424 229 458 259
rect 458 229 467 259
rect 415 207 467 229
<< metal2 >>
rect 14 501 656 507
rect 14 449 309 501
rect 361 449 656 501
rect 14 437 656 449
rect 14 385 309 437
rect 361 385 656 437
rect 14 379 656 385
rect 14 323 656 329
rect 14 271 203 323
rect 255 271 415 323
rect 467 271 656 323
rect 14 259 656 271
rect 14 207 203 259
rect 255 207 415 259
rect 467 207 656 259
rect 14 201 656 207
<< labels >>
flabel comment s 184 358 184 358 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 481 356 481 356 0 FreeSans 180 90 0 0 dummy_poly
flabel metal1 s 255 608 414 659 0 FreeSans 200 0 0 0 GATE
port 1 nsew
flabel metal1 s 255 44 414 95 0 FreeSans 200 0 0 0 GATE
port 1 nsew
flabel metal1 s 41 339 87 369 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal1 s 583 339 629 369 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal2 s 14 201 35 329 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 14 379 35 507 7 FreeSans 300 180 0 0 DRAIN
port 4 nsew
<< properties >>
string GDS_END 3927222
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 3917270
<< end >>
