magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 315 157 1193 203
rect 1 21 1193 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 393 47 423 177
rect 477 47 507 177
rect 561 47 591 177
rect 645 47 675 177
rect 833 47 863 177
rect 917 47 947 177
rect 1001 47 1031 177
rect 1085 47 1115 177
<< scpmoshvt >>
rect 79 413 109 497
rect 163 413 193 497
rect 393 297 423 497
rect 477 297 507 497
rect 561 297 591 497
rect 645 297 675 497
rect 833 297 863 497
rect 917 297 947 497
rect 1001 297 1031 497
rect 1085 297 1115 497
<< ndiff >>
rect 27 109 79 131
rect 27 75 35 109
rect 69 75 79 109
rect 27 47 79 75
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 109 287 131
rect 193 75 203 109
rect 237 75 287 109
rect 193 47 287 75
rect 341 101 393 177
rect 341 67 349 101
rect 383 67 393 101
rect 341 47 393 67
rect 423 165 477 177
rect 423 131 433 165
rect 467 131 477 165
rect 423 47 477 131
rect 507 97 561 177
rect 507 63 517 97
rect 551 63 561 97
rect 507 47 561 63
rect 591 165 645 177
rect 591 131 601 165
rect 635 131 645 165
rect 591 47 645 131
rect 675 97 727 177
rect 675 63 685 97
rect 719 63 727 97
rect 675 47 727 63
rect 781 97 833 177
rect 781 63 789 97
rect 823 63 833 97
rect 781 47 833 63
rect 863 165 917 177
rect 863 131 873 165
rect 907 131 917 165
rect 863 47 917 131
rect 947 165 1001 177
rect 947 131 957 165
rect 991 131 1001 165
rect 947 97 1001 131
rect 947 63 957 97
rect 991 63 1001 97
rect 947 47 1001 63
rect 1031 97 1085 177
rect 1031 63 1041 97
rect 1075 63 1085 97
rect 1031 47 1085 63
rect 1115 165 1167 177
rect 1115 131 1125 165
rect 1159 131 1167 165
rect 1115 97 1167 131
rect 1115 63 1125 97
rect 1159 63 1167 97
rect 1115 47 1167 63
<< pdiff >>
rect 27 472 79 497
rect 27 438 35 472
rect 69 438 79 472
rect 27 413 79 438
rect 109 489 163 497
rect 109 455 119 489
rect 153 455 163 489
rect 109 413 163 455
rect 193 483 287 497
rect 193 449 203 483
rect 237 449 287 483
rect 193 413 287 449
rect 341 485 393 497
rect 341 451 349 485
rect 383 451 393 485
rect 341 417 393 451
rect 341 383 349 417
rect 383 383 393 417
rect 341 349 393 383
rect 341 315 349 349
rect 383 315 393 349
rect 341 297 393 315
rect 423 477 477 497
rect 423 443 433 477
rect 467 443 477 477
rect 423 374 477 443
rect 423 340 433 374
rect 467 340 477 374
rect 423 297 477 340
rect 507 485 561 497
rect 507 451 517 485
rect 551 451 561 485
rect 507 417 561 451
rect 507 383 517 417
rect 551 383 561 417
rect 507 297 561 383
rect 591 485 645 497
rect 591 451 601 485
rect 635 451 645 485
rect 591 417 645 451
rect 591 383 601 417
rect 635 383 645 417
rect 591 349 645 383
rect 591 315 601 349
rect 635 315 645 349
rect 591 297 645 315
rect 675 485 833 497
rect 675 451 701 485
rect 735 451 773 485
rect 807 451 833 485
rect 675 417 833 451
rect 675 383 701 417
rect 735 383 773 417
rect 807 383 833 417
rect 675 297 833 383
rect 863 485 917 497
rect 863 451 873 485
rect 907 451 917 485
rect 863 417 917 451
rect 863 383 873 417
rect 907 383 917 417
rect 863 349 917 383
rect 863 315 873 349
rect 907 315 917 349
rect 863 297 917 315
rect 947 485 1001 497
rect 947 451 957 485
rect 991 451 1001 485
rect 947 417 1001 451
rect 947 383 957 417
rect 991 383 1001 417
rect 947 297 1001 383
rect 1031 485 1085 497
rect 1031 451 1041 485
rect 1075 451 1085 485
rect 1031 417 1085 451
rect 1031 383 1041 417
rect 1075 383 1085 417
rect 1031 349 1085 383
rect 1031 315 1041 349
rect 1075 315 1085 349
rect 1031 297 1085 315
rect 1115 485 1167 497
rect 1115 451 1125 485
rect 1159 451 1167 485
rect 1115 417 1167 451
rect 1115 383 1125 417
rect 1159 383 1167 417
rect 1115 349 1167 383
rect 1115 315 1125 349
rect 1159 315 1167 349
rect 1115 297 1167 315
<< ndiffc >>
rect 35 75 69 109
rect 119 59 153 93
rect 203 75 237 109
rect 349 67 383 101
rect 433 131 467 165
rect 517 63 551 97
rect 601 131 635 165
rect 685 63 719 97
rect 789 63 823 97
rect 873 131 907 165
rect 957 131 991 165
rect 957 63 991 97
rect 1041 63 1075 97
rect 1125 131 1159 165
rect 1125 63 1159 97
<< pdiffc >>
rect 35 438 69 472
rect 119 455 153 489
rect 203 449 237 483
rect 349 451 383 485
rect 349 383 383 417
rect 349 315 383 349
rect 433 443 467 477
rect 433 340 467 374
rect 517 451 551 485
rect 517 383 551 417
rect 601 451 635 485
rect 601 383 635 417
rect 601 315 635 349
rect 701 451 735 485
rect 773 451 807 485
rect 701 383 735 417
rect 773 383 807 417
rect 873 451 907 485
rect 873 383 907 417
rect 873 315 907 349
rect 957 451 991 485
rect 957 383 991 417
rect 1041 451 1075 485
rect 1041 383 1075 417
rect 1041 315 1075 349
rect 1125 451 1159 485
rect 1125 383 1159 417
rect 1125 315 1159 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 393 497 423 523
rect 477 497 507 523
rect 561 497 591 523
rect 645 497 675 523
rect 833 497 863 523
rect 917 497 947 523
rect 1001 497 1031 523
rect 1085 497 1115 523
rect 79 387 109 413
rect 46 357 109 387
rect 46 280 76 357
rect 163 284 193 413
rect 21 264 76 280
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 268 193 284
rect 118 234 128 268
rect 162 234 193 268
rect 393 265 423 297
rect 118 218 193 234
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 218
rect 272 259 423 265
rect 477 259 507 297
rect 561 259 591 297
rect 645 259 675 297
rect 833 259 863 297
rect 917 259 947 297
rect 1001 259 1031 297
rect 1085 261 1115 297
rect 1085 259 1175 261
rect 272 249 507 259
rect 272 215 282 249
rect 316 215 507 249
rect 272 205 507 215
rect 549 249 675 259
rect 549 215 565 249
rect 599 215 675 249
rect 549 205 675 215
rect 767 249 947 259
rect 767 215 783 249
rect 817 215 873 249
rect 907 215 947 249
rect 767 205 947 215
rect 989 249 1175 259
rect 989 215 1005 249
rect 1039 215 1125 249
rect 1159 215 1175 249
rect 989 205 1175 215
rect 272 199 423 205
rect 393 177 423 199
rect 477 177 507 205
rect 561 177 591 205
rect 645 177 675 205
rect 833 177 863 205
rect 917 177 947 205
rect 1001 177 1031 205
rect 1085 203 1175 205
rect 1085 177 1115 203
rect 79 21 109 47
rect 163 21 193 47
rect 393 21 423 47
rect 477 21 507 47
rect 561 21 591 47
rect 645 21 675 47
rect 833 21 863 47
rect 917 21 947 47
rect 1001 21 1031 47
rect 1085 21 1115 47
<< polycont >>
rect 32 230 66 264
rect 128 234 162 268
rect 282 215 316 249
rect 565 215 599 249
rect 783 215 817 249
rect 873 215 907 249
rect 1005 215 1039 249
rect 1125 215 1159 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 108 489 153 527
rect 17 472 74 488
rect 17 438 35 472
rect 69 438 74 472
rect 108 455 119 489
rect 108 439 153 455
rect 187 483 315 493
rect 187 449 203 483
rect 237 449 315 483
rect 17 396 74 438
rect 187 430 315 449
rect 17 357 246 396
rect 17 264 66 323
rect 122 268 178 323
rect 17 230 32 264
rect 112 234 128 268
rect 162 234 178 268
rect 17 214 66 230
rect 122 214 178 234
rect 212 255 246 357
rect 212 180 246 221
rect 17 146 246 180
rect 280 282 315 430
rect 349 485 383 527
rect 349 417 383 451
rect 349 349 383 383
rect 349 299 383 315
rect 417 477 467 493
rect 417 443 433 477
rect 417 374 467 443
rect 417 340 433 374
rect 501 485 551 527
rect 501 451 517 485
rect 501 417 551 451
rect 501 383 517 417
rect 501 367 551 383
rect 585 485 651 493
rect 585 451 601 485
rect 635 451 651 485
rect 585 417 651 451
rect 585 383 601 417
rect 635 383 651 417
rect 417 333 467 340
rect 585 349 651 383
rect 685 485 823 527
rect 685 451 701 485
rect 735 451 773 485
rect 807 451 823 485
rect 685 417 823 451
rect 685 383 701 417
rect 735 383 773 417
rect 807 383 823 417
rect 685 367 823 383
rect 857 485 923 493
rect 857 451 873 485
rect 907 451 923 485
rect 857 417 923 451
rect 857 383 873 417
rect 907 383 923 417
rect 585 333 601 349
rect 417 315 601 333
rect 635 333 651 349
rect 857 349 923 383
rect 957 485 991 527
rect 957 417 991 451
rect 957 367 991 383
rect 1025 485 1091 493
rect 1025 451 1041 485
rect 1075 451 1091 485
rect 1025 417 1091 451
rect 1025 383 1041 417
rect 1075 383 1091 417
rect 857 333 873 349
rect 635 315 873 333
rect 907 333 923 349
rect 1025 349 1091 383
rect 1025 333 1041 349
rect 907 315 1041 333
rect 1075 315 1091 349
rect 417 289 1091 315
rect 1125 485 1179 527
rect 1159 451 1179 485
rect 1125 417 1179 451
rect 1159 383 1179 417
rect 1125 349 1179 383
rect 1159 315 1179 349
rect 1125 289 1179 315
rect 280 249 316 282
rect 280 215 282 249
rect 17 109 69 146
rect 280 143 316 215
rect 417 165 483 289
rect 549 249 581 255
rect 549 215 565 249
rect 599 215 615 221
rect 649 215 710 289
rect 744 249 923 255
rect 744 215 783 249
rect 817 215 873 249
rect 907 215 923 249
rect 989 249 1175 255
rect 989 215 1005 249
rect 1039 215 1125 249
rect 1159 215 1175 249
rect 280 112 315 143
rect 417 131 433 165
rect 467 131 483 165
rect 585 165 923 181
rect 585 131 601 165
rect 635 131 873 165
rect 907 131 923 165
rect 957 165 1179 181
rect 991 147 1125 165
rect 991 131 1007 147
rect 187 109 315 112
rect 17 75 35 109
rect 17 51 69 75
rect 103 93 153 109
rect 103 59 119 93
rect 103 17 153 59
rect 187 75 203 109
rect 237 75 315 109
rect 187 51 315 75
rect 349 101 383 117
rect 957 97 1007 131
rect 1109 131 1125 147
rect 1159 131 1179 165
rect 383 67 517 97
rect 349 63 517 67
rect 551 63 685 97
rect 719 63 735 97
rect 349 51 735 63
rect 773 63 789 97
rect 823 63 957 97
rect 991 63 1007 97
rect 773 51 1007 63
rect 1041 97 1075 113
rect 1041 17 1075 63
rect 1109 97 1179 131
rect 1109 63 1125 97
rect 1159 63 1179 97
rect 1109 51 1179 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 212 221 246 255
rect 581 249 615 255
rect 581 221 599 249
rect 599 221 615 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 200 255 627 261
rect 200 221 212 255
rect 246 221 581 255
rect 615 221 627 255
rect 200 215 627 221
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 1137 221 1171 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 1045 221 1079 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 769 221 803 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 B_N
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 B_N
port 2 nsew signal input
flabel locali s 122 289 156 323 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 673 289 707 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 673 221 707 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 861 221 895 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nand4bb_2
rlabel metal1 s 0 -48 1196 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 1943734
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1933346
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 29.900 0.000 
<< end >>
