magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 182 157 456 203
rect 1 21 456 157
rect 30 -17 64 21
<< locali >>
rect 288 401 354 493
rect 288 367 443 401
rect 30 153 69 265
rect 173 153 255 265
rect 357 165 443 367
rect 304 131 443 165
rect 304 77 338 131
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 31 333 103 368
rect 220 367 254 527
rect 388 435 422 527
rect 31 299 323 333
rect 103 119 139 299
rect 289 199 323 299
rect 21 17 69 119
rect 103 51 161 119
rect 207 17 270 119
rect 372 17 438 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 173 153 255 265 6 A
port 1 nsew signal input
rlabel locali s 30 153 69 265 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 460 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 456 157 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 182 157 456 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 304 77 338 131 6 X
port 7 nsew signal output
rlabel locali s 304 131 443 165 6 X
port 7 nsew signal output
rlabel locali s 357 165 443 367 6 X
port 7 nsew signal output
rlabel locali s 288 367 443 401 6 X
port 7 nsew signal output
rlabel locali s 288 401 354 493 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 460 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 988668
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 984310
<< end >>
