magic
tech sky130B
magscale 1 2
timestamp 1666464484
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_0
timestamp 1666464484
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_1
timestamp 1666464484
transform 1 0 296 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808370  sky130_fd_pr__hvdfl1sd__example_55959141808370_0
timestamp 1666464484
transform -1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 30055428
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30053790
<< end >>
