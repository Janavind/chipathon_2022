magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< pwell >>
rect 10 10 806 392
<< nmoslvt >>
rect 92 36 122 366
rect 178 36 208 366
rect 264 36 294 366
rect 350 36 380 366
rect 436 36 466 366
rect 522 36 552 366
rect 608 36 638 366
rect 694 36 724 366
<< ndiff >>
rect 36 329 92 366
rect 36 295 47 329
rect 81 295 92 329
rect 36 257 92 295
rect 36 223 47 257
rect 81 223 92 257
rect 36 185 92 223
rect 36 151 47 185
rect 81 151 92 185
rect 36 113 92 151
rect 36 79 47 113
rect 81 79 92 113
rect 36 36 92 79
rect 122 329 178 366
rect 122 295 133 329
rect 167 295 178 329
rect 122 257 178 295
rect 122 223 133 257
rect 167 223 178 257
rect 122 185 178 223
rect 122 151 133 185
rect 167 151 178 185
rect 122 113 178 151
rect 122 79 133 113
rect 167 79 178 113
rect 122 36 178 79
rect 208 329 264 366
rect 208 295 219 329
rect 253 295 264 329
rect 208 257 264 295
rect 208 223 219 257
rect 253 223 264 257
rect 208 185 264 223
rect 208 151 219 185
rect 253 151 264 185
rect 208 113 264 151
rect 208 79 219 113
rect 253 79 264 113
rect 208 36 264 79
rect 294 329 350 366
rect 294 295 305 329
rect 339 295 350 329
rect 294 257 350 295
rect 294 223 305 257
rect 339 223 350 257
rect 294 185 350 223
rect 294 151 305 185
rect 339 151 350 185
rect 294 113 350 151
rect 294 79 305 113
rect 339 79 350 113
rect 294 36 350 79
rect 380 329 436 366
rect 380 295 391 329
rect 425 295 436 329
rect 380 257 436 295
rect 380 223 391 257
rect 425 223 436 257
rect 380 185 436 223
rect 380 151 391 185
rect 425 151 436 185
rect 380 113 436 151
rect 380 79 391 113
rect 425 79 436 113
rect 380 36 436 79
rect 466 329 522 366
rect 466 295 477 329
rect 511 295 522 329
rect 466 257 522 295
rect 466 223 477 257
rect 511 223 522 257
rect 466 185 522 223
rect 466 151 477 185
rect 511 151 522 185
rect 466 113 522 151
rect 466 79 477 113
rect 511 79 522 113
rect 466 36 522 79
rect 552 329 608 366
rect 552 295 563 329
rect 597 295 608 329
rect 552 257 608 295
rect 552 223 563 257
rect 597 223 608 257
rect 552 185 608 223
rect 552 151 563 185
rect 597 151 608 185
rect 552 113 608 151
rect 552 79 563 113
rect 597 79 608 113
rect 552 36 608 79
rect 638 329 694 366
rect 638 295 649 329
rect 683 295 694 329
rect 638 257 694 295
rect 638 223 649 257
rect 683 223 694 257
rect 638 185 694 223
rect 638 151 649 185
rect 683 151 694 185
rect 638 113 694 151
rect 638 79 649 113
rect 683 79 694 113
rect 638 36 694 79
rect 724 329 780 366
rect 724 295 735 329
rect 769 295 780 329
rect 724 257 780 295
rect 724 223 735 257
rect 769 223 780 257
rect 724 185 780 223
rect 724 151 735 185
rect 769 151 780 185
rect 724 113 780 151
rect 724 79 735 113
rect 769 79 780 113
rect 724 36 780 79
<< ndiffc >>
rect 47 295 81 329
rect 47 223 81 257
rect 47 151 81 185
rect 47 79 81 113
rect 133 295 167 329
rect 133 223 167 257
rect 133 151 167 185
rect 133 79 167 113
rect 219 295 253 329
rect 219 223 253 257
rect 219 151 253 185
rect 219 79 253 113
rect 305 295 339 329
rect 305 223 339 257
rect 305 151 339 185
rect 305 79 339 113
rect 391 295 425 329
rect 391 223 425 257
rect 391 151 425 185
rect 391 79 425 113
rect 477 295 511 329
rect 477 223 511 257
rect 477 151 511 185
rect 477 79 511 113
rect 563 295 597 329
rect 563 223 597 257
rect 563 151 597 185
rect 563 79 597 113
rect 649 295 683 329
rect 649 223 683 257
rect 649 151 683 185
rect 649 79 683 113
rect 735 295 769 329
rect 735 223 769 257
rect 735 151 769 185
rect 735 79 769 113
<< poly >>
rect 92 447 724 463
rect 92 413 153 447
rect 187 413 221 447
rect 255 413 289 447
rect 323 413 357 447
rect 391 413 425 447
rect 459 413 493 447
rect 527 413 561 447
rect 595 413 629 447
rect 663 413 724 447
rect 92 392 724 413
rect 92 366 122 392
rect 178 366 208 392
rect 264 366 294 392
rect 350 366 380 392
rect 436 366 466 392
rect 522 366 552 392
rect 608 366 638 392
rect 694 366 724 392
rect 92 10 122 36
rect 178 10 208 36
rect 264 10 294 36
rect 350 10 380 36
rect 436 10 466 36
rect 522 10 552 36
rect 608 10 638 36
rect 694 10 724 36
<< polycont >>
rect 153 413 187 447
rect 221 413 255 447
rect 289 413 323 447
rect 357 413 391 447
rect 425 413 459 447
rect 493 413 527 447
rect 561 413 595 447
rect 629 413 663 447
<< locali >>
rect 137 447 679 463
rect 137 413 139 447
rect 187 413 211 447
rect 255 413 283 447
rect 323 413 355 447
rect 391 413 425 447
rect 461 413 493 447
rect 533 413 561 447
rect 605 413 629 447
rect 677 413 679 447
rect 137 397 679 413
rect 47 329 81 357
rect 47 257 81 295
rect 47 185 81 223
rect 47 113 81 151
rect 47 51 81 79
rect 133 329 167 357
rect 133 257 167 295
rect 133 185 167 223
rect 133 113 167 151
rect 133 51 167 79
rect 219 329 253 357
rect 219 257 253 295
rect 219 185 253 223
rect 219 113 253 151
rect 219 51 253 79
rect 305 329 339 357
rect 305 257 339 295
rect 305 185 339 223
rect 305 113 339 151
rect 305 51 339 79
rect 391 329 425 357
rect 391 257 425 295
rect 391 185 425 223
rect 391 113 425 151
rect 391 51 425 79
rect 477 329 511 357
rect 477 257 511 295
rect 477 185 511 223
rect 477 113 511 151
rect 477 51 511 79
rect 563 329 597 357
rect 563 257 597 295
rect 563 185 597 223
rect 563 113 597 151
rect 563 51 597 79
rect 649 329 683 357
rect 649 257 683 295
rect 649 185 683 223
rect 649 113 683 151
rect 649 51 683 79
rect 735 329 769 357
rect 735 257 769 295
rect 735 185 769 223
rect 735 113 769 151
rect 735 51 769 79
<< viali >>
rect 139 413 153 447
rect 153 413 173 447
rect 211 413 221 447
rect 221 413 245 447
rect 283 413 289 447
rect 289 413 317 447
rect 355 413 357 447
rect 357 413 389 447
rect 427 413 459 447
rect 459 413 461 447
rect 499 413 527 447
rect 527 413 533 447
rect 571 413 595 447
rect 595 413 605 447
rect 643 413 663 447
rect 663 413 677 447
rect 47 295 81 329
rect 47 223 81 257
rect 47 151 81 185
rect 47 79 81 113
rect 133 295 167 329
rect 133 223 167 257
rect 133 151 167 185
rect 133 79 167 113
rect 219 295 253 329
rect 219 223 253 257
rect 219 151 253 185
rect 219 79 253 113
rect 305 295 339 329
rect 305 223 339 257
rect 305 151 339 185
rect 305 79 339 113
rect 391 295 425 329
rect 391 223 425 257
rect 391 151 425 185
rect 391 79 425 113
rect 477 295 511 329
rect 477 223 511 257
rect 477 151 511 185
rect 477 79 511 113
rect 563 295 597 329
rect 563 223 597 257
rect 563 151 597 185
rect 563 79 597 113
rect 649 295 683 329
rect 649 223 683 257
rect 649 151 683 185
rect 649 79 683 113
rect 735 295 769 329
rect 735 223 769 257
rect 735 151 769 185
rect 735 79 769 113
<< metal1 >>
rect 127 447 689 459
rect 127 413 139 447
rect 173 413 211 447
rect 245 413 283 447
rect 317 413 355 447
rect 389 413 427 447
rect 461 413 499 447
rect 533 413 571 447
rect 605 413 643 447
rect 677 413 689 447
rect 127 401 689 413
rect 41 329 87 357
rect 41 295 47 329
rect 81 295 87 329
rect 41 257 87 295
rect 41 223 47 257
rect 81 223 87 257
rect 41 185 87 223
rect 41 151 47 185
rect 81 151 87 185
rect 41 113 87 151
rect 41 79 47 113
rect 81 79 87 113
rect 41 -29 87 79
rect 124 338 176 357
rect 124 274 176 286
rect 124 185 176 222
rect 124 151 133 185
rect 167 151 176 185
rect 124 113 176 151
rect 124 79 133 113
rect 167 79 176 113
rect 124 51 176 79
rect 213 329 259 357
rect 213 295 219 329
rect 253 295 259 329
rect 213 257 259 295
rect 213 223 219 257
rect 253 223 259 257
rect 213 185 259 223
rect 213 151 219 185
rect 253 151 259 185
rect 213 113 259 151
rect 213 79 219 113
rect 253 79 259 113
rect 213 -29 259 79
rect 296 338 348 357
rect 296 274 348 286
rect 296 185 348 222
rect 296 151 305 185
rect 339 151 348 185
rect 296 113 348 151
rect 296 79 305 113
rect 339 79 348 113
rect 296 51 348 79
rect 385 329 431 357
rect 385 295 391 329
rect 425 295 431 329
rect 385 257 431 295
rect 385 223 391 257
rect 425 223 431 257
rect 385 185 431 223
rect 385 151 391 185
rect 425 151 431 185
rect 385 113 431 151
rect 385 79 391 113
rect 425 79 431 113
rect 385 -29 431 79
rect 468 338 520 357
rect 468 274 520 286
rect 468 185 520 222
rect 468 151 477 185
rect 511 151 520 185
rect 468 113 520 151
rect 468 79 477 113
rect 511 79 520 113
rect 468 51 520 79
rect 557 329 603 357
rect 557 295 563 329
rect 597 295 603 329
rect 557 257 603 295
rect 557 223 563 257
rect 597 223 603 257
rect 557 185 603 223
rect 557 151 563 185
rect 597 151 603 185
rect 557 113 603 151
rect 557 79 563 113
rect 597 79 603 113
rect 557 -29 603 79
rect 640 338 692 357
rect 640 274 692 286
rect 640 185 692 222
rect 640 151 649 185
rect 683 151 692 185
rect 640 113 692 151
rect 640 79 649 113
rect 683 79 692 113
rect 640 51 692 79
rect 729 329 775 357
rect 729 295 735 329
rect 769 295 775 329
rect 729 257 775 295
rect 729 223 735 257
rect 769 223 775 257
rect 729 185 775 223
rect 729 151 735 185
rect 769 151 775 185
rect 729 113 775 151
rect 729 79 735 113
rect 769 79 775 113
rect 729 -29 775 79
rect 41 -89 775 -29
<< via1 >>
rect 124 329 176 338
rect 124 295 133 329
rect 133 295 167 329
rect 167 295 176 329
rect 124 286 176 295
rect 124 257 176 274
rect 124 223 133 257
rect 133 223 167 257
rect 167 223 176 257
rect 124 222 176 223
rect 296 329 348 338
rect 296 295 305 329
rect 305 295 339 329
rect 339 295 348 329
rect 296 286 348 295
rect 296 257 348 274
rect 296 223 305 257
rect 305 223 339 257
rect 339 223 348 257
rect 296 222 348 223
rect 468 329 520 338
rect 468 295 477 329
rect 477 295 511 329
rect 511 295 520 329
rect 468 286 520 295
rect 468 257 520 274
rect 468 223 477 257
rect 477 223 511 257
rect 511 223 520 257
rect 468 222 520 223
rect 640 329 692 338
rect 640 295 649 329
rect 649 295 683 329
rect 683 295 692 329
rect 640 286 692 295
rect 640 257 692 274
rect 640 223 649 257
rect 649 223 683 257
rect 683 223 692 257
rect 640 222 692 223
<< metal2 >>
rect 117 348 183 357
rect 117 292 122 348
rect 178 292 183 348
rect 117 286 124 292
rect 176 286 183 292
rect 117 274 183 286
rect 117 268 124 274
rect 176 268 183 274
rect 117 212 122 268
rect 178 212 183 268
rect 117 203 183 212
rect 289 348 355 357
rect 289 292 294 348
rect 350 292 355 348
rect 289 286 296 292
rect 348 286 355 292
rect 289 274 355 286
rect 289 268 296 274
rect 348 268 355 274
rect 289 212 294 268
rect 350 212 355 268
rect 289 203 355 212
rect 461 348 527 357
rect 461 292 466 348
rect 522 292 527 348
rect 461 286 468 292
rect 520 286 527 292
rect 461 274 527 286
rect 461 268 468 274
rect 520 268 527 274
rect 461 212 466 268
rect 522 212 527 268
rect 461 203 527 212
rect 633 348 699 357
rect 633 292 638 348
rect 694 292 699 348
rect 633 286 640 292
rect 692 286 699 292
rect 633 274 699 286
rect 633 268 640 274
rect 692 268 699 274
rect 633 212 638 268
rect 694 212 699 268
rect 633 203 699 212
<< via2 >>
rect 122 338 178 348
rect 122 292 124 338
rect 124 292 176 338
rect 176 292 178 338
rect 122 222 124 268
rect 124 222 176 268
rect 176 222 178 268
rect 122 212 178 222
rect 294 338 350 348
rect 294 292 296 338
rect 296 292 348 338
rect 348 292 350 338
rect 294 222 296 268
rect 296 222 348 268
rect 348 222 350 268
rect 294 212 350 222
rect 466 338 522 348
rect 466 292 468 338
rect 468 292 520 338
rect 520 292 522 338
rect 466 222 468 268
rect 468 222 520 268
rect 520 222 522 268
rect 466 212 522 222
rect 638 338 694 348
rect 638 292 640 338
rect 640 292 692 338
rect 692 292 694 338
rect 638 222 640 268
rect 640 222 692 268
rect 692 222 694 268
rect 638 212 694 222
<< metal3 >>
rect 117 348 699 357
rect 117 292 122 348
rect 178 292 294 348
rect 350 292 466 348
rect 522 292 638 348
rect 694 292 699 348
rect 117 291 699 292
rect 117 268 183 291
rect 117 212 122 268
rect 178 212 183 268
rect 117 203 183 212
rect 289 268 355 291
rect 289 212 294 268
rect 350 212 355 268
rect 289 203 355 212
rect 461 268 527 291
rect 461 212 466 268
rect 522 212 527 268
rect 461 203 527 212
rect 633 268 699 291
rect 633 212 638 268
rect 694 212 699 268
rect 633 203 699 212
<< labels >>
flabel metal3 s 117 291 699 357 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 127 401 689 459 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel metal1 s 41 -89 775 -29 0 FreeSans 400 0 0 0 SOURCE
port 3 nsew
flabel pwell s 78 371 89 386 0 FreeSans 200 0 0 0 SUBSTRATE
port 4 nsew
<< properties >>
string GDS_END 3349294
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 3335312
string path 14.500 8.925 14.500 -2.225 
<< end >>
