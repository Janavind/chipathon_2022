magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1103 203
rect 29 -17 63 21
<< locali >>
rect 121 333 173 493
rect 307 333 345 493
rect 479 333 515 493
rect 763 333 801 421
rect 121 299 801 333
rect 17 215 85 271
rect 121 181 173 299
rect 209 215 358 265
rect 440 215 637 265
rect 673 215 891 265
rect 927 215 1087 265
rect 121 123 187 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 35 305 85 527
rect 207 367 273 527
rect 379 368 445 527
rect 551 367 617 527
rect 662 455 900 493
rect 662 367 714 455
rect 848 337 900 455
rect 934 371 986 527
rect 1020 337 1072 493
rect 848 303 1072 337
rect 35 89 87 173
rect 223 147 455 181
rect 223 89 260 147
rect 385 124 455 147
rect 490 131 1087 168
rect 35 52 260 89
rect 294 106 352 113
rect 294 89 355 106
rect 576 89 642 97
rect 294 51 642 89
rect 676 73 714 131
rect 848 130 1087 131
rect 748 17 814 97
rect 848 73 886 130
rect 920 17 986 96
rect 1020 73 1087 130
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 927 215 1087 265 6 A1
port 1 nsew signal input
rlabel locali s 673 215 891 265 6 A2
port 2 nsew signal input
rlabel locali s 440 215 637 265 6 B1
port 3 nsew signal input
rlabel locali s 209 215 358 265 6 C1
port 4 nsew signal input
rlabel locali s 17 215 85 271 6 D1
port 5 nsew signal input
rlabel metal1 s 0 -48 1104 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 1103 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 121 123 187 181 6 Y
port 10 nsew signal output
rlabel locali s 121 181 173 299 6 Y
port 10 nsew signal output
rlabel locali s 121 299 801 333 6 Y
port 10 nsew signal output
rlabel locali s 763 333 801 421 6 Y
port 10 nsew signal output
rlabel locali s 479 333 515 493 6 Y
port 10 nsew signal output
rlabel locali s 307 333 345 493 6 Y
port 10 nsew signal output
rlabel locali s 121 333 173 493 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 960620
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 951156
<< end >>
