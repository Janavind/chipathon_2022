magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -42 415 710 1116
<< pwell >>
rect 40 118 494 310
<< mvnmos >>
rect 119 144 239 284
rect 295 144 415 284
<< mvpmos >>
rect 119 750 239 950
rect 295 750 415 950
rect 471 750 591 950
rect 119 482 239 682
rect 295 482 415 682
rect 471 482 591 682
<< mvndiff >>
rect 66 272 119 284
rect 66 238 74 272
rect 108 238 119 272
rect 66 204 119 238
rect 66 170 74 204
rect 108 170 119 204
rect 66 144 119 170
rect 239 144 295 284
rect 415 272 468 284
rect 415 238 426 272
rect 460 238 468 272
rect 415 204 468 238
rect 415 170 426 204
rect 460 170 468 204
rect 415 144 468 170
<< mvpdiff >>
rect 66 932 119 950
rect 66 898 74 932
rect 108 898 119 932
rect 66 864 119 898
rect 66 830 74 864
rect 108 830 119 864
rect 66 796 119 830
rect 66 762 74 796
rect 108 762 119 796
rect 66 750 119 762
rect 239 932 295 950
rect 239 898 250 932
rect 284 898 295 932
rect 239 864 295 898
rect 239 830 250 864
rect 284 830 295 864
rect 239 796 295 830
rect 239 762 250 796
rect 284 762 295 796
rect 239 750 295 762
rect 415 932 471 950
rect 415 898 426 932
rect 460 898 471 932
rect 415 864 471 898
rect 415 830 426 864
rect 460 830 471 864
rect 415 796 471 830
rect 415 762 426 796
rect 460 762 471 796
rect 415 750 471 762
rect 591 932 644 950
rect 591 898 602 932
rect 636 898 644 932
rect 591 864 644 898
rect 591 830 602 864
rect 636 830 644 864
rect 591 796 644 830
rect 591 762 602 796
rect 636 762 644 796
rect 591 750 644 762
rect 66 670 119 682
rect 66 636 74 670
rect 108 636 119 670
rect 66 602 119 636
rect 66 568 74 602
rect 108 568 119 602
rect 66 534 119 568
rect 66 500 74 534
rect 108 500 119 534
rect 66 482 119 500
rect 239 670 295 682
rect 239 636 250 670
rect 284 636 295 670
rect 239 602 295 636
rect 239 568 250 602
rect 284 568 295 602
rect 239 534 295 568
rect 239 500 250 534
rect 284 500 295 534
rect 239 482 295 500
rect 415 670 471 682
rect 415 636 426 670
rect 460 636 471 670
rect 415 602 471 636
rect 415 568 426 602
rect 460 568 471 602
rect 415 534 471 568
rect 415 500 426 534
rect 460 500 471 534
rect 415 482 471 500
rect 591 670 644 682
rect 591 636 602 670
rect 636 636 644 670
rect 591 602 644 636
rect 591 568 602 602
rect 636 568 644 602
rect 591 534 644 568
rect 591 500 602 534
rect 636 500 644 534
rect 591 482 644 500
<< mvndiffc >>
rect 74 238 108 272
rect 74 170 108 204
rect 426 238 460 272
rect 426 170 460 204
<< mvpdiffc >>
rect 74 898 108 932
rect 74 830 108 864
rect 74 762 108 796
rect 250 898 284 932
rect 250 830 284 864
rect 250 762 284 796
rect 426 898 460 932
rect 426 830 460 864
rect 426 762 460 796
rect 602 898 636 932
rect 602 830 636 864
rect 602 762 636 796
rect 74 636 108 670
rect 74 568 108 602
rect 74 500 108 534
rect 250 636 284 670
rect 250 568 284 602
rect 250 500 284 534
rect 426 636 460 670
rect 426 568 460 602
rect 426 500 460 534
rect 602 636 636 670
rect 602 568 636 602
rect 602 500 636 534
<< poly >>
rect 119 950 239 976
rect 295 950 415 976
rect 471 950 591 976
rect 119 682 239 750
rect 295 682 415 750
rect 471 682 591 750
rect 119 434 239 482
rect 119 400 165 434
rect 199 400 239 434
rect 119 366 239 400
rect 119 332 165 366
rect 199 332 239 366
rect 119 284 239 332
rect 295 434 415 482
rect 295 400 336 434
rect 370 400 415 434
rect 295 366 415 400
rect 295 332 336 366
rect 370 332 415 366
rect 295 284 415 332
rect 471 434 591 482
rect 471 400 517 434
rect 551 400 591 434
rect 471 366 591 400
rect 471 332 517 366
rect 551 332 591 366
rect 471 316 591 332
rect 119 118 239 144
rect 295 118 415 144
<< polycont >>
rect 165 400 199 434
rect 165 332 199 366
rect 336 400 370 434
rect 336 332 370 366
rect 517 400 551 434
rect 517 332 551 366
<< locali >>
rect 74 932 108 944
rect 74 864 108 872
rect 74 796 108 830
rect 74 670 108 762
rect 74 602 108 636
rect 74 534 108 568
rect 74 484 108 500
rect 250 932 284 950
rect 250 864 284 898
rect 250 796 284 830
rect 250 670 284 762
rect 250 602 284 636
rect 250 534 284 568
rect 149 400 165 434
rect 199 400 215 434
rect 149 366 215 400
rect 149 332 165 366
rect 199 332 215 366
rect 74 272 108 288
rect 74 227 108 238
rect 250 261 284 500
rect 426 932 460 944
rect 426 864 460 872
rect 426 796 460 830
rect 426 670 460 762
rect 426 602 460 636
rect 426 534 460 568
rect 426 484 460 500
rect 602 932 636 948
rect 602 864 636 898
rect 602 796 636 830
rect 602 670 636 762
rect 602 602 636 636
rect 602 534 636 568
rect 320 400 336 434
rect 370 400 386 434
rect 320 366 386 400
rect 320 332 336 366
rect 370 332 386 366
rect 501 400 517 434
rect 551 400 567 434
rect 501 366 567 400
rect 501 332 517 366
rect 551 332 567 366
rect 426 272 460 288
rect 250 238 426 261
rect 602 238 636 500
rect 250 227 636 238
rect 74 155 108 170
rect 421 204 636 227
rect 421 170 426 204
rect 421 154 460 170
<< viali >>
rect 74 944 108 978
rect 74 898 108 906
rect 74 872 108 898
rect 426 944 460 978
rect 426 898 460 906
rect 426 872 460 898
rect 74 204 108 227
rect 74 193 108 204
rect 74 121 108 155
<< metal1 >>
rect 25 978 644 1062
rect 25 944 74 978
rect 108 944 426 978
rect 460 944 644 978
rect 25 906 644 944
rect 25 872 74 906
rect 108 872 426 906
rect 460 872 644 906
rect 25 859 644 872
rect 24 227 503 239
rect 24 193 74 227
rect 108 193 503 227
rect 24 155 503 193
rect 24 121 74 155
rect 108 121 503 155
rect 24 24 503 121
use sky130_fd_pr__nfet_01v8__example_559591418087  sky130_fd_pr__nfet_01v8__example_559591418087_0
timestamp 1666199351
transform 1 0 295 0 -1 284
box 120 0 121 1
use sky130_fd_pr__nfet_01v8__example_559591418089  sky130_fd_pr__nfet_01v8__example_559591418089_0
timestamp 1666199351
transform 1 0 119 0 -1 284
box -1 0 0 1
use sky130_fd_pr__pfet_01v8__example_559591418085  sky130_fd_pr__pfet_01v8__example_559591418085_0
timestamp 1666199351
transform 1 0 119 0 1 750
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_559591418085  sky130_fd_pr__pfet_01v8__example_559591418085_1
timestamp 1666199351
transform 1 0 295 0 1 750
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_559591418085  sky130_fd_pr__pfet_01v8__example_559591418085_2
timestamp 1666199351
transform 1 0 119 0 -1 682
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_559591418085  sky130_fd_pr__pfet_01v8__example_559591418085_3
timestamp 1666199351
transform 1 0 471 0 -1 682
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_559591418085  sky130_fd_pr__pfet_01v8__example_559591418085_4
timestamp 1666199351
transform 1 0 471 0 1 750
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_559591418085  sky130_fd_pr__pfet_01v8__example_559591418085_5
timestamp 1666199351
transform 1 0 295 0 -1 682
box -1 0 121 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1666199351
transform 0 -1 108 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1666199351
transform 0 -1 460 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1666199351
transform 0 -1 108 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1666199351
transform 0 -1 567 1 0 316
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1666199351
transform 0 -1 386 1 0 316
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_2
timestamp 1666199351
transform 0 -1 215 1 0 316
box 0 0 1 1
<< labels >>
flabel locali s 321 352 383 391 0 FreeSans 400 0 0 0 IN1
port 1 nsew
flabel locali s 156 353 207 394 0 FreeSans 400 0 0 0 IN0
port 2 nsew
flabel locali s 250 256 284 532 0 FreeSans 200 0 0 0 OUT
port 3 nsew
flabel metal1 s 24 24 107 238 0 FreeSans 320 0 0 0 VGND
port 4 nsew
flabel metal1 s 561 859 644 1062 0 FreeSans 320 0 0 0 VPWR
port 5 nsew
<< properties >>
string GDS_END 31883450
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31880436
<< end >>
