magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< dnwell >>
rect 20601 -14836 22062 -7928
<< nwell >>
rect 0 0 6792 494
rect 20750 -4052 21244 -3320
rect 20403 -7832 20707 -7470
rect 20403 -8134 22147 -7832
rect 20403 -14630 20707 -8134
rect 21845 -14630 22147 -8134
rect 20403 -14932 22147 -14630
rect 20403 -17308 20707 -14932
<< pwell >>
rect 21007 -8369 21785 -8215
rect 21007 -9914 21161 -8369
rect 21631 -9914 21785 -8369
rect 21007 -10566 21785 -9914
rect 21007 -14416 21161 -10566
rect 21631 -14416 21785 -10566
rect 21007 -14570 21785 -14416
<< mvnmos >>
rect 21268 -10540 21368 -9940
rect 21424 -10540 21524 -9940
<< mvpmos >>
rect 66 275 1066 375
rect 1198 275 2198 375
rect 2330 275 3330 375
rect 3462 275 4462 375
rect 4594 275 5594 375
rect 5726 275 6726 375
rect 66 119 1066 219
rect 1198 119 2198 219
rect 2330 119 3330 219
rect 3462 119 4462 219
rect 4594 119 5594 219
rect 5726 119 6726 219
rect 20869 -3986 20969 -3386
rect 21025 -3986 21125 -3386
<< mvndiff >>
rect 21215 -10018 21268 -9940
rect 21215 -10052 21223 -10018
rect 21257 -10052 21268 -10018
rect 21215 -10086 21268 -10052
rect 21215 -10120 21223 -10086
rect 21257 -10120 21268 -10086
rect 21215 -10154 21268 -10120
rect 21215 -10188 21223 -10154
rect 21257 -10188 21268 -10154
rect 21215 -10222 21268 -10188
rect 21215 -10256 21223 -10222
rect 21257 -10256 21268 -10222
rect 21215 -10290 21268 -10256
rect 21215 -10324 21223 -10290
rect 21257 -10324 21268 -10290
rect 21215 -10358 21268 -10324
rect 21215 -10392 21223 -10358
rect 21257 -10392 21268 -10358
rect 21215 -10426 21268 -10392
rect 21215 -10460 21223 -10426
rect 21257 -10460 21268 -10426
rect 21215 -10494 21268 -10460
rect 21215 -10528 21223 -10494
rect 21257 -10528 21268 -10494
rect 21215 -10540 21268 -10528
rect 21368 -10018 21424 -9940
rect 21368 -10052 21379 -10018
rect 21413 -10052 21424 -10018
rect 21368 -10086 21424 -10052
rect 21368 -10120 21379 -10086
rect 21413 -10120 21424 -10086
rect 21368 -10154 21424 -10120
rect 21368 -10188 21379 -10154
rect 21413 -10188 21424 -10154
rect 21368 -10222 21424 -10188
rect 21368 -10256 21379 -10222
rect 21413 -10256 21424 -10222
rect 21368 -10290 21424 -10256
rect 21368 -10324 21379 -10290
rect 21413 -10324 21424 -10290
rect 21368 -10358 21424 -10324
rect 21368 -10392 21379 -10358
rect 21413 -10392 21424 -10358
rect 21368 -10426 21424 -10392
rect 21368 -10460 21379 -10426
rect 21413 -10460 21424 -10426
rect 21368 -10494 21424 -10460
rect 21368 -10528 21379 -10494
rect 21413 -10528 21424 -10494
rect 21368 -10540 21424 -10528
rect 21524 -10018 21577 -9940
rect 21524 -10052 21535 -10018
rect 21569 -10052 21577 -10018
rect 21524 -10086 21577 -10052
rect 21524 -10120 21535 -10086
rect 21569 -10120 21577 -10086
rect 21524 -10154 21577 -10120
rect 21524 -10188 21535 -10154
rect 21569 -10188 21577 -10154
rect 21524 -10222 21577 -10188
rect 21524 -10256 21535 -10222
rect 21569 -10256 21577 -10222
rect 21524 -10290 21577 -10256
rect 21524 -10324 21535 -10290
rect 21569 -10324 21577 -10290
rect 21524 -10358 21577 -10324
rect 21524 -10392 21535 -10358
rect 21569 -10392 21577 -10358
rect 21524 -10426 21577 -10392
rect 21524 -10460 21535 -10426
rect 21569 -10460 21577 -10426
rect 21524 -10494 21577 -10460
rect 21524 -10528 21535 -10494
rect 21569 -10528 21577 -10494
rect 21524 -10540 21577 -10528
<< mvpdiff >>
rect 66 420 1066 428
rect 66 386 136 420
rect 170 386 204 420
rect 238 386 272 420
rect 306 386 340 420
rect 374 386 408 420
rect 442 386 476 420
rect 510 386 544 420
rect 578 386 612 420
rect 646 386 680 420
rect 714 386 748 420
rect 782 386 816 420
rect 850 386 884 420
rect 918 386 952 420
rect 986 386 1020 420
rect 1054 386 1066 420
rect 66 375 1066 386
rect 1198 420 2198 428
rect 1198 386 1210 420
rect 1244 386 1278 420
rect 1312 386 1346 420
rect 1380 386 1414 420
rect 1448 386 1482 420
rect 1516 386 1550 420
rect 1584 386 1618 420
rect 1652 386 1686 420
rect 1720 386 1754 420
rect 1788 386 1822 420
rect 1856 386 1890 420
rect 1924 386 1958 420
rect 1992 386 2026 420
rect 2060 386 2094 420
rect 2128 386 2198 420
rect 1198 375 2198 386
rect 2330 420 3330 428
rect 2330 386 2400 420
rect 2434 386 2468 420
rect 2502 386 2536 420
rect 2570 386 2604 420
rect 2638 386 2672 420
rect 2706 386 2740 420
rect 2774 386 2808 420
rect 2842 386 2876 420
rect 2910 386 2944 420
rect 2978 386 3012 420
rect 3046 386 3080 420
rect 3114 386 3148 420
rect 3182 386 3216 420
rect 3250 386 3284 420
rect 3318 386 3330 420
rect 2330 375 3330 386
rect 3462 420 4462 428
rect 3462 386 3474 420
rect 3508 386 3542 420
rect 3576 386 3610 420
rect 3644 386 3678 420
rect 3712 386 3746 420
rect 3780 386 3814 420
rect 3848 386 3882 420
rect 3916 386 3950 420
rect 3984 386 4018 420
rect 4052 386 4086 420
rect 4120 386 4154 420
rect 4188 386 4222 420
rect 4256 386 4290 420
rect 4324 386 4358 420
rect 4392 386 4462 420
rect 3462 375 4462 386
rect 4594 420 5594 428
rect 4594 386 4664 420
rect 4698 386 4732 420
rect 4766 386 4800 420
rect 4834 386 4868 420
rect 4902 386 4936 420
rect 4970 386 5004 420
rect 5038 386 5072 420
rect 5106 386 5140 420
rect 5174 386 5208 420
rect 5242 386 5276 420
rect 5310 386 5344 420
rect 5378 386 5412 420
rect 5446 386 5480 420
rect 5514 386 5548 420
rect 5582 386 5594 420
rect 4594 375 5594 386
rect 5726 420 6726 428
rect 5726 386 5738 420
rect 5772 386 5806 420
rect 5840 386 5874 420
rect 5908 386 5942 420
rect 5976 386 6010 420
rect 6044 386 6078 420
rect 6112 386 6146 420
rect 6180 386 6214 420
rect 6248 386 6282 420
rect 6316 386 6350 420
rect 6384 386 6418 420
rect 6452 386 6486 420
rect 6520 386 6554 420
rect 6588 386 6622 420
rect 6656 386 6726 420
rect 5726 375 6726 386
rect 66 264 1066 275
rect 66 230 136 264
rect 170 230 204 264
rect 238 230 272 264
rect 306 230 340 264
rect 374 230 408 264
rect 442 230 476 264
rect 510 230 544 264
rect 578 230 612 264
rect 646 230 680 264
rect 714 230 748 264
rect 782 230 816 264
rect 850 230 884 264
rect 918 230 952 264
rect 986 230 1020 264
rect 1054 230 1066 264
rect 66 219 1066 230
rect 1198 264 2198 275
rect 1198 230 1210 264
rect 1244 230 1278 264
rect 1312 230 1346 264
rect 1380 230 1414 264
rect 1448 230 1482 264
rect 1516 230 1550 264
rect 1584 230 1618 264
rect 1652 230 1686 264
rect 1720 230 1754 264
rect 1788 230 1822 264
rect 1856 230 1890 264
rect 1924 230 1958 264
rect 1992 230 2026 264
rect 2060 230 2094 264
rect 2128 230 2198 264
rect 1198 219 2198 230
rect 2330 264 3330 275
rect 2330 230 2400 264
rect 2434 230 2468 264
rect 2502 230 2536 264
rect 2570 230 2604 264
rect 2638 230 2672 264
rect 2706 230 2740 264
rect 2774 230 2808 264
rect 2842 230 2876 264
rect 2910 230 2944 264
rect 2978 230 3012 264
rect 3046 230 3080 264
rect 3114 230 3148 264
rect 3182 230 3216 264
rect 3250 230 3284 264
rect 3318 230 3330 264
rect 2330 219 3330 230
rect 3462 264 4462 275
rect 3462 230 3474 264
rect 3508 230 3542 264
rect 3576 230 3610 264
rect 3644 230 3678 264
rect 3712 230 3746 264
rect 3780 230 3814 264
rect 3848 230 3882 264
rect 3916 230 3950 264
rect 3984 230 4018 264
rect 4052 230 4086 264
rect 4120 230 4154 264
rect 4188 230 4222 264
rect 4256 230 4290 264
rect 4324 230 4358 264
rect 4392 230 4462 264
rect 3462 219 4462 230
rect 4594 264 5594 275
rect 4594 230 4664 264
rect 4698 230 4732 264
rect 4766 230 4800 264
rect 4834 230 4868 264
rect 4902 230 4936 264
rect 4970 230 5004 264
rect 5038 230 5072 264
rect 5106 230 5140 264
rect 5174 230 5208 264
rect 5242 230 5276 264
rect 5310 230 5344 264
rect 5378 230 5412 264
rect 5446 230 5480 264
rect 5514 230 5548 264
rect 5582 230 5594 264
rect 4594 219 5594 230
rect 5726 264 6726 275
rect 5726 230 5738 264
rect 5772 230 5806 264
rect 5840 230 5874 264
rect 5908 230 5942 264
rect 5976 230 6010 264
rect 6044 230 6078 264
rect 6112 230 6146 264
rect 6180 230 6214 264
rect 6248 230 6282 264
rect 6316 230 6350 264
rect 6384 230 6418 264
rect 6452 230 6486 264
rect 6520 230 6554 264
rect 6588 230 6622 264
rect 6656 230 6726 264
rect 5726 219 6726 230
rect 66 108 1066 119
rect 66 74 136 108
rect 170 74 204 108
rect 238 74 272 108
rect 306 74 340 108
rect 374 74 408 108
rect 442 74 476 108
rect 510 74 544 108
rect 578 74 612 108
rect 646 74 680 108
rect 714 74 748 108
rect 782 74 816 108
rect 850 74 884 108
rect 918 74 952 108
rect 986 74 1020 108
rect 1054 74 1066 108
rect 66 66 1066 74
rect 1198 108 2198 119
rect 1198 74 1210 108
rect 1244 74 1278 108
rect 1312 74 1346 108
rect 1380 74 1414 108
rect 1448 74 1482 108
rect 1516 74 1550 108
rect 1584 74 1618 108
rect 1652 74 1686 108
rect 1720 74 1754 108
rect 1788 74 1822 108
rect 1856 74 1890 108
rect 1924 74 1958 108
rect 1992 74 2026 108
rect 2060 74 2094 108
rect 2128 74 2198 108
rect 1198 66 2198 74
rect 2330 108 3330 119
rect 2330 74 2400 108
rect 2434 74 2468 108
rect 2502 74 2536 108
rect 2570 74 2604 108
rect 2638 74 2672 108
rect 2706 74 2740 108
rect 2774 74 2808 108
rect 2842 74 2876 108
rect 2910 74 2944 108
rect 2978 74 3012 108
rect 3046 74 3080 108
rect 3114 74 3148 108
rect 3182 74 3216 108
rect 3250 74 3284 108
rect 3318 74 3330 108
rect 2330 66 3330 74
rect 3462 108 4462 119
rect 3462 74 3474 108
rect 3508 74 3542 108
rect 3576 74 3610 108
rect 3644 74 3678 108
rect 3712 74 3746 108
rect 3780 74 3814 108
rect 3848 74 3882 108
rect 3916 74 3950 108
rect 3984 74 4018 108
rect 4052 74 4086 108
rect 4120 74 4154 108
rect 4188 74 4222 108
rect 4256 74 4290 108
rect 4324 74 4358 108
rect 4392 74 4462 108
rect 3462 66 4462 74
rect 4594 108 5594 119
rect 4594 74 4664 108
rect 4698 74 4732 108
rect 4766 74 4800 108
rect 4834 74 4868 108
rect 4902 74 4936 108
rect 4970 74 5004 108
rect 5038 74 5072 108
rect 5106 74 5140 108
rect 5174 74 5208 108
rect 5242 74 5276 108
rect 5310 74 5344 108
rect 5378 74 5412 108
rect 5446 74 5480 108
rect 5514 74 5548 108
rect 5582 74 5594 108
rect 4594 66 5594 74
rect 5726 108 6726 119
rect 5726 74 5738 108
rect 5772 74 5806 108
rect 5840 74 5874 108
rect 5908 74 5942 108
rect 5976 74 6010 108
rect 6044 74 6078 108
rect 6112 74 6146 108
rect 6180 74 6214 108
rect 6248 74 6282 108
rect 6316 74 6350 108
rect 6384 74 6418 108
rect 6452 74 6486 108
rect 6520 74 6554 108
rect 6588 74 6622 108
rect 6656 74 6726 108
rect 5726 66 6726 74
rect 20816 -3464 20869 -3386
rect 20816 -3498 20824 -3464
rect 20858 -3498 20869 -3464
rect 20816 -3532 20869 -3498
rect 20816 -3566 20824 -3532
rect 20858 -3566 20869 -3532
rect 20816 -3600 20869 -3566
rect 20816 -3634 20824 -3600
rect 20858 -3634 20869 -3600
rect 20816 -3668 20869 -3634
rect 20816 -3702 20824 -3668
rect 20858 -3702 20869 -3668
rect 20816 -3736 20869 -3702
rect 20816 -3770 20824 -3736
rect 20858 -3770 20869 -3736
rect 20816 -3804 20869 -3770
rect 20816 -3838 20824 -3804
rect 20858 -3838 20869 -3804
rect 20816 -3872 20869 -3838
rect 20816 -3906 20824 -3872
rect 20858 -3906 20869 -3872
rect 20816 -3940 20869 -3906
rect 20816 -3974 20824 -3940
rect 20858 -3974 20869 -3940
rect 20816 -3986 20869 -3974
rect 20969 -3464 21025 -3386
rect 20969 -3498 20980 -3464
rect 21014 -3498 21025 -3464
rect 20969 -3532 21025 -3498
rect 20969 -3566 20980 -3532
rect 21014 -3566 21025 -3532
rect 20969 -3600 21025 -3566
rect 20969 -3634 20980 -3600
rect 21014 -3634 21025 -3600
rect 20969 -3668 21025 -3634
rect 20969 -3702 20980 -3668
rect 21014 -3702 21025 -3668
rect 20969 -3736 21025 -3702
rect 20969 -3770 20980 -3736
rect 21014 -3770 21025 -3736
rect 20969 -3804 21025 -3770
rect 20969 -3838 20980 -3804
rect 21014 -3838 21025 -3804
rect 20969 -3872 21025 -3838
rect 20969 -3906 20980 -3872
rect 21014 -3906 21025 -3872
rect 20969 -3940 21025 -3906
rect 20969 -3974 20980 -3940
rect 21014 -3974 21025 -3940
rect 20969 -3986 21025 -3974
rect 21125 -3464 21178 -3386
rect 21125 -3498 21136 -3464
rect 21170 -3498 21178 -3464
rect 21125 -3532 21178 -3498
rect 21125 -3566 21136 -3532
rect 21170 -3566 21178 -3532
rect 21125 -3600 21178 -3566
rect 21125 -3634 21136 -3600
rect 21170 -3634 21178 -3600
rect 21125 -3668 21178 -3634
rect 21125 -3702 21136 -3668
rect 21170 -3702 21178 -3668
rect 21125 -3736 21178 -3702
rect 21125 -3770 21136 -3736
rect 21170 -3770 21178 -3736
rect 21125 -3804 21178 -3770
rect 21125 -3838 21136 -3804
rect 21170 -3838 21178 -3804
rect 21125 -3872 21178 -3838
rect 21125 -3906 21136 -3872
rect 21170 -3906 21178 -3872
rect 21125 -3940 21178 -3906
rect 21125 -3974 21136 -3940
rect 21170 -3974 21178 -3940
rect 21125 -3986 21178 -3974
<< mvndiffc >>
rect 21223 -10052 21257 -10018
rect 21223 -10120 21257 -10086
rect 21223 -10188 21257 -10154
rect 21223 -10256 21257 -10222
rect 21223 -10324 21257 -10290
rect 21223 -10392 21257 -10358
rect 21223 -10460 21257 -10426
rect 21223 -10528 21257 -10494
rect 21379 -10052 21413 -10018
rect 21379 -10120 21413 -10086
rect 21379 -10188 21413 -10154
rect 21379 -10256 21413 -10222
rect 21379 -10324 21413 -10290
rect 21379 -10392 21413 -10358
rect 21379 -10460 21413 -10426
rect 21379 -10528 21413 -10494
rect 21535 -10052 21569 -10018
rect 21535 -10120 21569 -10086
rect 21535 -10188 21569 -10154
rect 21535 -10256 21569 -10222
rect 21535 -10324 21569 -10290
rect 21535 -10392 21569 -10358
rect 21535 -10460 21569 -10426
rect 21535 -10528 21569 -10494
<< mvpdiffc >>
rect 136 386 170 420
rect 204 386 238 420
rect 272 386 306 420
rect 340 386 374 420
rect 408 386 442 420
rect 476 386 510 420
rect 544 386 578 420
rect 612 386 646 420
rect 680 386 714 420
rect 748 386 782 420
rect 816 386 850 420
rect 884 386 918 420
rect 952 386 986 420
rect 1020 386 1054 420
rect 1210 386 1244 420
rect 1278 386 1312 420
rect 1346 386 1380 420
rect 1414 386 1448 420
rect 1482 386 1516 420
rect 1550 386 1584 420
rect 1618 386 1652 420
rect 1686 386 1720 420
rect 1754 386 1788 420
rect 1822 386 1856 420
rect 1890 386 1924 420
rect 1958 386 1992 420
rect 2026 386 2060 420
rect 2094 386 2128 420
rect 2400 386 2434 420
rect 2468 386 2502 420
rect 2536 386 2570 420
rect 2604 386 2638 420
rect 2672 386 2706 420
rect 2740 386 2774 420
rect 2808 386 2842 420
rect 2876 386 2910 420
rect 2944 386 2978 420
rect 3012 386 3046 420
rect 3080 386 3114 420
rect 3148 386 3182 420
rect 3216 386 3250 420
rect 3284 386 3318 420
rect 3474 386 3508 420
rect 3542 386 3576 420
rect 3610 386 3644 420
rect 3678 386 3712 420
rect 3746 386 3780 420
rect 3814 386 3848 420
rect 3882 386 3916 420
rect 3950 386 3984 420
rect 4018 386 4052 420
rect 4086 386 4120 420
rect 4154 386 4188 420
rect 4222 386 4256 420
rect 4290 386 4324 420
rect 4358 386 4392 420
rect 4664 386 4698 420
rect 4732 386 4766 420
rect 4800 386 4834 420
rect 4868 386 4902 420
rect 4936 386 4970 420
rect 5004 386 5038 420
rect 5072 386 5106 420
rect 5140 386 5174 420
rect 5208 386 5242 420
rect 5276 386 5310 420
rect 5344 386 5378 420
rect 5412 386 5446 420
rect 5480 386 5514 420
rect 5548 386 5582 420
rect 5738 386 5772 420
rect 5806 386 5840 420
rect 5874 386 5908 420
rect 5942 386 5976 420
rect 6010 386 6044 420
rect 6078 386 6112 420
rect 6146 386 6180 420
rect 6214 386 6248 420
rect 6282 386 6316 420
rect 6350 386 6384 420
rect 6418 386 6452 420
rect 6486 386 6520 420
rect 6554 386 6588 420
rect 6622 386 6656 420
rect 136 230 170 264
rect 204 230 238 264
rect 272 230 306 264
rect 340 230 374 264
rect 408 230 442 264
rect 476 230 510 264
rect 544 230 578 264
rect 612 230 646 264
rect 680 230 714 264
rect 748 230 782 264
rect 816 230 850 264
rect 884 230 918 264
rect 952 230 986 264
rect 1020 230 1054 264
rect 1210 230 1244 264
rect 1278 230 1312 264
rect 1346 230 1380 264
rect 1414 230 1448 264
rect 1482 230 1516 264
rect 1550 230 1584 264
rect 1618 230 1652 264
rect 1686 230 1720 264
rect 1754 230 1788 264
rect 1822 230 1856 264
rect 1890 230 1924 264
rect 1958 230 1992 264
rect 2026 230 2060 264
rect 2094 230 2128 264
rect 2400 230 2434 264
rect 2468 230 2502 264
rect 2536 230 2570 264
rect 2604 230 2638 264
rect 2672 230 2706 264
rect 2740 230 2774 264
rect 2808 230 2842 264
rect 2876 230 2910 264
rect 2944 230 2978 264
rect 3012 230 3046 264
rect 3080 230 3114 264
rect 3148 230 3182 264
rect 3216 230 3250 264
rect 3284 230 3318 264
rect 3474 230 3508 264
rect 3542 230 3576 264
rect 3610 230 3644 264
rect 3678 230 3712 264
rect 3746 230 3780 264
rect 3814 230 3848 264
rect 3882 230 3916 264
rect 3950 230 3984 264
rect 4018 230 4052 264
rect 4086 230 4120 264
rect 4154 230 4188 264
rect 4222 230 4256 264
rect 4290 230 4324 264
rect 4358 230 4392 264
rect 4664 230 4698 264
rect 4732 230 4766 264
rect 4800 230 4834 264
rect 4868 230 4902 264
rect 4936 230 4970 264
rect 5004 230 5038 264
rect 5072 230 5106 264
rect 5140 230 5174 264
rect 5208 230 5242 264
rect 5276 230 5310 264
rect 5344 230 5378 264
rect 5412 230 5446 264
rect 5480 230 5514 264
rect 5548 230 5582 264
rect 5738 230 5772 264
rect 5806 230 5840 264
rect 5874 230 5908 264
rect 5942 230 5976 264
rect 6010 230 6044 264
rect 6078 230 6112 264
rect 6146 230 6180 264
rect 6214 230 6248 264
rect 6282 230 6316 264
rect 6350 230 6384 264
rect 6418 230 6452 264
rect 6486 230 6520 264
rect 6554 230 6588 264
rect 6622 230 6656 264
rect 136 74 170 108
rect 204 74 238 108
rect 272 74 306 108
rect 340 74 374 108
rect 408 74 442 108
rect 476 74 510 108
rect 544 74 578 108
rect 612 74 646 108
rect 680 74 714 108
rect 748 74 782 108
rect 816 74 850 108
rect 884 74 918 108
rect 952 74 986 108
rect 1020 74 1054 108
rect 1210 74 1244 108
rect 1278 74 1312 108
rect 1346 74 1380 108
rect 1414 74 1448 108
rect 1482 74 1516 108
rect 1550 74 1584 108
rect 1618 74 1652 108
rect 1686 74 1720 108
rect 1754 74 1788 108
rect 1822 74 1856 108
rect 1890 74 1924 108
rect 1958 74 1992 108
rect 2026 74 2060 108
rect 2094 74 2128 108
rect 2400 74 2434 108
rect 2468 74 2502 108
rect 2536 74 2570 108
rect 2604 74 2638 108
rect 2672 74 2706 108
rect 2740 74 2774 108
rect 2808 74 2842 108
rect 2876 74 2910 108
rect 2944 74 2978 108
rect 3012 74 3046 108
rect 3080 74 3114 108
rect 3148 74 3182 108
rect 3216 74 3250 108
rect 3284 74 3318 108
rect 3474 74 3508 108
rect 3542 74 3576 108
rect 3610 74 3644 108
rect 3678 74 3712 108
rect 3746 74 3780 108
rect 3814 74 3848 108
rect 3882 74 3916 108
rect 3950 74 3984 108
rect 4018 74 4052 108
rect 4086 74 4120 108
rect 4154 74 4188 108
rect 4222 74 4256 108
rect 4290 74 4324 108
rect 4358 74 4392 108
rect 4664 74 4698 108
rect 4732 74 4766 108
rect 4800 74 4834 108
rect 4868 74 4902 108
rect 4936 74 4970 108
rect 5004 74 5038 108
rect 5072 74 5106 108
rect 5140 74 5174 108
rect 5208 74 5242 108
rect 5276 74 5310 108
rect 5344 74 5378 108
rect 5412 74 5446 108
rect 5480 74 5514 108
rect 5548 74 5582 108
rect 5738 74 5772 108
rect 5806 74 5840 108
rect 5874 74 5908 108
rect 5942 74 5976 108
rect 6010 74 6044 108
rect 6078 74 6112 108
rect 6146 74 6180 108
rect 6214 74 6248 108
rect 6282 74 6316 108
rect 6350 74 6384 108
rect 6418 74 6452 108
rect 6486 74 6520 108
rect 6554 74 6588 108
rect 6622 74 6656 108
rect 20824 -3498 20858 -3464
rect 20824 -3566 20858 -3532
rect 20824 -3634 20858 -3600
rect 20824 -3702 20858 -3668
rect 20824 -3770 20858 -3736
rect 20824 -3838 20858 -3804
rect 20824 -3906 20858 -3872
rect 20824 -3974 20858 -3940
rect 20980 -3498 21014 -3464
rect 20980 -3566 21014 -3532
rect 20980 -3634 21014 -3600
rect 20980 -3702 21014 -3668
rect 20980 -3770 21014 -3736
rect 20980 -3838 21014 -3804
rect 20980 -3906 21014 -3872
rect 20980 -3974 21014 -3940
rect 21136 -3498 21170 -3464
rect 21136 -3566 21170 -3532
rect 21136 -3634 21170 -3600
rect 21136 -3702 21170 -3668
rect 21136 -3770 21170 -3736
rect 21136 -3838 21170 -3804
rect 21136 -3906 21170 -3872
rect 21136 -3974 21170 -3940
<< psubdiff >>
rect 21033 -8275 21113 -8241
rect 21147 -8275 21181 -8241
rect 21033 -8309 21181 -8275
rect 21135 -8343 21181 -8309
rect 21691 -8322 21759 -8241
rect 21691 -8343 21725 -8322
rect 21657 -8356 21725 -8343
rect 21657 -8390 21759 -8356
rect 21033 -14429 21135 -14395
rect 21067 -14442 21135 -14429
rect 21067 -14463 21101 -14442
rect 21033 -14544 21101 -14463
rect 21543 -14476 21657 -14442
rect 21543 -14510 21759 -14476
rect 21543 -14544 21649 -14510
rect 21683 -14544 21759 -14510
<< mvnsubdiff >>
rect 20470 -7504 20640 -7470
rect 20504 -7538 20538 -7504
rect 20572 -7538 20606 -7504
rect 20470 -7573 20640 -7538
rect 20504 -7607 20538 -7573
rect 20572 -7607 20606 -7573
rect 20470 -7642 20640 -7607
rect 20504 -7676 20538 -7642
rect 20572 -7676 20606 -7642
rect 20470 -7711 20640 -7676
rect 20504 -7745 20538 -7711
rect 20572 -7745 20606 -7711
rect 20470 -7780 20640 -7745
rect 20504 -7814 20538 -7780
rect 20572 -7814 20606 -7780
rect 20470 -7849 20640 -7814
rect 20504 -7883 20538 -7849
rect 20572 -7883 20606 -7849
rect 20470 -7898 20640 -7883
rect 20470 -7918 20674 -7898
rect 20504 -7952 20538 -7918
rect 20572 -7952 20606 -7918
rect 20640 -7952 20674 -7918
rect 20470 -7987 20674 -7952
rect 20504 -8021 20538 -7987
rect 20572 -8021 20606 -7987
rect 20640 -8021 20674 -7987
rect 21116 -7932 21151 -7898
rect 21185 -7932 21220 -7898
rect 21254 -7932 21289 -7898
rect 21323 -7932 21358 -7898
rect 21392 -7932 21427 -7898
rect 21461 -7932 21496 -7898
rect 21530 -7932 21565 -7898
rect 21599 -7932 21634 -7898
rect 21668 -7932 21703 -7898
rect 21737 -7932 21772 -7898
rect 21806 -7932 21841 -7898
rect 21875 -7932 21910 -7898
rect 21944 -7932 21979 -7898
rect 22013 -7932 22081 -7898
rect 21116 -7966 22081 -7932
rect 21116 -8000 21151 -7966
rect 21185 -8000 21220 -7966
rect 21254 -8000 21289 -7966
rect 21323 -8000 21358 -7966
rect 21392 -8000 21427 -7966
rect 21461 -8000 21496 -7966
rect 21530 -8000 21565 -7966
rect 21599 -8000 21634 -7966
rect 21668 -8000 21703 -7966
rect 21737 -8000 21772 -7966
rect 21806 -8000 21841 -7966
rect 21875 -8000 21910 -7966
rect 21944 -8000 21979 -7966
rect 20470 -8056 20674 -8021
rect 20504 -8090 20538 -8056
rect 20572 -8090 20606 -8056
rect 20640 -8068 20674 -8056
rect 21048 -8034 21979 -8000
rect 21048 -8068 21083 -8034
rect 21117 -8068 21152 -8034
rect 21186 -8068 21221 -8034
rect 21255 -8068 21290 -8034
rect 21324 -8068 21359 -8034
rect 21393 -8068 21428 -8034
rect 21462 -8068 21497 -8034
rect 21531 -8068 21566 -8034
rect 21600 -8068 21635 -8034
rect 21669 -8068 21704 -8034
rect 21738 -8068 21773 -8034
rect 21807 -8068 21842 -8034
rect 21876 -8068 21911 -8034
rect 20470 -8125 20640 -8090
rect 20504 -8159 20538 -8125
rect 20572 -8159 20606 -8125
rect 20470 -8194 20640 -8159
rect 20504 -8228 20538 -8194
rect 20572 -8228 20606 -8194
rect 20470 -8263 20640 -8228
rect 20504 -8297 20538 -8263
rect 20572 -8297 20606 -8263
rect 20470 -8332 20640 -8297
rect 21911 -10211 21979 -10176
rect 21945 -10244 21979 -10211
rect 21945 -10245 22081 -10244
rect 21911 -10279 22081 -10245
rect 21911 -10280 21979 -10279
rect 21945 -10313 21979 -10280
rect 22013 -10313 22047 -10279
rect 21945 -10314 22081 -10313
rect 21911 -10348 22081 -10314
rect 21911 -10349 21979 -10348
rect 21945 -10382 21979 -10349
rect 22013 -10382 22047 -10348
rect 21945 -10383 22081 -10382
rect 21911 -10417 22081 -10383
rect 21911 -10418 21979 -10417
rect 21945 -10451 21979 -10418
rect 22013 -10451 22047 -10417
rect 21945 -10452 22081 -10451
rect 21911 -10486 22081 -10452
rect 21911 -10487 21979 -10486
rect 21945 -10520 21979 -10487
rect 22013 -10520 22047 -10486
rect 21945 -10521 22081 -10520
rect 21911 -10555 22081 -10521
rect 21911 -10556 21979 -10555
rect 21945 -10589 21979 -10556
rect 22013 -10589 22047 -10555
rect 21945 -10590 22081 -10589
rect 21911 -10624 22081 -10590
rect 21911 -10625 21979 -10624
rect 21945 -10658 21979 -10625
rect 22013 -10658 22047 -10624
rect 21945 -10659 22081 -10658
rect 21911 -10693 22081 -10659
rect 21911 -10694 21979 -10693
rect 21945 -10727 21979 -10694
rect 22013 -10727 22047 -10693
rect 21945 -10728 22081 -10727
rect 21911 -10762 22081 -10728
rect 21911 -10763 21979 -10762
rect 21945 -10796 21979 -10763
rect 22013 -10796 22047 -10762
rect 21945 -10797 22081 -10796
rect 21911 -10831 22081 -10797
rect 21911 -10832 21979 -10831
rect 21945 -10865 21979 -10832
rect 22013 -10865 22047 -10831
rect 21945 -10866 22081 -10865
rect 21911 -10900 22081 -10866
rect 21911 -10901 21979 -10900
rect 21945 -10934 21979 -10901
rect 22013 -10934 22047 -10900
rect 21945 -10935 22081 -10934
rect 21911 -10969 22081 -10935
rect 21911 -10970 21979 -10969
rect 21945 -11003 21979 -10970
rect 22013 -11003 22047 -10969
rect 21945 -11004 22081 -11003
rect 21911 -11038 22081 -11004
rect 21911 -11039 21979 -11038
rect 21945 -11072 21979 -11039
rect 22013 -11072 22047 -11038
rect 21945 -11073 22081 -11072
rect 21911 -11107 22081 -11073
rect 21911 -11108 21979 -11107
rect 21945 -11141 21979 -11108
rect 22013 -11141 22047 -11107
rect 21945 -11142 22081 -11141
rect 21911 -11176 22081 -11142
rect 21911 -11177 21979 -11176
rect 21945 -11210 21979 -11177
rect 22013 -11210 22047 -11176
rect 21945 -11211 22081 -11210
rect 21911 -11245 22081 -11211
rect 21911 -11246 21979 -11245
rect 21945 -11279 21979 -11246
rect 22013 -11279 22047 -11245
rect 21945 -11280 22081 -11279
rect 21911 -11314 22081 -11280
rect 21911 -11315 21979 -11314
rect 21945 -11348 21979 -11315
rect 22013 -11348 22047 -11314
rect 21945 -11349 22081 -11348
rect 21911 -11383 22081 -11349
rect 21911 -11384 21979 -11383
rect 21945 -11417 21979 -11384
rect 22013 -11417 22047 -11383
rect 21945 -11418 22081 -11417
rect 21911 -11452 22081 -11418
rect 21911 -11453 21979 -11452
rect 21945 -11486 21979 -11453
rect 22013 -11486 22047 -11452
rect 21945 -11487 22081 -11486
rect 21911 -11521 22081 -11487
rect 21911 -11522 21979 -11521
rect 21945 -11555 21979 -11522
rect 22013 -11555 22047 -11521
rect 21945 -11556 22081 -11555
rect 21911 -11590 22081 -11556
rect 21911 -11591 21979 -11590
rect 21945 -11624 21979 -11591
rect 22013 -11624 22047 -11590
rect 21945 -11625 22081 -11624
rect 21911 -11659 22081 -11625
rect 21911 -11660 21979 -11659
rect 21945 -11693 21979 -11660
rect 22013 -11693 22047 -11659
rect 21945 -11694 22081 -11693
rect 21911 -11728 22081 -11694
rect 21911 -11729 21979 -11728
rect 21945 -11762 21979 -11729
rect 22013 -11762 22047 -11728
rect 21945 -11763 22081 -11762
rect 21911 -11797 22081 -11763
rect 21911 -11798 21979 -11797
rect 21945 -11831 21979 -11798
rect 22013 -11831 22047 -11797
rect 21945 -11832 22081 -11831
rect 21911 -11866 22081 -11832
rect 21911 -11867 21979 -11866
rect 21945 -11900 21979 -11867
rect 22013 -11900 22047 -11866
rect 21945 -11901 22081 -11900
rect 21911 -11935 22081 -11901
rect 21911 -11936 21979 -11935
rect 21945 -11969 21979 -11936
rect 22013 -11969 22047 -11935
rect 21945 -11970 22081 -11969
rect 21911 -12004 22081 -11970
rect 21911 -12005 21979 -12004
rect 21945 -12038 21979 -12005
rect 22013 -12038 22047 -12004
rect 21945 -12039 22081 -12038
rect 21911 -12073 22081 -12039
rect 21911 -12074 21979 -12073
rect 21945 -12107 21979 -12074
rect 22013 -12107 22047 -12073
rect 21945 -12108 22081 -12107
rect 21911 -12142 22081 -12108
rect 21911 -12143 21979 -12142
rect 21945 -12176 21979 -12143
rect 22013 -12176 22047 -12142
rect 21945 -12177 22081 -12176
rect 21911 -12211 22081 -12177
rect 21911 -12212 21979 -12211
rect 21945 -12245 21979 -12212
rect 22013 -12245 22047 -12211
rect 21945 -12246 22081 -12245
rect 21911 -12280 22081 -12246
rect 21911 -12281 21979 -12280
rect 21945 -12314 21979 -12281
rect 22013 -12314 22047 -12280
rect 21945 -12315 22081 -12314
rect 21911 -12349 22081 -12315
rect 21911 -12350 21979 -12349
rect 21945 -12383 21979 -12350
rect 22013 -12383 22047 -12349
rect 21945 -12384 22081 -12383
rect 21911 -12418 22081 -12384
rect 21911 -12419 21979 -12418
rect 21945 -12452 21979 -12419
rect 22013 -12452 22047 -12418
rect 21945 -12453 22081 -12452
rect 21911 -12487 22081 -12453
rect 21911 -12488 21979 -12487
rect 21945 -12521 21979 -12488
rect 22013 -12521 22047 -12487
rect 21945 -12522 22081 -12521
rect 21911 -12556 22081 -12522
rect 21911 -12557 21979 -12556
rect 21945 -12590 21979 -12557
rect 22013 -12590 22047 -12556
rect 21945 -12591 22081 -12590
rect 21911 -12625 22081 -12591
rect 21911 -12626 21979 -12625
rect 21945 -12659 21979 -12626
rect 22013 -12659 22047 -12625
rect 21945 -12660 22081 -12659
rect 21911 -12694 22081 -12660
rect 21911 -12695 21979 -12694
rect 21945 -12728 21979 -12695
rect 22013 -12728 22047 -12694
rect 21945 -12729 22081 -12728
rect 21911 -12763 22081 -12729
rect 21911 -12764 21979 -12763
rect 21945 -12797 21979 -12764
rect 22013 -12797 22047 -12763
rect 21945 -12798 22081 -12797
rect 21911 -12832 22081 -12798
rect 21911 -12833 21979 -12832
rect 21945 -12866 21979 -12833
rect 22013 -12866 22047 -12832
rect 21945 -12867 22081 -12866
rect 21911 -12901 22081 -12867
rect 21911 -12902 21979 -12901
rect 21945 -12935 21979 -12902
rect 22013 -12935 22047 -12901
rect 21945 -12936 22081 -12935
rect 21911 -12970 22081 -12936
rect 21911 -12971 21979 -12970
rect 21945 -13004 21979 -12971
rect 22013 -13004 22047 -12970
rect 21945 -13005 22081 -13004
rect 21911 -13039 22081 -13005
rect 21911 -13040 21979 -13039
rect 21945 -13073 21979 -13040
rect 22013 -13073 22047 -13039
rect 21945 -13074 22081 -13073
rect 21911 -13108 22081 -13074
rect 21911 -13109 21979 -13108
rect 21945 -13142 21979 -13109
rect 22013 -13142 22047 -13108
rect 21945 -13143 22081 -13142
rect 21911 -13177 22081 -13143
rect 21911 -13178 21979 -13177
rect 21945 -13211 21979 -13178
rect 22013 -13211 22047 -13177
rect 21945 -13212 22081 -13211
rect 21911 -13246 22081 -13212
rect 21911 -13247 21979 -13246
rect 21945 -13280 21979 -13247
rect 22013 -13280 22047 -13246
rect 21945 -13281 22081 -13280
rect 21911 -13315 22081 -13281
rect 21911 -13316 21979 -13315
rect 21945 -13349 21979 -13316
rect 22013 -13349 22047 -13315
rect 21945 -13350 22081 -13349
rect 21911 -13384 22081 -13350
rect 21911 -13385 21979 -13384
rect 21945 -13418 21979 -13385
rect 22013 -13418 22047 -13384
rect 21945 -13419 22081 -13418
rect 21911 -13453 22081 -13419
rect 21911 -13454 21979 -13453
rect 21945 -13487 21979 -13454
rect 22013 -13487 22047 -13453
rect 21945 -13488 22081 -13487
rect 21911 -13522 22081 -13488
rect 21911 -13523 21979 -13522
rect 21945 -13556 21979 -13523
rect 22013 -13556 22047 -13522
rect 21945 -13557 22081 -13556
rect 21911 -13591 22081 -13557
rect 21911 -13592 21979 -13591
rect 21945 -13625 21979 -13592
rect 22013 -13625 22047 -13591
rect 21945 -13626 22081 -13625
rect 21911 -13660 22081 -13626
rect 21911 -13661 21979 -13660
rect 21945 -13694 21979 -13661
rect 22013 -13694 22047 -13660
rect 21945 -13695 22081 -13694
rect 21911 -13729 22081 -13695
rect 21911 -13730 21979 -13729
rect 21945 -13763 21979 -13730
rect 22013 -13763 22047 -13729
rect 21945 -13764 22081 -13763
rect 21911 -13798 22081 -13764
rect 21911 -13799 21979 -13798
rect 21945 -13832 21979 -13799
rect 22013 -13832 22047 -13798
rect 21945 -13833 22081 -13832
rect 21911 -13867 22081 -13833
rect 21911 -13868 21979 -13867
rect 21945 -13901 21979 -13868
rect 22013 -13901 22047 -13867
rect 21945 -13902 22081 -13901
rect 21911 -13936 22081 -13902
rect 21911 -13937 21979 -13936
rect 21945 -13970 21979 -13937
rect 22013 -13970 22047 -13936
rect 21945 -13971 22081 -13970
rect 21911 -14005 22081 -13971
rect 21911 -14006 21979 -14005
rect 21945 -14039 21979 -14006
rect 22013 -14039 22047 -14005
rect 21945 -14040 22081 -14039
rect 21911 -14074 22081 -14040
rect 21911 -14075 21979 -14074
rect 21945 -14108 21979 -14075
rect 22013 -14108 22047 -14074
rect 21945 -14109 22081 -14108
rect 21911 -14143 22081 -14109
rect 21911 -14144 21979 -14143
rect 21945 -14177 21979 -14144
rect 22013 -14177 22047 -14143
rect 21945 -14178 22081 -14177
rect 21911 -14212 22081 -14178
rect 21911 -14213 21979 -14212
rect 21945 -14246 21979 -14213
rect 22013 -14246 22047 -14212
rect 21945 -14247 22081 -14246
rect 21911 -14281 22081 -14247
rect 21911 -14282 21979 -14281
rect 21945 -14315 21979 -14282
rect 22013 -14315 22047 -14281
rect 21945 -14316 22081 -14315
rect 21911 -14350 22081 -14316
rect 21911 -14351 21979 -14350
rect 21945 -14384 21979 -14351
rect 22013 -14384 22047 -14350
rect 21945 -14385 22081 -14384
rect 21911 -14419 22081 -14385
rect 21911 -14420 21979 -14419
rect 21945 -14453 21979 -14420
rect 22013 -14453 22047 -14419
rect 21945 -14454 22081 -14453
rect 21911 -14488 22081 -14454
rect 21911 -14489 21979 -14488
rect 21945 -14522 21979 -14489
rect 22013 -14522 22047 -14488
rect 21945 -14523 22081 -14522
rect 21911 -14557 22081 -14523
rect 21911 -14558 21979 -14557
rect 21945 -14591 21979 -14558
rect 22013 -14591 22047 -14557
rect 21945 -14592 22081 -14591
rect 21911 -14626 22081 -14592
rect 21911 -14627 21979 -14626
rect 21945 -14660 21979 -14627
rect 22013 -14660 22047 -14626
rect 21945 -14661 22081 -14660
rect 21911 -14695 22081 -14661
rect 21911 -14696 21979 -14695
rect 20708 -14730 20743 -14696
rect 20777 -14730 20812 -14696
rect 20846 -14730 20881 -14696
rect 20915 -14730 20950 -14696
rect 20984 -14730 21019 -14696
rect 21053 -14730 21088 -14696
rect 21122 -14730 21157 -14696
rect 21191 -14730 21226 -14696
rect 21260 -14730 21295 -14696
rect 21329 -14730 21364 -14696
rect 21398 -14730 21433 -14696
rect 21467 -14730 21502 -14696
rect 21536 -14730 21571 -14696
rect 20708 -14764 21571 -14730
rect 21945 -14729 21979 -14696
rect 22013 -14729 22047 -14695
rect 21945 -14764 22081 -14729
rect 20708 -14798 20743 -14764
rect 20777 -14798 20812 -14764
rect 20846 -14798 20881 -14764
rect 20915 -14798 20950 -14764
rect 20984 -14798 21019 -14764
rect 21053 -14798 21088 -14764
rect 21122 -14798 21157 -14764
rect 21191 -14798 21226 -14764
rect 21260 -14798 21295 -14764
rect 21329 -14798 21364 -14764
rect 21398 -14798 21433 -14764
rect 21467 -14798 21502 -14764
rect 21536 -14798 21571 -14764
rect 20708 -14832 21571 -14798
rect 20708 -14866 20743 -14832
rect 20777 -14866 20812 -14832
rect 20846 -14866 20881 -14832
rect 20915 -14866 20950 -14832
rect 20984 -14866 21019 -14832
rect 21053 -14866 21088 -14832
rect 21122 -14866 21157 -14832
rect 21191 -14866 21226 -14832
rect 21260 -14866 21295 -14832
rect 21329 -14866 21364 -14832
rect 21398 -14866 21433 -14832
rect 21467 -14866 21502 -14832
rect 21536 -14866 21571 -14832
rect 22013 -14798 22047 -14764
rect 22013 -14866 22081 -14798
rect 20470 -17308 20640 -17274
<< psubdiffcont >>
rect 21113 -8275 21147 -8241
rect 21033 -14395 21135 -8309
rect 21181 -8343 21691 -8241
rect 21725 -8356 21759 -8322
rect 21033 -14463 21067 -14429
rect 21101 -14544 21543 -14442
rect 21657 -14476 21759 -8390
rect 21649 -14544 21683 -14510
<< mvnsubdiffcont >>
rect 20470 -7538 20504 -7504
rect 20538 -7538 20572 -7504
rect 20606 -7538 20640 -7504
rect 20470 -7607 20504 -7573
rect 20538 -7607 20572 -7573
rect 20606 -7607 20640 -7573
rect 20470 -7676 20504 -7642
rect 20538 -7676 20572 -7642
rect 20606 -7676 20640 -7642
rect 20470 -7745 20504 -7711
rect 20538 -7745 20572 -7711
rect 20606 -7745 20640 -7711
rect 20470 -7814 20504 -7780
rect 20538 -7814 20572 -7780
rect 20606 -7814 20640 -7780
rect 20470 -7883 20504 -7849
rect 20538 -7883 20572 -7849
rect 20606 -7883 20640 -7849
rect 20470 -7952 20504 -7918
rect 20538 -7952 20572 -7918
rect 20606 -7952 20640 -7918
rect 20470 -8021 20504 -7987
rect 20538 -8021 20572 -7987
rect 20606 -8021 20640 -7987
rect 20674 -8000 21116 -7898
rect 21151 -7932 21185 -7898
rect 21220 -7932 21254 -7898
rect 21289 -7932 21323 -7898
rect 21358 -7932 21392 -7898
rect 21427 -7932 21461 -7898
rect 21496 -7932 21530 -7898
rect 21565 -7932 21599 -7898
rect 21634 -7932 21668 -7898
rect 21703 -7932 21737 -7898
rect 21772 -7932 21806 -7898
rect 21841 -7932 21875 -7898
rect 21910 -7932 21944 -7898
rect 21979 -7932 22013 -7898
rect 21151 -8000 21185 -7966
rect 21220 -8000 21254 -7966
rect 21289 -8000 21323 -7966
rect 21358 -8000 21392 -7966
rect 21427 -8000 21461 -7966
rect 21496 -8000 21530 -7966
rect 21565 -8000 21599 -7966
rect 21634 -8000 21668 -7966
rect 21703 -8000 21737 -7966
rect 21772 -8000 21806 -7966
rect 21841 -8000 21875 -7966
rect 21910 -8000 21944 -7966
rect 20470 -8090 20504 -8056
rect 20538 -8090 20572 -8056
rect 20606 -8090 20640 -8056
rect 20674 -8068 21048 -8000
rect 21979 -8034 22081 -7966
rect 21083 -8068 21117 -8034
rect 21152 -8068 21186 -8034
rect 21221 -8068 21255 -8034
rect 21290 -8068 21324 -8034
rect 21359 -8068 21393 -8034
rect 21428 -8068 21462 -8034
rect 21497 -8068 21531 -8034
rect 21566 -8068 21600 -8034
rect 21635 -8068 21669 -8034
rect 21704 -8068 21738 -8034
rect 21773 -8068 21807 -8034
rect 21842 -8068 21876 -8034
rect 20470 -8159 20504 -8125
rect 20538 -8159 20572 -8125
rect 20606 -8159 20640 -8125
rect 20470 -8228 20504 -8194
rect 20538 -8228 20572 -8194
rect 20606 -8228 20640 -8194
rect 20470 -8297 20504 -8263
rect 20538 -8297 20572 -8263
rect 20606 -8297 20640 -8263
rect 20470 -14696 20640 -8332
rect 21911 -10176 22081 -8034
rect 21911 -10245 21945 -10211
rect 21979 -10244 22081 -10176
rect 21911 -10314 21945 -10280
rect 21979 -10313 22013 -10279
rect 22047 -10313 22081 -10279
rect 21911 -10383 21945 -10349
rect 21979 -10382 22013 -10348
rect 22047 -10382 22081 -10348
rect 21911 -10452 21945 -10418
rect 21979 -10451 22013 -10417
rect 22047 -10451 22081 -10417
rect 21911 -10521 21945 -10487
rect 21979 -10520 22013 -10486
rect 22047 -10520 22081 -10486
rect 21911 -10590 21945 -10556
rect 21979 -10589 22013 -10555
rect 22047 -10589 22081 -10555
rect 21911 -10659 21945 -10625
rect 21979 -10658 22013 -10624
rect 22047 -10658 22081 -10624
rect 21911 -10728 21945 -10694
rect 21979 -10727 22013 -10693
rect 22047 -10727 22081 -10693
rect 21911 -10797 21945 -10763
rect 21979 -10796 22013 -10762
rect 22047 -10796 22081 -10762
rect 21911 -10866 21945 -10832
rect 21979 -10865 22013 -10831
rect 22047 -10865 22081 -10831
rect 21911 -10935 21945 -10901
rect 21979 -10934 22013 -10900
rect 22047 -10934 22081 -10900
rect 21911 -11004 21945 -10970
rect 21979 -11003 22013 -10969
rect 22047 -11003 22081 -10969
rect 21911 -11073 21945 -11039
rect 21979 -11072 22013 -11038
rect 22047 -11072 22081 -11038
rect 21911 -11142 21945 -11108
rect 21979 -11141 22013 -11107
rect 22047 -11141 22081 -11107
rect 21911 -11211 21945 -11177
rect 21979 -11210 22013 -11176
rect 22047 -11210 22081 -11176
rect 21911 -11280 21945 -11246
rect 21979 -11279 22013 -11245
rect 22047 -11279 22081 -11245
rect 21911 -11349 21945 -11315
rect 21979 -11348 22013 -11314
rect 22047 -11348 22081 -11314
rect 21911 -11418 21945 -11384
rect 21979 -11417 22013 -11383
rect 22047 -11417 22081 -11383
rect 21911 -11487 21945 -11453
rect 21979 -11486 22013 -11452
rect 22047 -11486 22081 -11452
rect 21911 -11556 21945 -11522
rect 21979 -11555 22013 -11521
rect 22047 -11555 22081 -11521
rect 21911 -11625 21945 -11591
rect 21979 -11624 22013 -11590
rect 22047 -11624 22081 -11590
rect 21911 -11694 21945 -11660
rect 21979 -11693 22013 -11659
rect 22047 -11693 22081 -11659
rect 21911 -11763 21945 -11729
rect 21979 -11762 22013 -11728
rect 22047 -11762 22081 -11728
rect 21911 -11832 21945 -11798
rect 21979 -11831 22013 -11797
rect 22047 -11831 22081 -11797
rect 21911 -11901 21945 -11867
rect 21979 -11900 22013 -11866
rect 22047 -11900 22081 -11866
rect 21911 -11970 21945 -11936
rect 21979 -11969 22013 -11935
rect 22047 -11969 22081 -11935
rect 21911 -12039 21945 -12005
rect 21979 -12038 22013 -12004
rect 22047 -12038 22081 -12004
rect 21911 -12108 21945 -12074
rect 21979 -12107 22013 -12073
rect 22047 -12107 22081 -12073
rect 21911 -12177 21945 -12143
rect 21979 -12176 22013 -12142
rect 22047 -12176 22081 -12142
rect 21911 -12246 21945 -12212
rect 21979 -12245 22013 -12211
rect 22047 -12245 22081 -12211
rect 21911 -12315 21945 -12281
rect 21979 -12314 22013 -12280
rect 22047 -12314 22081 -12280
rect 21911 -12384 21945 -12350
rect 21979 -12383 22013 -12349
rect 22047 -12383 22081 -12349
rect 21911 -12453 21945 -12419
rect 21979 -12452 22013 -12418
rect 22047 -12452 22081 -12418
rect 21911 -12522 21945 -12488
rect 21979 -12521 22013 -12487
rect 22047 -12521 22081 -12487
rect 21911 -12591 21945 -12557
rect 21979 -12590 22013 -12556
rect 22047 -12590 22081 -12556
rect 21911 -12660 21945 -12626
rect 21979 -12659 22013 -12625
rect 22047 -12659 22081 -12625
rect 21911 -12729 21945 -12695
rect 21979 -12728 22013 -12694
rect 22047 -12728 22081 -12694
rect 21911 -12798 21945 -12764
rect 21979 -12797 22013 -12763
rect 22047 -12797 22081 -12763
rect 21911 -12867 21945 -12833
rect 21979 -12866 22013 -12832
rect 22047 -12866 22081 -12832
rect 21911 -12936 21945 -12902
rect 21979 -12935 22013 -12901
rect 22047 -12935 22081 -12901
rect 21911 -13005 21945 -12971
rect 21979 -13004 22013 -12970
rect 22047 -13004 22081 -12970
rect 21911 -13074 21945 -13040
rect 21979 -13073 22013 -13039
rect 22047 -13073 22081 -13039
rect 21911 -13143 21945 -13109
rect 21979 -13142 22013 -13108
rect 22047 -13142 22081 -13108
rect 21911 -13212 21945 -13178
rect 21979 -13211 22013 -13177
rect 22047 -13211 22081 -13177
rect 21911 -13281 21945 -13247
rect 21979 -13280 22013 -13246
rect 22047 -13280 22081 -13246
rect 21911 -13350 21945 -13316
rect 21979 -13349 22013 -13315
rect 22047 -13349 22081 -13315
rect 21911 -13419 21945 -13385
rect 21979 -13418 22013 -13384
rect 22047 -13418 22081 -13384
rect 21911 -13488 21945 -13454
rect 21979 -13487 22013 -13453
rect 22047 -13487 22081 -13453
rect 21911 -13557 21945 -13523
rect 21979 -13556 22013 -13522
rect 22047 -13556 22081 -13522
rect 21911 -13626 21945 -13592
rect 21979 -13625 22013 -13591
rect 22047 -13625 22081 -13591
rect 21911 -13695 21945 -13661
rect 21979 -13694 22013 -13660
rect 22047 -13694 22081 -13660
rect 21911 -13764 21945 -13730
rect 21979 -13763 22013 -13729
rect 22047 -13763 22081 -13729
rect 21911 -13833 21945 -13799
rect 21979 -13832 22013 -13798
rect 22047 -13832 22081 -13798
rect 21911 -13902 21945 -13868
rect 21979 -13901 22013 -13867
rect 22047 -13901 22081 -13867
rect 21911 -13971 21945 -13937
rect 21979 -13970 22013 -13936
rect 22047 -13970 22081 -13936
rect 21911 -14040 21945 -14006
rect 21979 -14039 22013 -14005
rect 22047 -14039 22081 -14005
rect 21911 -14109 21945 -14075
rect 21979 -14108 22013 -14074
rect 22047 -14108 22081 -14074
rect 21911 -14178 21945 -14144
rect 21979 -14177 22013 -14143
rect 22047 -14177 22081 -14143
rect 21911 -14247 21945 -14213
rect 21979 -14246 22013 -14212
rect 22047 -14246 22081 -14212
rect 21911 -14316 21945 -14282
rect 21979 -14315 22013 -14281
rect 22047 -14315 22081 -14281
rect 21911 -14385 21945 -14351
rect 21979 -14384 22013 -14350
rect 22047 -14384 22081 -14350
rect 21911 -14454 21945 -14420
rect 21979 -14453 22013 -14419
rect 22047 -14453 22081 -14419
rect 21911 -14523 21945 -14489
rect 21979 -14522 22013 -14488
rect 22047 -14522 22081 -14488
rect 21911 -14592 21945 -14558
rect 21979 -14591 22013 -14557
rect 22047 -14591 22081 -14557
rect 21911 -14661 21945 -14627
rect 21979 -14660 22013 -14626
rect 22047 -14660 22081 -14626
rect 20470 -14866 20708 -14696
rect 20743 -14730 20777 -14696
rect 20812 -14730 20846 -14696
rect 20881 -14730 20915 -14696
rect 20950 -14730 20984 -14696
rect 21019 -14730 21053 -14696
rect 21088 -14730 21122 -14696
rect 21157 -14730 21191 -14696
rect 21226 -14730 21260 -14696
rect 21295 -14730 21329 -14696
rect 21364 -14730 21398 -14696
rect 21433 -14730 21467 -14696
rect 21502 -14730 21536 -14696
rect 21571 -14764 21945 -14696
rect 21979 -14729 22013 -14695
rect 22047 -14729 22081 -14695
rect 20743 -14798 20777 -14764
rect 20812 -14798 20846 -14764
rect 20881 -14798 20915 -14764
rect 20950 -14798 20984 -14764
rect 21019 -14798 21053 -14764
rect 21088 -14798 21122 -14764
rect 21157 -14798 21191 -14764
rect 21226 -14798 21260 -14764
rect 21295 -14798 21329 -14764
rect 21364 -14798 21398 -14764
rect 21433 -14798 21467 -14764
rect 21502 -14798 21536 -14764
rect 20743 -14866 20777 -14832
rect 20812 -14866 20846 -14832
rect 20881 -14866 20915 -14832
rect 20950 -14866 20984 -14832
rect 21019 -14866 21053 -14832
rect 21088 -14866 21122 -14832
rect 21157 -14866 21191 -14832
rect 21226 -14866 21260 -14832
rect 21295 -14866 21329 -14832
rect 21364 -14866 21398 -14832
rect 21433 -14866 21467 -14832
rect 21502 -14866 21536 -14832
rect 21571 -14866 22013 -14764
rect 22047 -14798 22081 -14764
rect 20470 -17274 20640 -14866
<< poly >>
rect -40 342 66 375
rect -40 308 -17 342
rect 17 308 66 342
rect -40 275 66 308
rect 1066 342 1198 375
rect 1066 308 1115 342
rect 1149 308 1198 342
rect 1066 275 1198 308
rect 2198 342 2330 375
rect 2198 308 2247 342
rect 2281 308 2330 342
rect 2198 275 2330 308
rect 3330 342 3462 375
rect 3330 308 3379 342
rect 3413 308 3462 342
rect 3330 275 3462 308
rect 4462 342 4594 375
rect 4462 308 4511 342
rect 4545 308 4594 342
rect 4462 275 4594 308
rect 5594 342 5726 375
rect 5594 308 5643 342
rect 5677 308 5726 342
rect 5594 275 5726 308
rect 6726 342 6832 375
rect 6726 308 6775 342
rect 6809 308 6832 342
rect 6726 275 6832 308
rect -40 187 66 219
rect -40 153 -17 187
rect 17 153 66 187
rect -40 119 66 153
rect 1066 187 1198 219
rect 1066 153 1115 187
rect 1149 153 1198 187
rect 1066 119 1198 153
rect 2198 187 2330 219
rect 2198 153 2247 187
rect 2281 153 2330 187
rect 2198 119 2330 153
rect 3330 187 3462 219
rect 3330 153 3379 187
rect 3413 153 3462 187
rect 3330 119 3462 153
rect 4462 187 4594 219
rect 4462 153 4511 187
rect 4545 153 4594 187
rect 4462 119 4594 153
rect 5594 187 5726 219
rect 5594 153 5643 187
rect 5677 153 5726 187
rect 5594 119 5726 153
rect 6726 187 6832 219
rect 6726 153 6775 187
rect 6809 153 6832 187
rect 6726 119 6832 153
rect -40 85 -17 119
rect 17 85 40 119
rect -40 69 40 85
rect 1092 85 1115 119
rect 1149 85 1172 119
rect 1092 69 1172 85
rect 2224 85 2247 119
rect 2281 85 2304 119
rect 2224 69 2304 85
rect 3356 85 3379 119
rect 3413 85 3436 119
rect 3356 69 3436 85
rect 4488 85 4511 119
rect 4545 85 4568 119
rect 4488 69 4568 85
rect 5620 85 5643 119
rect 5677 85 5700 119
rect 5620 69 5700 85
rect 6752 85 6775 119
rect 6809 85 6832 119
rect 6752 69 6832 85
rect 20869 -3386 20969 -3354
rect 21025 -3386 21125 -3354
rect 20869 -4018 20969 -3986
rect 21025 -4018 21125 -3986
rect 20869 -4034 21125 -4018
rect 20869 -4068 20885 -4034
rect 20919 -4068 20980 -4034
rect 21014 -4068 21075 -4034
rect 21109 -4068 21125 -4034
rect 20869 -4084 21125 -4068
rect 21268 -9940 21368 -9914
rect 21424 -9940 21524 -9914
rect 21268 -10589 21368 -10540
rect 21268 -10623 21301 -10589
rect 21335 -10623 21368 -10589
rect 21268 -10646 21368 -10623
rect 21424 -10589 21524 -10540
rect 21424 -10623 21457 -10589
rect 21491 -10623 21524 -10589
rect 21424 -10646 21524 -10623
<< polycont >>
rect -17 308 17 342
rect 1115 308 1149 342
rect 2247 308 2281 342
rect 3379 308 3413 342
rect 4511 308 4545 342
rect 5643 308 5677 342
rect 6775 308 6809 342
rect -17 153 17 187
rect 1115 153 1149 187
rect 2247 153 2281 187
rect 3379 153 3413 187
rect 4511 153 4545 187
rect 5643 153 5677 187
rect 6775 153 6809 187
rect -17 85 17 119
rect 1115 85 1149 119
rect 2247 85 2281 119
rect 3379 85 3413 119
rect 4511 85 4545 119
rect 5643 85 5677 119
rect 6775 85 6809 119
rect 20885 -4068 20919 -4034
rect 20980 -4068 21014 -4034
rect 21075 -4068 21109 -4034
rect 21301 -10623 21335 -10589
rect 21457 -10623 21491 -10589
<< locali >>
rect 134 386 136 420
rect 170 386 172 420
rect 238 386 244 420
rect 306 386 316 420
rect 374 386 388 420
rect 442 386 460 420
rect 510 386 532 420
rect 578 386 604 420
rect 646 386 676 420
rect 714 386 748 420
rect 782 386 816 420
rect 854 386 884 420
rect 926 386 952 420
rect 998 386 1020 420
rect 1244 386 1266 420
rect 1312 386 1338 420
rect 1380 386 1410 420
rect 1448 386 1482 420
rect 1516 386 1550 420
rect 1588 386 1618 420
rect 1660 386 1686 420
rect 1732 386 1754 420
rect 1804 386 1822 420
rect 1876 386 1890 420
rect 1948 386 1958 420
rect 2020 386 2026 420
rect 2092 386 2094 420
rect 2128 386 2130 420
rect 2398 386 2400 420
rect 2434 386 2436 420
rect 2502 386 2508 420
rect 2570 386 2580 420
rect 2638 386 2652 420
rect 2706 386 2724 420
rect 2774 386 2796 420
rect 2842 386 2868 420
rect 2910 386 2940 420
rect 2978 386 3012 420
rect 3046 386 3080 420
rect 3118 386 3148 420
rect 3190 386 3216 420
rect 3262 386 3284 420
rect 3508 386 3530 420
rect 3576 386 3602 420
rect 3644 386 3674 420
rect 3712 386 3746 420
rect 3780 386 3814 420
rect 3852 386 3882 420
rect 3924 386 3950 420
rect 3996 386 4018 420
rect 4068 386 4086 420
rect 4140 386 4154 420
rect 4212 386 4222 420
rect 4284 386 4290 420
rect 4356 386 4358 420
rect 4392 386 4394 420
rect 4662 386 4664 420
rect 4698 386 4700 420
rect 4766 386 4772 420
rect 4834 386 4844 420
rect 4902 386 4916 420
rect 4970 386 4988 420
rect 5038 386 5060 420
rect 5106 386 5132 420
rect 5174 386 5204 420
rect 5242 386 5276 420
rect 5310 386 5344 420
rect 5382 386 5412 420
rect 5454 386 5480 420
rect 5526 386 5548 420
rect 5772 386 5794 420
rect 5840 386 5866 420
rect 5908 386 5938 420
rect 5976 386 6010 420
rect 6044 386 6078 420
rect 6116 386 6146 420
rect 6188 386 6214 420
rect 6260 386 6282 420
rect 6332 386 6350 420
rect 6404 386 6418 420
rect 6476 386 6486 420
rect 6548 386 6554 420
rect 6620 386 6622 420
rect 6656 386 6658 420
rect -26 351 26 359
rect 1106 351 1158 359
rect 2238 351 2290 359
rect 3370 351 3422 359
rect 4502 351 4554 359
rect 5634 351 5686 359
rect 6766 351 6818 359
rect -26 342 6818 351
rect -26 308 -17 342
rect 17 308 1115 342
rect 1149 308 2247 342
rect 2281 308 3379 342
rect 3413 308 4511 342
rect 4545 308 5643 342
rect 5677 308 6775 342
rect 6809 308 6818 342
rect -26 299 6818 308
rect -26 187 26 299
rect 134 230 136 264
rect 170 230 172 264
rect 238 230 244 264
rect 306 230 316 264
rect 374 230 388 264
rect 442 230 460 264
rect 510 230 532 264
rect 578 230 604 264
rect 646 230 676 264
rect 714 230 748 264
rect 782 230 816 264
rect 854 230 884 264
rect 926 230 952 264
rect 998 230 1020 264
rect -26 186 -17 187
rect -19 153 -17 186
rect 17 186 26 187
rect 1106 187 1158 299
rect 1244 230 1266 264
rect 1312 230 1338 264
rect 1380 230 1410 264
rect 1448 230 1482 264
rect 1516 230 1550 264
rect 1588 230 1618 264
rect 1660 230 1686 264
rect 1732 230 1754 264
rect 1804 230 1822 264
rect 1876 230 1890 264
rect 1948 230 1958 264
rect 2020 230 2026 264
rect 2092 230 2094 264
rect 2128 230 2130 264
rect 1106 186 1115 187
rect 17 153 19 186
rect -19 152 19 153
rect 1113 153 1115 186
rect 1149 186 1158 187
rect 2238 187 2290 299
rect 2398 230 2400 264
rect 2434 230 2436 264
rect 2502 230 2508 264
rect 2570 230 2580 264
rect 2638 230 2652 264
rect 2706 230 2724 264
rect 2774 230 2796 264
rect 2842 230 2868 264
rect 2910 230 2940 264
rect 2978 230 3012 264
rect 3046 230 3080 264
rect 3118 230 3148 264
rect 3190 230 3216 264
rect 3262 230 3284 264
rect 2238 186 2247 187
rect 1149 153 1151 186
rect 1113 152 1151 153
rect 2245 153 2247 186
rect 2281 186 2290 187
rect 3370 187 3422 299
rect 3508 230 3530 264
rect 3576 230 3602 264
rect 3644 230 3674 264
rect 3712 230 3746 264
rect 3780 230 3814 264
rect 3852 230 3882 264
rect 3924 230 3950 264
rect 3996 230 4018 264
rect 4068 230 4086 264
rect 4140 230 4154 264
rect 4212 230 4222 264
rect 4284 230 4290 264
rect 4356 230 4358 264
rect 4392 230 4394 264
rect 3370 186 3379 187
rect 2281 153 2283 186
rect 2245 152 2283 153
rect 3377 153 3379 186
rect 3413 186 3422 187
rect 4502 187 4554 299
rect 4662 230 4664 264
rect 4698 230 4700 264
rect 4766 230 4772 264
rect 4834 230 4844 264
rect 4902 230 4916 264
rect 4970 230 4988 264
rect 5038 230 5060 264
rect 5106 230 5132 264
rect 5174 230 5204 264
rect 5242 230 5276 264
rect 5310 230 5344 264
rect 5382 230 5412 264
rect 5454 230 5480 264
rect 5526 230 5548 264
rect 4502 186 4511 187
rect 3413 153 3415 186
rect 3377 152 3415 153
rect 4509 153 4511 186
rect 4545 186 4554 187
rect 5634 187 5686 299
rect 5772 230 5794 264
rect 5840 230 5866 264
rect 5908 230 5938 264
rect 5976 230 6010 264
rect 6044 230 6078 264
rect 6116 230 6146 264
rect 6188 230 6214 264
rect 6260 230 6282 264
rect 6332 230 6350 264
rect 6404 230 6418 264
rect 6476 230 6486 264
rect 6548 230 6554 264
rect 6620 230 6622 264
rect 6656 230 6658 264
rect 5634 186 5643 187
rect 4545 153 4547 186
rect 4509 152 4547 153
rect 5641 153 5643 186
rect 5677 186 5686 187
rect 6766 187 6818 299
rect 6766 186 6775 187
rect 5677 153 5679 186
rect 5641 152 5679 153
rect 6773 153 6775 186
rect 6809 186 6818 187
rect 6809 153 6811 186
rect 6773 152 6811 153
rect -26 136 26 152
rect 1106 136 1158 152
rect 2238 136 2290 152
rect 3370 136 3422 152
rect 4502 136 4554 152
rect 5634 136 5686 152
rect 6766 136 6818 152
rect -24 119 24 136
rect -24 85 -17 119
rect 17 85 24 119
rect 1108 119 1156 136
rect -24 69 24 85
rect 134 74 136 108
rect 170 74 172 108
rect 238 74 244 108
rect 306 74 316 108
rect 374 74 388 108
rect 442 74 460 108
rect 510 74 532 108
rect 578 74 604 108
rect 646 74 676 108
rect 714 74 748 108
rect 782 74 816 108
rect 854 74 884 108
rect 926 74 952 108
rect 998 74 1020 108
rect 1108 85 1115 119
rect 1149 85 1156 119
rect 2240 119 2288 136
rect 1108 69 1156 85
rect 1244 74 1266 108
rect 1312 74 1338 108
rect 1380 74 1410 108
rect 1448 74 1482 108
rect 1516 74 1550 108
rect 1588 74 1618 108
rect 1660 74 1686 108
rect 1732 74 1754 108
rect 1804 74 1822 108
rect 1876 74 1890 108
rect 1948 74 1958 108
rect 2020 74 2026 108
rect 2092 74 2094 108
rect 2128 74 2130 108
rect 2240 85 2247 119
rect 2281 85 2288 119
rect 3372 119 3420 136
rect 2240 69 2288 85
rect 2398 74 2400 108
rect 2434 74 2436 108
rect 2502 74 2508 108
rect 2570 74 2580 108
rect 2638 74 2652 108
rect 2706 74 2724 108
rect 2774 74 2796 108
rect 2842 74 2868 108
rect 2910 74 2940 108
rect 2978 74 3012 108
rect 3046 74 3080 108
rect 3118 74 3148 108
rect 3190 74 3216 108
rect 3262 74 3284 108
rect 3372 85 3379 119
rect 3413 85 3420 119
rect 4504 119 4552 136
rect 3372 69 3420 85
rect 3508 74 3530 108
rect 3576 74 3602 108
rect 3644 74 3674 108
rect 3712 74 3746 108
rect 3780 74 3814 108
rect 3852 74 3882 108
rect 3924 74 3950 108
rect 3996 74 4018 108
rect 4068 74 4086 108
rect 4140 74 4154 108
rect 4212 74 4222 108
rect 4284 74 4290 108
rect 4356 74 4358 108
rect 4392 74 4394 108
rect 4504 85 4511 119
rect 4545 85 4552 119
rect 5636 119 5684 136
rect 4504 69 4552 85
rect 4662 74 4664 108
rect 4698 74 4700 108
rect 4766 74 4772 108
rect 4834 74 4844 108
rect 4902 74 4916 108
rect 4970 74 4988 108
rect 5038 74 5060 108
rect 5106 74 5132 108
rect 5174 74 5204 108
rect 5242 74 5276 108
rect 5310 74 5344 108
rect 5382 74 5412 108
rect 5454 74 5480 108
rect 5526 74 5548 108
rect 5636 85 5643 119
rect 5677 85 5684 119
rect 6768 119 6816 136
rect 5636 69 5684 85
rect 5772 74 5794 108
rect 5840 74 5866 108
rect 5908 74 5938 108
rect 5976 74 6010 108
rect 6044 74 6078 108
rect 6116 74 6146 108
rect 6188 74 6214 108
rect 6260 74 6282 108
rect 6332 74 6350 108
rect 6404 74 6418 108
rect 6476 74 6486 108
rect 6548 74 6554 108
rect 6620 74 6622 108
rect 6656 74 6658 108
rect 6768 85 6775 119
rect 6809 85 6816 119
rect 6768 69 6816 85
rect 20824 -3464 20858 -3448
rect 20824 -3532 20858 -3498
rect 20824 -3600 20858 -3566
rect 20824 -3668 20858 -3634
rect 20824 -3736 20858 -3719
rect 20824 -3794 20858 -3770
rect 20824 -3872 20858 -3838
rect 20824 -3940 20858 -3906
rect 20824 -3990 20858 -3974
rect 20980 -3464 21014 -3459
rect 20980 -3532 21014 -3531
rect 20980 -3600 21014 -3566
rect 20980 -3668 21014 -3634
rect 20980 -3736 21014 -3702
rect 20980 -3804 21014 -3770
rect 20980 -3872 21014 -3838
rect 20980 -3940 21014 -3906
rect 20980 -3990 21014 -3974
rect 21136 -3464 21170 -3448
rect 21136 -3532 21170 -3498
rect 21136 -3600 21170 -3566
rect 21136 -3668 21170 -3634
rect 21136 -3736 21170 -3719
rect 21136 -3794 21170 -3770
rect 21136 -3872 21170 -3838
rect 21136 -3940 21170 -3906
rect 21136 -3990 21170 -3974
rect 20869 -4068 20885 -4034
rect 20919 -4068 20980 -4034
rect 21014 -4068 21075 -4034
rect 21109 -4068 21125 -4034
rect 20470 -7504 20640 -7470
rect 20504 -7538 20538 -7504
rect 20572 -7538 20606 -7504
rect 20470 -7573 20640 -7538
rect 20504 -7607 20538 -7573
rect 20572 -7607 20606 -7573
rect 20470 -7642 20640 -7607
rect 20504 -7676 20538 -7642
rect 20572 -7676 20606 -7642
rect 20470 -7711 20640 -7676
rect 20504 -7745 20538 -7711
rect 20572 -7745 20606 -7711
rect 20470 -7780 20640 -7745
rect 20504 -7814 20538 -7780
rect 20572 -7814 20606 -7780
rect 20470 -7849 20640 -7814
rect 20504 -7883 20538 -7849
rect 20572 -7883 20606 -7849
rect 20470 -7887 20640 -7883
rect 20470 -7893 22091 -7887
rect 20470 -7918 20651 -7893
rect 20685 -7898 20724 -7893
rect 20758 -7898 20797 -7893
rect 20831 -7898 20870 -7893
rect 20904 -7898 20943 -7893
rect 20977 -7898 21017 -7893
rect 21051 -7898 21091 -7893
rect 21125 -7898 21165 -7893
rect 21199 -7898 21239 -7893
rect 21273 -7898 21313 -7893
rect 21347 -7898 21387 -7893
rect 21421 -7898 21461 -7893
rect 20504 -7952 20538 -7918
rect 20572 -7952 20606 -7918
rect 20640 -7927 20651 -7918
rect 21125 -7927 21151 -7898
rect 21199 -7927 21220 -7898
rect 21273 -7927 21289 -7898
rect 21347 -7927 21358 -7898
rect 21421 -7927 21427 -7898
rect 20640 -7952 20674 -7927
rect 20470 -7965 20674 -7952
rect 21116 -7932 21151 -7927
rect 21185 -7932 21220 -7927
rect 21254 -7932 21289 -7927
rect 21323 -7932 21358 -7927
rect 21392 -7932 21427 -7927
rect 21495 -7898 21535 -7893
rect 21569 -7898 21609 -7893
rect 21643 -7898 21683 -7893
rect 21717 -7898 21757 -7893
rect 21791 -7898 21831 -7893
rect 21865 -7898 21905 -7893
rect 21939 -7898 21979 -7893
rect 21495 -7927 21496 -7898
rect 21461 -7932 21496 -7927
rect 21530 -7927 21535 -7898
rect 21599 -7927 21609 -7898
rect 21668 -7927 21683 -7898
rect 21737 -7927 21757 -7898
rect 21806 -7927 21831 -7898
rect 21875 -7927 21905 -7898
rect 21530 -7932 21565 -7927
rect 21599 -7932 21634 -7927
rect 21668 -7932 21703 -7927
rect 21737 -7932 21772 -7927
rect 21806 -7932 21841 -7927
rect 21875 -7932 21910 -7927
rect 21944 -7932 21979 -7898
rect 22013 -7932 22091 -7893
rect 21116 -7965 22091 -7932
rect 20470 -7987 20651 -7965
rect 20504 -8021 20538 -7987
rect 20572 -8021 20606 -7987
rect 20640 -7999 20651 -7987
rect 21125 -7966 21165 -7965
rect 21199 -7966 21239 -7965
rect 21273 -7966 21313 -7965
rect 21347 -7966 21387 -7965
rect 21421 -7966 21461 -7965
rect 21125 -7999 21151 -7966
rect 21199 -7999 21220 -7966
rect 21273 -7999 21289 -7966
rect 21347 -7999 21358 -7966
rect 21421 -7999 21427 -7966
rect 20640 -8021 20674 -7999
rect 21116 -8000 21151 -7999
rect 21185 -8000 21220 -7999
rect 21254 -8000 21289 -7999
rect 21323 -8000 21358 -7999
rect 21392 -8000 21427 -7999
rect 21495 -7966 21535 -7965
rect 21569 -7966 21609 -7965
rect 21643 -7966 21683 -7965
rect 21717 -7966 21757 -7965
rect 21791 -7966 21831 -7965
rect 21865 -7966 21905 -7965
rect 21939 -7966 21979 -7965
rect 21495 -7999 21496 -7966
rect 21461 -8000 21496 -7999
rect 21530 -7999 21535 -7966
rect 21599 -7999 21609 -7966
rect 21668 -7999 21683 -7966
rect 21737 -7999 21757 -7966
rect 21806 -7999 21831 -7966
rect 21875 -7999 21905 -7966
rect 21530 -8000 21565 -7999
rect 21599 -8000 21634 -7999
rect 21668 -8000 21703 -7999
rect 21737 -8000 21772 -7999
rect 21806 -8000 21841 -7999
rect 21875 -8000 21910 -7999
rect 21944 -8000 21979 -7966
rect 20470 -8037 20674 -8021
rect 21048 -8034 21979 -8000
rect 21048 -8037 21083 -8034
rect 21117 -8037 21152 -8034
rect 21186 -8037 21221 -8034
rect 21255 -8037 21290 -8034
rect 21324 -8037 21359 -8034
rect 21393 -8037 21428 -8034
rect 20470 -8056 20651 -8037
rect 20504 -8090 20538 -8056
rect 20572 -8090 20606 -8056
rect 20640 -8071 20651 -8056
rect 21053 -8068 21083 -8037
rect 21127 -8068 21152 -8037
rect 21201 -8068 21221 -8037
rect 21275 -8068 21290 -8037
rect 21349 -8068 21359 -8037
rect 21423 -8068 21428 -8037
rect 21462 -8037 21497 -8034
rect 21462 -8068 21463 -8037
rect 20685 -8071 20724 -8068
rect 20758 -8071 20797 -8068
rect 20831 -8071 20871 -8068
rect 20905 -8071 20945 -8068
rect 20979 -8071 21019 -8068
rect 21053 -8071 21093 -8068
rect 21127 -8071 21167 -8068
rect 21201 -8071 21241 -8068
rect 21275 -8071 21315 -8068
rect 21349 -8071 21389 -8068
rect 21423 -8071 21463 -8068
rect 21531 -8037 21566 -8034
rect 21600 -8037 21635 -8034
rect 21669 -8037 21704 -8034
rect 21738 -8037 21773 -8034
rect 21807 -8037 21842 -8034
rect 21876 -8037 21911 -8034
rect 21531 -8068 21537 -8037
rect 21600 -8068 21611 -8037
rect 21669 -8068 21685 -8037
rect 21738 -8068 21759 -8037
rect 21807 -8068 21833 -8037
rect 21876 -8068 21907 -8037
rect 21497 -8071 21537 -8068
rect 21571 -8071 21611 -8068
rect 21645 -8071 21685 -8068
rect 21719 -8071 21759 -8068
rect 21793 -8071 21833 -8068
rect 21867 -8071 21907 -8068
rect 20640 -8077 21907 -8071
rect 20470 -8125 20640 -8090
rect 20504 -8159 20538 -8125
rect 20572 -8159 20606 -8125
rect 20470 -8194 20640 -8159
rect 20504 -8228 20538 -8194
rect 20572 -8228 20606 -8194
rect 20470 -8263 20640 -8228
rect 20504 -8297 20538 -8263
rect 20572 -8297 20606 -8263
rect 20470 -8332 20640 -8297
rect 21033 -8275 21113 -8241
rect 21147 -8275 21181 -8241
rect 21033 -8309 21181 -8275
rect 21135 -8343 21181 -8309
rect 21691 -8322 21759 -8241
rect 21691 -8343 21725 -8322
rect 21657 -8356 21725 -8343
rect 21657 -8390 21759 -8356
rect 21223 -10006 21257 -10002
rect 21223 -10078 21257 -10052
rect 21223 -10150 21257 -10120
rect 21223 -10222 21257 -10188
rect 21223 -10290 21257 -10256
rect 21223 -10358 21257 -10328
rect 21223 -10426 21257 -10400
rect 21223 -10494 21257 -10472
rect 21379 -10006 21413 -10002
rect 21379 -10078 21413 -10052
rect 21379 -10150 21413 -10120
rect 21379 -10222 21413 -10188
rect 21379 -10290 21413 -10256
rect 21379 -10358 21413 -10328
rect 21379 -10426 21413 -10400
rect 21379 -10494 21413 -10472
rect 21535 -10006 21569 -10002
rect 21535 -10078 21569 -10052
rect 21535 -10150 21569 -10120
rect 21535 -10222 21569 -10188
rect 21535 -10290 21569 -10256
rect 21535 -10358 21569 -10328
rect 21535 -10426 21569 -10400
rect 21535 -10494 21569 -10472
rect 21284 -10587 21301 -10582
rect 21335 -10587 21507 -10582
rect 21284 -10589 21507 -10587
rect 21284 -10623 21301 -10589
rect 21335 -10623 21457 -10589
rect 21491 -10623 21507 -10589
rect 21284 -10625 21507 -10623
rect 21284 -10630 21301 -10625
rect 21335 -10630 21507 -10625
rect 21033 -14429 21135 -14395
rect 21067 -14442 21135 -14429
rect 21067 -14463 21101 -14442
rect 21033 -14544 21101 -14463
rect 21543 -14476 21657 -14442
rect 21543 -14510 21759 -14476
rect 21543 -14544 21649 -14510
rect 21683 -14544 21759 -14510
rect 21901 -12463 21907 -8077
rect 21901 -12488 21979 -12463
rect 21901 -12502 21911 -12488
rect 21901 -12536 21907 -12502
rect 21945 -12522 21979 -12488
rect 21941 -12535 21979 -12522
rect 22085 -12535 22091 -7965
rect 21941 -12536 22091 -12535
rect 21901 -12556 22091 -12536
rect 21901 -12557 21979 -12556
rect 21901 -12575 21911 -12557
rect 21901 -12609 21907 -12575
rect 21945 -12591 21979 -12557
rect 22013 -12590 22047 -12556
rect 22081 -12574 22091 -12556
rect 21941 -12608 21979 -12591
rect 22013 -12608 22051 -12590
rect 22085 -12608 22091 -12574
rect 21941 -12609 22091 -12608
rect 21901 -12625 22091 -12609
rect 21901 -12626 21979 -12625
rect 21901 -12648 21911 -12626
rect 21901 -12682 21907 -12648
rect 21945 -12660 21979 -12626
rect 22013 -12659 22047 -12625
rect 22081 -12647 22091 -12625
rect 21941 -12681 21979 -12660
rect 22013 -12681 22051 -12659
rect 22085 -12681 22091 -12647
rect 21941 -12682 22091 -12681
rect 21901 -12694 22091 -12682
rect 21901 -12695 21979 -12694
rect 21901 -12721 21911 -12695
rect 21901 -12755 21907 -12721
rect 21945 -12729 21979 -12695
rect 22013 -12728 22047 -12694
rect 22081 -12720 22091 -12694
rect 21941 -12754 21979 -12729
rect 22013 -12754 22051 -12728
rect 22085 -12754 22091 -12720
rect 21941 -12755 22091 -12754
rect 21901 -12763 22091 -12755
rect 21901 -12764 21979 -12763
rect 21901 -12794 21911 -12764
rect 21901 -12828 21907 -12794
rect 21945 -12798 21979 -12764
rect 22013 -12797 22047 -12763
rect 22081 -12793 22091 -12763
rect 21941 -12827 21979 -12798
rect 22013 -12827 22051 -12797
rect 22085 -12827 22091 -12793
rect 21941 -12828 22091 -12827
rect 21901 -12832 22091 -12828
rect 21901 -12833 21979 -12832
rect 21901 -12867 21911 -12833
rect 21945 -12867 21979 -12833
rect 22013 -12866 22047 -12832
rect 22081 -12866 22091 -12832
rect 21901 -12901 21907 -12867
rect 21941 -12900 21979 -12867
rect 22013 -12900 22051 -12866
rect 22085 -12900 22091 -12866
rect 21941 -12901 22091 -12900
rect 21901 -12902 21979 -12901
rect 21901 -12936 21911 -12902
rect 21945 -12935 21979 -12902
rect 22013 -12935 22047 -12901
rect 22081 -12935 22091 -12901
rect 21945 -12936 22091 -12935
rect 21901 -12939 22091 -12936
rect 21901 -12940 21979 -12939
rect 21901 -12974 21907 -12940
rect 21941 -12971 21979 -12940
rect 22013 -12970 22051 -12939
rect 21901 -13005 21911 -12974
rect 21945 -13004 21979 -12971
rect 22013 -13004 22047 -12970
rect 22085 -12973 22091 -12939
rect 22081 -13004 22091 -12973
rect 21945 -13005 22091 -13004
rect 21901 -13012 22091 -13005
rect 21901 -13013 21979 -13012
rect 21901 -13047 21907 -13013
rect 21941 -13040 21979 -13013
rect 22013 -13039 22051 -13012
rect 21901 -13074 21911 -13047
rect 21945 -13073 21979 -13040
rect 22013 -13073 22047 -13039
rect 22085 -13046 22091 -13012
rect 22081 -13073 22091 -13046
rect 21945 -13074 22091 -13073
rect 21901 -13085 22091 -13074
rect 21901 -13086 21979 -13085
rect 21901 -13120 21907 -13086
rect 21941 -13109 21979 -13086
rect 22013 -13108 22051 -13085
rect 21901 -13143 21911 -13120
rect 21945 -13142 21979 -13109
rect 22013 -13142 22047 -13108
rect 22085 -13119 22091 -13085
rect 22081 -13142 22091 -13119
rect 21945 -13143 22091 -13142
rect 21901 -13158 22091 -13143
rect 21901 -13159 21979 -13158
rect 21901 -13193 21907 -13159
rect 21941 -13178 21979 -13159
rect 22013 -13177 22051 -13158
rect 21901 -13212 21911 -13193
rect 21945 -13211 21979 -13178
rect 22013 -13211 22047 -13177
rect 22085 -13192 22091 -13158
rect 22081 -13211 22091 -13192
rect 21945 -13212 22091 -13211
rect 21901 -13231 22091 -13212
rect 21901 -13232 21979 -13231
rect 21901 -13266 21907 -13232
rect 21941 -13247 21979 -13232
rect 22013 -13246 22051 -13231
rect 21901 -13281 21911 -13266
rect 21945 -13280 21979 -13247
rect 22013 -13280 22047 -13246
rect 22085 -13265 22091 -13231
rect 22081 -13280 22091 -13265
rect 21945 -13281 22091 -13280
rect 21901 -13304 22091 -13281
rect 21901 -13305 21979 -13304
rect 21901 -13339 21907 -13305
rect 21941 -13316 21979 -13305
rect 22013 -13315 22051 -13304
rect 21901 -13350 21911 -13339
rect 21945 -13349 21979 -13316
rect 22013 -13349 22047 -13315
rect 22085 -13338 22091 -13304
rect 22081 -13349 22091 -13338
rect 21945 -13350 22091 -13349
rect 21901 -13377 22091 -13350
rect 21901 -13378 21979 -13377
rect 21901 -13412 21907 -13378
rect 21941 -13385 21979 -13378
rect 22013 -13384 22051 -13377
rect 21901 -13419 21911 -13412
rect 21945 -13418 21979 -13385
rect 22013 -13418 22047 -13384
rect 22085 -13411 22091 -13377
rect 22081 -13418 22091 -13411
rect 21945 -13419 22091 -13418
rect 21901 -13450 22091 -13419
rect 21901 -13451 21979 -13450
rect 21901 -13485 21907 -13451
rect 21941 -13454 21979 -13451
rect 22013 -13453 22051 -13450
rect 21901 -13488 21911 -13485
rect 21945 -13487 21979 -13454
rect 22013 -13487 22047 -13453
rect 22085 -13484 22091 -13450
rect 22081 -13487 22091 -13484
rect 21945 -13488 22091 -13487
rect 21901 -13522 22091 -13488
rect 21901 -13523 21979 -13522
rect 21901 -13524 21911 -13523
rect 21901 -13558 21907 -13524
rect 21945 -13557 21979 -13523
rect 22013 -13556 22047 -13522
rect 22081 -13523 22091 -13522
rect 22013 -13557 22051 -13556
rect 22085 -13557 22091 -13523
rect 21941 -13558 22091 -13557
rect 21901 -13591 22091 -13558
rect 21901 -13592 21979 -13591
rect 21901 -13597 21911 -13592
rect 21901 -13631 21907 -13597
rect 21945 -13626 21979 -13592
rect 22013 -13625 22047 -13591
rect 22081 -13596 22091 -13591
rect 21941 -13630 21979 -13626
rect 22013 -13630 22051 -13625
rect 22085 -13630 22091 -13596
rect 21941 -13631 22091 -13630
rect 21901 -13660 22091 -13631
rect 21901 -13661 21979 -13660
rect 21901 -13670 21911 -13661
rect 21901 -13704 21907 -13670
rect 21945 -13695 21979 -13661
rect 22013 -13694 22047 -13660
rect 22081 -13669 22091 -13660
rect 21941 -13703 21979 -13695
rect 22013 -13703 22051 -13694
rect 22085 -13703 22091 -13669
rect 21941 -13704 22091 -13703
rect 21901 -13729 22091 -13704
rect 21901 -13730 21979 -13729
rect 21901 -13743 21911 -13730
rect 21901 -13777 21907 -13743
rect 21945 -13764 21979 -13730
rect 22013 -13763 22047 -13729
rect 22081 -13742 22091 -13729
rect 21941 -13776 21979 -13764
rect 22013 -13776 22051 -13763
rect 22085 -13776 22091 -13742
rect 21941 -13777 22091 -13776
rect 21901 -13798 22091 -13777
rect 21901 -13799 21979 -13798
rect 21901 -13816 21911 -13799
rect 21901 -13850 21907 -13816
rect 21945 -13833 21979 -13799
rect 22013 -13832 22047 -13798
rect 22081 -13815 22091 -13798
rect 21941 -13849 21979 -13833
rect 22013 -13849 22051 -13832
rect 22085 -13849 22091 -13815
rect 21941 -13850 22091 -13849
rect 21901 -13867 22091 -13850
rect 21901 -13868 21979 -13867
rect 21901 -13889 21911 -13868
rect 21901 -13923 21907 -13889
rect 21945 -13902 21979 -13868
rect 22013 -13901 22047 -13867
rect 22081 -13888 22091 -13867
rect 21941 -13922 21979 -13902
rect 22013 -13922 22051 -13901
rect 22085 -13922 22091 -13888
rect 21941 -13923 22091 -13922
rect 21901 -13936 22091 -13923
rect 21901 -13937 21979 -13936
rect 21901 -13962 21911 -13937
rect 21901 -13996 21907 -13962
rect 21945 -13971 21979 -13937
rect 22013 -13970 22047 -13936
rect 22081 -13961 22091 -13936
rect 21941 -13995 21979 -13971
rect 22013 -13995 22051 -13970
rect 22085 -13995 22091 -13961
rect 21941 -13996 22091 -13995
rect 21901 -14005 22091 -13996
rect 21901 -14006 21979 -14005
rect 21901 -14035 21911 -14006
rect 21901 -14069 21907 -14035
rect 21945 -14040 21979 -14006
rect 22013 -14039 22047 -14005
rect 22081 -14034 22091 -14005
rect 21941 -14068 21979 -14040
rect 22013 -14068 22051 -14039
rect 22085 -14068 22091 -14034
rect 21941 -14069 22091 -14068
rect 21901 -14074 22091 -14069
rect 21901 -14075 21979 -14074
rect 21901 -14108 21911 -14075
rect 21901 -14142 21907 -14108
rect 21945 -14109 21979 -14075
rect 22013 -14108 22047 -14074
rect 22081 -14107 22091 -14074
rect 21941 -14141 21979 -14109
rect 22013 -14141 22051 -14108
rect 22085 -14141 22091 -14107
rect 21941 -14142 22091 -14141
rect 21901 -14143 22091 -14142
rect 21901 -14144 21979 -14143
rect 21901 -14178 21911 -14144
rect 21945 -14177 21979 -14144
rect 22013 -14177 22047 -14143
rect 22081 -14177 22091 -14143
rect 21945 -14178 22091 -14177
rect 21901 -14180 22091 -14178
rect 21901 -14181 21979 -14180
rect 21901 -14215 21907 -14181
rect 21941 -14213 21979 -14181
rect 22013 -14212 22051 -14180
rect 21901 -14247 21911 -14215
rect 21945 -14246 21979 -14213
rect 22013 -14246 22047 -14212
rect 22085 -14214 22091 -14180
rect 22081 -14246 22091 -14214
rect 21945 -14247 22091 -14246
rect 21901 -14253 22091 -14247
rect 21901 -14254 21979 -14253
rect 21901 -14288 21907 -14254
rect 21941 -14282 21979 -14254
rect 22013 -14281 22051 -14253
rect 21901 -14316 21911 -14288
rect 21945 -14315 21979 -14282
rect 22013 -14315 22047 -14281
rect 22085 -14287 22091 -14253
rect 22081 -14315 22091 -14287
rect 21945 -14316 22091 -14315
rect 21901 -14326 22091 -14316
rect 21901 -14327 21979 -14326
rect 21901 -14361 21907 -14327
rect 21941 -14351 21979 -14327
rect 22013 -14350 22051 -14326
rect 21901 -14385 21911 -14361
rect 21945 -14384 21979 -14351
rect 22013 -14384 22047 -14350
rect 22085 -14360 22091 -14326
rect 22081 -14384 22091 -14360
rect 21945 -14385 22091 -14384
rect 21901 -14399 22091 -14385
rect 21901 -14400 21979 -14399
rect 21901 -14434 21907 -14400
rect 21941 -14420 21979 -14400
rect 22013 -14419 22051 -14399
rect 21901 -14454 21911 -14434
rect 21945 -14453 21979 -14420
rect 22013 -14453 22047 -14419
rect 22085 -14433 22091 -14399
rect 22081 -14453 22091 -14433
rect 21945 -14454 22091 -14453
rect 21901 -14472 22091 -14454
rect 21901 -14473 21979 -14472
rect 21901 -14507 21907 -14473
rect 21941 -14489 21979 -14473
rect 22013 -14488 22051 -14472
rect 21901 -14523 21911 -14507
rect 21945 -14522 21979 -14489
rect 22013 -14522 22047 -14488
rect 22085 -14506 22091 -14472
rect 22081 -14522 22091 -14506
rect 21945 -14523 22091 -14522
rect 21901 -14545 22091 -14523
rect 21901 -14546 21979 -14545
rect 21901 -14580 21907 -14546
rect 21941 -14558 21979 -14546
rect 22013 -14557 22051 -14545
rect 21901 -14592 21911 -14580
rect 21945 -14591 21979 -14558
rect 22013 -14591 22047 -14557
rect 22085 -14579 22091 -14545
rect 22081 -14591 22091 -14579
rect 21945 -14592 22091 -14591
rect 21901 -14618 22091 -14592
rect 21901 -14619 21979 -14618
rect 21901 -14653 21907 -14619
rect 21941 -14627 21979 -14619
rect 22013 -14626 22051 -14618
rect 21901 -14661 21911 -14653
rect 21945 -14660 21979 -14627
rect 22013 -14660 22047 -14626
rect 22085 -14652 22091 -14618
rect 22081 -14660 22091 -14652
rect 21945 -14661 22091 -14660
rect 21901 -14686 22091 -14661
rect 20640 -14691 22091 -14686
rect 20640 -14692 21979 -14691
rect 20640 -14696 20651 -14692
rect 20685 -14696 20725 -14692
rect 20759 -14696 20799 -14692
rect 20833 -14696 20873 -14692
rect 20907 -14696 20947 -14692
rect 20981 -14696 21021 -14692
rect 21055 -14696 21095 -14692
rect 21129 -14696 21169 -14692
rect 21203 -14696 21243 -14692
rect 21277 -14696 21317 -14692
rect 21351 -14696 21391 -14692
rect 21425 -14696 21465 -14692
rect 21499 -14696 21539 -14692
rect 21573 -14696 21613 -14692
rect 21647 -14696 21687 -14692
rect 21721 -14696 21761 -14692
rect 21795 -14696 21834 -14692
rect 21868 -14696 21907 -14692
rect 21941 -14696 21979 -14692
rect 22013 -14695 22051 -14691
rect 20708 -14726 20725 -14696
rect 20777 -14726 20799 -14696
rect 20846 -14726 20873 -14696
rect 20915 -14726 20947 -14696
rect 20708 -14730 20743 -14726
rect 20777 -14730 20812 -14726
rect 20846 -14730 20881 -14726
rect 20915 -14730 20950 -14726
rect 20984 -14730 21019 -14696
rect 21055 -14726 21088 -14696
rect 21129 -14726 21157 -14696
rect 21203 -14726 21226 -14696
rect 21277 -14726 21295 -14696
rect 21351 -14726 21364 -14696
rect 21425 -14726 21433 -14696
rect 21499 -14726 21502 -14696
rect 21053 -14730 21088 -14726
rect 21122 -14730 21157 -14726
rect 21191 -14730 21226 -14726
rect 21260 -14730 21295 -14726
rect 21329 -14730 21364 -14726
rect 21398 -14730 21433 -14726
rect 21467 -14730 21502 -14726
rect 21536 -14726 21539 -14696
rect 21536 -14730 21571 -14726
rect 20708 -14764 21571 -14730
rect 21945 -14729 21979 -14696
rect 22013 -14729 22047 -14695
rect 22085 -14725 22091 -14691
rect 22081 -14729 22091 -14725
rect 21945 -14764 22091 -14729
rect 20708 -14798 20725 -14764
rect 20777 -14798 20799 -14764
rect 20846 -14798 20873 -14764
rect 20915 -14798 20947 -14764
rect 20984 -14798 21019 -14764
rect 21055 -14798 21088 -14764
rect 21129 -14798 21157 -14764
rect 21203 -14798 21226 -14764
rect 21277 -14798 21295 -14764
rect 21351 -14798 21364 -14764
rect 21425 -14798 21433 -14764
rect 21499 -14798 21502 -14764
rect 21536 -14798 21539 -14764
rect 22013 -14798 22047 -14764
rect 22085 -14798 22091 -14764
rect 20708 -14832 21571 -14798
rect 20708 -14836 20743 -14832
rect 20777 -14836 20812 -14832
rect 20846 -14836 20881 -14832
rect 20915 -14836 20950 -14832
rect 20708 -14866 20725 -14836
rect 20777 -14866 20799 -14836
rect 20846 -14866 20873 -14836
rect 20915 -14866 20947 -14836
rect 20984 -14866 21019 -14832
rect 21053 -14836 21088 -14832
rect 21122 -14836 21157 -14832
rect 21191 -14836 21226 -14832
rect 21260 -14836 21295 -14832
rect 21329 -14836 21364 -14832
rect 21398 -14836 21433 -14832
rect 21467 -14836 21502 -14832
rect 21055 -14866 21088 -14836
rect 21129 -14866 21157 -14836
rect 21203 -14866 21226 -14836
rect 21277 -14866 21295 -14836
rect 21351 -14866 21364 -14836
rect 21425 -14866 21433 -14836
rect 21499 -14866 21502 -14836
rect 21536 -14836 21571 -14832
rect 21536 -14866 21539 -14836
rect 22013 -14866 22091 -14798
rect 20640 -14870 20651 -14866
rect 20685 -14870 20725 -14866
rect 20759 -14870 20799 -14866
rect 20833 -14870 20873 -14866
rect 20907 -14870 20947 -14866
rect 20981 -14870 21021 -14866
rect 21055 -14870 21095 -14866
rect 21129 -14870 21169 -14866
rect 21203 -14870 21243 -14866
rect 21277 -14870 21317 -14866
rect 21351 -14870 21391 -14866
rect 21425 -14870 21465 -14866
rect 21499 -14870 21539 -14866
rect 21573 -14870 21613 -14866
rect 21647 -14870 21686 -14866
rect 21720 -14870 21759 -14866
rect 21793 -14870 21832 -14866
rect 21866 -14870 21905 -14866
rect 21939 -14870 21978 -14866
rect 22012 -14870 22091 -14866
rect 20640 -14876 22091 -14870
rect 20470 -17308 20640 -17274
<< viali >>
rect 100 386 134 420
rect 172 386 204 420
rect 204 386 206 420
rect 244 386 272 420
rect 272 386 278 420
rect 316 386 340 420
rect 340 386 350 420
rect 388 386 408 420
rect 408 386 422 420
rect 460 386 476 420
rect 476 386 494 420
rect 532 386 544 420
rect 544 386 566 420
rect 604 386 612 420
rect 612 386 638 420
rect 676 386 680 420
rect 680 386 710 420
rect 748 386 782 420
rect 820 386 850 420
rect 850 386 854 420
rect 892 386 918 420
rect 918 386 926 420
rect 964 386 986 420
rect 986 386 998 420
rect 1036 386 1054 420
rect 1054 386 1070 420
rect 1194 386 1210 420
rect 1210 386 1228 420
rect 1266 386 1278 420
rect 1278 386 1300 420
rect 1338 386 1346 420
rect 1346 386 1372 420
rect 1410 386 1414 420
rect 1414 386 1444 420
rect 1482 386 1516 420
rect 1554 386 1584 420
rect 1584 386 1588 420
rect 1626 386 1652 420
rect 1652 386 1660 420
rect 1698 386 1720 420
rect 1720 386 1732 420
rect 1770 386 1788 420
rect 1788 386 1804 420
rect 1842 386 1856 420
rect 1856 386 1876 420
rect 1914 386 1924 420
rect 1924 386 1948 420
rect 1986 386 1992 420
rect 1992 386 2020 420
rect 2058 386 2060 420
rect 2060 386 2092 420
rect 2130 386 2164 420
rect 2364 386 2398 420
rect 2436 386 2468 420
rect 2468 386 2470 420
rect 2508 386 2536 420
rect 2536 386 2542 420
rect 2580 386 2604 420
rect 2604 386 2614 420
rect 2652 386 2672 420
rect 2672 386 2686 420
rect 2724 386 2740 420
rect 2740 386 2758 420
rect 2796 386 2808 420
rect 2808 386 2830 420
rect 2868 386 2876 420
rect 2876 386 2902 420
rect 2940 386 2944 420
rect 2944 386 2974 420
rect 3012 386 3046 420
rect 3084 386 3114 420
rect 3114 386 3118 420
rect 3156 386 3182 420
rect 3182 386 3190 420
rect 3228 386 3250 420
rect 3250 386 3262 420
rect 3300 386 3318 420
rect 3318 386 3334 420
rect 3458 386 3474 420
rect 3474 386 3492 420
rect 3530 386 3542 420
rect 3542 386 3564 420
rect 3602 386 3610 420
rect 3610 386 3636 420
rect 3674 386 3678 420
rect 3678 386 3708 420
rect 3746 386 3780 420
rect 3818 386 3848 420
rect 3848 386 3852 420
rect 3890 386 3916 420
rect 3916 386 3924 420
rect 3962 386 3984 420
rect 3984 386 3996 420
rect 4034 386 4052 420
rect 4052 386 4068 420
rect 4106 386 4120 420
rect 4120 386 4140 420
rect 4178 386 4188 420
rect 4188 386 4212 420
rect 4250 386 4256 420
rect 4256 386 4284 420
rect 4322 386 4324 420
rect 4324 386 4356 420
rect 4394 386 4428 420
rect 4628 386 4662 420
rect 4700 386 4732 420
rect 4732 386 4734 420
rect 4772 386 4800 420
rect 4800 386 4806 420
rect 4844 386 4868 420
rect 4868 386 4878 420
rect 4916 386 4936 420
rect 4936 386 4950 420
rect 4988 386 5004 420
rect 5004 386 5022 420
rect 5060 386 5072 420
rect 5072 386 5094 420
rect 5132 386 5140 420
rect 5140 386 5166 420
rect 5204 386 5208 420
rect 5208 386 5238 420
rect 5276 386 5310 420
rect 5348 386 5378 420
rect 5378 386 5382 420
rect 5420 386 5446 420
rect 5446 386 5454 420
rect 5492 386 5514 420
rect 5514 386 5526 420
rect 5564 386 5582 420
rect 5582 386 5598 420
rect 5722 386 5738 420
rect 5738 386 5756 420
rect 5794 386 5806 420
rect 5806 386 5828 420
rect 5866 386 5874 420
rect 5874 386 5900 420
rect 5938 386 5942 420
rect 5942 386 5972 420
rect 6010 386 6044 420
rect 6082 386 6112 420
rect 6112 386 6116 420
rect 6154 386 6180 420
rect 6180 386 6188 420
rect 6226 386 6248 420
rect 6248 386 6260 420
rect 6298 386 6316 420
rect 6316 386 6332 420
rect 6370 386 6384 420
rect 6384 386 6404 420
rect 6442 386 6452 420
rect 6452 386 6476 420
rect 6514 386 6520 420
rect 6520 386 6548 420
rect 6586 386 6588 420
rect 6588 386 6620 420
rect 6658 386 6692 420
rect 100 230 134 264
rect 172 230 204 264
rect 204 230 206 264
rect 244 230 272 264
rect 272 230 278 264
rect 316 230 340 264
rect 340 230 350 264
rect 388 230 408 264
rect 408 230 422 264
rect 460 230 476 264
rect 476 230 494 264
rect 532 230 544 264
rect 544 230 566 264
rect 604 230 612 264
rect 612 230 638 264
rect 676 230 680 264
rect 680 230 710 264
rect 748 230 782 264
rect 820 230 850 264
rect 850 230 854 264
rect 892 230 918 264
rect 918 230 926 264
rect 964 230 986 264
rect 986 230 998 264
rect 1036 230 1054 264
rect 1054 230 1070 264
rect -53 152 -19 186
rect 1194 230 1210 264
rect 1210 230 1228 264
rect 1266 230 1278 264
rect 1278 230 1300 264
rect 1338 230 1346 264
rect 1346 230 1372 264
rect 1410 230 1414 264
rect 1414 230 1444 264
rect 1482 230 1516 264
rect 1554 230 1584 264
rect 1584 230 1588 264
rect 1626 230 1652 264
rect 1652 230 1660 264
rect 1698 230 1720 264
rect 1720 230 1732 264
rect 1770 230 1788 264
rect 1788 230 1804 264
rect 1842 230 1856 264
rect 1856 230 1876 264
rect 1914 230 1924 264
rect 1924 230 1948 264
rect 1986 230 1992 264
rect 1992 230 2020 264
rect 2058 230 2060 264
rect 2060 230 2092 264
rect 2130 230 2164 264
rect 19 152 53 186
rect 1079 152 1113 186
rect 2364 230 2398 264
rect 2436 230 2468 264
rect 2468 230 2470 264
rect 2508 230 2536 264
rect 2536 230 2542 264
rect 2580 230 2604 264
rect 2604 230 2614 264
rect 2652 230 2672 264
rect 2672 230 2686 264
rect 2724 230 2740 264
rect 2740 230 2758 264
rect 2796 230 2808 264
rect 2808 230 2830 264
rect 2868 230 2876 264
rect 2876 230 2902 264
rect 2940 230 2944 264
rect 2944 230 2974 264
rect 3012 230 3046 264
rect 3084 230 3114 264
rect 3114 230 3118 264
rect 3156 230 3182 264
rect 3182 230 3190 264
rect 3228 230 3250 264
rect 3250 230 3262 264
rect 3300 230 3318 264
rect 3318 230 3334 264
rect 1151 152 1185 186
rect 2211 152 2245 186
rect 3458 230 3474 264
rect 3474 230 3492 264
rect 3530 230 3542 264
rect 3542 230 3564 264
rect 3602 230 3610 264
rect 3610 230 3636 264
rect 3674 230 3678 264
rect 3678 230 3708 264
rect 3746 230 3780 264
rect 3818 230 3848 264
rect 3848 230 3852 264
rect 3890 230 3916 264
rect 3916 230 3924 264
rect 3962 230 3984 264
rect 3984 230 3996 264
rect 4034 230 4052 264
rect 4052 230 4068 264
rect 4106 230 4120 264
rect 4120 230 4140 264
rect 4178 230 4188 264
rect 4188 230 4212 264
rect 4250 230 4256 264
rect 4256 230 4284 264
rect 4322 230 4324 264
rect 4324 230 4356 264
rect 4394 230 4428 264
rect 2283 152 2317 186
rect 3343 152 3377 186
rect 4628 230 4662 264
rect 4700 230 4732 264
rect 4732 230 4734 264
rect 4772 230 4800 264
rect 4800 230 4806 264
rect 4844 230 4868 264
rect 4868 230 4878 264
rect 4916 230 4936 264
rect 4936 230 4950 264
rect 4988 230 5004 264
rect 5004 230 5022 264
rect 5060 230 5072 264
rect 5072 230 5094 264
rect 5132 230 5140 264
rect 5140 230 5166 264
rect 5204 230 5208 264
rect 5208 230 5238 264
rect 5276 230 5310 264
rect 5348 230 5378 264
rect 5378 230 5382 264
rect 5420 230 5446 264
rect 5446 230 5454 264
rect 5492 230 5514 264
rect 5514 230 5526 264
rect 5564 230 5582 264
rect 5582 230 5598 264
rect 3415 152 3449 186
rect 4475 152 4509 186
rect 5722 230 5738 264
rect 5738 230 5756 264
rect 5794 230 5806 264
rect 5806 230 5828 264
rect 5866 230 5874 264
rect 5874 230 5900 264
rect 5938 230 5942 264
rect 5942 230 5972 264
rect 6010 230 6044 264
rect 6082 230 6112 264
rect 6112 230 6116 264
rect 6154 230 6180 264
rect 6180 230 6188 264
rect 6226 230 6248 264
rect 6248 230 6260 264
rect 6298 230 6316 264
rect 6316 230 6332 264
rect 6370 230 6384 264
rect 6384 230 6404 264
rect 6442 230 6452 264
rect 6452 230 6476 264
rect 6514 230 6520 264
rect 6520 230 6548 264
rect 6586 230 6588 264
rect 6588 230 6620 264
rect 6658 230 6692 264
rect 4547 152 4581 186
rect 5607 152 5641 186
rect 5679 152 5713 186
rect 6739 152 6773 186
rect 6811 152 6845 186
rect 100 74 134 108
rect 172 74 204 108
rect 204 74 206 108
rect 244 74 272 108
rect 272 74 278 108
rect 316 74 340 108
rect 340 74 350 108
rect 388 74 408 108
rect 408 74 422 108
rect 460 74 476 108
rect 476 74 494 108
rect 532 74 544 108
rect 544 74 566 108
rect 604 74 612 108
rect 612 74 638 108
rect 676 74 680 108
rect 680 74 710 108
rect 748 74 782 108
rect 820 74 850 108
rect 850 74 854 108
rect 892 74 918 108
rect 918 74 926 108
rect 964 74 986 108
rect 986 74 998 108
rect 1036 74 1054 108
rect 1054 74 1070 108
rect 1194 74 1210 108
rect 1210 74 1228 108
rect 1266 74 1278 108
rect 1278 74 1300 108
rect 1338 74 1346 108
rect 1346 74 1372 108
rect 1410 74 1414 108
rect 1414 74 1444 108
rect 1482 74 1516 108
rect 1554 74 1584 108
rect 1584 74 1588 108
rect 1626 74 1652 108
rect 1652 74 1660 108
rect 1698 74 1720 108
rect 1720 74 1732 108
rect 1770 74 1788 108
rect 1788 74 1804 108
rect 1842 74 1856 108
rect 1856 74 1876 108
rect 1914 74 1924 108
rect 1924 74 1948 108
rect 1986 74 1992 108
rect 1992 74 2020 108
rect 2058 74 2060 108
rect 2060 74 2092 108
rect 2130 74 2164 108
rect 2364 74 2398 108
rect 2436 74 2468 108
rect 2468 74 2470 108
rect 2508 74 2536 108
rect 2536 74 2542 108
rect 2580 74 2604 108
rect 2604 74 2614 108
rect 2652 74 2672 108
rect 2672 74 2686 108
rect 2724 74 2740 108
rect 2740 74 2758 108
rect 2796 74 2808 108
rect 2808 74 2830 108
rect 2868 74 2876 108
rect 2876 74 2902 108
rect 2940 74 2944 108
rect 2944 74 2974 108
rect 3012 74 3046 108
rect 3084 74 3114 108
rect 3114 74 3118 108
rect 3156 74 3182 108
rect 3182 74 3190 108
rect 3228 74 3250 108
rect 3250 74 3262 108
rect 3300 74 3318 108
rect 3318 74 3334 108
rect 3458 74 3474 108
rect 3474 74 3492 108
rect 3530 74 3542 108
rect 3542 74 3564 108
rect 3602 74 3610 108
rect 3610 74 3636 108
rect 3674 74 3678 108
rect 3678 74 3708 108
rect 3746 74 3780 108
rect 3818 74 3848 108
rect 3848 74 3852 108
rect 3890 74 3916 108
rect 3916 74 3924 108
rect 3962 74 3984 108
rect 3984 74 3996 108
rect 4034 74 4052 108
rect 4052 74 4068 108
rect 4106 74 4120 108
rect 4120 74 4140 108
rect 4178 74 4188 108
rect 4188 74 4212 108
rect 4250 74 4256 108
rect 4256 74 4284 108
rect 4322 74 4324 108
rect 4324 74 4356 108
rect 4394 74 4428 108
rect 4628 74 4662 108
rect 4700 74 4732 108
rect 4732 74 4734 108
rect 4772 74 4800 108
rect 4800 74 4806 108
rect 4844 74 4868 108
rect 4868 74 4878 108
rect 4916 74 4936 108
rect 4936 74 4950 108
rect 4988 74 5004 108
rect 5004 74 5022 108
rect 5060 74 5072 108
rect 5072 74 5094 108
rect 5132 74 5140 108
rect 5140 74 5166 108
rect 5204 74 5208 108
rect 5208 74 5238 108
rect 5276 74 5310 108
rect 5348 74 5378 108
rect 5378 74 5382 108
rect 5420 74 5446 108
rect 5446 74 5454 108
rect 5492 74 5514 108
rect 5514 74 5526 108
rect 5564 74 5582 108
rect 5582 74 5598 108
rect 5722 74 5738 108
rect 5738 74 5756 108
rect 5794 74 5806 108
rect 5806 74 5828 108
rect 5866 74 5874 108
rect 5874 74 5900 108
rect 5938 74 5942 108
rect 5942 74 5972 108
rect 6010 74 6044 108
rect 6082 74 6112 108
rect 6112 74 6116 108
rect 6154 74 6180 108
rect 6180 74 6188 108
rect 6226 74 6248 108
rect 6248 74 6260 108
rect 6298 74 6316 108
rect 6316 74 6332 108
rect 6370 74 6384 108
rect 6384 74 6404 108
rect 6442 74 6452 108
rect 6452 74 6476 108
rect 6514 74 6520 108
rect 6520 74 6548 108
rect 6586 74 6588 108
rect 6588 74 6620 108
rect 6658 74 6692 108
rect 20824 -3702 20858 -3685
rect 20824 -3719 20858 -3702
rect 20824 -3804 20858 -3794
rect 20824 -3828 20858 -3804
rect 20980 -3459 21014 -3425
rect 20980 -3498 21014 -3497
rect 20980 -3531 21014 -3498
rect 21136 -3702 21170 -3685
rect 21136 -3719 21170 -3702
rect 21136 -3804 21170 -3794
rect 21136 -3828 21170 -3804
rect 20651 -7898 20685 -7893
rect 20724 -7898 20758 -7893
rect 20797 -7898 20831 -7893
rect 20870 -7898 20904 -7893
rect 20943 -7898 20977 -7893
rect 21017 -7898 21051 -7893
rect 21091 -7898 21125 -7893
rect 21165 -7898 21199 -7893
rect 21239 -7898 21273 -7893
rect 21313 -7898 21347 -7893
rect 21387 -7898 21421 -7893
rect 20651 -7927 20674 -7898
rect 20674 -7927 20685 -7898
rect 20724 -7927 20758 -7898
rect 20797 -7927 20831 -7898
rect 20870 -7927 20904 -7898
rect 20943 -7927 20977 -7898
rect 21017 -7927 21051 -7898
rect 21091 -7927 21116 -7898
rect 21116 -7927 21125 -7898
rect 21165 -7927 21185 -7898
rect 21185 -7927 21199 -7898
rect 21239 -7927 21254 -7898
rect 21254 -7927 21273 -7898
rect 21313 -7927 21323 -7898
rect 21323 -7927 21347 -7898
rect 21387 -7927 21392 -7898
rect 21392 -7927 21421 -7898
rect 21461 -7927 21495 -7893
rect 21535 -7898 21569 -7893
rect 21609 -7898 21643 -7893
rect 21683 -7898 21717 -7893
rect 21757 -7898 21791 -7893
rect 21831 -7898 21865 -7893
rect 21905 -7898 21939 -7893
rect 21979 -7898 22013 -7893
rect 21535 -7927 21565 -7898
rect 21565 -7927 21569 -7898
rect 21609 -7927 21634 -7898
rect 21634 -7927 21643 -7898
rect 21683 -7927 21703 -7898
rect 21703 -7927 21717 -7898
rect 21757 -7927 21772 -7898
rect 21772 -7927 21791 -7898
rect 21831 -7927 21841 -7898
rect 21841 -7927 21865 -7898
rect 21905 -7927 21910 -7898
rect 21910 -7927 21939 -7898
rect 21979 -7927 22013 -7898
rect 20651 -7999 20674 -7965
rect 20674 -7999 20685 -7965
rect 20724 -7999 20758 -7965
rect 20797 -7999 20831 -7965
rect 20870 -7999 20904 -7965
rect 20943 -7999 20977 -7965
rect 21017 -7999 21051 -7965
rect 21091 -7999 21116 -7965
rect 21116 -7999 21125 -7965
rect 21165 -7966 21199 -7965
rect 21239 -7966 21273 -7965
rect 21313 -7966 21347 -7965
rect 21387 -7966 21421 -7965
rect 21165 -7999 21185 -7966
rect 21185 -7999 21199 -7966
rect 21239 -7999 21254 -7966
rect 21254 -7999 21273 -7966
rect 21313 -7999 21323 -7966
rect 21323 -7999 21347 -7966
rect 21387 -7999 21392 -7966
rect 21392 -7999 21421 -7966
rect 21461 -7999 21495 -7965
rect 21535 -7966 21569 -7965
rect 21609 -7966 21643 -7965
rect 21683 -7966 21717 -7965
rect 21757 -7966 21791 -7965
rect 21831 -7966 21865 -7965
rect 21905 -7966 21939 -7965
rect 21979 -7966 22085 -7965
rect 21535 -7999 21565 -7966
rect 21565 -7999 21569 -7966
rect 21609 -7999 21634 -7966
rect 21634 -7999 21643 -7966
rect 21683 -7999 21703 -7966
rect 21703 -7999 21717 -7966
rect 21757 -7999 21772 -7966
rect 21772 -7999 21791 -7966
rect 21831 -7999 21841 -7966
rect 21841 -7999 21865 -7966
rect 21905 -7999 21910 -7966
rect 21910 -7999 21939 -7966
rect 20651 -8068 20674 -8037
rect 20674 -8068 20685 -8037
rect 20724 -8068 20758 -8037
rect 20797 -8068 20831 -8037
rect 20871 -8068 20905 -8037
rect 20945 -8068 20979 -8037
rect 21019 -8068 21048 -8037
rect 21048 -8068 21053 -8037
rect 21093 -8068 21117 -8037
rect 21117 -8068 21127 -8037
rect 21167 -8068 21186 -8037
rect 21186 -8068 21201 -8037
rect 21241 -8068 21255 -8037
rect 21255 -8068 21275 -8037
rect 21315 -8068 21324 -8037
rect 21324 -8068 21349 -8037
rect 21389 -8068 21393 -8037
rect 21393 -8068 21423 -8037
rect 20651 -8071 20685 -8068
rect 20724 -8071 20758 -8068
rect 20797 -8071 20831 -8068
rect 20871 -8071 20905 -8068
rect 20945 -8071 20979 -8068
rect 21019 -8071 21053 -8068
rect 21093 -8071 21127 -8068
rect 21167 -8071 21201 -8068
rect 21241 -8071 21275 -8068
rect 21315 -8071 21349 -8068
rect 21389 -8071 21423 -8068
rect 21463 -8071 21497 -8037
rect 21979 -8037 22081 -7966
rect 21537 -8068 21566 -8037
rect 21566 -8068 21571 -8037
rect 21611 -8068 21635 -8037
rect 21635 -8068 21645 -8037
rect 21685 -8068 21704 -8037
rect 21704 -8068 21719 -8037
rect 21759 -8068 21773 -8037
rect 21773 -8068 21793 -8037
rect 21833 -8068 21842 -8037
rect 21842 -8068 21867 -8037
rect 21537 -8071 21571 -8068
rect 21611 -8071 21645 -8068
rect 21685 -8071 21719 -8068
rect 21759 -8071 21793 -8068
rect 21833 -8071 21867 -8068
rect 21223 -10018 21257 -10006
rect 21223 -10040 21257 -10018
rect 21223 -10086 21257 -10078
rect 21223 -10112 21257 -10086
rect 21223 -10154 21257 -10150
rect 21223 -10184 21257 -10154
rect 21223 -10256 21257 -10222
rect 21223 -10324 21257 -10294
rect 21223 -10328 21257 -10324
rect 21223 -10392 21257 -10366
rect 21223 -10400 21257 -10392
rect 21223 -10460 21257 -10438
rect 21223 -10472 21257 -10460
rect 21223 -10528 21257 -10510
rect 21223 -10544 21257 -10528
rect 21379 -10018 21413 -10006
rect 21379 -10040 21413 -10018
rect 21379 -10086 21413 -10078
rect 21379 -10112 21413 -10086
rect 21379 -10154 21413 -10150
rect 21379 -10184 21413 -10154
rect 21379 -10256 21413 -10222
rect 21379 -10324 21413 -10294
rect 21379 -10328 21413 -10324
rect 21379 -10392 21413 -10366
rect 21379 -10400 21413 -10392
rect 21379 -10460 21413 -10438
rect 21379 -10472 21413 -10460
rect 21379 -10528 21413 -10510
rect 21379 -10544 21413 -10528
rect 21535 -10018 21569 -10006
rect 21535 -10040 21569 -10018
rect 21535 -10086 21569 -10078
rect 21535 -10112 21569 -10086
rect 21535 -10154 21569 -10150
rect 21535 -10184 21569 -10154
rect 21535 -10256 21569 -10222
rect 21535 -10324 21569 -10294
rect 21535 -10328 21569 -10324
rect 21535 -10392 21569 -10366
rect 21535 -10400 21569 -10392
rect 21535 -10460 21569 -10438
rect 21535 -10472 21569 -10460
rect 21535 -10528 21569 -10510
rect 21535 -10544 21569 -10528
rect 21301 -10587 21335 -10553
rect 21301 -10659 21335 -10625
rect 21907 -10176 21911 -8037
rect 21911 -10176 22081 -8037
rect 21907 -10211 21979 -10176
rect 21907 -10245 21911 -10211
rect 21911 -10245 21945 -10211
rect 21945 -10244 21979 -10211
rect 21979 -10244 22081 -10176
rect 22081 -10244 22085 -7966
rect 21945 -10245 22085 -10244
rect 21907 -10279 22085 -10245
rect 21907 -10280 21979 -10279
rect 21907 -10314 21911 -10280
rect 21911 -10314 21945 -10280
rect 21945 -10313 21979 -10280
rect 21979 -10313 22013 -10279
rect 22013 -10313 22047 -10279
rect 22047 -10313 22081 -10279
rect 22081 -10313 22085 -10279
rect 21945 -10314 22085 -10313
rect 21907 -10348 22085 -10314
rect 21907 -10349 21979 -10348
rect 21907 -10383 21911 -10349
rect 21911 -10383 21945 -10349
rect 21945 -10382 21979 -10349
rect 21979 -10382 22013 -10348
rect 22013 -10382 22047 -10348
rect 22047 -10382 22081 -10348
rect 22081 -10382 22085 -10348
rect 21945 -10383 22085 -10382
rect 21907 -10417 22085 -10383
rect 21907 -10418 21979 -10417
rect 21907 -10452 21911 -10418
rect 21911 -10452 21945 -10418
rect 21945 -10451 21979 -10418
rect 21979 -10451 22013 -10417
rect 22013 -10451 22047 -10417
rect 22047 -10451 22081 -10417
rect 22081 -10451 22085 -10417
rect 21945 -10452 22085 -10451
rect 21907 -10486 22085 -10452
rect 21907 -10487 21979 -10486
rect 21907 -10521 21911 -10487
rect 21911 -10521 21945 -10487
rect 21945 -10520 21979 -10487
rect 21979 -10520 22013 -10486
rect 22013 -10520 22047 -10486
rect 22047 -10520 22081 -10486
rect 22081 -10520 22085 -10486
rect 21945 -10521 22085 -10520
rect 21907 -10555 22085 -10521
rect 21907 -10556 21979 -10555
rect 21907 -10590 21911 -10556
rect 21911 -10590 21945 -10556
rect 21945 -10589 21979 -10556
rect 21979 -10589 22013 -10555
rect 22013 -10589 22047 -10555
rect 22047 -10589 22081 -10555
rect 22081 -10589 22085 -10555
rect 21945 -10590 22085 -10589
rect 21907 -10624 22085 -10590
rect 21907 -10625 21979 -10624
rect 21907 -10659 21911 -10625
rect 21911 -10659 21945 -10625
rect 21945 -10658 21979 -10625
rect 21979 -10658 22013 -10624
rect 22013 -10658 22047 -10624
rect 22047 -10658 22081 -10624
rect 22081 -10658 22085 -10624
rect 21945 -10659 22085 -10658
rect 21907 -10693 22085 -10659
rect 21907 -10694 21979 -10693
rect 21907 -10728 21911 -10694
rect 21911 -10728 21945 -10694
rect 21945 -10727 21979 -10694
rect 21979 -10727 22013 -10693
rect 22013 -10727 22047 -10693
rect 22047 -10727 22081 -10693
rect 22081 -10727 22085 -10693
rect 21945 -10728 22085 -10727
rect 21907 -10762 22085 -10728
rect 21907 -10763 21979 -10762
rect 21907 -10797 21911 -10763
rect 21911 -10797 21945 -10763
rect 21945 -10796 21979 -10763
rect 21979 -10796 22013 -10762
rect 22013 -10796 22047 -10762
rect 22047 -10796 22081 -10762
rect 22081 -10796 22085 -10762
rect 21945 -10797 22085 -10796
rect 21907 -10831 22085 -10797
rect 21907 -10832 21979 -10831
rect 21907 -10866 21911 -10832
rect 21911 -10866 21945 -10832
rect 21945 -10865 21979 -10832
rect 21979 -10865 22013 -10831
rect 22013 -10865 22047 -10831
rect 22047 -10865 22081 -10831
rect 22081 -10865 22085 -10831
rect 21945 -10866 22085 -10865
rect 21907 -10900 22085 -10866
rect 21907 -10901 21979 -10900
rect 21907 -10935 21911 -10901
rect 21911 -10935 21945 -10901
rect 21945 -10934 21979 -10901
rect 21979 -10934 22013 -10900
rect 22013 -10934 22047 -10900
rect 22047 -10934 22081 -10900
rect 22081 -10934 22085 -10900
rect 21945 -10935 22085 -10934
rect 21907 -10969 22085 -10935
rect 21907 -10970 21979 -10969
rect 21907 -11004 21911 -10970
rect 21911 -11004 21945 -10970
rect 21945 -11003 21979 -10970
rect 21979 -11003 22013 -10969
rect 22013 -11003 22047 -10969
rect 22047 -11003 22081 -10969
rect 22081 -11003 22085 -10969
rect 21945 -11004 22085 -11003
rect 21907 -11038 22085 -11004
rect 21907 -11039 21979 -11038
rect 21907 -11073 21911 -11039
rect 21911 -11073 21945 -11039
rect 21945 -11072 21979 -11039
rect 21979 -11072 22013 -11038
rect 22013 -11072 22047 -11038
rect 22047 -11072 22081 -11038
rect 22081 -11072 22085 -11038
rect 21945 -11073 22085 -11072
rect 21907 -11107 22085 -11073
rect 21907 -11108 21979 -11107
rect 21907 -11142 21911 -11108
rect 21911 -11142 21945 -11108
rect 21945 -11141 21979 -11108
rect 21979 -11141 22013 -11107
rect 22013 -11141 22047 -11107
rect 22047 -11141 22081 -11107
rect 22081 -11141 22085 -11107
rect 21945 -11142 22085 -11141
rect 21907 -11176 22085 -11142
rect 21907 -11177 21979 -11176
rect 21907 -11211 21911 -11177
rect 21911 -11211 21945 -11177
rect 21945 -11210 21979 -11177
rect 21979 -11210 22013 -11176
rect 22013 -11210 22047 -11176
rect 22047 -11210 22081 -11176
rect 22081 -11210 22085 -11176
rect 21945 -11211 22085 -11210
rect 21907 -11245 22085 -11211
rect 21907 -11246 21979 -11245
rect 21907 -11280 21911 -11246
rect 21911 -11280 21945 -11246
rect 21945 -11279 21979 -11246
rect 21979 -11279 22013 -11245
rect 22013 -11279 22047 -11245
rect 22047 -11279 22081 -11245
rect 22081 -11279 22085 -11245
rect 21945 -11280 22085 -11279
rect 21907 -11314 22085 -11280
rect 21907 -11315 21979 -11314
rect 21907 -11349 21911 -11315
rect 21911 -11349 21945 -11315
rect 21945 -11348 21979 -11315
rect 21979 -11348 22013 -11314
rect 22013 -11348 22047 -11314
rect 22047 -11348 22081 -11314
rect 22081 -11348 22085 -11314
rect 21945 -11349 22085 -11348
rect 21907 -11383 22085 -11349
rect 21907 -11384 21979 -11383
rect 21907 -11418 21911 -11384
rect 21911 -11418 21945 -11384
rect 21945 -11417 21979 -11384
rect 21979 -11417 22013 -11383
rect 22013 -11417 22047 -11383
rect 22047 -11417 22081 -11383
rect 22081 -11417 22085 -11383
rect 21945 -11418 22085 -11417
rect 21907 -11452 22085 -11418
rect 21907 -11453 21979 -11452
rect 21907 -11487 21911 -11453
rect 21911 -11487 21945 -11453
rect 21945 -11486 21979 -11453
rect 21979 -11486 22013 -11452
rect 22013 -11486 22047 -11452
rect 22047 -11486 22081 -11452
rect 22081 -11486 22085 -11452
rect 21945 -11487 22085 -11486
rect 21907 -11521 22085 -11487
rect 21907 -11522 21979 -11521
rect 21907 -11556 21911 -11522
rect 21911 -11556 21945 -11522
rect 21945 -11555 21979 -11522
rect 21979 -11555 22013 -11521
rect 22013 -11555 22047 -11521
rect 22047 -11555 22081 -11521
rect 22081 -11555 22085 -11521
rect 21945 -11556 22085 -11555
rect 21907 -11590 22085 -11556
rect 21907 -11591 21979 -11590
rect 21907 -11625 21911 -11591
rect 21911 -11625 21945 -11591
rect 21945 -11624 21979 -11591
rect 21979 -11624 22013 -11590
rect 22013 -11624 22047 -11590
rect 22047 -11624 22081 -11590
rect 22081 -11624 22085 -11590
rect 21945 -11625 22085 -11624
rect 21907 -11659 22085 -11625
rect 21907 -11660 21979 -11659
rect 21907 -11694 21911 -11660
rect 21911 -11694 21945 -11660
rect 21945 -11693 21979 -11660
rect 21979 -11693 22013 -11659
rect 22013 -11693 22047 -11659
rect 22047 -11693 22081 -11659
rect 22081 -11693 22085 -11659
rect 21945 -11694 22085 -11693
rect 21907 -11728 22085 -11694
rect 21907 -11729 21979 -11728
rect 21907 -11763 21911 -11729
rect 21911 -11763 21945 -11729
rect 21945 -11762 21979 -11729
rect 21979 -11762 22013 -11728
rect 22013 -11762 22047 -11728
rect 22047 -11762 22081 -11728
rect 22081 -11762 22085 -11728
rect 21945 -11763 22085 -11762
rect 21907 -11797 22085 -11763
rect 21907 -11798 21979 -11797
rect 21907 -11832 21911 -11798
rect 21911 -11832 21945 -11798
rect 21945 -11831 21979 -11798
rect 21979 -11831 22013 -11797
rect 22013 -11831 22047 -11797
rect 22047 -11831 22081 -11797
rect 22081 -11831 22085 -11797
rect 21945 -11832 22085 -11831
rect 21907 -11866 22085 -11832
rect 21907 -11867 21979 -11866
rect 21907 -11901 21911 -11867
rect 21911 -11901 21945 -11867
rect 21945 -11900 21979 -11867
rect 21979 -11900 22013 -11866
rect 22013 -11900 22047 -11866
rect 22047 -11900 22081 -11866
rect 22081 -11900 22085 -11866
rect 21945 -11901 22085 -11900
rect 21907 -11935 22085 -11901
rect 21907 -11936 21979 -11935
rect 21907 -11970 21911 -11936
rect 21911 -11970 21945 -11936
rect 21945 -11969 21979 -11936
rect 21979 -11969 22013 -11935
rect 22013 -11969 22047 -11935
rect 22047 -11969 22081 -11935
rect 22081 -11969 22085 -11935
rect 21945 -11970 22085 -11969
rect 21907 -12004 22085 -11970
rect 21907 -12005 21979 -12004
rect 21907 -12039 21911 -12005
rect 21911 -12039 21945 -12005
rect 21945 -12038 21979 -12005
rect 21979 -12038 22013 -12004
rect 22013 -12038 22047 -12004
rect 22047 -12038 22081 -12004
rect 22081 -12038 22085 -12004
rect 21945 -12039 22085 -12038
rect 21907 -12073 22085 -12039
rect 21907 -12074 21979 -12073
rect 21907 -12108 21911 -12074
rect 21911 -12108 21945 -12074
rect 21945 -12107 21979 -12074
rect 21979 -12107 22013 -12073
rect 22013 -12107 22047 -12073
rect 22047 -12107 22081 -12073
rect 22081 -12107 22085 -12073
rect 21945 -12108 22085 -12107
rect 21907 -12142 22085 -12108
rect 21907 -12143 21979 -12142
rect 21907 -12177 21911 -12143
rect 21911 -12177 21945 -12143
rect 21945 -12176 21979 -12143
rect 21979 -12176 22013 -12142
rect 22013 -12176 22047 -12142
rect 22047 -12176 22081 -12142
rect 22081 -12176 22085 -12142
rect 21945 -12177 22085 -12176
rect 21907 -12211 22085 -12177
rect 21907 -12212 21979 -12211
rect 21907 -12246 21911 -12212
rect 21911 -12246 21945 -12212
rect 21945 -12245 21979 -12212
rect 21979 -12245 22013 -12211
rect 22013 -12245 22047 -12211
rect 22047 -12245 22081 -12211
rect 22081 -12245 22085 -12211
rect 21945 -12246 22085 -12245
rect 21907 -12280 22085 -12246
rect 21907 -12281 21979 -12280
rect 21907 -12315 21911 -12281
rect 21911 -12315 21945 -12281
rect 21945 -12314 21979 -12281
rect 21979 -12314 22013 -12280
rect 22013 -12314 22047 -12280
rect 22047 -12314 22081 -12280
rect 22081 -12314 22085 -12280
rect 21945 -12315 22085 -12314
rect 21907 -12349 22085 -12315
rect 21907 -12350 21979 -12349
rect 21907 -12384 21911 -12350
rect 21911 -12384 21945 -12350
rect 21945 -12383 21979 -12350
rect 21979 -12383 22013 -12349
rect 22013 -12383 22047 -12349
rect 22047 -12383 22081 -12349
rect 22081 -12383 22085 -12349
rect 21945 -12384 22085 -12383
rect 21907 -12418 22085 -12384
rect 21907 -12419 21979 -12418
rect 21907 -12453 21911 -12419
rect 21911 -12453 21945 -12419
rect 21945 -12452 21979 -12419
rect 21979 -12452 22013 -12418
rect 22013 -12452 22047 -12418
rect 22047 -12452 22081 -12418
rect 22081 -12452 22085 -12418
rect 21945 -12453 22085 -12452
rect 21907 -12463 22085 -12453
rect 21979 -12487 22085 -12463
rect 21907 -12522 21911 -12502
rect 21911 -12522 21941 -12502
rect 21979 -12521 22013 -12487
rect 22013 -12521 22047 -12487
rect 22047 -12521 22081 -12487
rect 22081 -12521 22085 -12487
rect 21907 -12536 21941 -12522
rect 21979 -12535 22085 -12521
rect 21907 -12591 21911 -12575
rect 21911 -12591 21941 -12575
rect 21979 -12590 22013 -12574
rect 22051 -12590 22081 -12574
rect 22081 -12590 22085 -12574
rect 21907 -12609 21941 -12591
rect 21979 -12608 22013 -12590
rect 22051 -12608 22085 -12590
rect 21907 -12660 21911 -12648
rect 21911 -12660 21941 -12648
rect 21979 -12659 22013 -12647
rect 22051 -12659 22081 -12647
rect 22081 -12659 22085 -12647
rect 21907 -12682 21941 -12660
rect 21979 -12681 22013 -12659
rect 22051 -12681 22085 -12659
rect 21907 -12729 21911 -12721
rect 21911 -12729 21941 -12721
rect 21979 -12728 22013 -12720
rect 22051 -12728 22081 -12720
rect 22081 -12728 22085 -12720
rect 21907 -12755 21941 -12729
rect 21979 -12754 22013 -12728
rect 22051 -12754 22085 -12728
rect 21907 -12798 21911 -12794
rect 21911 -12798 21941 -12794
rect 21979 -12797 22013 -12793
rect 22051 -12797 22081 -12793
rect 22081 -12797 22085 -12793
rect 21907 -12828 21941 -12798
rect 21979 -12827 22013 -12797
rect 22051 -12827 22085 -12797
rect 21907 -12901 21941 -12867
rect 21979 -12900 22013 -12866
rect 22051 -12900 22085 -12866
rect 21907 -12971 21941 -12940
rect 21979 -12970 22013 -12939
rect 22051 -12970 22085 -12939
rect 21907 -12974 21911 -12971
rect 21911 -12974 21941 -12971
rect 21979 -12973 22013 -12970
rect 22051 -12973 22081 -12970
rect 22081 -12973 22085 -12970
rect 21907 -13040 21941 -13013
rect 21979 -13039 22013 -13012
rect 22051 -13039 22085 -13012
rect 21907 -13047 21911 -13040
rect 21911 -13047 21941 -13040
rect 21979 -13046 22013 -13039
rect 22051 -13046 22081 -13039
rect 22081 -13046 22085 -13039
rect 21907 -13109 21941 -13086
rect 21979 -13108 22013 -13085
rect 22051 -13108 22085 -13085
rect 21907 -13120 21911 -13109
rect 21911 -13120 21941 -13109
rect 21979 -13119 22013 -13108
rect 22051 -13119 22081 -13108
rect 22081 -13119 22085 -13108
rect 21907 -13178 21941 -13159
rect 21979 -13177 22013 -13158
rect 22051 -13177 22085 -13158
rect 21907 -13193 21911 -13178
rect 21911 -13193 21941 -13178
rect 21979 -13192 22013 -13177
rect 22051 -13192 22081 -13177
rect 22081 -13192 22085 -13177
rect 21907 -13247 21941 -13232
rect 21979 -13246 22013 -13231
rect 22051 -13246 22085 -13231
rect 21907 -13266 21911 -13247
rect 21911 -13266 21941 -13247
rect 21979 -13265 22013 -13246
rect 22051 -13265 22081 -13246
rect 22081 -13265 22085 -13246
rect 21907 -13316 21941 -13305
rect 21979 -13315 22013 -13304
rect 22051 -13315 22085 -13304
rect 21907 -13339 21911 -13316
rect 21911 -13339 21941 -13316
rect 21979 -13338 22013 -13315
rect 22051 -13338 22081 -13315
rect 22081 -13338 22085 -13315
rect 21907 -13385 21941 -13378
rect 21979 -13384 22013 -13377
rect 22051 -13384 22085 -13377
rect 21907 -13412 21911 -13385
rect 21911 -13412 21941 -13385
rect 21979 -13411 22013 -13384
rect 22051 -13411 22081 -13384
rect 22081 -13411 22085 -13384
rect 21907 -13454 21941 -13451
rect 21979 -13453 22013 -13450
rect 22051 -13453 22085 -13450
rect 21907 -13485 21911 -13454
rect 21911 -13485 21941 -13454
rect 21979 -13484 22013 -13453
rect 22051 -13484 22081 -13453
rect 22081 -13484 22085 -13453
rect 21907 -13557 21911 -13524
rect 21911 -13557 21941 -13524
rect 21979 -13556 22013 -13523
rect 22051 -13556 22081 -13523
rect 22081 -13556 22085 -13523
rect 21979 -13557 22013 -13556
rect 22051 -13557 22085 -13556
rect 21907 -13558 21941 -13557
rect 21907 -13626 21911 -13597
rect 21911 -13626 21941 -13597
rect 21979 -13625 22013 -13596
rect 22051 -13625 22081 -13596
rect 22081 -13625 22085 -13596
rect 21907 -13631 21941 -13626
rect 21979 -13630 22013 -13625
rect 22051 -13630 22085 -13625
rect 21907 -13695 21911 -13670
rect 21911 -13695 21941 -13670
rect 21979 -13694 22013 -13669
rect 22051 -13694 22081 -13669
rect 22081 -13694 22085 -13669
rect 21907 -13704 21941 -13695
rect 21979 -13703 22013 -13694
rect 22051 -13703 22085 -13694
rect 21907 -13764 21911 -13743
rect 21911 -13764 21941 -13743
rect 21979 -13763 22013 -13742
rect 22051 -13763 22081 -13742
rect 22081 -13763 22085 -13742
rect 21907 -13777 21941 -13764
rect 21979 -13776 22013 -13763
rect 22051 -13776 22085 -13763
rect 21907 -13833 21911 -13816
rect 21911 -13833 21941 -13816
rect 21979 -13832 22013 -13815
rect 22051 -13832 22081 -13815
rect 22081 -13832 22085 -13815
rect 21907 -13850 21941 -13833
rect 21979 -13849 22013 -13832
rect 22051 -13849 22085 -13832
rect 21907 -13902 21911 -13889
rect 21911 -13902 21941 -13889
rect 21979 -13901 22013 -13888
rect 22051 -13901 22081 -13888
rect 22081 -13901 22085 -13888
rect 21907 -13923 21941 -13902
rect 21979 -13922 22013 -13901
rect 22051 -13922 22085 -13901
rect 21907 -13971 21911 -13962
rect 21911 -13971 21941 -13962
rect 21979 -13970 22013 -13961
rect 22051 -13970 22081 -13961
rect 22081 -13970 22085 -13961
rect 21907 -13996 21941 -13971
rect 21979 -13995 22013 -13970
rect 22051 -13995 22085 -13970
rect 21907 -14040 21911 -14035
rect 21911 -14040 21941 -14035
rect 21979 -14039 22013 -14034
rect 22051 -14039 22081 -14034
rect 22081 -14039 22085 -14034
rect 21907 -14069 21941 -14040
rect 21979 -14068 22013 -14039
rect 22051 -14068 22085 -14039
rect 21907 -14109 21911 -14108
rect 21911 -14109 21941 -14108
rect 21979 -14108 22013 -14107
rect 22051 -14108 22081 -14107
rect 22081 -14108 22085 -14107
rect 21907 -14142 21941 -14109
rect 21979 -14141 22013 -14108
rect 22051 -14141 22085 -14108
rect 21907 -14213 21941 -14181
rect 21979 -14212 22013 -14180
rect 22051 -14212 22085 -14180
rect 21907 -14215 21911 -14213
rect 21911 -14215 21941 -14213
rect 21979 -14214 22013 -14212
rect 22051 -14214 22081 -14212
rect 22081 -14214 22085 -14212
rect 21907 -14282 21941 -14254
rect 21979 -14281 22013 -14253
rect 22051 -14281 22085 -14253
rect 21907 -14288 21911 -14282
rect 21911 -14288 21941 -14282
rect 21979 -14287 22013 -14281
rect 22051 -14287 22081 -14281
rect 22081 -14287 22085 -14281
rect 21907 -14351 21941 -14327
rect 21979 -14350 22013 -14326
rect 22051 -14350 22085 -14326
rect 21907 -14361 21911 -14351
rect 21911 -14361 21941 -14351
rect 21979 -14360 22013 -14350
rect 22051 -14360 22081 -14350
rect 22081 -14360 22085 -14350
rect 21907 -14420 21941 -14400
rect 21979 -14419 22013 -14399
rect 22051 -14419 22085 -14399
rect 21907 -14434 21911 -14420
rect 21911 -14434 21941 -14420
rect 21979 -14433 22013 -14419
rect 22051 -14433 22081 -14419
rect 22081 -14433 22085 -14419
rect 21907 -14489 21941 -14473
rect 21979 -14488 22013 -14472
rect 22051 -14488 22085 -14472
rect 21907 -14507 21911 -14489
rect 21911 -14507 21941 -14489
rect 21979 -14506 22013 -14488
rect 22051 -14506 22081 -14488
rect 22081 -14506 22085 -14488
rect 21907 -14558 21941 -14546
rect 21979 -14557 22013 -14545
rect 22051 -14557 22085 -14545
rect 21907 -14580 21911 -14558
rect 21911 -14580 21941 -14558
rect 21979 -14579 22013 -14557
rect 22051 -14579 22081 -14557
rect 22081 -14579 22085 -14557
rect 21907 -14627 21941 -14619
rect 21979 -14626 22013 -14618
rect 22051 -14626 22085 -14618
rect 21907 -14653 21911 -14627
rect 21911 -14653 21941 -14627
rect 21979 -14652 22013 -14626
rect 22051 -14652 22081 -14626
rect 22081 -14652 22085 -14626
rect 20651 -14696 20685 -14692
rect 20725 -14696 20759 -14692
rect 20799 -14696 20833 -14692
rect 20873 -14696 20907 -14692
rect 20947 -14696 20981 -14692
rect 21021 -14696 21055 -14692
rect 21095 -14696 21129 -14692
rect 21169 -14696 21203 -14692
rect 21243 -14696 21277 -14692
rect 21317 -14696 21351 -14692
rect 21391 -14696 21425 -14692
rect 21465 -14696 21499 -14692
rect 21539 -14696 21573 -14692
rect 21613 -14696 21647 -14692
rect 21687 -14696 21721 -14692
rect 21761 -14696 21795 -14692
rect 21834 -14696 21868 -14692
rect 21907 -14696 21941 -14692
rect 21979 -14695 22013 -14691
rect 22051 -14695 22085 -14691
rect 20651 -14726 20685 -14696
rect 20725 -14726 20743 -14696
rect 20743 -14726 20759 -14696
rect 20799 -14726 20812 -14696
rect 20812 -14726 20833 -14696
rect 20873 -14726 20881 -14696
rect 20881 -14726 20907 -14696
rect 20947 -14726 20950 -14696
rect 20950 -14726 20981 -14696
rect 21021 -14726 21053 -14696
rect 21053 -14726 21055 -14696
rect 21095 -14726 21122 -14696
rect 21122 -14726 21129 -14696
rect 21169 -14726 21191 -14696
rect 21191 -14726 21203 -14696
rect 21243 -14726 21260 -14696
rect 21260 -14726 21277 -14696
rect 21317 -14726 21329 -14696
rect 21329 -14726 21351 -14696
rect 21391 -14726 21398 -14696
rect 21398 -14726 21425 -14696
rect 21465 -14726 21467 -14696
rect 21467 -14726 21499 -14696
rect 21539 -14726 21571 -14696
rect 21571 -14726 21573 -14696
rect 21613 -14726 21647 -14696
rect 21687 -14726 21721 -14696
rect 21761 -14726 21795 -14696
rect 21834 -14726 21868 -14696
rect 21907 -14726 21941 -14696
rect 21979 -14725 22013 -14695
rect 22051 -14725 22081 -14695
rect 22081 -14725 22085 -14695
rect 20651 -14798 20685 -14764
rect 20725 -14798 20743 -14764
rect 20743 -14798 20759 -14764
rect 20799 -14798 20812 -14764
rect 20812 -14798 20833 -14764
rect 20873 -14798 20881 -14764
rect 20881 -14798 20907 -14764
rect 20947 -14798 20950 -14764
rect 20950 -14798 20981 -14764
rect 21021 -14798 21053 -14764
rect 21053 -14798 21055 -14764
rect 21095 -14798 21122 -14764
rect 21122 -14798 21129 -14764
rect 21169 -14798 21191 -14764
rect 21191 -14798 21203 -14764
rect 21243 -14798 21260 -14764
rect 21260 -14798 21277 -14764
rect 21317 -14798 21329 -14764
rect 21329 -14798 21351 -14764
rect 21391 -14798 21398 -14764
rect 21398 -14798 21425 -14764
rect 21465 -14798 21467 -14764
rect 21467 -14798 21499 -14764
rect 21539 -14798 21571 -14764
rect 21571 -14798 21573 -14764
rect 21613 -14798 21647 -14764
rect 21686 -14798 21720 -14764
rect 21759 -14798 21793 -14764
rect 21832 -14798 21866 -14764
rect 21905 -14798 21939 -14764
rect 21979 -14798 22013 -14764
rect 22051 -14798 22081 -14764
rect 22081 -14798 22085 -14764
rect 20651 -14866 20685 -14836
rect 20725 -14866 20743 -14836
rect 20743 -14866 20759 -14836
rect 20799 -14866 20812 -14836
rect 20812 -14866 20833 -14836
rect 20873 -14866 20881 -14836
rect 20881 -14866 20907 -14836
rect 20947 -14866 20950 -14836
rect 20950 -14866 20981 -14836
rect 21021 -14866 21053 -14836
rect 21053 -14866 21055 -14836
rect 21095 -14866 21122 -14836
rect 21122 -14866 21129 -14836
rect 21169 -14866 21191 -14836
rect 21191 -14866 21203 -14836
rect 21243 -14866 21260 -14836
rect 21260 -14866 21277 -14836
rect 21317 -14866 21329 -14836
rect 21329 -14866 21351 -14836
rect 21391 -14866 21398 -14836
rect 21398 -14866 21425 -14836
rect 21465 -14866 21467 -14836
rect 21467 -14866 21499 -14836
rect 21539 -14866 21571 -14836
rect 21571 -14866 21573 -14836
rect 21613 -14866 21647 -14836
rect 21686 -14866 21720 -14836
rect 21759 -14866 21793 -14836
rect 21832 -14866 21866 -14836
rect 21905 -14866 21939 -14836
rect 21978 -14866 22012 -14836
rect 20651 -14870 20685 -14866
rect 20725 -14870 20759 -14866
rect 20799 -14870 20833 -14866
rect 20873 -14870 20907 -14866
rect 20947 -14870 20981 -14866
rect 21021 -14870 21055 -14866
rect 21095 -14870 21129 -14866
rect 21169 -14870 21203 -14866
rect 21243 -14870 21277 -14866
rect 21317 -14870 21351 -14866
rect 21391 -14870 21425 -14866
rect 21465 -14870 21499 -14866
rect 21539 -14870 21573 -14866
rect 21613 -14870 21647 -14866
rect 21686 -14870 21720 -14866
rect 21759 -14870 21793 -14866
rect 21832 -14870 21866 -14866
rect 21905 -14870 21939 -14866
rect 21978 -14870 22012 -14866
<< metal1 >>
rect 3655 2027 3661 2079
rect 3713 2027 3742 2079
rect 3794 2027 3823 2079
rect 3875 2027 3905 2079
rect 3957 2027 3963 2079
rect 3655 2001 3963 2027
rect 3655 1949 3661 2001
rect 3713 1949 3742 2001
rect 3794 1949 3823 2001
rect 3875 1949 3905 2001
rect 3957 1949 3963 2001
rect 88 380 94 432
rect 146 380 158 432
rect 210 380 222 432
rect 274 420 286 432
rect 338 420 350 432
rect 402 420 414 432
rect 466 420 478 432
rect 530 420 542 432
rect 594 420 606 432
rect 278 386 286 420
rect 530 386 532 420
rect 594 386 604 420
rect 274 380 286 386
rect 338 380 350 386
rect 402 380 414 386
rect 466 380 478 386
rect 530 380 542 386
rect 594 380 606 386
rect 658 380 670 432
rect 722 380 734 432
rect 786 380 798 432
rect 850 420 862 432
rect 914 420 926 432
rect 978 420 990 432
rect 1042 420 1054 432
rect 854 386 862 420
rect 850 380 862 386
rect 914 380 926 386
rect 978 380 990 386
rect 1042 380 1054 386
rect 1106 380 1118 432
rect 1170 380 1182 432
rect 1234 380 1246 432
rect 1298 420 1310 432
rect 1362 420 1374 432
rect 1426 420 1438 432
rect 1490 420 1502 432
rect 1554 420 1566 432
rect 1618 420 1630 432
rect 1300 386 1310 420
rect 1372 386 1374 420
rect 1618 386 1626 420
rect 1298 380 1310 386
rect 1362 380 1374 386
rect 1426 380 1438 386
rect 1490 380 1502 386
rect 1554 380 1566 386
rect 1618 380 1630 386
rect 1682 380 1694 432
rect 1746 380 1758 432
rect 1810 380 1822 432
rect 1874 420 1886 432
rect 1938 420 1950 432
rect 2002 420 2014 432
rect 2066 420 2078 432
rect 2130 420 2142 432
rect 1876 386 1886 420
rect 1948 386 1950 420
rect 1874 380 1886 386
rect 1938 380 1950 386
rect 2002 380 2014 386
rect 2066 380 2078 386
rect 2130 380 2142 386
rect 2194 380 2206 432
rect 2258 380 2270 432
rect 2322 380 2334 432
rect 2386 420 2398 432
rect 2450 420 2462 432
rect 2514 420 2526 432
rect 2578 420 2590 432
rect 2642 420 2654 432
rect 2578 386 2580 420
rect 2642 386 2652 420
rect 2386 380 2398 386
rect 2450 380 2462 386
rect 2514 380 2526 386
rect 2578 380 2590 386
rect 2642 380 2654 386
rect 2706 380 2718 432
rect 2770 380 2782 432
rect 2834 380 2846 432
rect 2898 420 2910 432
rect 2962 420 2974 432
rect 3026 420 3039 432
rect 3091 420 3104 432
rect 3156 420 3169 432
rect 3221 420 3234 432
rect 2902 386 2910 420
rect 3221 386 3228 420
rect 2898 380 2910 386
rect 2962 380 2974 386
rect 3026 380 3039 386
rect 3091 380 3104 386
rect 3156 380 3169 386
rect 3221 380 3234 386
rect 3286 380 3299 432
rect 3351 380 3364 432
rect 3416 380 3429 432
rect 3481 420 3494 432
rect 3546 420 3559 432
rect 3611 420 3624 432
rect 3676 420 3689 432
rect 3741 420 3754 432
rect 3806 420 3819 432
rect 3492 386 3494 420
rect 3741 386 3746 420
rect 3806 386 3818 420
rect 3481 380 3494 386
rect 3546 380 3559 386
rect 3611 380 3624 386
rect 3676 380 3689 386
rect 3741 380 3754 386
rect 3806 380 3819 386
rect 3871 380 3884 432
rect 3936 380 3949 432
rect 4001 380 4014 432
rect 4066 420 4079 432
rect 4131 420 4144 432
rect 4196 420 4209 432
rect 4261 420 4274 432
rect 4326 420 4339 432
rect 4391 420 4404 432
rect 4068 386 4079 420
rect 4140 386 4144 420
rect 4391 386 4394 420
rect 4066 380 4079 386
rect 4131 380 4144 386
rect 4196 380 4209 386
rect 4261 380 4274 386
rect 4326 380 4339 386
rect 4391 380 4404 386
rect 4456 380 4469 432
rect 4521 380 4534 432
rect 4586 380 4599 432
rect 4651 420 4664 432
rect 4716 420 4729 432
rect 4781 420 4794 432
rect 4846 420 4859 432
rect 4911 420 4924 432
rect 4976 420 4989 432
rect 4662 386 4664 420
rect 4911 386 4916 420
rect 4976 386 4988 420
rect 4651 380 4664 386
rect 4716 380 4729 386
rect 4781 380 4794 386
rect 4846 380 4859 386
rect 4911 380 4924 386
rect 4976 380 4989 386
rect 5041 380 5054 432
rect 5106 380 5119 432
rect 5171 380 5184 432
rect 5236 420 5249 432
rect 5301 420 5314 432
rect 5366 420 5379 432
rect 5431 420 5444 432
rect 5496 420 5509 432
rect 5561 420 5574 432
rect 5238 386 5249 420
rect 5310 386 5314 420
rect 5561 386 5564 420
rect 5236 380 5249 386
rect 5301 380 5314 386
rect 5366 380 5379 386
rect 5431 380 5444 386
rect 5496 380 5509 386
rect 5561 380 5574 386
rect 5626 380 5639 432
rect 5691 380 5704 432
rect 5756 380 5769 432
rect 5821 420 5834 432
rect 5886 420 5899 432
rect 5951 420 5964 432
rect 6016 420 6029 432
rect 6081 420 6094 432
rect 6146 420 6159 432
rect 5828 386 5834 420
rect 6081 386 6082 420
rect 6146 386 6154 420
rect 5821 380 5834 386
rect 5886 380 5899 386
rect 5951 380 5964 386
rect 6016 380 6029 386
rect 6081 380 6094 386
rect 6146 380 6159 386
rect 6211 380 6224 432
rect 6276 380 6289 432
rect 6341 380 6354 432
rect 6406 380 6419 432
rect 6471 420 6484 432
rect 6536 420 6549 432
rect 6601 420 6614 432
rect 6666 420 6679 432
rect 6476 386 6484 420
rect 6548 386 6549 420
rect 6471 380 6484 386
rect 6536 380 6549 386
rect 6601 380 6614 386
rect 6666 380 6679 386
rect 6731 380 6737 432
rect 330 297 6737 312
rect 330 296 4051 297
rect 330 270 2210 296
rect 88 264 2210 270
rect 88 230 100 264
rect 134 230 172 264
rect 206 230 244 264
rect 278 230 316 264
rect 350 230 388 264
rect 422 230 460 264
rect 494 230 532 264
rect 566 230 604 264
rect 638 230 676 264
rect 710 230 748 264
rect 782 230 820 264
rect 854 230 892 264
rect 926 230 964 264
rect 998 230 1036 264
rect 1070 230 1194 264
rect 1228 230 1266 264
rect 1300 230 1338 264
rect 1372 230 1410 264
rect 1444 230 1482 264
rect 1516 230 1554 264
rect 1588 230 1626 264
rect 1660 230 1698 264
rect 1732 230 1770 264
rect 1804 230 1842 264
rect 1876 230 1914 264
rect 1948 230 1986 264
rect 2020 230 2058 264
rect 2092 230 2130 264
rect 2164 244 2210 264
rect 2262 244 2279 296
rect 2331 244 2348 296
rect 2400 244 2417 296
rect 2469 264 2486 296
rect 2538 264 2555 296
rect 2607 264 2624 296
rect 2676 264 2693 296
rect 2745 264 2762 296
rect 2814 264 2831 296
rect 2883 264 2899 296
rect 2951 264 2967 296
rect 3019 264 3035 296
rect 3087 264 4051 296
rect 4103 264 4120 297
rect 4172 264 4189 297
rect 4241 264 4258 297
rect 4310 264 4327 297
rect 4379 264 4396 297
rect 2470 244 2486 264
rect 2542 244 2555 264
rect 2614 244 2624 264
rect 2686 244 2693 264
rect 2758 244 2762 264
rect 2830 244 2831 264
rect 2164 230 2364 244
rect 2398 230 2436 244
rect 2470 230 2508 244
rect 2542 230 2580 244
rect 2614 230 2652 244
rect 2686 230 2724 244
rect 2758 230 2796 244
rect 2830 230 2868 244
rect 2902 230 2940 244
rect 2974 230 3012 244
rect 3046 230 3084 244
rect 3118 230 3156 264
rect 3190 230 3228 264
rect 3262 230 3300 264
rect 3334 230 3458 264
rect 3492 230 3530 264
rect 3564 230 3602 264
rect 3636 230 3674 264
rect 3708 230 3746 264
rect 3780 230 3818 264
rect 3852 230 3890 264
rect 3924 230 3962 264
rect 3996 230 4034 264
rect 4103 245 4106 264
rect 4172 245 4178 264
rect 4241 245 4250 264
rect 4310 245 4322 264
rect 4379 245 4394 264
rect 4448 245 4465 297
rect 4517 245 4534 297
rect 4586 245 4603 297
rect 4655 264 4672 297
rect 4724 264 4740 297
rect 4792 264 4808 297
rect 4860 264 4876 297
rect 4928 264 6737 297
rect 4662 245 4672 264
rect 4734 245 4740 264
rect 4806 245 4808 264
rect 4068 230 4106 245
rect 4140 230 4178 245
rect 4212 230 4250 245
rect 4284 230 4322 245
rect 4356 230 4394 245
rect 4428 230 4628 245
rect 4662 230 4700 245
rect 4734 230 4772 245
rect 4806 230 4844 245
rect 4878 230 4916 245
rect 4950 230 4988 264
rect 5022 230 5060 264
rect 5094 230 5132 264
rect 5166 230 5204 264
rect 5238 230 5276 264
rect 5310 230 5348 264
rect 5382 230 5420 264
rect 5454 230 5492 264
rect 5526 230 5564 264
rect 5598 230 5722 264
rect 5756 230 5794 264
rect 5828 230 5866 264
rect 5900 230 5938 264
rect 5972 230 6010 264
rect 6044 230 6082 264
rect 6116 230 6154 264
rect 6188 230 6226 264
rect 6260 230 6298 264
rect 6332 230 6370 264
rect 6404 230 6442 264
rect 6476 230 6514 264
rect 6548 230 6586 264
rect 6620 230 6658 264
rect 6692 230 6737 264
rect 88 224 6737 230
rect -65 140 -59 192
rect -7 140 5 192
rect 57 186 6857 192
rect 57 152 1079 186
rect 1113 152 1151 186
rect 1185 152 2211 186
rect 2245 152 2283 186
rect 2317 152 3343 186
rect 3377 152 3415 186
rect 3449 152 4475 186
rect 4509 152 4547 186
rect 4581 152 5607 186
rect 5641 152 5679 186
rect 5713 152 6739 186
rect 6773 152 6811 186
rect 6845 152 6857 186
rect 57 146 6857 152
rect 57 140 63 146
rect 88 62 94 114
rect 146 62 158 114
rect 210 62 222 114
rect 274 108 286 114
rect 338 108 350 114
rect 402 108 414 114
rect 466 108 478 114
rect 530 108 542 114
rect 594 108 606 114
rect 278 74 286 108
rect 530 74 532 108
rect 594 74 604 108
rect 274 62 286 74
rect 338 62 350 74
rect 402 62 414 74
rect 466 62 478 74
rect 530 62 542 74
rect 594 62 606 74
rect 658 62 670 114
rect 722 62 734 114
rect 786 62 798 114
rect 850 108 862 114
rect 914 108 926 114
rect 978 108 990 114
rect 1042 108 1054 114
rect 854 74 862 108
rect 850 62 862 74
rect 914 62 926 74
rect 978 62 990 74
rect 1042 62 1054 74
rect 1106 62 1118 114
rect 1170 62 1182 114
rect 1234 62 1246 114
rect 1298 108 1310 114
rect 1362 108 1374 114
rect 1426 108 1438 114
rect 1490 108 1502 114
rect 1554 108 1566 114
rect 1618 108 1630 114
rect 1300 74 1310 108
rect 1372 74 1374 108
rect 1618 74 1626 108
rect 1298 62 1310 74
rect 1362 62 1374 74
rect 1426 62 1438 74
rect 1490 62 1502 74
rect 1554 62 1566 74
rect 1618 62 1630 74
rect 1682 62 1694 114
rect 1746 62 1758 114
rect 1810 62 1822 114
rect 1874 108 1886 114
rect 1938 108 1950 114
rect 2002 108 2014 114
rect 2066 108 2078 114
rect 2130 108 2142 114
rect 1876 74 1886 108
rect 1948 74 1950 108
rect 1874 62 1886 74
rect 1938 62 1950 74
rect 2002 62 2014 74
rect 2066 62 2078 74
rect 2130 62 2142 74
rect 2194 62 2206 114
rect 2258 62 2270 114
rect 2322 62 2334 114
rect 2386 108 2398 114
rect 2450 108 2462 114
rect 2514 108 2526 114
rect 2578 108 2590 114
rect 2642 108 2654 114
rect 2578 74 2580 108
rect 2642 74 2652 108
rect 2386 62 2398 74
rect 2450 62 2462 74
rect 2514 62 2526 74
rect 2578 62 2590 74
rect 2642 62 2654 74
rect 2706 62 2718 114
rect 2770 62 2782 114
rect 2834 62 2846 114
rect 2898 108 2910 114
rect 2962 108 2974 114
rect 3026 108 3039 114
rect 3091 108 3104 114
rect 3156 108 3169 114
rect 3221 108 3234 114
rect 2902 74 2910 108
rect 3221 74 3228 108
rect 2898 62 2910 74
rect 2962 62 2974 74
rect 3026 62 3039 74
rect 3091 62 3104 74
rect 3156 62 3169 74
rect 3221 62 3234 74
rect 3286 62 3299 114
rect 3351 62 3364 114
rect 3416 62 3429 114
rect 3481 108 3494 114
rect 3546 108 3559 114
rect 3611 108 3624 114
rect 3676 108 3689 114
rect 3741 108 3754 114
rect 3806 108 3819 114
rect 3492 74 3494 108
rect 3741 74 3746 108
rect 3806 74 3818 108
rect 3481 62 3494 74
rect 3546 62 3559 74
rect 3611 62 3624 74
rect 3676 62 3689 74
rect 3741 62 3754 74
rect 3806 62 3819 74
rect 3871 62 3884 114
rect 3936 62 3949 114
rect 4001 62 4014 114
rect 4066 108 4079 114
rect 4131 108 4144 114
rect 4196 108 4209 114
rect 4261 108 4274 114
rect 4326 108 4339 114
rect 4391 108 4404 114
rect 4068 74 4079 108
rect 4140 74 4144 108
rect 4391 74 4394 108
rect 4066 62 4079 74
rect 4131 62 4144 74
rect 4196 62 4209 74
rect 4261 62 4274 74
rect 4326 62 4339 74
rect 4391 62 4404 74
rect 4456 62 4469 114
rect 4521 62 4534 114
rect 4586 62 4599 114
rect 4651 108 4664 114
rect 4716 108 4729 114
rect 4781 108 4794 114
rect 4846 108 4859 114
rect 4911 108 4924 114
rect 4976 108 4989 114
rect 4662 74 4664 108
rect 4911 74 4916 108
rect 4976 74 4988 108
rect 4651 62 4664 74
rect 4716 62 4729 74
rect 4781 62 4794 74
rect 4846 62 4859 74
rect 4911 62 4924 74
rect 4976 62 4989 74
rect 5041 62 5054 114
rect 5106 62 5119 114
rect 5171 62 5184 114
rect 5236 108 5249 114
rect 5301 108 5314 114
rect 5366 108 5379 114
rect 5431 108 5444 114
rect 5496 108 5509 114
rect 5561 108 5574 114
rect 5238 74 5249 108
rect 5310 74 5314 108
rect 5561 74 5564 108
rect 5236 62 5249 74
rect 5301 62 5314 74
rect 5366 62 5379 74
rect 5431 62 5444 74
rect 5496 62 5509 74
rect 5561 62 5574 74
rect 5626 62 5639 114
rect 5691 62 5704 114
rect 5756 62 5769 114
rect 5821 108 5834 114
rect 5886 108 5899 114
rect 5951 108 5964 114
rect 6016 108 6029 114
rect 6081 108 6094 114
rect 6146 108 6159 114
rect 5828 74 5834 108
rect 6081 74 6082 108
rect 6146 74 6154 108
rect 5821 62 5834 74
rect 5886 62 5899 74
rect 5951 62 5964 74
rect 6016 62 6029 74
rect 6081 62 6094 74
rect 6146 62 6159 74
rect 6211 62 6224 114
rect 6276 62 6289 114
rect 6341 62 6354 114
rect 6406 62 6419 114
rect 6471 108 6484 114
rect 6536 108 6549 114
rect 6601 108 6614 114
rect 6666 108 6679 114
rect 6476 74 6484 108
rect 6548 74 6549 108
rect 6471 62 6484 74
rect 6536 62 6549 74
rect 6601 62 6614 74
rect 6666 62 6679 74
rect 6731 62 6737 114
rect -182 -88 -130 -82
rect -182 -152 -130 -140
rect -182 -3457 -130 -204
rect 20974 -3425 21020 -3413
rect -182 -3482 445 -3457
rect 20974 -3459 20980 -3425
rect 21014 -3459 21020 -3425
rect -182 -3489 20509 -3482
rect 413 -3497 20509 -3489
tri 20509 -3497 20524 -3482 sw
rect 20974 -3497 21020 -3459
rect 413 -3511 20524 -3497
tri 20524 -3511 20538 -3497 sw
rect 20974 -3511 20980 -3497
rect 413 -3514 20980 -3511
tri 20486 -3531 20503 -3514 ne
rect 20503 -3531 20980 -3514
rect 21014 -3511 21020 -3497
rect 21657 -3421 21709 -3415
rect 21657 -3485 21709 -3473
rect 21014 -3531 21657 -3511
tri 20503 -3543 20515 -3531 ne
rect 20515 -3537 21657 -3531
rect 20515 -3543 21709 -3537
rect 20818 -3679 21240 -3673
rect 20818 -3685 21188 -3679
rect 20818 -3719 20824 -3685
rect 20858 -3719 21136 -3685
rect 21170 -3719 21188 -3685
rect 20818 -3731 21188 -3719
rect 20818 -3782 21240 -3731
rect 20818 -3794 21188 -3782
rect 20818 -3828 20824 -3794
rect 20858 -3828 21136 -3794
rect 21170 -3828 21188 -3794
rect 20818 -3834 21188 -3828
rect 20818 -3840 21240 -3834
rect -2935 -4716 -2763 -4547
rect -3365 -5079 -3205 -4949
rect 21111 -5194 21117 -5142
rect 21169 -5194 21181 -5142
rect 21233 -5194 21239 -5142
rect 20619 -7893 22091 -7887
rect 20619 -7927 20651 -7893
rect 20685 -7927 20724 -7893
rect 20758 -7927 20797 -7893
rect 20831 -7927 20870 -7893
rect 20904 -7927 20943 -7893
rect 20977 -7927 21017 -7893
rect 21051 -7927 21091 -7893
rect 21125 -7927 21165 -7893
rect 21199 -7927 21239 -7893
rect 21273 -7927 21313 -7893
rect 21347 -7927 21387 -7893
rect 21421 -7927 21461 -7893
rect 21495 -7927 21535 -7893
rect 21569 -7927 21609 -7893
rect 21643 -7927 21683 -7893
rect 21717 -7927 21757 -7893
rect 21791 -7927 21831 -7893
rect 21865 -7927 21905 -7893
rect 21939 -7927 21979 -7893
rect 22013 -7927 22091 -7893
rect 20619 -7965 22091 -7927
rect 20619 -7999 20651 -7965
rect 20685 -7999 20724 -7965
rect 20758 -7999 20797 -7965
rect 20831 -7999 20870 -7965
rect 20904 -7999 20943 -7965
rect 20977 -7999 21017 -7965
rect 21051 -7999 21091 -7965
rect 21125 -7999 21165 -7965
rect 21199 -7999 21239 -7965
rect 21273 -7999 21313 -7965
rect 21347 -7999 21387 -7965
rect 21421 -7999 21461 -7965
rect 21495 -7999 21535 -7965
rect 21569 -7999 21609 -7965
rect 21643 -7999 21683 -7965
rect 21717 -7999 21757 -7965
rect 21791 -7999 21831 -7965
rect 21865 -7999 21905 -7965
rect 21939 -7999 21979 -7965
rect 20619 -8037 21979 -7999
rect 20619 -8071 20651 -8037
rect 20685 -8071 20724 -8037
rect 20758 -8071 20797 -8037
rect 20831 -8071 20871 -8037
rect 20905 -8071 20945 -8037
rect 20979 -8071 21019 -8037
rect 21053 -8071 21093 -8037
rect 21127 -8071 21167 -8037
rect 21201 -8071 21241 -8037
rect 21275 -8071 21315 -8037
rect 21349 -8071 21389 -8037
rect 21423 -8071 21463 -8037
rect 21497 -8071 21537 -8037
rect 21571 -8071 21611 -8037
rect 21645 -8071 21685 -8037
rect 21719 -8071 21759 -8037
rect 21793 -8071 21833 -8037
rect 21867 -8071 21907 -8037
rect 20619 -8077 21907 -8071
rect 21217 -10006 21263 -9994
rect 21217 -10040 21223 -10006
rect 21257 -10040 21263 -10006
rect 21217 -10078 21263 -10040
rect 21217 -10112 21223 -10078
rect 21257 -10112 21263 -10078
rect 21217 -10150 21263 -10112
rect 21217 -10184 21223 -10150
rect 21257 -10184 21263 -10150
rect 21217 -10222 21263 -10184
rect 21370 -10006 21422 -9994
rect 21370 -10016 21379 -10006
rect 21413 -10016 21422 -10006
rect 21370 -10078 21422 -10068
rect 21370 -10080 21379 -10078
rect 21413 -10080 21422 -10078
rect 21370 -10144 21422 -10132
rect 21370 -10202 21422 -10196
tri 21370 -10205 21373 -10202 ne
rect 21217 -10256 21223 -10222
rect 21257 -10256 21263 -10222
rect 21217 -10294 21263 -10256
rect 21217 -10328 21223 -10294
rect 21257 -10328 21263 -10294
rect 21217 -10348 21263 -10328
rect 21373 -10222 21419 -10202
tri 21419 -10205 21422 -10202 nw
rect 21529 -10006 21575 -9994
rect 21529 -10040 21535 -10006
rect 21569 -10040 21575 -10006
rect 21529 -10078 21575 -10040
rect 21529 -10112 21535 -10078
rect 21569 -10112 21575 -10078
rect 21529 -10150 21575 -10112
rect 21529 -10184 21535 -10150
rect 21569 -10184 21575 -10150
rect 21373 -10256 21379 -10222
rect 21413 -10256 21419 -10222
rect 21373 -10294 21419 -10256
rect 21373 -10328 21379 -10294
rect 21413 -10328 21419 -10294
rect 21214 -10354 21266 -10348
rect 21214 -10418 21266 -10406
rect 21214 -10472 21223 -10470
rect 21257 -10472 21266 -10470
rect 21214 -10482 21266 -10472
rect 21214 -10540 21223 -10534
rect 21217 -10544 21223 -10540
rect 21257 -10540 21266 -10534
rect 21373 -10366 21419 -10328
rect 21529 -10222 21575 -10184
rect 21529 -10256 21535 -10222
rect 21569 -10256 21575 -10222
rect 21529 -10294 21575 -10256
rect 21529 -10328 21535 -10294
rect 21569 -10328 21575 -10294
rect 21529 -10348 21575 -10328
rect 21373 -10400 21379 -10366
rect 21413 -10400 21419 -10366
rect 21373 -10438 21419 -10400
rect 21373 -10472 21379 -10438
rect 21413 -10472 21419 -10438
rect 21373 -10510 21419 -10472
rect 21257 -10544 21263 -10540
rect 21217 -10556 21263 -10544
rect 21295 -10553 21341 -10541
rect 21295 -10587 21301 -10553
rect 21335 -10587 21341 -10553
rect 21373 -10544 21379 -10510
rect 21413 -10544 21419 -10510
rect 21526 -10354 21578 -10348
rect 21526 -10418 21578 -10406
rect 21526 -10472 21535 -10470
rect 21569 -10472 21578 -10470
rect 21526 -10482 21578 -10472
rect 21526 -10540 21535 -10534
rect 21373 -10556 21419 -10544
rect 21529 -10544 21535 -10540
rect 21569 -10540 21578 -10534
rect 21569 -10544 21575 -10540
rect 21529 -10556 21575 -10544
rect 21295 -10625 21341 -10587
rect 21295 -10659 21301 -10625
rect 21335 -10659 21341 -10625
rect 21295 -10671 21341 -10659
rect 21901 -12463 21907 -8077
rect 21901 -12502 21979 -12463
rect 21901 -12536 21907 -12502
rect 21941 -12535 21979 -12502
rect 22085 -12535 22091 -7965
rect 21941 -12536 22091 -12535
rect 21901 -12574 22091 -12536
rect 21901 -12575 21979 -12574
rect 21901 -12609 21907 -12575
rect 21941 -12608 21979 -12575
rect 22013 -12608 22051 -12574
rect 22085 -12608 22091 -12574
rect 21941 -12609 22091 -12608
rect 21901 -12647 22091 -12609
rect 21901 -12648 21979 -12647
rect 21901 -12682 21907 -12648
rect 21941 -12681 21979 -12648
rect 22013 -12681 22051 -12647
rect 22085 -12681 22091 -12647
rect 21941 -12682 22091 -12681
rect 21901 -12720 22091 -12682
rect 21901 -12721 21979 -12720
rect 21901 -12755 21907 -12721
rect 21941 -12754 21979 -12721
rect 22013 -12754 22051 -12720
rect 22085 -12754 22091 -12720
rect 21941 -12755 22091 -12754
rect 21901 -12793 22091 -12755
rect 21901 -12794 21979 -12793
rect 21901 -12828 21907 -12794
rect 21941 -12827 21979 -12794
rect 22013 -12827 22051 -12793
rect 22085 -12827 22091 -12793
rect 21941 -12828 22091 -12827
rect 21901 -12866 22091 -12828
rect 21901 -12867 21979 -12866
rect 21901 -12901 21907 -12867
rect 21941 -12900 21979 -12867
rect 22013 -12900 22051 -12866
rect 22085 -12900 22091 -12866
rect 21941 -12901 22091 -12900
rect 21901 -12939 22091 -12901
rect 21901 -12940 21979 -12939
rect 21901 -12974 21907 -12940
rect 21941 -12973 21979 -12940
rect 22013 -12973 22051 -12939
rect 22085 -12973 22091 -12939
rect 21941 -12974 22091 -12973
rect 21901 -13012 22091 -12974
rect 21901 -13013 21979 -13012
rect 21901 -13047 21907 -13013
rect 21941 -13046 21979 -13013
rect 22013 -13046 22051 -13012
rect 22085 -13046 22091 -13012
rect 21941 -13047 22091 -13046
rect 21901 -13085 22091 -13047
rect 21901 -13086 21979 -13085
rect 21901 -13120 21907 -13086
rect 21941 -13119 21979 -13086
rect 22013 -13119 22051 -13085
rect 22085 -13119 22091 -13085
rect 21941 -13120 22091 -13119
rect 21901 -13158 22091 -13120
rect 21901 -13159 21979 -13158
rect 21901 -13193 21907 -13159
rect 21941 -13192 21979 -13159
rect 22013 -13192 22051 -13158
rect 22085 -13192 22091 -13158
rect 21941 -13193 22091 -13192
rect 21901 -13231 22091 -13193
rect 21901 -13232 21979 -13231
rect 21901 -13266 21907 -13232
rect 21941 -13265 21979 -13232
rect 22013 -13265 22051 -13231
rect 22085 -13265 22091 -13231
rect 21941 -13266 22091 -13265
rect 21901 -13304 22091 -13266
rect 21901 -13305 21979 -13304
rect 21901 -13339 21907 -13305
rect 21941 -13338 21979 -13305
rect 22013 -13338 22051 -13304
rect 22085 -13338 22091 -13304
rect 21941 -13339 22091 -13338
rect 21901 -13377 22091 -13339
rect 21901 -13378 21979 -13377
rect 21901 -13412 21907 -13378
rect 21941 -13411 21979 -13378
rect 22013 -13411 22051 -13377
rect 22085 -13411 22091 -13377
rect 21941 -13412 22091 -13411
rect 21901 -13450 22091 -13412
rect 21901 -13451 21979 -13450
rect 21901 -13485 21907 -13451
rect 21941 -13484 21979 -13451
rect 22013 -13484 22051 -13450
rect 22085 -13484 22091 -13450
rect 21941 -13485 22091 -13484
rect 21901 -13523 22091 -13485
rect 21901 -13524 21979 -13523
rect 21901 -13558 21907 -13524
rect 21941 -13557 21979 -13524
rect 22013 -13557 22051 -13523
rect 22085 -13557 22091 -13523
rect 21941 -13558 22091 -13557
rect 21901 -13596 22091 -13558
rect 21901 -13597 21979 -13596
rect 21901 -13631 21907 -13597
rect 21941 -13630 21979 -13597
rect 22013 -13630 22051 -13596
rect 22085 -13630 22091 -13596
rect 21941 -13631 22091 -13630
rect 21901 -13669 22091 -13631
rect 21901 -13670 21979 -13669
rect 21901 -13704 21907 -13670
rect 21941 -13703 21979 -13670
rect 22013 -13703 22051 -13669
rect 22085 -13703 22091 -13669
rect 21941 -13704 22091 -13703
rect 21901 -13742 22091 -13704
rect 21901 -13743 21979 -13742
rect 21901 -13777 21907 -13743
rect 21941 -13776 21979 -13743
rect 22013 -13776 22051 -13742
rect 22085 -13776 22091 -13742
rect 21941 -13777 22091 -13776
rect 21901 -13815 22091 -13777
rect 21901 -13816 21979 -13815
rect 21901 -13850 21907 -13816
rect 21941 -13849 21979 -13816
rect 22013 -13849 22051 -13815
rect 22085 -13849 22091 -13815
rect 21941 -13850 22091 -13849
rect 21901 -13888 22091 -13850
rect 21901 -13889 21979 -13888
rect 21901 -13923 21907 -13889
rect 21941 -13922 21979 -13889
rect 22013 -13922 22051 -13888
rect 22085 -13922 22091 -13888
rect 21941 -13923 22091 -13922
rect 21901 -13961 22091 -13923
rect 21901 -13962 21979 -13961
rect 21901 -13996 21907 -13962
rect 21941 -13995 21979 -13962
rect 22013 -13995 22051 -13961
rect 22085 -13995 22091 -13961
rect 21941 -13996 22091 -13995
rect 21901 -14034 22091 -13996
rect 21901 -14035 21979 -14034
rect 21901 -14069 21907 -14035
rect 21941 -14068 21979 -14035
rect 22013 -14068 22051 -14034
rect 22085 -14068 22091 -14034
rect 21941 -14069 22091 -14068
rect 21901 -14107 22091 -14069
rect 21901 -14108 21979 -14107
rect 21901 -14142 21907 -14108
rect 21941 -14141 21979 -14108
rect 22013 -14141 22051 -14107
rect 22085 -14141 22091 -14107
rect 21941 -14142 22091 -14141
rect 21901 -14180 22091 -14142
rect 21901 -14181 21979 -14180
rect 21901 -14215 21907 -14181
rect 21941 -14214 21979 -14181
rect 22013 -14214 22051 -14180
rect 22085 -14214 22091 -14180
rect 21941 -14215 22091 -14214
rect 21901 -14253 22091 -14215
rect 21901 -14254 21979 -14253
rect 21901 -14288 21907 -14254
rect 21941 -14287 21979 -14254
rect 22013 -14287 22051 -14253
rect 22085 -14287 22091 -14253
rect 21941 -14288 22091 -14287
rect 21901 -14326 22091 -14288
rect 21901 -14327 21979 -14326
rect 21901 -14361 21907 -14327
rect 21941 -14360 21979 -14327
rect 22013 -14360 22051 -14326
rect 22085 -14360 22091 -14326
rect 21941 -14361 22091 -14360
rect 21901 -14399 22091 -14361
rect 21901 -14400 21979 -14399
rect 21901 -14434 21907 -14400
rect 21941 -14433 21979 -14400
rect 22013 -14433 22051 -14399
rect 22085 -14433 22091 -14399
rect 21941 -14434 22091 -14433
rect 21332 -14466 21582 -14436
rect 21332 -14518 21338 -14466
rect 21390 -14518 21431 -14466
rect 21483 -14518 21524 -14466
rect 21576 -14518 21582 -14466
rect 21332 -14548 21582 -14518
rect 21901 -14472 22091 -14434
rect 21901 -14473 21979 -14472
rect 21901 -14507 21907 -14473
rect 21941 -14506 21979 -14473
rect 22013 -14506 22051 -14472
rect 22085 -14506 22091 -14472
rect 21941 -14507 22091 -14506
rect 21901 -14545 22091 -14507
rect 21901 -14546 21979 -14545
rect 21901 -14580 21907 -14546
rect 21941 -14579 21979 -14546
rect 22013 -14579 22051 -14545
rect 22085 -14579 22091 -14545
rect 21941 -14580 22091 -14579
rect 21901 -14618 22091 -14580
rect 21901 -14619 21979 -14618
rect 21901 -14653 21907 -14619
rect 21941 -14652 21979 -14619
rect 22013 -14652 22051 -14618
rect 22085 -14652 22091 -14618
rect 21941 -14653 22091 -14652
rect 21901 -14686 22091 -14653
rect 20619 -14691 22091 -14686
rect 20619 -14692 21979 -14691
rect 20619 -14726 20651 -14692
rect 20685 -14726 20725 -14692
rect 20759 -14726 20799 -14692
rect 20833 -14726 20873 -14692
rect 20907 -14726 20947 -14692
rect 20981 -14726 21021 -14692
rect 21055 -14726 21095 -14692
rect 21129 -14726 21169 -14692
rect 21203 -14726 21243 -14692
rect 21277 -14726 21317 -14692
rect 21351 -14726 21391 -14692
rect 21425 -14726 21465 -14692
rect 21499 -14726 21539 -14692
rect 21573 -14726 21613 -14692
rect 21647 -14726 21687 -14692
rect 21721 -14726 21761 -14692
rect 21795 -14726 21834 -14692
rect 21868 -14726 21907 -14692
rect 21941 -14725 21979 -14692
rect 22013 -14725 22051 -14691
rect 22085 -14725 22091 -14691
rect 21941 -14726 22091 -14725
rect 20619 -14764 22091 -14726
rect 20619 -14798 20651 -14764
rect 20685 -14798 20725 -14764
rect 20759 -14798 20799 -14764
rect 20833 -14798 20873 -14764
rect 20907 -14798 20947 -14764
rect 20981 -14798 21021 -14764
rect 21055 -14798 21095 -14764
rect 21129 -14798 21169 -14764
rect 21203 -14798 21243 -14764
rect 21277 -14798 21317 -14764
rect 21351 -14798 21391 -14764
rect 21425 -14798 21465 -14764
rect 21499 -14798 21539 -14764
rect 21573 -14798 21613 -14764
rect 21647 -14798 21686 -14764
rect 21720 -14798 21759 -14764
rect 21793 -14798 21832 -14764
rect 21866 -14798 21905 -14764
rect 21939 -14798 21979 -14764
rect 22013 -14798 22051 -14764
rect 22085 -14798 22091 -14764
rect 20619 -14836 22091 -14798
rect 20619 -14870 20651 -14836
rect 20685 -14870 20725 -14836
rect 20759 -14870 20799 -14836
rect 20833 -14870 20873 -14836
rect 20907 -14870 20947 -14836
rect 20981 -14870 21021 -14836
rect 21055 -14870 21095 -14836
rect 21129 -14870 21169 -14836
rect 21203 -14870 21243 -14836
rect 21277 -14870 21317 -14836
rect 21351 -14870 21391 -14836
rect 21425 -14870 21465 -14836
rect 21499 -14870 21539 -14836
rect 21573 -14870 21613 -14836
rect 21647 -14870 21686 -14836
rect 21720 -14870 21759 -14836
rect 21793 -14870 21832 -14836
rect 21866 -14870 21905 -14836
rect 21939 -14870 21978 -14836
rect 22012 -14870 22091 -14836
rect 20619 -14876 22091 -14870
<< via1 >>
rect 3661 2027 3713 2079
rect 3742 2027 3794 2079
rect 3823 2027 3875 2079
rect 3905 2027 3957 2079
rect 3661 1949 3713 2001
rect 3742 1949 3794 2001
rect 3823 1949 3875 2001
rect 3905 1949 3957 2001
rect 94 420 146 432
rect 94 386 100 420
rect 100 386 134 420
rect 134 386 146 420
rect 94 380 146 386
rect 158 420 210 432
rect 158 386 172 420
rect 172 386 206 420
rect 206 386 210 420
rect 158 380 210 386
rect 222 420 274 432
rect 286 420 338 432
rect 350 420 402 432
rect 414 420 466 432
rect 478 420 530 432
rect 542 420 594 432
rect 606 420 658 432
rect 222 386 244 420
rect 244 386 274 420
rect 286 386 316 420
rect 316 386 338 420
rect 350 386 388 420
rect 388 386 402 420
rect 414 386 422 420
rect 422 386 460 420
rect 460 386 466 420
rect 478 386 494 420
rect 494 386 530 420
rect 542 386 566 420
rect 566 386 594 420
rect 606 386 638 420
rect 638 386 658 420
rect 222 380 274 386
rect 286 380 338 386
rect 350 380 402 386
rect 414 380 466 386
rect 478 380 530 386
rect 542 380 594 386
rect 606 380 658 386
rect 670 420 722 432
rect 670 386 676 420
rect 676 386 710 420
rect 710 386 722 420
rect 670 380 722 386
rect 734 420 786 432
rect 734 386 748 420
rect 748 386 782 420
rect 782 386 786 420
rect 734 380 786 386
rect 798 420 850 432
rect 862 420 914 432
rect 926 420 978 432
rect 990 420 1042 432
rect 1054 420 1106 432
rect 798 386 820 420
rect 820 386 850 420
rect 862 386 892 420
rect 892 386 914 420
rect 926 386 964 420
rect 964 386 978 420
rect 990 386 998 420
rect 998 386 1036 420
rect 1036 386 1042 420
rect 1054 386 1070 420
rect 1070 386 1106 420
rect 798 380 850 386
rect 862 380 914 386
rect 926 380 978 386
rect 990 380 1042 386
rect 1054 380 1106 386
rect 1118 380 1170 432
rect 1182 420 1234 432
rect 1182 386 1194 420
rect 1194 386 1228 420
rect 1228 386 1234 420
rect 1182 380 1234 386
rect 1246 420 1298 432
rect 1310 420 1362 432
rect 1374 420 1426 432
rect 1438 420 1490 432
rect 1502 420 1554 432
rect 1566 420 1618 432
rect 1630 420 1682 432
rect 1246 386 1266 420
rect 1266 386 1298 420
rect 1310 386 1338 420
rect 1338 386 1362 420
rect 1374 386 1410 420
rect 1410 386 1426 420
rect 1438 386 1444 420
rect 1444 386 1482 420
rect 1482 386 1490 420
rect 1502 386 1516 420
rect 1516 386 1554 420
rect 1566 386 1588 420
rect 1588 386 1618 420
rect 1630 386 1660 420
rect 1660 386 1682 420
rect 1246 380 1298 386
rect 1310 380 1362 386
rect 1374 380 1426 386
rect 1438 380 1490 386
rect 1502 380 1554 386
rect 1566 380 1618 386
rect 1630 380 1682 386
rect 1694 420 1746 432
rect 1694 386 1698 420
rect 1698 386 1732 420
rect 1732 386 1746 420
rect 1694 380 1746 386
rect 1758 420 1810 432
rect 1758 386 1770 420
rect 1770 386 1804 420
rect 1804 386 1810 420
rect 1758 380 1810 386
rect 1822 420 1874 432
rect 1886 420 1938 432
rect 1950 420 2002 432
rect 2014 420 2066 432
rect 2078 420 2130 432
rect 2142 420 2194 432
rect 1822 386 1842 420
rect 1842 386 1874 420
rect 1886 386 1914 420
rect 1914 386 1938 420
rect 1950 386 1986 420
rect 1986 386 2002 420
rect 2014 386 2020 420
rect 2020 386 2058 420
rect 2058 386 2066 420
rect 2078 386 2092 420
rect 2092 386 2130 420
rect 2142 386 2164 420
rect 2164 386 2194 420
rect 1822 380 1874 386
rect 1886 380 1938 386
rect 1950 380 2002 386
rect 2014 380 2066 386
rect 2078 380 2130 386
rect 2142 380 2194 386
rect 2206 380 2258 432
rect 2270 380 2322 432
rect 2334 420 2386 432
rect 2398 420 2450 432
rect 2462 420 2514 432
rect 2526 420 2578 432
rect 2590 420 2642 432
rect 2654 420 2706 432
rect 2334 386 2364 420
rect 2364 386 2386 420
rect 2398 386 2436 420
rect 2436 386 2450 420
rect 2462 386 2470 420
rect 2470 386 2508 420
rect 2508 386 2514 420
rect 2526 386 2542 420
rect 2542 386 2578 420
rect 2590 386 2614 420
rect 2614 386 2642 420
rect 2654 386 2686 420
rect 2686 386 2706 420
rect 2334 380 2386 386
rect 2398 380 2450 386
rect 2462 380 2514 386
rect 2526 380 2578 386
rect 2590 380 2642 386
rect 2654 380 2706 386
rect 2718 420 2770 432
rect 2718 386 2724 420
rect 2724 386 2758 420
rect 2758 386 2770 420
rect 2718 380 2770 386
rect 2782 420 2834 432
rect 2782 386 2796 420
rect 2796 386 2830 420
rect 2830 386 2834 420
rect 2782 380 2834 386
rect 2846 420 2898 432
rect 2910 420 2962 432
rect 2974 420 3026 432
rect 3039 420 3091 432
rect 3104 420 3156 432
rect 3169 420 3221 432
rect 3234 420 3286 432
rect 2846 386 2868 420
rect 2868 386 2898 420
rect 2910 386 2940 420
rect 2940 386 2962 420
rect 2974 386 3012 420
rect 3012 386 3026 420
rect 3039 386 3046 420
rect 3046 386 3084 420
rect 3084 386 3091 420
rect 3104 386 3118 420
rect 3118 386 3156 420
rect 3169 386 3190 420
rect 3190 386 3221 420
rect 3234 386 3262 420
rect 3262 386 3286 420
rect 2846 380 2898 386
rect 2910 380 2962 386
rect 2974 380 3026 386
rect 3039 380 3091 386
rect 3104 380 3156 386
rect 3169 380 3221 386
rect 3234 380 3286 386
rect 3299 420 3351 432
rect 3299 386 3300 420
rect 3300 386 3334 420
rect 3334 386 3351 420
rect 3299 380 3351 386
rect 3364 380 3416 432
rect 3429 420 3481 432
rect 3494 420 3546 432
rect 3559 420 3611 432
rect 3624 420 3676 432
rect 3689 420 3741 432
rect 3754 420 3806 432
rect 3819 420 3871 432
rect 3429 386 3458 420
rect 3458 386 3481 420
rect 3494 386 3530 420
rect 3530 386 3546 420
rect 3559 386 3564 420
rect 3564 386 3602 420
rect 3602 386 3611 420
rect 3624 386 3636 420
rect 3636 386 3674 420
rect 3674 386 3676 420
rect 3689 386 3708 420
rect 3708 386 3741 420
rect 3754 386 3780 420
rect 3780 386 3806 420
rect 3819 386 3852 420
rect 3852 386 3871 420
rect 3429 380 3481 386
rect 3494 380 3546 386
rect 3559 380 3611 386
rect 3624 380 3676 386
rect 3689 380 3741 386
rect 3754 380 3806 386
rect 3819 380 3871 386
rect 3884 420 3936 432
rect 3884 386 3890 420
rect 3890 386 3924 420
rect 3924 386 3936 420
rect 3884 380 3936 386
rect 3949 420 4001 432
rect 3949 386 3962 420
rect 3962 386 3996 420
rect 3996 386 4001 420
rect 3949 380 4001 386
rect 4014 420 4066 432
rect 4079 420 4131 432
rect 4144 420 4196 432
rect 4209 420 4261 432
rect 4274 420 4326 432
rect 4339 420 4391 432
rect 4404 420 4456 432
rect 4014 386 4034 420
rect 4034 386 4066 420
rect 4079 386 4106 420
rect 4106 386 4131 420
rect 4144 386 4178 420
rect 4178 386 4196 420
rect 4209 386 4212 420
rect 4212 386 4250 420
rect 4250 386 4261 420
rect 4274 386 4284 420
rect 4284 386 4322 420
rect 4322 386 4326 420
rect 4339 386 4356 420
rect 4356 386 4391 420
rect 4404 386 4428 420
rect 4428 386 4456 420
rect 4014 380 4066 386
rect 4079 380 4131 386
rect 4144 380 4196 386
rect 4209 380 4261 386
rect 4274 380 4326 386
rect 4339 380 4391 386
rect 4404 380 4456 386
rect 4469 380 4521 432
rect 4534 380 4586 432
rect 4599 420 4651 432
rect 4664 420 4716 432
rect 4729 420 4781 432
rect 4794 420 4846 432
rect 4859 420 4911 432
rect 4924 420 4976 432
rect 4989 420 5041 432
rect 4599 386 4628 420
rect 4628 386 4651 420
rect 4664 386 4700 420
rect 4700 386 4716 420
rect 4729 386 4734 420
rect 4734 386 4772 420
rect 4772 386 4781 420
rect 4794 386 4806 420
rect 4806 386 4844 420
rect 4844 386 4846 420
rect 4859 386 4878 420
rect 4878 386 4911 420
rect 4924 386 4950 420
rect 4950 386 4976 420
rect 4989 386 5022 420
rect 5022 386 5041 420
rect 4599 380 4651 386
rect 4664 380 4716 386
rect 4729 380 4781 386
rect 4794 380 4846 386
rect 4859 380 4911 386
rect 4924 380 4976 386
rect 4989 380 5041 386
rect 5054 420 5106 432
rect 5054 386 5060 420
rect 5060 386 5094 420
rect 5094 386 5106 420
rect 5054 380 5106 386
rect 5119 420 5171 432
rect 5119 386 5132 420
rect 5132 386 5166 420
rect 5166 386 5171 420
rect 5119 380 5171 386
rect 5184 420 5236 432
rect 5249 420 5301 432
rect 5314 420 5366 432
rect 5379 420 5431 432
rect 5444 420 5496 432
rect 5509 420 5561 432
rect 5574 420 5626 432
rect 5184 386 5204 420
rect 5204 386 5236 420
rect 5249 386 5276 420
rect 5276 386 5301 420
rect 5314 386 5348 420
rect 5348 386 5366 420
rect 5379 386 5382 420
rect 5382 386 5420 420
rect 5420 386 5431 420
rect 5444 386 5454 420
rect 5454 386 5492 420
rect 5492 386 5496 420
rect 5509 386 5526 420
rect 5526 386 5561 420
rect 5574 386 5598 420
rect 5598 386 5626 420
rect 5184 380 5236 386
rect 5249 380 5301 386
rect 5314 380 5366 386
rect 5379 380 5431 386
rect 5444 380 5496 386
rect 5509 380 5561 386
rect 5574 380 5626 386
rect 5639 380 5691 432
rect 5704 420 5756 432
rect 5704 386 5722 420
rect 5722 386 5756 420
rect 5704 380 5756 386
rect 5769 420 5821 432
rect 5834 420 5886 432
rect 5899 420 5951 432
rect 5964 420 6016 432
rect 6029 420 6081 432
rect 6094 420 6146 432
rect 6159 420 6211 432
rect 5769 386 5794 420
rect 5794 386 5821 420
rect 5834 386 5866 420
rect 5866 386 5886 420
rect 5899 386 5900 420
rect 5900 386 5938 420
rect 5938 386 5951 420
rect 5964 386 5972 420
rect 5972 386 6010 420
rect 6010 386 6016 420
rect 6029 386 6044 420
rect 6044 386 6081 420
rect 6094 386 6116 420
rect 6116 386 6146 420
rect 6159 386 6188 420
rect 6188 386 6211 420
rect 5769 380 5821 386
rect 5834 380 5886 386
rect 5899 380 5951 386
rect 5964 380 6016 386
rect 6029 380 6081 386
rect 6094 380 6146 386
rect 6159 380 6211 386
rect 6224 420 6276 432
rect 6224 386 6226 420
rect 6226 386 6260 420
rect 6260 386 6276 420
rect 6224 380 6276 386
rect 6289 420 6341 432
rect 6289 386 6298 420
rect 6298 386 6332 420
rect 6332 386 6341 420
rect 6289 380 6341 386
rect 6354 420 6406 432
rect 6354 386 6370 420
rect 6370 386 6404 420
rect 6404 386 6406 420
rect 6354 380 6406 386
rect 6419 420 6471 432
rect 6484 420 6536 432
rect 6549 420 6601 432
rect 6614 420 6666 432
rect 6679 420 6731 432
rect 6419 386 6442 420
rect 6442 386 6471 420
rect 6484 386 6514 420
rect 6514 386 6536 420
rect 6549 386 6586 420
rect 6586 386 6601 420
rect 6614 386 6620 420
rect 6620 386 6658 420
rect 6658 386 6666 420
rect 6679 386 6692 420
rect 6692 386 6731 420
rect 6419 380 6471 386
rect 6484 380 6536 386
rect 6549 380 6601 386
rect 6614 380 6666 386
rect 6679 380 6731 386
rect 2210 244 2262 296
rect 2279 244 2331 296
rect 2348 264 2400 296
rect 2348 244 2364 264
rect 2364 244 2398 264
rect 2398 244 2400 264
rect 2417 264 2469 296
rect 2486 264 2538 296
rect 2555 264 2607 296
rect 2624 264 2676 296
rect 2693 264 2745 296
rect 2762 264 2814 296
rect 2831 264 2883 296
rect 2899 264 2951 296
rect 2967 264 3019 296
rect 3035 264 3087 296
rect 4051 264 4103 297
rect 4120 264 4172 297
rect 4189 264 4241 297
rect 4258 264 4310 297
rect 4327 264 4379 297
rect 4396 264 4448 297
rect 2417 244 2436 264
rect 2436 244 2469 264
rect 2486 244 2508 264
rect 2508 244 2538 264
rect 2555 244 2580 264
rect 2580 244 2607 264
rect 2624 244 2652 264
rect 2652 244 2676 264
rect 2693 244 2724 264
rect 2724 244 2745 264
rect 2762 244 2796 264
rect 2796 244 2814 264
rect 2831 244 2868 264
rect 2868 244 2883 264
rect 2899 244 2902 264
rect 2902 244 2940 264
rect 2940 244 2951 264
rect 2967 244 2974 264
rect 2974 244 3012 264
rect 3012 244 3019 264
rect 3035 244 3046 264
rect 3046 244 3084 264
rect 3084 244 3087 264
rect 4051 245 4068 264
rect 4068 245 4103 264
rect 4120 245 4140 264
rect 4140 245 4172 264
rect 4189 245 4212 264
rect 4212 245 4241 264
rect 4258 245 4284 264
rect 4284 245 4310 264
rect 4327 245 4356 264
rect 4356 245 4379 264
rect 4396 245 4428 264
rect 4428 245 4448 264
rect 4465 245 4517 297
rect 4534 245 4586 297
rect 4603 264 4655 297
rect 4672 264 4724 297
rect 4740 264 4792 297
rect 4808 264 4860 297
rect 4876 264 4928 297
rect 4603 245 4628 264
rect 4628 245 4655 264
rect 4672 245 4700 264
rect 4700 245 4724 264
rect 4740 245 4772 264
rect 4772 245 4792 264
rect 4808 245 4844 264
rect 4844 245 4860 264
rect 4876 245 4878 264
rect 4878 245 4916 264
rect 4916 245 4928 264
rect -59 186 -7 192
rect -59 152 -53 186
rect -53 152 -19 186
rect -19 152 -7 186
rect -59 140 -7 152
rect 5 186 57 192
rect 5 152 19 186
rect 19 152 53 186
rect 53 152 57 186
rect 5 140 57 152
rect 94 108 146 114
rect 94 74 100 108
rect 100 74 134 108
rect 134 74 146 108
rect 94 62 146 74
rect 158 108 210 114
rect 158 74 172 108
rect 172 74 206 108
rect 206 74 210 108
rect 158 62 210 74
rect 222 108 274 114
rect 286 108 338 114
rect 350 108 402 114
rect 414 108 466 114
rect 478 108 530 114
rect 542 108 594 114
rect 606 108 658 114
rect 222 74 244 108
rect 244 74 274 108
rect 286 74 316 108
rect 316 74 338 108
rect 350 74 388 108
rect 388 74 402 108
rect 414 74 422 108
rect 422 74 460 108
rect 460 74 466 108
rect 478 74 494 108
rect 494 74 530 108
rect 542 74 566 108
rect 566 74 594 108
rect 606 74 638 108
rect 638 74 658 108
rect 222 62 274 74
rect 286 62 338 74
rect 350 62 402 74
rect 414 62 466 74
rect 478 62 530 74
rect 542 62 594 74
rect 606 62 658 74
rect 670 108 722 114
rect 670 74 676 108
rect 676 74 710 108
rect 710 74 722 108
rect 670 62 722 74
rect 734 108 786 114
rect 734 74 748 108
rect 748 74 782 108
rect 782 74 786 108
rect 734 62 786 74
rect 798 108 850 114
rect 862 108 914 114
rect 926 108 978 114
rect 990 108 1042 114
rect 1054 108 1106 114
rect 798 74 820 108
rect 820 74 850 108
rect 862 74 892 108
rect 892 74 914 108
rect 926 74 964 108
rect 964 74 978 108
rect 990 74 998 108
rect 998 74 1036 108
rect 1036 74 1042 108
rect 1054 74 1070 108
rect 1070 74 1106 108
rect 798 62 850 74
rect 862 62 914 74
rect 926 62 978 74
rect 990 62 1042 74
rect 1054 62 1106 74
rect 1118 62 1170 114
rect 1182 108 1234 114
rect 1182 74 1194 108
rect 1194 74 1228 108
rect 1228 74 1234 108
rect 1182 62 1234 74
rect 1246 108 1298 114
rect 1310 108 1362 114
rect 1374 108 1426 114
rect 1438 108 1490 114
rect 1502 108 1554 114
rect 1566 108 1618 114
rect 1630 108 1682 114
rect 1246 74 1266 108
rect 1266 74 1298 108
rect 1310 74 1338 108
rect 1338 74 1362 108
rect 1374 74 1410 108
rect 1410 74 1426 108
rect 1438 74 1444 108
rect 1444 74 1482 108
rect 1482 74 1490 108
rect 1502 74 1516 108
rect 1516 74 1554 108
rect 1566 74 1588 108
rect 1588 74 1618 108
rect 1630 74 1660 108
rect 1660 74 1682 108
rect 1246 62 1298 74
rect 1310 62 1362 74
rect 1374 62 1426 74
rect 1438 62 1490 74
rect 1502 62 1554 74
rect 1566 62 1618 74
rect 1630 62 1682 74
rect 1694 108 1746 114
rect 1694 74 1698 108
rect 1698 74 1732 108
rect 1732 74 1746 108
rect 1694 62 1746 74
rect 1758 108 1810 114
rect 1758 74 1770 108
rect 1770 74 1804 108
rect 1804 74 1810 108
rect 1758 62 1810 74
rect 1822 108 1874 114
rect 1886 108 1938 114
rect 1950 108 2002 114
rect 2014 108 2066 114
rect 2078 108 2130 114
rect 2142 108 2194 114
rect 1822 74 1842 108
rect 1842 74 1874 108
rect 1886 74 1914 108
rect 1914 74 1938 108
rect 1950 74 1986 108
rect 1986 74 2002 108
rect 2014 74 2020 108
rect 2020 74 2058 108
rect 2058 74 2066 108
rect 2078 74 2092 108
rect 2092 74 2130 108
rect 2142 74 2164 108
rect 2164 74 2194 108
rect 1822 62 1874 74
rect 1886 62 1938 74
rect 1950 62 2002 74
rect 2014 62 2066 74
rect 2078 62 2130 74
rect 2142 62 2194 74
rect 2206 62 2258 114
rect 2270 62 2322 114
rect 2334 108 2386 114
rect 2398 108 2450 114
rect 2462 108 2514 114
rect 2526 108 2578 114
rect 2590 108 2642 114
rect 2654 108 2706 114
rect 2334 74 2364 108
rect 2364 74 2386 108
rect 2398 74 2436 108
rect 2436 74 2450 108
rect 2462 74 2470 108
rect 2470 74 2508 108
rect 2508 74 2514 108
rect 2526 74 2542 108
rect 2542 74 2578 108
rect 2590 74 2614 108
rect 2614 74 2642 108
rect 2654 74 2686 108
rect 2686 74 2706 108
rect 2334 62 2386 74
rect 2398 62 2450 74
rect 2462 62 2514 74
rect 2526 62 2578 74
rect 2590 62 2642 74
rect 2654 62 2706 74
rect 2718 108 2770 114
rect 2718 74 2724 108
rect 2724 74 2758 108
rect 2758 74 2770 108
rect 2718 62 2770 74
rect 2782 108 2834 114
rect 2782 74 2796 108
rect 2796 74 2830 108
rect 2830 74 2834 108
rect 2782 62 2834 74
rect 2846 108 2898 114
rect 2910 108 2962 114
rect 2974 108 3026 114
rect 3039 108 3091 114
rect 3104 108 3156 114
rect 3169 108 3221 114
rect 3234 108 3286 114
rect 2846 74 2868 108
rect 2868 74 2898 108
rect 2910 74 2940 108
rect 2940 74 2962 108
rect 2974 74 3012 108
rect 3012 74 3026 108
rect 3039 74 3046 108
rect 3046 74 3084 108
rect 3084 74 3091 108
rect 3104 74 3118 108
rect 3118 74 3156 108
rect 3169 74 3190 108
rect 3190 74 3221 108
rect 3234 74 3262 108
rect 3262 74 3286 108
rect 2846 62 2898 74
rect 2910 62 2962 74
rect 2974 62 3026 74
rect 3039 62 3091 74
rect 3104 62 3156 74
rect 3169 62 3221 74
rect 3234 62 3286 74
rect 3299 108 3351 114
rect 3299 74 3300 108
rect 3300 74 3334 108
rect 3334 74 3351 108
rect 3299 62 3351 74
rect 3364 62 3416 114
rect 3429 108 3481 114
rect 3494 108 3546 114
rect 3559 108 3611 114
rect 3624 108 3676 114
rect 3689 108 3741 114
rect 3754 108 3806 114
rect 3819 108 3871 114
rect 3429 74 3458 108
rect 3458 74 3481 108
rect 3494 74 3530 108
rect 3530 74 3546 108
rect 3559 74 3564 108
rect 3564 74 3602 108
rect 3602 74 3611 108
rect 3624 74 3636 108
rect 3636 74 3674 108
rect 3674 74 3676 108
rect 3689 74 3708 108
rect 3708 74 3741 108
rect 3754 74 3780 108
rect 3780 74 3806 108
rect 3819 74 3852 108
rect 3852 74 3871 108
rect 3429 62 3481 74
rect 3494 62 3546 74
rect 3559 62 3611 74
rect 3624 62 3676 74
rect 3689 62 3741 74
rect 3754 62 3806 74
rect 3819 62 3871 74
rect 3884 108 3936 114
rect 3884 74 3890 108
rect 3890 74 3924 108
rect 3924 74 3936 108
rect 3884 62 3936 74
rect 3949 108 4001 114
rect 3949 74 3962 108
rect 3962 74 3996 108
rect 3996 74 4001 108
rect 3949 62 4001 74
rect 4014 108 4066 114
rect 4079 108 4131 114
rect 4144 108 4196 114
rect 4209 108 4261 114
rect 4274 108 4326 114
rect 4339 108 4391 114
rect 4404 108 4456 114
rect 4014 74 4034 108
rect 4034 74 4066 108
rect 4079 74 4106 108
rect 4106 74 4131 108
rect 4144 74 4178 108
rect 4178 74 4196 108
rect 4209 74 4212 108
rect 4212 74 4250 108
rect 4250 74 4261 108
rect 4274 74 4284 108
rect 4284 74 4322 108
rect 4322 74 4326 108
rect 4339 74 4356 108
rect 4356 74 4391 108
rect 4404 74 4428 108
rect 4428 74 4456 108
rect 4014 62 4066 74
rect 4079 62 4131 74
rect 4144 62 4196 74
rect 4209 62 4261 74
rect 4274 62 4326 74
rect 4339 62 4391 74
rect 4404 62 4456 74
rect 4469 62 4521 114
rect 4534 62 4586 114
rect 4599 108 4651 114
rect 4664 108 4716 114
rect 4729 108 4781 114
rect 4794 108 4846 114
rect 4859 108 4911 114
rect 4924 108 4976 114
rect 4989 108 5041 114
rect 4599 74 4628 108
rect 4628 74 4651 108
rect 4664 74 4700 108
rect 4700 74 4716 108
rect 4729 74 4734 108
rect 4734 74 4772 108
rect 4772 74 4781 108
rect 4794 74 4806 108
rect 4806 74 4844 108
rect 4844 74 4846 108
rect 4859 74 4878 108
rect 4878 74 4911 108
rect 4924 74 4950 108
rect 4950 74 4976 108
rect 4989 74 5022 108
rect 5022 74 5041 108
rect 4599 62 4651 74
rect 4664 62 4716 74
rect 4729 62 4781 74
rect 4794 62 4846 74
rect 4859 62 4911 74
rect 4924 62 4976 74
rect 4989 62 5041 74
rect 5054 108 5106 114
rect 5054 74 5060 108
rect 5060 74 5094 108
rect 5094 74 5106 108
rect 5054 62 5106 74
rect 5119 108 5171 114
rect 5119 74 5132 108
rect 5132 74 5166 108
rect 5166 74 5171 108
rect 5119 62 5171 74
rect 5184 108 5236 114
rect 5249 108 5301 114
rect 5314 108 5366 114
rect 5379 108 5431 114
rect 5444 108 5496 114
rect 5509 108 5561 114
rect 5574 108 5626 114
rect 5184 74 5204 108
rect 5204 74 5236 108
rect 5249 74 5276 108
rect 5276 74 5301 108
rect 5314 74 5348 108
rect 5348 74 5366 108
rect 5379 74 5382 108
rect 5382 74 5420 108
rect 5420 74 5431 108
rect 5444 74 5454 108
rect 5454 74 5492 108
rect 5492 74 5496 108
rect 5509 74 5526 108
rect 5526 74 5561 108
rect 5574 74 5598 108
rect 5598 74 5626 108
rect 5184 62 5236 74
rect 5249 62 5301 74
rect 5314 62 5366 74
rect 5379 62 5431 74
rect 5444 62 5496 74
rect 5509 62 5561 74
rect 5574 62 5626 74
rect 5639 62 5691 114
rect 5704 108 5756 114
rect 5704 74 5722 108
rect 5722 74 5756 108
rect 5704 62 5756 74
rect 5769 108 5821 114
rect 5834 108 5886 114
rect 5899 108 5951 114
rect 5964 108 6016 114
rect 6029 108 6081 114
rect 6094 108 6146 114
rect 6159 108 6211 114
rect 5769 74 5794 108
rect 5794 74 5821 108
rect 5834 74 5866 108
rect 5866 74 5886 108
rect 5899 74 5900 108
rect 5900 74 5938 108
rect 5938 74 5951 108
rect 5964 74 5972 108
rect 5972 74 6010 108
rect 6010 74 6016 108
rect 6029 74 6044 108
rect 6044 74 6081 108
rect 6094 74 6116 108
rect 6116 74 6146 108
rect 6159 74 6188 108
rect 6188 74 6211 108
rect 5769 62 5821 74
rect 5834 62 5886 74
rect 5899 62 5951 74
rect 5964 62 6016 74
rect 6029 62 6081 74
rect 6094 62 6146 74
rect 6159 62 6211 74
rect 6224 108 6276 114
rect 6224 74 6226 108
rect 6226 74 6260 108
rect 6260 74 6276 108
rect 6224 62 6276 74
rect 6289 108 6341 114
rect 6289 74 6298 108
rect 6298 74 6332 108
rect 6332 74 6341 108
rect 6289 62 6341 74
rect 6354 108 6406 114
rect 6354 74 6370 108
rect 6370 74 6404 108
rect 6404 74 6406 108
rect 6354 62 6406 74
rect 6419 108 6471 114
rect 6484 108 6536 114
rect 6549 108 6601 114
rect 6614 108 6666 114
rect 6679 108 6731 114
rect 6419 74 6442 108
rect 6442 74 6471 108
rect 6484 74 6514 108
rect 6514 74 6536 108
rect 6549 74 6586 108
rect 6586 74 6601 108
rect 6614 74 6620 108
rect 6620 74 6658 108
rect 6658 74 6666 108
rect 6679 74 6692 108
rect 6692 74 6731 108
rect 6419 62 6471 74
rect 6484 62 6536 74
rect 6549 62 6601 74
rect 6614 62 6666 74
rect 6679 62 6731 74
rect -182 -140 -130 -88
rect -182 -204 -130 -152
rect 21657 -3473 21709 -3421
rect 21657 -3537 21709 -3485
rect 21188 -3731 21240 -3679
rect 21188 -3834 21240 -3782
rect 21117 -5194 21169 -5142
rect 21181 -5194 21233 -5142
rect 21370 -10040 21379 -10016
rect 21379 -10040 21413 -10016
rect 21413 -10040 21422 -10016
rect 21370 -10068 21422 -10040
rect 21370 -10112 21379 -10080
rect 21379 -10112 21413 -10080
rect 21413 -10112 21422 -10080
rect 21370 -10132 21422 -10112
rect 21370 -10150 21422 -10144
rect 21370 -10184 21379 -10150
rect 21379 -10184 21413 -10150
rect 21413 -10184 21422 -10150
rect 21370 -10196 21422 -10184
rect 21214 -10366 21266 -10354
rect 21214 -10400 21223 -10366
rect 21223 -10400 21257 -10366
rect 21257 -10400 21266 -10366
rect 21214 -10406 21266 -10400
rect 21214 -10438 21266 -10418
rect 21214 -10470 21223 -10438
rect 21223 -10470 21257 -10438
rect 21257 -10470 21266 -10438
rect 21214 -10510 21266 -10482
rect 21214 -10534 21223 -10510
rect 21223 -10534 21257 -10510
rect 21257 -10534 21266 -10510
rect 21526 -10366 21578 -10354
rect 21526 -10400 21535 -10366
rect 21535 -10400 21569 -10366
rect 21569 -10400 21578 -10366
rect 21526 -10406 21578 -10400
rect 21526 -10438 21578 -10418
rect 21526 -10470 21535 -10438
rect 21535 -10470 21569 -10438
rect 21569 -10470 21578 -10438
rect 21526 -10510 21578 -10482
rect 21526 -10534 21535 -10510
rect 21535 -10534 21569 -10510
rect 21569 -10534 21578 -10510
rect 21338 -14518 21390 -14466
rect 21431 -14518 21483 -14466
rect 21524 -14518 21576 -14466
<< metal2 >>
rect 3651 1949 3660 2085
rect 3796 2029 3821 2085
rect 3877 2029 3902 2085
rect 3958 2029 3967 2085
rect 3796 2027 3823 2029
rect 3875 2027 3905 2029
rect 3957 2027 3967 2029
rect 3796 2005 3967 2027
rect 3796 1949 3821 2005
rect 3877 1949 3902 2005
rect 3958 1949 3967 2005
rect 3651 432 3660 434
rect 3716 432 3740 434
rect 3796 432 3821 434
rect 3877 432 3902 434
rect 3958 432 3967 434
rect 88 380 94 432
rect 146 380 158 432
rect 210 380 222 432
rect 274 380 286 432
rect 338 380 350 432
rect 402 380 414 432
rect 466 380 478 432
rect 530 380 542 432
rect 594 380 606 432
rect 658 380 670 432
rect 722 380 734 432
rect 786 380 798 432
rect 850 380 862 432
rect 914 380 926 432
rect 978 380 990 432
rect 1042 380 1054 432
rect 1106 380 1118 432
rect 1170 380 1182 432
rect 1234 380 1246 432
rect 1298 380 1310 432
rect 1362 380 1374 432
rect 1426 380 1438 432
rect 1490 380 1502 432
rect 1554 380 1566 432
rect 1618 380 1630 432
rect 1682 380 1694 432
rect 1746 380 1758 432
rect 1810 380 1822 432
rect 1874 380 1886 432
rect 1938 380 1950 432
rect 2002 380 2014 432
rect 2066 380 2078 432
rect 2130 380 2142 432
rect 2194 380 2206 432
rect 2258 380 2270 432
rect 2322 380 2334 432
rect 2386 380 2398 432
rect 2450 380 2462 432
rect 2514 380 2526 432
rect 2578 380 2590 432
rect 2642 380 2654 432
rect 2706 380 2718 432
rect 2770 380 2782 432
rect 2834 380 2846 432
rect 2898 380 2910 432
rect 2962 380 2974 432
rect 3026 380 3039 432
rect 3091 380 3104 432
rect 3156 380 3169 432
rect 3221 380 3234 432
rect 3286 380 3299 432
rect 3351 380 3364 432
rect 3416 380 3429 432
rect 3481 380 3494 432
rect 3546 380 3559 432
rect 3611 380 3624 432
rect 3806 380 3819 432
rect 3877 380 3884 432
rect 4001 380 4014 432
rect 4066 380 4079 432
rect 4131 380 4144 432
rect 4196 380 4209 432
rect 4261 380 4274 432
rect 4326 380 4339 432
rect 4391 380 4404 432
rect 4456 380 4469 432
rect 4521 380 4534 432
rect 4586 380 4599 432
rect 4651 380 4664 432
rect 4716 380 4729 432
rect 4781 380 4794 432
rect 4846 380 4859 432
rect 4911 380 4924 432
rect 4976 380 4989 432
rect 5041 380 5054 432
rect 5106 380 5119 432
rect 5171 380 5184 432
rect 5236 380 5249 432
rect 5301 380 5314 432
rect 5366 380 5379 432
rect 5431 380 5444 432
rect 5496 380 5509 432
rect 5561 380 5574 432
rect 5626 380 5639 432
rect 5691 380 5704 432
rect 5756 380 5769 432
rect 5821 380 5834 432
rect 5886 380 5899 432
rect 5951 380 5964 432
rect 6016 380 6029 432
rect 6081 380 6094 432
rect 6146 380 6159 432
rect 6211 380 6224 432
rect 6276 380 6289 432
rect 6341 380 6354 432
rect 6406 380 6419 432
rect 6471 380 6484 432
rect 6536 380 6549 432
rect 6601 380 6614 432
rect 6666 380 6679 432
rect 6731 380 6737 432
rect 3651 378 3660 380
rect 3716 378 3740 380
rect 3796 378 3821 380
rect 3877 378 3902 380
rect 3958 378 3967 380
rect 2204 296 2213 298
rect 2269 296 2295 298
rect 2351 296 2377 298
rect 2433 296 2459 298
rect 2515 296 2541 298
rect 2597 296 2623 298
rect 2679 296 2704 298
rect 2760 296 2785 298
rect 2841 296 2866 298
rect 2922 296 2947 298
rect 3003 296 3028 298
rect 3084 296 3093 298
rect 2204 244 2210 296
rect 2269 244 2279 296
rect 2538 244 2541 296
rect 2607 244 2623 296
rect 2679 244 2693 296
rect 2760 244 2762 296
rect 3019 244 3028 296
rect 3087 244 3093 296
rect 2204 242 2213 244
rect 2269 242 2295 244
rect 2351 242 2377 244
rect 2433 242 2459 244
rect 2515 242 2541 244
rect 2597 242 2623 244
rect 2679 242 2704 244
rect 2760 242 2785 244
rect 2841 242 2866 244
rect 2922 242 2947 244
rect 3003 242 3028 244
rect 3084 242 3093 244
rect 4045 297 4054 299
rect 4110 297 4136 299
rect 4192 297 4218 299
rect 4274 297 4300 299
rect 4356 297 4382 299
rect 4438 297 4464 299
rect 4520 297 4545 299
rect 4601 297 4626 299
rect 4682 297 4707 299
rect 4763 297 4788 299
rect 4844 297 4869 299
rect 4925 297 4934 299
rect 4045 245 4051 297
rect 4110 245 4120 297
rect 4379 245 4382 297
rect 4448 245 4464 297
rect 4520 245 4534 297
rect 4601 245 4603 297
rect 4860 245 4869 297
rect 4928 245 4934 297
rect 4045 243 4054 245
rect 4110 243 4136 245
rect 4192 243 4218 245
rect 4274 243 4300 245
rect 4356 243 4382 245
rect 4438 243 4464 245
rect 4520 243 4545 245
rect 4601 243 4626 245
rect 4682 243 4707 245
rect 4763 243 4788 245
rect 4844 243 4869 245
rect 4925 243 4934 245
rect -185 140 -59 192
rect -7 140 5 192
rect 57 140 63 192
rect -185 116 -107 140
tri -107 116 -83 140 nw
rect -185 114 -109 116
tri -109 114 -107 116 nw
rect 3651 114 3660 116
rect 3716 114 3740 116
rect 3796 114 3821 116
rect 3877 114 3902 116
rect 3958 114 3967 116
rect -185 -88 -130 114
tri -130 93 -109 114 nw
rect 88 62 94 114
rect 146 62 158 114
rect 210 62 222 114
rect 274 62 286 114
rect 338 62 350 114
rect 402 62 414 114
rect 466 62 478 114
rect 530 62 542 114
rect 594 62 606 114
rect 658 62 670 114
rect 722 62 734 114
rect 786 62 798 114
rect 850 62 862 114
rect 914 62 926 114
rect 978 62 990 114
rect 1042 62 1054 114
rect 1106 62 1118 114
rect 1170 62 1182 114
rect 1234 62 1246 114
rect 1298 62 1310 114
rect 1362 62 1374 114
rect 1426 62 1438 114
rect 1490 62 1502 114
rect 1554 62 1566 114
rect 1618 62 1630 114
rect 1682 62 1694 114
rect 1746 62 1758 114
rect 1810 62 1822 114
rect 1874 62 1886 114
rect 1938 62 1950 114
rect 2002 62 2014 114
rect 2066 62 2078 114
rect 2130 62 2142 114
rect 2194 62 2206 114
rect 2258 62 2270 114
rect 2322 62 2334 114
rect 2386 62 2398 114
rect 2450 62 2462 114
rect 2514 62 2526 114
rect 2578 62 2590 114
rect 2642 62 2654 114
rect 2706 62 2718 114
rect 2770 62 2782 114
rect 2834 62 2846 114
rect 2898 62 2910 114
rect 2962 62 2974 114
rect 3026 62 3039 114
rect 3091 62 3104 114
rect 3156 62 3169 114
rect 3221 62 3234 114
rect 3286 62 3299 114
rect 3351 62 3364 114
rect 3416 62 3429 114
rect 3481 62 3494 114
rect 3546 62 3559 114
rect 3611 62 3624 114
rect 3806 62 3819 114
rect 3877 62 3884 114
rect 4001 62 4014 114
rect 4066 62 4079 114
rect 4131 62 4144 114
rect 4196 62 4209 114
rect 4261 62 4274 114
rect 4326 62 4339 114
rect 4391 62 4404 114
rect 4456 62 4469 114
rect 4521 62 4534 114
rect 4586 62 4599 114
rect 4651 62 4664 114
rect 4716 62 4729 114
rect 4781 62 4794 114
rect 4846 62 4859 114
rect 4911 62 4924 114
rect 4976 62 4989 114
rect 5041 62 5054 114
rect 5106 62 5119 114
rect 5171 62 5184 114
rect 5236 62 5249 114
rect 5301 62 5314 114
rect 5366 62 5379 114
rect 5431 62 5444 114
rect 5496 62 5509 114
rect 5561 62 5574 114
rect 5626 62 5639 114
rect 5691 62 5704 114
rect 5756 62 5769 114
rect 5821 62 5834 114
rect 5886 62 5899 114
rect 5951 62 5964 114
rect 6016 62 6029 114
rect 6081 62 6094 114
rect 6146 62 6159 114
rect 6211 62 6224 114
rect 6276 62 6289 114
rect 6341 62 6354 114
rect 6406 62 6419 114
rect 6471 62 6484 114
rect 6536 62 6549 114
rect 6601 62 6614 114
rect 6666 62 6679 114
rect 6731 62 6737 114
rect 3651 60 3660 62
rect 3716 60 3740 62
rect 3796 60 3821 62
rect 3877 60 3902 62
rect 3958 60 3967 62
rect -185 -140 -182 -88
rect -185 -152 -130 -140
rect -185 -204 -182 -152
rect -185 -207 -130 -204
tri -185 -210 -182 -207 ne
rect -182 -210 -130 -207
rect 21657 -3421 21709 -3415
rect 21657 -3485 21709 -3473
rect 21709 -3537 21972 -3491
rect 21657 -3543 21972 -3537
rect 21188 -3679 21240 -3673
rect 21188 -3782 21240 -3731
rect 21188 -5142 21240 -3834
rect 21111 -5194 21117 -5142
rect 21169 -5194 21181 -5142
rect 21233 -5194 21240 -5142
rect 21188 -10348 21240 -5194
rect 21370 -10016 21422 -10010
tri 21422 -10026 21424 -10024 sw
rect 21422 -10055 21424 -10026
tri 21424 -10055 21453 -10026 sw
tri 21891 -10055 21920 -10026 se
rect 21920 -10055 21972 -3543
rect 21422 -10068 21972 -10055
rect 21370 -10080 21972 -10068
rect 21422 -10107 21972 -10080
rect 21370 -10144 21422 -10132
tri 21422 -10137 21452 -10107 nw
rect 21370 -10202 21422 -10196
rect 21188 -10354 21578 -10348
rect 21188 -10406 21214 -10354
rect 21266 -10406 21526 -10354
rect 21188 -10418 21578 -10406
rect 21188 -10470 21214 -10418
rect 21266 -10470 21526 -10418
rect 21188 -10482 21578 -10470
rect 21188 -10534 21214 -10482
rect 21266 -10534 21526 -10482
rect 21188 -10540 21578 -10534
rect 21332 -14466 21582 -14436
rect 21332 -14518 21338 -14466
rect 21390 -14518 21431 -14466
rect 21483 -14518 21524 -14466
rect 21576 -14518 21582 -14466
rect 21332 -14548 21582 -14518
<< via2 >>
rect 3660 2079 3796 2085
rect 3660 2027 3661 2079
rect 3661 2027 3713 2079
rect 3713 2027 3742 2079
rect 3742 2027 3794 2079
rect 3794 2027 3796 2079
rect 3821 2079 3877 2085
rect 3821 2029 3823 2079
rect 3823 2029 3875 2079
rect 3875 2029 3877 2079
rect 3902 2079 3958 2085
rect 3902 2029 3905 2079
rect 3905 2029 3957 2079
rect 3957 2029 3958 2079
rect 3660 2001 3796 2027
rect 3660 1949 3661 2001
rect 3661 1949 3713 2001
rect 3713 1949 3742 2001
rect 3742 1949 3794 2001
rect 3794 1949 3796 2001
rect 3821 2001 3877 2005
rect 3821 1949 3823 2001
rect 3823 1949 3875 2001
rect 3875 1949 3877 2001
rect 3902 2001 3958 2005
rect 3902 1949 3905 2001
rect 3905 1949 3957 2001
rect 3957 1949 3958 2001
rect 3660 432 3716 434
rect 3740 432 3796 434
rect 3821 432 3877 434
rect 3902 432 3958 434
rect 3660 380 3676 432
rect 3676 380 3689 432
rect 3689 380 3716 432
rect 3740 380 3741 432
rect 3741 380 3754 432
rect 3754 380 3796 432
rect 3821 380 3871 432
rect 3871 380 3877 432
rect 3902 380 3936 432
rect 3936 380 3949 432
rect 3949 380 3958 432
rect 3660 378 3716 380
rect 3740 378 3796 380
rect 3821 378 3877 380
rect 3902 378 3958 380
rect 2213 296 2269 298
rect 2295 296 2351 298
rect 2377 296 2433 298
rect 2459 296 2515 298
rect 2541 296 2597 298
rect 2623 296 2679 298
rect 2704 296 2760 298
rect 2785 296 2841 298
rect 2866 296 2922 298
rect 2947 296 3003 298
rect 3028 296 3084 298
rect 2213 244 2262 296
rect 2262 244 2269 296
rect 2295 244 2331 296
rect 2331 244 2348 296
rect 2348 244 2351 296
rect 2377 244 2400 296
rect 2400 244 2417 296
rect 2417 244 2433 296
rect 2459 244 2469 296
rect 2469 244 2486 296
rect 2486 244 2515 296
rect 2541 244 2555 296
rect 2555 244 2597 296
rect 2623 244 2624 296
rect 2624 244 2676 296
rect 2676 244 2679 296
rect 2704 244 2745 296
rect 2745 244 2760 296
rect 2785 244 2814 296
rect 2814 244 2831 296
rect 2831 244 2841 296
rect 2866 244 2883 296
rect 2883 244 2899 296
rect 2899 244 2922 296
rect 2947 244 2951 296
rect 2951 244 2967 296
rect 2967 244 3003 296
rect 3028 244 3035 296
rect 3035 244 3084 296
rect 2213 242 2269 244
rect 2295 242 2351 244
rect 2377 242 2433 244
rect 2459 242 2515 244
rect 2541 242 2597 244
rect 2623 242 2679 244
rect 2704 242 2760 244
rect 2785 242 2841 244
rect 2866 242 2922 244
rect 2947 242 3003 244
rect 3028 242 3084 244
rect 4054 297 4110 299
rect 4136 297 4192 299
rect 4218 297 4274 299
rect 4300 297 4356 299
rect 4382 297 4438 299
rect 4464 297 4520 299
rect 4545 297 4601 299
rect 4626 297 4682 299
rect 4707 297 4763 299
rect 4788 297 4844 299
rect 4869 297 4925 299
rect 4054 245 4103 297
rect 4103 245 4110 297
rect 4136 245 4172 297
rect 4172 245 4189 297
rect 4189 245 4192 297
rect 4218 245 4241 297
rect 4241 245 4258 297
rect 4258 245 4274 297
rect 4300 245 4310 297
rect 4310 245 4327 297
rect 4327 245 4356 297
rect 4382 245 4396 297
rect 4396 245 4438 297
rect 4464 245 4465 297
rect 4465 245 4517 297
rect 4517 245 4520 297
rect 4545 245 4586 297
rect 4586 245 4601 297
rect 4626 245 4655 297
rect 4655 245 4672 297
rect 4672 245 4682 297
rect 4707 245 4724 297
rect 4724 245 4740 297
rect 4740 245 4763 297
rect 4788 245 4792 297
rect 4792 245 4808 297
rect 4808 245 4844 297
rect 4869 245 4876 297
rect 4876 245 4925 297
rect 4054 243 4110 245
rect 4136 243 4192 245
rect 4218 243 4274 245
rect 4300 243 4356 245
rect 4382 243 4438 245
rect 4464 243 4520 245
rect 4545 243 4601 245
rect 4626 243 4682 245
rect 4707 243 4763 245
rect 4788 243 4844 245
rect 4869 243 4925 245
rect 3660 114 3716 116
rect 3740 114 3796 116
rect 3821 114 3877 116
rect 3902 114 3958 116
rect 3660 62 3676 114
rect 3676 62 3689 114
rect 3689 62 3716 114
rect 3740 62 3741 114
rect 3741 62 3754 114
rect 3754 62 3796 114
rect 3821 62 3871 114
rect 3871 62 3877 114
rect 3902 62 3936 114
rect 3936 62 3949 114
rect 3949 62 3958 114
rect 3660 60 3716 62
rect 3740 60 3796 62
rect 3821 60 3877 62
rect 3902 60 3958 62
<< metal3 >>
rect 3655 2085 3963 2090
rect 3655 1949 3660 2085
rect 3796 2029 3821 2085
rect 3877 2029 3902 2085
rect 3958 2029 3963 2085
rect 3796 2005 3963 2029
rect 3796 1949 3821 2005
rect 3877 1949 3902 2005
rect 3958 1949 3963 2005
rect 3655 434 3963 1949
rect 3655 378 3660 434
rect 3716 378 3740 434
rect 3796 378 3821 434
rect 3877 378 3902 434
rect 3958 378 3963 434
rect 2208 298 3089 303
rect 2208 242 2213 298
rect 2269 242 2295 298
rect 2351 242 2377 298
rect 2433 242 2459 298
rect 2515 242 2541 298
rect 2597 242 2623 298
rect 2679 242 2704 298
rect 2760 242 2785 298
rect 2841 242 2866 298
rect 2922 242 2947 298
rect 3003 242 3028 298
rect 3084 242 3089 298
rect 2208 237 3089 242
rect 3655 116 3963 378
rect 4049 299 4930 304
rect 4049 243 4054 299
rect 4110 243 4136 299
rect 4192 243 4218 299
rect 4274 243 4300 299
rect 4356 243 4382 299
rect 4438 243 4464 299
rect 4520 243 4545 299
rect 4601 243 4626 299
rect 4682 243 4707 299
rect 4763 243 4788 299
rect 4844 243 4869 299
rect 4925 243 4930 299
rect 4049 238 4930 243
rect 3655 60 3660 116
rect 3716 60 3740 116
rect 3796 60 3821 116
rect 3877 60 3902 116
rect 3958 60 3963 116
rect 3655 55 3963 60
use sky130_fd_io__gpio_ovtv2_hotswap_guardrings  sky130_fd_io__gpio_ovtv2_hotswap_guardrings_0
timestamp 1666199351
transform -1 0 22914 0 -1 3000
box 0 0 26980 8664
use sky130_fd_pr__nfet_01v8__example_5595914180834  sky130_fd_pr__nfet_01v8__example_5595914180834_0
timestamp 1666199351
transform -1 0 21524 0 1 -10540
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_5595914180837  sky130_fd_pr__pfet_01v8__example_5595914180837_0
timestamp 1666199351
transform -1 0 21125 0 1 -3986
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_5595914180847  sky130_fd_pr__pfet_01v8__example_5595914180847_0
timestamp 1666199351
transform 0 -1 1066 1 0 119
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_5595914180847  sky130_fd_pr__pfet_01v8__example_5595914180847_1
timestamp 1666199351
transform 0 1 1198 1 0 119
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_5595914180847  sky130_fd_pr__pfet_01v8__example_5595914180847_2
timestamp 1666199351
transform 0 1 3462 1 0 119
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_5595914180847  sky130_fd_pr__pfet_01v8__example_5595914180847_3
timestamp 1666199351
transform 0 -1 3330 1 0 119
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_5595914180847  sky130_fd_pr__pfet_01v8__example_5595914180847_4
timestamp 1666199351
transform 0 1 5726 1 0 119
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_5595914180847  sky130_fd_pr__pfet_01v8__example_5595914180847_5
timestamp 1666199351
transform 0 -1 5594 1 0 119
box -1 0 257 1
<< labels >>
flabel metal1 s -2935 -4716 -2763 -4547 3 FreeSans 520 0 0 0 VPB_DRVR
port 1 nsew
flabel metal1 s -3365 -5079 -3205 -4949 3 FreeSans 520 0 0 0 VSSD
port 2 nsew
flabel metal1 s 20670 -8075 20849 -7911 3 FreeSans 200 180 0 0 VDDIO
port 3 nsew
flabel metal2 s 21188 -4142 21240 -4102 3 FreeSans 520 0 0 0 PU_H_N
port 4 nsew
flabel metal2 s 4139 247 4197 299 3 FreeSans 520 0 0 0 VDDIO
port 3 nsew
flabel metal2 s 4469 380 4569 432 3 FreeSans 520 0 0 0 PAD
port 5 nsew
flabel metal2 s 21920 -3759 21972 -3681 3 FreeSans 520 0 0 0 PUG_H
port 6 nsew
flabel locali s 21377 -10630 21418 -10582 3 FreeSans 520 0 0 0 NGHS_H
port 7 nsew
flabel locali s 20963 -4067 21021 -4037 3 FreeSans 520 0 0 0 PGHS_H
port 8 nsew
flabel locali s 21665 -10335 21705 -10236 3 FreeSans 520 0 0 0 VSSIO
port 9 nsew
<< properties >>
string GDS_END 36449962
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 36309346
<< end >>
