magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 3 157 272 203
rect 3 21 808 157
rect 25 -17 59 21
<< scnmos >>
rect 82 47 112 177
rect 166 47 196 177
rect 283 47 313 131
rect 367 47 397 131
rect 532 47 562 131
rect 616 47 646 131
rect 700 47 730 131
<< scpmoshvt >>
rect 82 297 112 497
rect 166 297 196 497
rect 283 297 313 425
rect 355 297 385 425
rect 544 369 574 497
rect 635 369 665 497
rect 719 369 749 497
<< ndiff >>
rect 29 161 82 177
rect 29 127 37 161
rect 71 127 82 161
rect 29 93 82 127
rect 29 59 37 93
rect 71 59 82 93
rect 29 47 82 59
rect 112 129 166 177
rect 112 95 122 129
rect 156 95 166 129
rect 112 47 166 95
rect 196 131 246 177
rect 196 106 283 131
rect 196 72 206 106
rect 240 72 283 106
rect 196 47 283 72
rect 313 106 367 131
rect 313 72 323 106
rect 357 72 367 106
rect 313 47 367 72
rect 397 97 532 131
rect 397 63 407 97
rect 441 63 488 97
rect 522 63 532 97
rect 397 47 532 63
rect 562 106 616 131
rect 562 72 572 106
rect 606 72 616 106
rect 562 47 616 72
rect 646 47 700 131
rect 730 103 782 131
rect 730 69 740 103
rect 774 69 782 103
rect 730 47 782 69
<< pdiff >>
rect 29 481 82 497
rect 29 447 37 481
rect 71 447 82 481
rect 29 413 82 447
rect 29 379 37 413
rect 71 379 82 413
rect 29 345 82 379
rect 29 311 37 345
rect 71 311 82 345
rect 29 297 82 311
rect 112 458 166 497
rect 112 424 122 458
rect 156 424 166 458
rect 112 369 166 424
rect 112 335 122 369
rect 156 335 166 369
rect 112 297 166 335
rect 196 481 248 497
rect 196 447 206 481
rect 240 447 248 481
rect 492 472 544 497
rect 196 425 248 447
rect 492 438 500 472
rect 534 438 544 472
rect 196 297 283 425
rect 313 297 355 425
rect 385 359 438 425
rect 492 369 544 438
rect 574 485 635 497
rect 574 451 591 485
rect 625 451 635 485
rect 574 369 635 451
rect 665 485 719 497
rect 665 451 675 485
rect 709 451 719 485
rect 665 369 719 451
rect 749 472 801 497
rect 749 438 759 472
rect 793 438 801 472
rect 749 369 801 438
rect 385 325 395 359
rect 429 325 438 359
rect 385 297 438 325
<< ndiffc >>
rect 37 127 71 161
rect 37 59 71 93
rect 122 95 156 129
rect 206 72 240 106
rect 323 72 357 106
rect 407 63 441 97
rect 488 63 522 97
rect 572 72 606 106
rect 740 69 774 103
<< pdiffc >>
rect 37 447 71 481
rect 37 379 71 413
rect 37 311 71 345
rect 122 424 156 458
rect 122 335 156 369
rect 206 447 240 481
rect 500 438 534 472
rect 591 451 625 485
rect 675 451 709 485
rect 759 438 793 472
rect 395 325 429 359
<< poly >>
rect 82 497 112 523
rect 166 497 196 523
rect 544 497 574 523
rect 635 497 665 523
rect 719 497 749 523
rect 283 425 313 451
rect 355 425 385 451
rect 82 265 112 297
rect 166 265 196 297
rect 283 265 313 297
rect 82 249 217 265
rect 82 215 173 249
rect 207 215 217 249
rect 82 199 217 215
rect 259 249 313 265
rect 259 215 269 249
rect 303 215 313 249
rect 355 275 385 297
rect 544 287 574 369
rect 635 327 665 369
rect 355 265 397 275
rect 355 249 413 265
rect 355 242 369 249
rect 259 199 313 215
rect 359 215 369 242
rect 403 215 413 249
rect 359 199 413 215
rect 458 248 574 287
rect 458 214 468 248
rect 502 214 574 248
rect 458 211 574 214
rect 616 311 670 327
rect 616 277 626 311
rect 660 277 670 311
rect 616 261 670 277
rect 719 265 749 369
rect 82 177 112 199
rect 166 177 196 199
rect 283 131 313 199
rect 367 131 397 199
rect 458 153 562 211
rect 532 131 562 153
rect 616 131 646 261
rect 719 249 790 265
rect 719 229 746 249
rect 700 215 746 229
rect 780 215 790 249
rect 700 199 790 215
rect 700 131 730 199
rect 82 21 112 47
rect 166 21 196 47
rect 283 21 313 47
rect 367 21 397 47
rect 532 21 562 47
rect 616 21 646 47
rect 700 21 730 47
<< polycont >>
rect 173 215 207 249
rect 269 215 303 249
rect 369 215 403 249
rect 468 214 502 248
rect 626 277 660 311
rect 746 215 780 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 37 481 71 527
rect 37 413 71 447
rect 37 345 71 379
rect 37 289 71 311
rect 105 458 156 493
rect 105 424 122 458
rect 190 481 256 527
rect 190 447 206 481
rect 240 447 256 481
rect 500 474 534 493
rect 675 485 725 527
rect 308 472 534 474
rect 105 369 156 424
rect 308 440 500 472
rect 308 395 342 440
rect 105 335 122 369
rect 105 305 156 335
rect 190 361 342 395
rect 488 438 500 440
rect 575 451 591 485
rect 625 451 641 485
rect 488 413 534 438
rect 37 161 71 186
rect 37 93 71 127
rect 37 17 71 59
rect 105 162 139 305
rect 190 265 224 361
rect 395 359 429 381
rect 488 379 570 413
rect 429 325 502 343
rect 173 249 224 265
rect 207 215 224 249
rect 173 199 224 215
rect 269 249 335 323
rect 395 309 502 325
rect 303 215 335 249
rect 269 199 335 215
rect 369 249 427 275
rect 403 215 427 249
rect 369 199 427 215
rect 468 248 502 309
rect 468 165 502 214
rect 105 129 156 162
rect 105 95 122 129
rect 323 131 502 165
rect 536 174 570 379
rect 607 401 641 451
rect 709 451 725 485
rect 675 435 725 451
rect 759 472 793 493
rect 759 401 793 438
rect 607 367 793 401
rect 610 311 706 331
rect 610 277 626 311
rect 660 277 706 311
rect 610 271 706 277
rect 536 140 606 174
rect 654 153 706 271
rect 746 249 798 331
rect 780 215 798 249
rect 746 153 798 215
rect 323 106 357 131
rect 105 51 156 95
rect 190 72 206 106
rect 240 72 276 106
rect 190 17 276 72
rect 572 106 606 140
rect 323 51 357 72
rect 391 63 407 97
rect 441 63 488 97
rect 522 63 538 97
rect 391 17 538 63
rect 572 51 606 72
rect 721 103 801 119
rect 721 69 740 103
rect 774 69 801 103
rect 721 17 801 69
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel pwell s 25 -17 59 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 25 527 59 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 25 -17 59 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 25 527 59 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 25 527 59 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 25 -17 59 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 764 221 798 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 764 289 798 323 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 764 153 798 187 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 301 221 335 255 0 FreeSans 200 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 393 221 427 255 0 FreeSans 200 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 117 85 151 119 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 672 289 706 323 0 FreeSans 200 0 0 0 B2
port 4 nsew signal input
flabel locali s 301 289 335 323 0 FreeSans 200 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 117 425 151 459 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 117 357 151 391 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
rlabel comment s 0 0 0 0 4 a2bb2o_2
rlabel metal1 s 0 -48 828 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 3934450
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3926722
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 20.700 0.000 
<< end >>
