magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 832 157 1287 203
rect 1 21 1287 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 435 47 465 131
rect 530 47 560 119
rect 627 47 657 119
rect 722 47 752 131
rect 910 47 940 177
rect 1004 47 1034 177
rect 1095 47 1125 177
rect 1179 47 1209 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 435 369 465 497
rect 530 413 560 497
rect 614 413 644 497
rect 711 413 741 497
rect 910 297 940 497
rect 1004 297 1034 497
rect 1088 297 1118 497
rect 1179 297 1209 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 119 351 131
rect 299 85 307 119
rect 341 85 351 119
rect 299 47 351 85
rect 381 89 435 131
rect 381 55 391 89
rect 425 55 435 89
rect 381 47 435 55
rect 465 119 515 131
rect 858 165 910 177
rect 858 131 866 165
rect 900 131 910 165
rect 672 119 722 131
rect 465 47 530 119
rect 560 107 627 119
rect 560 73 570 107
rect 604 73 627 107
rect 560 47 627 73
rect 657 47 722 119
rect 752 106 804 131
rect 752 72 762 106
rect 796 72 804 106
rect 752 47 804 72
rect 858 97 910 131
rect 858 63 866 97
rect 900 63 910 97
rect 858 47 910 63
rect 940 47 1004 177
rect 1034 89 1095 177
rect 1034 55 1051 89
rect 1085 55 1095 89
rect 1034 47 1095 55
rect 1125 89 1179 177
rect 1125 55 1135 89
rect 1169 55 1179 89
rect 1125 47 1179 55
rect 1209 93 1261 177
rect 1209 59 1219 93
rect 1253 59 1261 93
rect 1209 47 1261 59
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 483 351 497
rect 299 449 307 483
rect 341 449 351 483
rect 299 415 351 449
rect 299 381 307 415
rect 341 381 351 415
rect 299 369 351 381
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 369 435 383
rect 465 413 530 497
rect 560 485 614 497
rect 560 451 570 485
rect 604 451 614 485
rect 560 413 614 451
rect 644 413 711 497
rect 741 485 793 497
rect 741 451 751 485
rect 785 451 793 485
rect 741 413 793 451
rect 856 485 910 497
rect 856 451 864 485
rect 898 451 910 485
rect 465 369 515 413
rect 856 297 910 451
rect 940 471 1004 497
rect 940 437 960 471
rect 994 437 1004 471
rect 940 368 1004 437
rect 940 334 960 368
rect 994 334 1004 368
rect 940 297 1004 334
rect 1034 489 1088 497
rect 1034 455 1044 489
rect 1078 455 1088 489
rect 1034 421 1088 455
rect 1034 387 1044 421
rect 1078 387 1088 421
rect 1034 297 1088 387
rect 1118 477 1179 497
rect 1118 443 1131 477
rect 1165 443 1179 477
rect 1118 297 1179 443
rect 1209 475 1261 497
rect 1209 441 1219 475
rect 1253 441 1261 475
rect 1209 384 1261 441
rect 1209 350 1219 384
rect 1253 350 1261 384
rect 1209 297 1261 350
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 85 341 119
rect 391 55 425 89
rect 866 131 900 165
rect 570 73 604 107
rect 762 72 796 106
rect 866 63 900 97
rect 1051 55 1085 89
rect 1135 55 1169 89
rect 1219 59 1253 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 449 341 483
rect 307 381 341 415
rect 391 451 425 485
rect 391 383 425 417
rect 570 451 604 485
rect 751 451 785 485
rect 864 451 898 485
rect 960 437 994 471
rect 960 334 994 368
rect 1044 455 1078 489
rect 1044 387 1078 421
rect 1131 443 1165 477
rect 1219 441 1253 475
rect 1219 350 1253 384
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 435 497 465 523
rect 530 497 560 523
rect 614 497 644 523
rect 711 497 741 523
rect 910 497 940 523
rect 1004 497 1034 523
rect 1088 497 1118 523
rect 1179 497 1209 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 22 264 76 280
rect 163 274 193 363
rect 22 230 32 264
rect 66 230 76 264
rect 22 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 351 241 381 369
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 294 225 381 241
rect 294 191 304 225
rect 338 191 381 225
rect 435 219 465 369
rect 530 337 560 413
rect 614 376 644 413
rect 603 366 669 376
rect 507 321 561 337
rect 603 332 619 366
rect 653 332 669 366
rect 603 322 669 332
rect 711 373 741 413
rect 711 357 799 373
rect 711 323 755 357
rect 789 323 799 357
rect 507 287 517 321
rect 551 287 561 321
rect 711 307 799 323
rect 507 280 561 287
rect 507 271 657 280
rect 527 250 657 271
rect 294 175 381 191
rect 351 131 381 175
rect 423 203 477 219
rect 423 169 433 203
rect 467 169 477 203
rect 423 153 477 169
rect 519 198 585 208
rect 519 164 535 198
rect 569 164 585 198
rect 519 154 585 164
rect 435 131 465 153
rect 530 119 560 154
rect 627 119 657 250
rect 722 131 752 307
rect 910 259 940 297
rect 1004 265 1034 297
rect 1088 265 1118 297
rect 1179 265 1209 297
rect 794 249 940 259
rect 794 215 810 249
rect 844 215 940 249
rect 794 205 940 215
rect 910 177 940 205
rect 982 249 1037 265
rect 982 215 993 249
rect 1027 215 1037 249
rect 982 199 1037 215
rect 1079 249 1209 265
rect 1079 215 1089 249
rect 1123 215 1209 249
rect 1079 199 1209 215
rect 1004 177 1034 199
rect 1095 177 1125 199
rect 1179 177 1209 199
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 435 21 465 47
rect 530 21 560 47
rect 627 21 657 47
rect 722 21 752 47
rect 910 21 940 47
rect 1004 21 1034 47
rect 1095 21 1125 47
rect 1179 21 1209 47
<< polycont >>
rect 32 230 66 264
rect 134 230 168 264
rect 304 191 338 225
rect 619 332 653 366
rect 755 323 789 357
rect 517 287 551 321
rect 433 169 467 203
rect 535 164 569 198
rect 810 215 844 249
rect 993 215 1027 249
rect 1089 215 1123 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 391 485 450 527
rect 750 485 818 527
rect 237 443 248 477
rect 203 409 248 443
rect 69 375 156 393
rect 35 359 156 375
rect 18 264 66 325
rect 18 230 32 264
rect 18 197 66 230
rect 122 323 156 359
rect 122 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 287 449 307 483
rect 341 449 357 483
rect 287 415 357 449
rect 287 381 307 415
rect 341 381 357 415
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 122 161 156 214
rect 17 127 156 161
rect 17 119 69 127
rect 17 85 35 119
rect 203 119 237 337
rect 287 333 357 381
rect 425 451 450 485
rect 554 451 570 485
rect 604 451 716 485
rect 391 417 450 451
rect 425 383 450 417
rect 682 417 716 451
rect 750 451 751 485
rect 785 451 818 485
rect 750 435 818 451
rect 856 485 912 527
rect 856 451 864 485
rect 898 451 912 485
rect 856 427 912 451
rect 960 471 994 493
rect 682 400 721 417
rect 683 399 721 400
rect 391 367 450 383
rect 581 391 635 399
rect 684 397 721 399
rect 581 357 585 391
rect 619 382 635 391
rect 619 366 653 382
rect 581 356 619 357
rect 287 299 424 333
rect 288 225 354 265
rect 288 191 304 225
rect 338 191 354 225
rect 390 219 424 299
rect 490 323 551 337
rect 524 321 551 323
rect 490 287 517 289
rect 490 271 551 287
rect 586 332 619 356
rect 586 314 653 332
rect 390 203 467 219
rect 586 208 620 314
rect 687 265 721 397
rect 960 373 994 437
rect 1028 489 1097 527
rect 1028 455 1044 489
rect 1078 455 1097 489
rect 1028 421 1097 455
rect 1028 387 1044 421
rect 1078 387 1097 421
rect 1028 375 1097 387
rect 1131 477 1185 493
rect 1165 443 1185 477
rect 1131 375 1185 443
rect 755 368 994 373
rect 755 357 960 368
rect 789 334 960 357
rect 994 334 1117 341
rect 789 323 1117 334
rect 755 307 1117 323
rect 1083 265 1117 307
rect 1151 300 1185 375
rect 1219 475 1271 527
rect 1253 441 1271 475
rect 1219 384 1271 441
rect 1253 350 1271 384
rect 1219 334 1271 350
rect 1151 285 1271 300
rect 1152 283 1271 285
rect 1153 282 1271 283
rect 1155 277 1271 282
rect 390 169 433 203
rect 390 157 467 169
rect 17 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 303 153 467 157
rect 517 198 620 208
rect 517 164 535 198
rect 569 164 620 198
rect 303 123 424 153
rect 517 147 620 164
rect 654 249 844 265
rect 654 215 810 249
rect 654 199 844 215
rect 896 249 1048 265
rect 896 215 993 249
rect 1027 215 1048 249
rect 896 207 1048 215
rect 1083 249 1123 265
rect 1083 215 1089 249
rect 896 199 963 207
rect 1083 199 1123 215
rect 303 119 341 123
rect 303 85 307 119
rect 654 107 689 199
rect 1083 173 1117 199
rect 1157 178 1271 277
rect 1154 173 1271 178
rect 991 165 1117 173
rect 303 69 341 85
rect 103 17 169 59
rect 375 55 391 89
rect 425 55 441 89
rect 554 73 570 107
rect 604 73 689 107
rect 848 131 866 165
rect 900 139 1117 165
rect 1151 153 1271 173
rect 900 131 1019 139
rect 375 17 441 55
rect 744 72 762 106
rect 796 72 812 106
rect 744 17 812 72
rect 848 97 916 131
rect 848 63 866 97
rect 900 63 916 97
rect 848 51 916 63
rect 1051 89 1085 105
rect 1151 97 1185 153
rect 1051 17 1085 55
rect 1119 89 1185 97
rect 1119 55 1135 89
rect 1169 55 1185 89
rect 1119 51 1185 55
rect 1219 93 1271 119
rect 1253 59 1271 93
rect 1219 17 1271 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 585 357 619 391
rect 490 321 524 323
rect 490 289 517 321
rect 517 289 524 321
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 573 391 631 397
rect 573 388 585 391
rect 248 360 585 388
rect 248 357 260 360
rect 202 351 260 357
rect 573 357 585 360
rect 619 357 631 391
rect 573 351 631 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 478 323 536 329
rect 478 320 490 323
rect 156 292 490 320
rect 156 289 168 292
rect 110 283 168 289
rect 478 289 490 292
rect 524 289 536 323
rect 478 283 536 289
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 954 221 988 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1138 425 1172 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1230 153 1264 187 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1230 221 1264 255 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 47 544 47 544 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 dlrtp_2
rlabel metal1 s 0 -48 1288 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1288 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_END 2798016
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2786822
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
