magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -47 1824 21 1825
rect -47 1716 965 1824
rect -47 1500 1013 1716
rect -47 1384 839 1500
<< pwell >>
rect 207 1128 1089 1254
rect 33 992 1089 1128
rect 207 796 1089 992
rect 33 635 1089 796
rect 27 202 1089 635
<< mvnmos >>
rect 112 1018 212 1102
rect 112 686 212 770
rect 286 228 386 1228
rect 442 228 542 1228
rect 598 228 698 1228
rect 754 228 854 1228
rect 910 228 1010 1228
<< mvpmos >>
rect 72 1450 192 1650
rect 248 1450 368 1650
rect 424 1450 544 1650
rect 600 1450 720 1650
rect 794 1566 894 1650
<< mvndiff >>
rect 233 1158 286 1228
rect 233 1124 241 1158
rect 275 1124 286 1158
rect 233 1102 286 1124
rect 59 1090 112 1102
rect 59 1056 67 1090
rect 101 1056 112 1090
rect 59 1018 112 1056
rect 212 1090 286 1102
rect 212 1056 241 1090
rect 275 1056 286 1090
rect 212 1022 286 1056
rect 212 1018 241 1022
rect 233 988 241 1018
rect 275 988 286 1022
rect 233 954 286 988
rect 233 920 241 954
rect 275 920 286 954
rect 233 886 286 920
rect 233 852 241 886
rect 275 852 286 886
rect 233 818 286 852
rect 233 784 241 818
rect 275 784 286 818
rect 233 770 286 784
rect 59 758 112 770
rect 59 724 67 758
rect 101 724 112 758
rect 59 686 112 724
rect 212 750 286 770
rect 212 716 241 750
rect 275 716 286 750
rect 212 686 286 716
rect 233 682 286 686
rect 233 648 241 682
rect 275 648 286 682
rect 233 614 286 648
rect 233 580 241 614
rect 275 580 286 614
rect 233 546 286 580
rect 233 512 241 546
rect 275 512 286 546
rect 233 478 286 512
rect 233 444 241 478
rect 275 444 286 478
rect 233 410 286 444
rect 233 376 241 410
rect 275 376 286 410
rect 233 342 286 376
rect 233 308 241 342
rect 275 308 286 342
rect 233 274 286 308
rect 233 240 241 274
rect 275 240 286 274
rect 233 228 286 240
rect 386 1158 442 1228
rect 386 1124 397 1158
rect 431 1124 442 1158
rect 386 1090 442 1124
rect 386 1056 397 1090
rect 431 1056 442 1090
rect 386 1022 442 1056
rect 386 988 397 1022
rect 431 988 442 1022
rect 386 954 442 988
rect 386 920 397 954
rect 431 920 442 954
rect 386 886 442 920
rect 386 852 397 886
rect 431 852 442 886
rect 386 818 442 852
rect 386 784 397 818
rect 431 784 442 818
rect 386 750 442 784
rect 386 716 397 750
rect 431 716 442 750
rect 386 682 442 716
rect 386 648 397 682
rect 431 648 442 682
rect 386 614 442 648
rect 386 580 397 614
rect 431 580 442 614
rect 386 546 442 580
rect 386 512 397 546
rect 431 512 442 546
rect 386 478 442 512
rect 386 444 397 478
rect 431 444 442 478
rect 386 410 442 444
rect 386 376 397 410
rect 431 376 442 410
rect 386 342 442 376
rect 386 308 397 342
rect 431 308 442 342
rect 386 274 442 308
rect 386 240 397 274
rect 431 240 442 274
rect 386 228 442 240
rect 542 1158 598 1228
rect 542 1124 553 1158
rect 587 1124 598 1158
rect 542 1090 598 1124
rect 542 1056 553 1090
rect 587 1056 598 1090
rect 542 1022 598 1056
rect 542 988 553 1022
rect 587 988 598 1022
rect 542 954 598 988
rect 542 920 553 954
rect 587 920 598 954
rect 542 886 598 920
rect 542 852 553 886
rect 587 852 598 886
rect 542 818 598 852
rect 542 784 553 818
rect 587 784 598 818
rect 542 750 598 784
rect 542 716 553 750
rect 587 716 598 750
rect 542 682 598 716
rect 542 648 553 682
rect 587 648 598 682
rect 542 614 598 648
rect 542 580 553 614
rect 587 580 598 614
rect 542 546 598 580
rect 542 512 553 546
rect 587 512 598 546
rect 542 478 598 512
rect 542 444 553 478
rect 587 444 598 478
rect 542 410 598 444
rect 542 376 553 410
rect 587 376 598 410
rect 542 342 598 376
rect 542 308 553 342
rect 587 308 598 342
rect 542 274 598 308
rect 542 240 553 274
rect 587 240 598 274
rect 542 228 598 240
rect 698 1158 754 1228
rect 698 1124 709 1158
rect 743 1124 754 1158
rect 698 1090 754 1124
rect 698 1056 709 1090
rect 743 1056 754 1090
rect 698 1022 754 1056
rect 698 988 709 1022
rect 743 988 754 1022
rect 698 954 754 988
rect 698 920 709 954
rect 743 920 754 954
rect 698 886 754 920
rect 698 852 709 886
rect 743 852 754 886
rect 698 818 754 852
rect 698 784 709 818
rect 743 784 754 818
rect 698 750 754 784
rect 698 716 709 750
rect 743 716 754 750
rect 698 682 754 716
rect 698 648 709 682
rect 743 648 754 682
rect 698 614 754 648
rect 698 580 709 614
rect 743 580 754 614
rect 698 546 754 580
rect 698 512 709 546
rect 743 512 754 546
rect 698 478 754 512
rect 698 444 709 478
rect 743 444 754 478
rect 698 410 754 444
rect 698 376 709 410
rect 743 376 754 410
rect 698 342 754 376
rect 698 308 709 342
rect 743 308 754 342
rect 698 274 754 308
rect 698 240 709 274
rect 743 240 754 274
rect 698 228 754 240
rect 854 1158 910 1228
rect 854 1124 865 1158
rect 899 1124 910 1158
rect 854 1090 910 1124
rect 854 1056 865 1090
rect 899 1056 910 1090
rect 854 1022 910 1056
rect 854 988 865 1022
rect 899 988 910 1022
rect 854 954 910 988
rect 854 920 865 954
rect 899 920 910 954
rect 854 886 910 920
rect 854 852 865 886
rect 899 852 910 886
rect 854 818 910 852
rect 854 784 865 818
rect 899 784 910 818
rect 854 750 910 784
rect 854 716 865 750
rect 899 716 910 750
rect 854 682 910 716
rect 854 648 865 682
rect 899 648 910 682
rect 854 614 910 648
rect 854 580 865 614
rect 899 580 910 614
rect 854 546 910 580
rect 854 512 865 546
rect 899 512 910 546
rect 854 478 910 512
rect 854 444 865 478
rect 899 444 910 478
rect 854 410 910 444
rect 854 376 865 410
rect 899 376 910 410
rect 854 342 910 376
rect 854 308 865 342
rect 899 308 910 342
rect 854 274 910 308
rect 854 240 865 274
rect 899 240 910 274
rect 854 228 910 240
rect 1010 1158 1063 1228
rect 1010 1124 1021 1158
rect 1055 1124 1063 1158
rect 1010 1090 1063 1124
rect 1010 1056 1021 1090
rect 1055 1056 1063 1090
rect 1010 1022 1063 1056
rect 1010 988 1021 1022
rect 1055 988 1063 1022
rect 1010 954 1063 988
rect 1010 920 1021 954
rect 1055 920 1063 954
rect 1010 886 1063 920
rect 1010 852 1021 886
rect 1055 852 1063 886
rect 1010 818 1063 852
rect 1010 784 1021 818
rect 1055 784 1063 818
rect 1010 750 1063 784
rect 1010 716 1021 750
rect 1055 716 1063 750
rect 1010 682 1063 716
rect 1010 648 1021 682
rect 1055 648 1063 682
rect 1010 614 1063 648
rect 1010 580 1021 614
rect 1055 580 1063 614
rect 1010 546 1063 580
rect 1010 512 1021 546
rect 1055 512 1063 546
rect 1010 478 1063 512
rect 1010 444 1021 478
rect 1055 444 1063 478
rect 1010 410 1063 444
rect 1010 376 1021 410
rect 1055 376 1063 410
rect 1010 342 1063 376
rect 1010 308 1021 342
rect 1055 308 1063 342
rect 1010 274 1063 308
rect 1010 240 1021 274
rect 1055 240 1063 274
rect 1010 228 1063 240
<< mvpdiff >>
rect 19 1638 72 1650
rect 19 1604 27 1638
rect 61 1604 72 1638
rect 19 1570 72 1604
rect 19 1536 27 1570
rect 61 1536 72 1570
rect 19 1502 72 1536
rect 19 1468 27 1502
rect 61 1468 72 1502
rect 19 1450 72 1468
rect 192 1638 248 1650
rect 192 1604 203 1638
rect 237 1604 248 1638
rect 192 1570 248 1604
rect 192 1536 203 1570
rect 237 1536 248 1570
rect 192 1502 248 1536
rect 192 1468 203 1502
rect 237 1468 248 1502
rect 192 1450 248 1468
rect 368 1638 424 1650
rect 368 1604 379 1638
rect 413 1604 424 1638
rect 368 1570 424 1604
rect 368 1536 379 1570
rect 413 1536 424 1570
rect 368 1502 424 1536
rect 368 1468 379 1502
rect 413 1468 424 1502
rect 368 1450 424 1468
rect 544 1638 600 1650
rect 544 1604 555 1638
rect 589 1604 600 1638
rect 544 1570 600 1604
rect 544 1536 555 1570
rect 589 1536 600 1570
rect 544 1502 600 1536
rect 544 1468 555 1502
rect 589 1468 600 1502
rect 544 1450 600 1468
rect 720 1638 794 1650
rect 720 1604 731 1638
rect 765 1604 794 1638
rect 720 1570 794 1604
rect 720 1536 731 1570
rect 765 1566 794 1570
rect 894 1638 947 1650
rect 894 1604 905 1638
rect 939 1604 947 1638
rect 894 1566 947 1604
rect 765 1536 773 1566
rect 720 1502 773 1536
rect 720 1468 731 1502
rect 765 1468 773 1502
rect 720 1450 773 1468
<< mvndiffc >>
rect 241 1124 275 1158
rect 67 1056 101 1090
rect 241 1056 275 1090
rect 241 988 275 1022
rect 241 920 275 954
rect 241 852 275 886
rect 241 784 275 818
rect 67 724 101 758
rect 241 716 275 750
rect 241 648 275 682
rect 241 580 275 614
rect 241 512 275 546
rect 241 444 275 478
rect 241 376 275 410
rect 241 308 275 342
rect 241 240 275 274
rect 397 1124 431 1158
rect 397 1056 431 1090
rect 397 988 431 1022
rect 397 920 431 954
rect 397 852 431 886
rect 397 784 431 818
rect 397 716 431 750
rect 397 648 431 682
rect 397 580 431 614
rect 397 512 431 546
rect 397 444 431 478
rect 397 376 431 410
rect 397 308 431 342
rect 397 240 431 274
rect 553 1124 587 1158
rect 553 1056 587 1090
rect 553 988 587 1022
rect 553 920 587 954
rect 553 852 587 886
rect 553 784 587 818
rect 553 716 587 750
rect 553 648 587 682
rect 553 580 587 614
rect 553 512 587 546
rect 553 444 587 478
rect 553 376 587 410
rect 553 308 587 342
rect 553 240 587 274
rect 709 1124 743 1158
rect 709 1056 743 1090
rect 709 988 743 1022
rect 709 920 743 954
rect 709 852 743 886
rect 709 784 743 818
rect 709 716 743 750
rect 709 648 743 682
rect 709 580 743 614
rect 709 512 743 546
rect 709 444 743 478
rect 709 376 743 410
rect 709 308 743 342
rect 709 240 743 274
rect 865 1124 899 1158
rect 865 1056 899 1090
rect 865 988 899 1022
rect 865 920 899 954
rect 865 852 899 886
rect 865 784 899 818
rect 865 716 899 750
rect 865 648 899 682
rect 865 580 899 614
rect 865 512 899 546
rect 865 444 899 478
rect 865 376 899 410
rect 865 308 899 342
rect 865 240 899 274
rect 1021 1124 1055 1158
rect 1021 1056 1055 1090
rect 1021 988 1055 1022
rect 1021 920 1055 954
rect 1021 852 1055 886
rect 1021 784 1055 818
rect 1021 716 1055 750
rect 1021 648 1055 682
rect 1021 580 1055 614
rect 1021 512 1055 546
rect 1021 444 1055 478
rect 1021 376 1055 410
rect 1021 308 1055 342
rect 1021 240 1055 274
<< mvpdiffc >>
rect 27 1604 61 1638
rect 27 1536 61 1570
rect 27 1468 61 1502
rect 203 1604 237 1638
rect 203 1536 237 1570
rect 203 1468 237 1502
rect 379 1604 413 1638
rect 379 1536 413 1570
rect 379 1468 413 1502
rect 555 1604 589 1638
rect 555 1536 589 1570
rect 555 1468 589 1502
rect 731 1604 765 1638
rect 731 1536 765 1570
rect 905 1604 939 1638
rect 731 1468 765 1502
<< psubdiff >>
rect 53 585 155 609
rect 87 551 121 585
rect 53 486 155 551
rect 87 452 121 486
rect 53 386 155 452
rect 87 352 121 386
rect 53 286 155 352
rect 87 252 121 286
rect 53 228 155 252
<< mvnsubdiff >>
rect 87 1724 111 1758
rect 145 1724 184 1758
rect 218 1724 257 1758
rect 291 1724 330 1758
rect 364 1724 403 1758
rect 437 1724 476 1758
rect 510 1724 549 1758
rect 583 1724 622 1758
rect 656 1724 695 1758
rect 729 1724 768 1758
rect 802 1724 841 1758
rect 875 1724 899 1758
<< psubdiffcont >>
rect 53 551 87 585
rect 121 551 155 585
rect 53 452 87 486
rect 121 452 155 486
rect 53 352 87 386
rect 121 352 155 386
rect 53 252 87 286
rect 121 252 155 286
<< mvnsubdiffcont >>
rect 111 1724 145 1758
rect 184 1724 218 1758
rect 257 1724 291 1758
rect 330 1724 364 1758
rect 403 1724 437 1758
rect 476 1724 510 1758
rect 549 1724 583 1758
rect 622 1724 656 1758
rect 695 1724 729 1758
rect 768 1724 802 1758
rect 841 1724 875 1758
<< poly >>
rect 72 1650 192 1682
rect 248 1650 368 1682
rect 424 1650 544 1682
rect 600 1650 720 1682
rect 794 1650 894 1682
rect 794 1517 894 1566
rect 794 1483 836 1517
rect 870 1483 894 1517
rect 72 1418 192 1450
rect 248 1418 368 1450
rect 112 1402 368 1418
rect 112 1368 128 1402
rect 162 1368 223 1402
rect 257 1368 318 1402
rect 352 1368 368 1402
rect 112 1352 368 1368
rect 424 1418 544 1450
rect 600 1418 720 1450
rect 424 1402 720 1418
rect 424 1368 440 1402
rect 474 1368 516 1402
rect 550 1368 593 1402
rect 627 1368 670 1402
rect 704 1368 720 1402
rect 794 1449 894 1483
rect 794 1415 836 1449
rect 870 1415 894 1449
rect 794 1399 894 1415
rect 424 1352 720 1368
rect 112 1271 212 1288
rect 112 1237 145 1271
rect 179 1237 212 1271
rect 112 1203 212 1237
rect 286 1228 386 1260
rect 442 1228 542 1260
rect 598 1228 698 1260
rect 754 1228 854 1260
rect 910 1228 1010 1260
rect 112 1169 145 1203
rect 179 1169 212 1203
rect 112 1102 212 1169
rect 112 986 212 1018
rect 112 928 212 944
rect 112 894 150 928
rect 184 894 212 928
rect 112 860 212 894
rect 112 826 150 860
rect 184 826 212 860
rect 112 770 212 826
rect 112 654 212 686
rect 286 158 386 228
rect 286 124 319 158
rect 353 124 386 158
rect 286 90 386 124
rect 286 56 319 90
rect 353 56 386 90
rect 286 40 386 56
rect 442 158 542 228
rect 442 124 479 158
rect 513 124 542 158
rect 442 90 542 124
rect 442 56 479 90
rect 513 56 542 90
rect 442 40 542 56
rect 598 158 698 228
rect 598 124 635 158
rect 669 124 698 158
rect 598 90 698 124
rect 598 56 635 90
rect 669 56 698 90
rect 598 40 698 56
rect 754 158 854 228
rect 754 124 785 158
rect 819 124 854 158
rect 754 90 854 124
rect 754 56 785 90
rect 819 56 854 90
rect 754 40 854 56
rect 910 156 1010 228
rect 910 122 940 156
rect 974 122 1010 156
rect 910 88 1010 122
rect 910 54 940 88
rect 974 54 1010 88
rect 910 38 1010 54
<< polycont >>
rect 836 1483 870 1517
rect 128 1368 162 1402
rect 223 1368 257 1402
rect 318 1368 352 1402
rect 440 1368 474 1402
rect 516 1368 550 1402
rect 593 1368 627 1402
rect 670 1368 704 1402
rect 836 1415 870 1449
rect 145 1237 179 1271
rect 145 1169 179 1203
rect 150 894 184 928
rect 150 826 184 860
rect 319 124 353 158
rect 319 56 353 90
rect 479 124 513 158
rect 479 56 513 90
rect 635 124 669 158
rect 635 56 669 90
rect 785 124 819 158
rect 785 56 819 90
rect 940 122 974 156
rect 940 54 974 88
<< locali >>
rect 87 1724 111 1758
rect 145 1724 146 1758
rect 180 1724 184 1758
rect 218 1724 222 1758
rect 256 1724 257 1758
rect 291 1724 298 1758
rect 364 1724 374 1758
rect 437 1724 450 1758
rect 510 1724 526 1758
rect 583 1724 602 1758
rect 656 1724 678 1758
rect 729 1724 754 1758
rect 802 1724 831 1758
rect 875 1724 899 1758
rect 27 1582 61 1604
rect 27 1510 61 1536
rect 27 1452 61 1468
rect 203 1582 237 1604
rect 203 1510 237 1536
rect 203 1452 237 1468
rect 379 1582 413 1604
rect 379 1510 413 1536
rect 379 1452 413 1468
rect 555 1582 589 1604
rect 555 1510 589 1536
rect 555 1452 589 1468
rect 731 1582 765 1604
rect 905 1582 939 1604
rect 731 1510 765 1536
rect 731 1452 765 1468
rect 816 1522 831 1556
rect 865 1522 870 1556
rect 816 1517 870 1522
rect 816 1484 836 1517
rect 816 1450 831 1484
rect 870 1483 939 1514
rect 865 1450 939 1483
rect 816 1449 939 1450
rect 816 1415 836 1449
rect 870 1415 939 1449
rect 112 1368 128 1402
rect 162 1368 223 1402
rect 257 1368 318 1402
rect 352 1368 368 1402
rect 424 1368 440 1402
rect 474 1368 516 1402
rect 550 1368 593 1402
rect 627 1368 670 1402
rect 704 1400 720 1402
rect 704 1368 722 1400
rect 153 1299 191 1333
rect 119 1271 225 1299
rect 119 1237 145 1271
rect 179 1237 225 1271
rect 119 1205 225 1237
rect 119 1203 203 1205
rect 119 1169 145 1203
rect 179 1169 203 1203
rect 309 1181 363 1368
rect 424 1356 722 1368
rect 424 1322 478 1356
rect 512 1322 568 1356
rect 602 1322 658 1356
rect 692 1322 722 1356
rect 424 1316 722 1322
rect 816 1282 939 1415
rect 732 1248 770 1282
rect 804 1248 939 1282
rect 698 1229 939 1248
rect 119 1153 203 1169
rect 241 1158 275 1174
rect 61 1090 166 1106
rect 61 1056 67 1090
rect 101 1072 166 1090
rect 101 1056 200 1072
rect 61 1032 200 1056
rect 61 998 166 1032
rect 61 959 200 998
rect 61 928 166 959
rect 61 894 150 928
rect 184 894 200 925
rect 61 886 200 894
rect 61 883 166 886
rect 138 860 166 883
rect 138 826 150 860
rect 184 826 200 852
rect 138 800 200 826
rect 241 1092 275 1124
rect 309 1147 320 1181
rect 354 1147 363 1181
rect 309 1109 363 1147
rect 309 1075 320 1109
rect 354 1075 363 1109
rect 309 1074 363 1075
rect 397 1158 431 1160
rect 397 1122 431 1124
rect 241 1022 275 1056
rect 241 954 275 985
rect 241 886 275 912
rect 241 818 275 839
rect 67 758 101 771
rect 241 750 275 766
rect 241 682 275 693
rect 241 614 275 620
rect 64 585 142 612
rect 30 551 53 578
rect 87 551 121 585
rect 155 551 176 578
rect 30 523 176 551
rect 64 489 142 523
rect 30 486 176 489
rect 30 452 53 486
rect 87 452 121 486
rect 155 452 176 486
rect 30 434 176 452
rect 64 400 142 434
rect 30 386 176 400
rect 30 352 53 386
rect 87 352 121 386
rect 155 352 176 386
rect 30 346 176 352
rect 64 312 142 346
rect 30 286 176 312
rect 30 258 53 286
rect 87 252 121 286
rect 155 258 176 286
rect 64 224 142 252
rect 241 506 275 512
rect 241 432 275 444
rect 241 358 275 376
rect 241 284 275 308
rect 241 224 275 240
rect 397 1050 431 1056
rect 397 978 431 988
rect 397 906 431 920
rect 397 834 431 852
rect 397 762 431 784
rect 397 690 431 716
rect 397 618 431 648
rect 397 546 431 580
rect 397 478 431 512
rect 397 410 431 440
rect 397 342 431 368
rect 397 274 431 296
rect 553 1158 587 1160
rect 553 1122 587 1124
rect 553 1050 587 1056
rect 553 978 587 988
rect 553 906 587 920
rect 553 834 587 852
rect 553 762 587 784
rect 553 690 587 716
rect 553 618 587 648
rect 553 546 587 580
rect 553 478 587 512
rect 553 410 587 440
rect 553 342 587 368
rect 553 274 587 296
rect 709 1158 743 1160
rect 709 1122 743 1124
rect 709 1050 743 1056
rect 709 978 743 988
rect 709 906 743 920
rect 709 834 743 852
rect 709 762 743 784
rect 709 690 743 716
rect 709 618 743 648
rect 709 546 743 580
rect 709 478 743 512
rect 709 410 743 440
rect 709 342 743 368
rect 709 274 743 296
rect 865 1158 899 1160
rect 865 1122 899 1124
rect 865 1050 899 1056
rect 865 978 899 988
rect 865 906 899 920
rect 865 834 899 852
rect 865 762 899 784
rect 865 690 899 716
rect 865 618 899 648
rect 865 546 899 580
rect 865 478 899 512
rect 865 410 899 440
rect 865 342 899 368
rect 865 274 899 296
rect 1021 1158 1055 1160
rect 1021 1122 1055 1124
rect 1021 1050 1055 1056
rect 1021 978 1055 988
rect 1021 906 1055 920
rect 1021 834 1055 852
rect 1021 762 1055 784
rect 1021 690 1055 716
rect 1021 618 1055 648
rect 1021 546 1055 580
rect 1021 478 1055 512
rect 1021 410 1055 440
rect 1021 342 1055 368
rect 1021 274 1055 296
rect 319 158 320 174
rect 353 124 354 147
rect 319 109 354 124
rect 319 90 320 109
rect 479 158 513 174
rect 479 90 513 124
rect 319 40 353 56
rect 479 40 513 56
rect 635 158 669 174
rect 635 90 669 124
rect 635 40 669 56
rect 785 158 819 174
rect 785 90 819 124
rect 785 40 819 56
rect 940 156 974 172
rect 940 88 974 122
rect 940 38 974 54
<< viali >>
rect 146 1724 180 1758
rect 222 1724 256 1758
rect 298 1724 330 1758
rect 330 1724 332 1758
rect 374 1724 403 1758
rect 403 1724 408 1758
rect 450 1724 476 1758
rect 476 1724 484 1758
rect 526 1724 549 1758
rect 549 1724 560 1758
rect 602 1724 622 1758
rect 622 1724 636 1758
rect 678 1724 695 1758
rect 695 1724 712 1758
rect 754 1724 768 1758
rect 768 1724 788 1758
rect 831 1724 841 1758
rect 841 1724 865 1758
rect 27 1638 61 1654
rect 27 1620 61 1638
rect 27 1570 61 1582
rect 27 1548 61 1570
rect 27 1502 61 1510
rect 27 1476 61 1502
rect 203 1638 237 1654
rect 203 1620 237 1638
rect 203 1570 237 1582
rect 203 1548 237 1570
rect 203 1502 237 1510
rect 203 1476 237 1502
rect 379 1638 413 1654
rect 379 1620 413 1638
rect 379 1570 413 1582
rect 379 1548 413 1570
rect 379 1502 413 1510
rect 379 1476 413 1502
rect 555 1638 589 1654
rect 555 1620 589 1638
rect 555 1570 589 1582
rect 555 1548 589 1570
rect 555 1502 589 1510
rect 555 1476 589 1502
rect 731 1638 765 1654
rect 731 1620 765 1638
rect 731 1570 765 1582
rect 731 1548 765 1570
rect 905 1638 939 1654
rect 905 1620 939 1638
rect 731 1502 765 1510
rect 731 1476 765 1502
rect 831 1522 865 1556
rect 905 1548 939 1582
rect 831 1483 836 1484
rect 836 1483 865 1484
rect 831 1450 865 1483
rect 119 1299 153 1333
rect 191 1299 225 1333
rect 478 1322 512 1356
rect 568 1322 602 1356
rect 658 1322 692 1356
rect 698 1248 732 1282
rect 770 1248 804 1282
rect 166 1072 200 1106
rect 166 998 200 1032
rect 166 928 200 959
rect 166 925 184 928
rect 184 925 200 928
rect 166 860 200 886
rect 166 852 184 860
rect 184 852 200 860
rect 67 771 101 805
rect 241 1090 275 1092
rect 241 1058 275 1090
rect 320 1147 354 1181
rect 320 1075 354 1109
rect 397 1160 431 1194
rect 397 1090 431 1122
rect 397 1088 431 1090
rect 241 988 275 1019
rect 241 985 275 988
rect 241 920 275 946
rect 241 912 275 920
rect 241 852 275 873
rect 241 839 275 852
rect 67 724 101 733
rect 67 699 101 724
rect 241 784 275 800
rect 241 766 275 784
rect 241 716 275 727
rect 241 693 275 716
rect 241 648 275 654
rect 241 620 275 648
rect 30 585 64 612
rect 142 585 176 612
rect 30 578 53 585
rect 53 578 64 585
rect 142 578 155 585
rect 155 578 176 585
rect 30 489 64 523
rect 142 489 176 523
rect 30 400 64 434
rect 142 400 176 434
rect 30 312 64 346
rect 142 312 176 346
rect 30 252 53 258
rect 53 252 64 258
rect 142 252 155 258
rect 155 252 176 258
rect 30 224 64 252
rect 142 224 176 252
rect 241 546 275 580
rect 241 478 275 506
rect 241 472 275 478
rect 241 410 275 432
rect 241 398 275 410
rect 241 342 275 358
rect 241 324 275 342
rect 241 274 275 284
rect 241 250 275 274
rect 397 1022 431 1050
rect 397 1016 431 1022
rect 397 954 431 978
rect 397 944 431 954
rect 397 886 431 906
rect 397 872 431 886
rect 397 818 431 834
rect 397 800 431 818
rect 397 750 431 762
rect 397 728 431 750
rect 397 682 431 690
rect 397 656 431 682
rect 397 614 431 618
rect 397 584 431 614
rect 397 512 431 546
rect 397 444 431 474
rect 397 440 431 444
rect 397 376 431 402
rect 397 368 431 376
rect 397 308 431 330
rect 397 296 431 308
rect 397 240 431 258
rect 397 224 431 240
rect 553 1160 587 1194
rect 553 1090 587 1122
rect 553 1088 587 1090
rect 553 1022 587 1050
rect 553 1016 587 1022
rect 553 954 587 978
rect 553 944 587 954
rect 553 886 587 906
rect 553 872 587 886
rect 553 818 587 834
rect 553 800 587 818
rect 553 750 587 762
rect 553 728 587 750
rect 553 682 587 690
rect 553 656 587 682
rect 553 614 587 618
rect 553 584 587 614
rect 553 512 587 546
rect 553 444 587 474
rect 553 440 587 444
rect 553 376 587 402
rect 553 368 587 376
rect 553 308 587 330
rect 553 296 587 308
rect 553 240 587 258
rect 553 224 587 240
rect 709 1160 743 1194
rect 709 1090 743 1122
rect 709 1088 743 1090
rect 709 1022 743 1050
rect 709 1016 743 1022
rect 709 954 743 978
rect 709 944 743 954
rect 709 886 743 906
rect 709 872 743 886
rect 709 818 743 834
rect 709 800 743 818
rect 709 750 743 762
rect 709 728 743 750
rect 709 682 743 690
rect 709 656 743 682
rect 709 614 743 618
rect 709 584 743 614
rect 709 512 743 546
rect 709 444 743 474
rect 709 440 743 444
rect 709 376 743 402
rect 709 368 743 376
rect 709 308 743 330
rect 709 296 743 308
rect 709 240 743 258
rect 709 224 743 240
rect 865 1160 899 1194
rect 865 1090 899 1122
rect 865 1088 899 1090
rect 865 1022 899 1050
rect 865 1016 899 1022
rect 865 954 899 978
rect 865 944 899 954
rect 865 886 899 906
rect 865 872 899 886
rect 865 818 899 834
rect 865 800 899 818
rect 865 750 899 762
rect 865 728 899 750
rect 865 682 899 690
rect 865 656 899 682
rect 865 614 899 618
rect 865 584 899 614
rect 865 512 899 546
rect 865 444 899 474
rect 865 440 899 444
rect 865 376 899 402
rect 865 368 899 376
rect 865 308 899 330
rect 865 296 899 308
rect 865 240 899 258
rect 865 224 899 240
rect 1021 1160 1055 1194
rect 1021 1090 1055 1122
rect 1021 1088 1055 1090
rect 1021 1022 1055 1050
rect 1021 1016 1055 1022
rect 1021 954 1055 978
rect 1021 944 1055 954
rect 1021 886 1055 906
rect 1021 872 1055 886
rect 1021 818 1055 834
rect 1021 800 1055 818
rect 1021 750 1055 762
rect 1021 728 1055 750
rect 1021 682 1055 690
rect 1021 656 1055 682
rect 1021 614 1055 618
rect 1021 584 1055 614
rect 1021 512 1055 546
rect 1021 444 1055 474
rect 1021 440 1055 444
rect 1021 376 1055 402
rect 1021 368 1055 376
rect 1021 308 1055 330
rect 1021 296 1055 308
rect 1021 240 1055 258
rect 1021 224 1055 240
rect 320 158 354 181
rect 320 147 353 158
rect 353 147 354 158
rect 320 90 354 109
rect 320 75 353 90
rect 353 75 354 90
<< metal1 >>
rect 21 1758 1014 1846
rect 21 1724 146 1758
rect 180 1724 222 1758
rect 256 1724 298 1758
rect 332 1724 374 1758
rect 408 1724 450 1758
rect 484 1724 526 1758
rect 560 1724 602 1758
rect 636 1724 678 1758
rect 712 1724 754 1758
rect 788 1724 831 1758
rect 865 1724 1014 1758
rect 21 1718 1014 1724
rect 21 1654 67 1718
tri 67 1685 100 1718 nw
tri 339 1685 372 1718 ne
rect 372 1685 420 1718
tri 420 1685 453 1718 nw
tri 691 1685 724 1718 ne
rect 724 1685 771 1718
tri 372 1684 373 1685 ne
rect 21 1620 27 1654
rect 61 1620 67 1654
rect 21 1582 67 1620
rect 21 1548 27 1582
rect 61 1548 67 1582
rect 21 1510 67 1548
rect 21 1476 27 1510
rect 61 1476 67 1510
rect 21 1464 67 1476
rect 197 1654 243 1666
rect 197 1620 203 1654
rect 237 1620 243 1654
rect 197 1582 243 1620
rect 197 1548 203 1582
rect 237 1548 243 1582
rect 197 1510 243 1548
rect 197 1476 203 1510
rect 237 1476 243 1510
tri 151 1362 197 1408 se
rect 197 1391 243 1476
rect 373 1654 419 1685
tri 419 1684 420 1685 nw
tri 724 1684 725 1685 ne
rect 373 1620 379 1654
rect 413 1620 419 1654
rect 373 1582 419 1620
rect 373 1548 379 1582
rect 413 1548 419 1582
rect 373 1510 419 1548
rect 373 1476 379 1510
rect 413 1476 419 1510
rect 373 1464 419 1476
rect 549 1654 595 1666
rect 549 1620 555 1654
rect 589 1620 595 1654
rect 549 1582 595 1620
rect 549 1548 555 1582
rect 589 1548 595 1582
rect 549 1510 595 1548
rect 549 1476 555 1510
rect 589 1476 595 1510
rect 549 1464 595 1476
rect 725 1654 771 1685
tri 771 1684 805 1718 nw
rect 725 1620 731 1654
rect 765 1620 771 1654
rect 725 1582 771 1620
rect 725 1548 731 1582
rect 765 1548 771 1582
rect 899 1654 945 1666
rect 899 1620 905 1654
rect 939 1620 945 1654
rect 899 1582 945 1620
rect 725 1510 771 1548
rect 725 1476 731 1510
rect 765 1476 771 1510
tri 595 1464 598 1467 sw
rect 725 1464 771 1476
rect 825 1556 871 1568
rect 825 1522 831 1556
rect 865 1522 871 1556
rect 825 1484 871 1522
tri 817 1464 825 1472 se
rect 825 1464 831 1484
rect 549 1450 598 1464
tri 598 1450 612 1464 sw
tri 803 1450 817 1464 se
rect 817 1450 831 1464
rect 865 1450 871 1484
rect 549 1438 612 1450
tri 612 1438 624 1450 sw
tri 791 1438 803 1450 se
rect 803 1438 871 1450
rect 549 1436 624 1438
tri 624 1436 626 1438 sw
tri 789 1436 791 1438 se
rect 791 1436 858 1438
rect 549 1425 858 1436
tri 858 1425 871 1438 nw
rect 899 1548 905 1582
rect 939 1548 945 1582
tri 549 1415 559 1425 ne
rect 559 1415 824 1425
tri 243 1391 267 1415 sw
tri 559 1391 583 1415 ne
rect 583 1391 824 1415
tri 824 1391 858 1425 nw
tri 890 1391 899 1400 se
rect 899 1391 945 1548
tri 945 1391 976 1422 sw
rect 197 1367 267 1391
tri 267 1367 291 1391 sw
tri 866 1367 890 1391 se
rect 890 1367 976 1391
tri 976 1367 1000 1391 sw
rect 197 1362 291 1367
tri 291 1362 296 1367 sw
tri 861 1362 866 1367 se
rect 866 1362 1000 1367
tri 1000 1362 1005 1367 sw
rect 107 1356 1005 1362
tri 100 1339 107 1346 se
rect 107 1339 478 1356
tri 94 1333 100 1339 se
rect 100 1333 478 1339
tri 61 1300 94 1333 se
rect 94 1300 119 1333
rect 61 1299 119 1300
rect 153 1299 191 1333
rect 225 1322 478 1333
rect 512 1322 568 1356
rect 602 1322 658 1356
rect 692 1322 1005 1356
rect 225 1316 1005 1322
tri 1005 1316 1051 1362 sw
rect 225 1306 250 1316
tri 250 1306 260 1316 nw
tri 990 1306 1000 1316 ne
rect 1000 1306 1051 1316
tri 1051 1306 1061 1316 sw
rect 225 1299 237 1306
rect 61 1293 237 1299
tri 237 1293 250 1306 nw
tri 1000 1293 1013 1306 ne
rect 1013 1293 1061 1306
rect 61 1288 147 1293
tri 147 1288 152 1293 nw
tri 1013 1291 1015 1293 ne
rect 61 1282 141 1288
tri 141 1282 147 1288 nw
tri 299 1282 305 1288 se
rect 305 1282 816 1288
rect 61 1243 107 1282
tri 107 1248 141 1282 nw
tri 265 1248 299 1282 se
rect 299 1248 698 1282
rect 732 1248 770 1282
rect 804 1248 816 1282
tri 260 1243 265 1248 se
rect 265 1243 816 1248
tri 246 1229 260 1243 se
rect 260 1242 816 1243
rect 260 1229 305 1242
tri 305 1229 318 1242 nw
tri 211 1194 246 1229 se
rect 246 1194 270 1229
tri 270 1194 305 1229 nw
rect 391 1194 437 1206
tri 210 1193 211 1194 se
rect 211 1193 269 1194
tri 269 1193 270 1194 nw
tri 198 1181 210 1193 se
rect 210 1181 257 1193
tri 257 1181 269 1193 nw
rect 309 1181 363 1193
tri 187 1170 198 1181 se
rect 198 1170 246 1181
tri 246 1170 257 1181 nw
tri 164 1147 187 1170 se
rect 187 1147 223 1170
tri 223 1147 246 1170 nw
rect 309 1147 320 1181
rect 354 1147 363 1181
tri 160 1143 164 1147 se
rect 164 1143 219 1147
tri 219 1143 223 1147 nw
rect 160 1106 206 1143
tri 206 1130 219 1143 nw
rect 160 1072 166 1106
rect 200 1072 206 1106
rect 309 1109 363 1147
rect 160 1032 206 1072
rect 160 998 166 1032
rect 200 998 206 1032
rect 160 959 206 998
rect 160 925 166 959
rect 200 925 206 959
rect 160 886 206 925
rect 160 852 166 886
rect 200 852 206 886
rect 160 840 206 852
rect 235 1092 281 1104
rect 235 1058 241 1092
rect 275 1058 281 1092
rect 235 1019 281 1058
rect 235 985 241 1019
rect 275 985 281 1019
rect 235 946 281 985
rect 235 912 241 946
rect 275 912 281 946
rect 235 873 281 912
rect 235 839 241 873
rect 275 839 281 873
rect 61 805 107 817
rect 61 771 67 805
rect 101 771 107 805
rect 61 733 107 771
rect 61 699 67 733
rect 101 699 107 733
tri 57 656 61 660 se
rect 61 656 107 699
rect 235 800 281 839
rect 235 766 241 800
rect 275 766 281 800
rect 235 727 281 766
rect 235 693 241 727
rect 275 693 281 727
tri 107 656 111 660 sw
tri 55 654 57 656 se
rect 57 654 111 656
tri 111 654 113 656 sw
rect 235 654 281 693
tri 25 624 55 654 se
rect 55 624 113 654
tri 113 624 143 654 sw
rect 235 624 241 654
rect 24 620 241 624
rect 275 620 281 654
rect 24 612 281 620
rect 24 578 30 612
rect 64 578 142 612
rect 176 580 281 612
rect 176 578 241 580
rect 24 546 241 578
rect 275 546 281 580
rect 24 523 281 546
rect 24 489 30 523
rect 64 489 142 523
rect 176 506 281 523
rect 176 489 241 506
rect 24 472 241 489
rect 275 472 281 506
rect 24 434 281 472
rect 24 400 30 434
rect 64 400 142 434
rect 176 432 281 434
rect 176 400 241 432
rect 24 398 241 400
rect 275 398 281 432
rect 24 358 281 398
rect 24 346 241 358
rect 24 312 30 346
rect 64 312 142 346
rect 176 324 241 346
rect 275 324 281 358
rect 176 312 281 324
rect 24 284 281 312
rect 24 258 241 284
rect 24 224 30 258
rect 64 224 142 258
rect 176 250 241 258
rect 275 250 281 284
rect 176 224 281 250
rect 24 212 281 224
rect 309 1075 320 1109
rect 354 1075 363 1109
rect 309 181 363 1075
rect 391 1160 397 1194
rect 431 1160 437 1194
rect 391 1122 437 1160
rect 391 1088 397 1122
rect 431 1088 437 1122
rect 391 1050 437 1088
rect 391 1016 397 1050
rect 431 1016 437 1050
rect 391 978 437 1016
rect 391 944 397 978
rect 431 944 437 978
rect 391 906 437 944
rect 391 872 397 906
rect 431 872 437 906
rect 391 834 437 872
rect 391 800 397 834
rect 431 800 437 834
rect 391 762 437 800
rect 391 728 397 762
rect 431 728 437 762
rect 391 690 437 728
rect 391 656 397 690
rect 431 656 437 690
rect 391 618 437 656
rect 391 584 397 618
rect 431 584 437 618
rect 391 546 437 584
rect 391 512 397 546
rect 431 512 437 546
rect 391 474 437 512
rect 391 440 397 474
rect 431 440 437 474
rect 391 402 437 440
rect 391 368 397 402
rect 431 368 437 402
rect 391 330 437 368
rect 391 296 397 330
rect 431 296 437 330
rect 391 258 437 296
rect 391 224 397 258
rect 431 224 437 258
rect 391 212 437 224
rect 547 1194 593 1206
rect 547 1160 553 1194
rect 587 1160 593 1194
rect 547 1122 593 1160
rect 547 1088 553 1122
rect 587 1088 593 1122
rect 547 1050 593 1088
rect 547 1016 553 1050
rect 587 1016 593 1050
rect 547 978 593 1016
rect 547 944 553 978
rect 587 944 593 978
rect 547 906 593 944
rect 547 872 553 906
rect 587 872 593 906
rect 547 834 593 872
rect 547 800 553 834
rect 587 800 593 834
rect 547 762 593 800
rect 547 728 553 762
rect 587 728 593 762
rect 547 690 593 728
rect 547 656 553 690
rect 587 656 593 690
rect 547 618 593 656
rect 547 584 553 618
rect 587 584 593 618
rect 547 546 593 584
rect 547 512 553 546
rect 587 512 593 546
rect 547 474 593 512
rect 547 440 553 474
rect 587 440 593 474
rect 547 402 593 440
rect 547 368 553 402
rect 587 368 593 402
rect 547 330 593 368
rect 547 296 553 330
rect 587 296 593 330
rect 547 258 593 296
rect 547 224 553 258
rect 587 224 593 258
rect 547 212 593 224
rect 703 1194 749 1206
rect 703 1160 709 1194
rect 743 1160 749 1194
rect 703 1122 749 1160
rect 703 1088 709 1122
rect 743 1088 749 1122
rect 703 1050 749 1088
rect 703 1016 709 1050
rect 743 1016 749 1050
rect 703 978 749 1016
rect 703 944 709 978
rect 743 944 749 978
rect 703 906 749 944
rect 703 872 709 906
rect 743 872 749 906
rect 703 834 749 872
rect 703 800 709 834
rect 743 800 749 834
rect 703 762 749 800
rect 703 728 709 762
rect 743 728 749 762
rect 703 690 749 728
rect 703 656 709 690
rect 743 656 749 690
rect 703 618 749 656
rect 703 584 709 618
rect 743 584 749 618
rect 703 546 749 584
rect 703 512 709 546
rect 743 512 749 546
rect 703 474 749 512
rect 703 440 709 474
rect 743 440 749 474
rect 703 402 749 440
rect 703 368 709 402
rect 743 368 749 402
rect 703 330 749 368
rect 703 296 709 330
rect 743 296 749 330
rect 703 258 749 296
rect 703 224 709 258
rect 743 224 749 258
rect 703 212 749 224
rect 859 1194 905 1206
rect 859 1160 865 1194
rect 899 1160 905 1194
rect 859 1122 905 1160
rect 859 1088 865 1122
rect 899 1088 905 1122
rect 859 1050 905 1088
rect 859 1016 865 1050
rect 899 1016 905 1050
rect 859 978 905 1016
rect 859 944 865 978
rect 899 944 905 978
rect 859 906 905 944
rect 859 872 865 906
rect 899 872 905 906
rect 859 834 905 872
rect 859 800 865 834
rect 899 800 905 834
rect 859 762 905 800
rect 859 728 865 762
rect 899 728 905 762
rect 859 690 905 728
rect 859 656 865 690
rect 899 656 905 690
rect 859 618 905 656
rect 859 584 865 618
rect 899 584 905 618
rect 859 546 905 584
rect 859 512 865 546
rect 899 512 905 546
rect 859 474 905 512
rect 859 440 865 474
rect 899 440 905 474
rect 859 402 905 440
rect 859 368 865 402
rect 899 368 905 402
rect 859 330 905 368
rect 859 296 865 330
rect 899 296 905 330
rect 859 258 905 296
rect 859 224 865 258
rect 899 224 905 258
rect 859 212 905 224
rect 1015 1194 1061 1293
rect 1015 1160 1021 1194
rect 1055 1160 1061 1194
rect 1015 1122 1061 1160
rect 1015 1088 1021 1122
rect 1055 1088 1061 1122
rect 1015 1050 1061 1088
rect 1015 1016 1021 1050
rect 1055 1016 1061 1050
rect 1015 978 1061 1016
rect 1015 944 1021 978
rect 1055 944 1061 978
rect 1015 906 1061 944
rect 1015 872 1021 906
rect 1055 872 1061 906
rect 1015 834 1061 872
rect 1015 800 1021 834
rect 1055 800 1061 834
rect 1015 762 1061 800
rect 1015 728 1021 762
rect 1055 728 1061 762
rect 1015 690 1061 728
rect 1015 656 1021 690
rect 1055 656 1061 690
rect 1015 618 1061 656
rect 1015 584 1021 618
rect 1055 584 1061 618
rect 1015 546 1061 584
rect 1015 512 1021 546
rect 1055 512 1061 546
rect 1015 474 1061 512
rect 1015 440 1021 474
rect 1055 440 1061 474
rect 1015 402 1061 440
rect 1015 368 1021 402
rect 1055 368 1061 402
rect 1015 330 1061 368
rect 1015 296 1021 330
rect 1055 296 1061 330
rect 1015 258 1061 296
rect 1015 224 1021 258
rect 1055 224 1061 258
rect 1015 212 1061 224
rect 309 147 320 181
rect 354 147 363 181
rect 309 109 363 147
rect 309 75 320 109
rect 354 75 363 109
rect 309 33 363 75
use sky130_fd_pr__nfet_01v8__example_55959141808248  sky130_fd_pr__nfet_01v8__example_55959141808248_0
timestamp 1666199351
transform 1 0 910 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808445  sky130_fd_pr__nfet_01v8__example_55959141808445_0
timestamp 1666199351
transform 1 0 286 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808447  sky130_fd_pr__nfet_01v8__example_55959141808447_0
timestamp 1666199351
transform 1 0 442 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808447  sky130_fd_pr__nfet_01v8__example_55959141808447_1
timestamp 1666199351
transform 1 0 598 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808447  sky130_fd_pr__nfet_01v8__example_55959141808447_2
timestamp 1666199351
transform 1 0 754 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808455  sky130_fd_pr__nfet_01v8__example_55959141808455_0
timestamp 1666199351
transform -1 0 212 0 -1 1102
box -19 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808584  sky130_fd_pr__nfet_01v8__example_55959141808584_0
timestamp 1666199351
transform -1 0 212 0 -1 770
box 100 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808450  sky130_fd_pr__pfet_01v8__example_55959141808450_0
timestamp 1666199351
transform -1 0 720 0 -1 1650
box -1 0 297 1
use sky130_fd_pr__pfet_01v8__example_55959141808451  sky130_fd_pr__pfet_01v8__example_55959141808451_0
timestamp 1666199351
transform 1 0 794 0 -1 1650
box -19 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808457  sky130_fd_pr__pfet_01v8__example_55959141808457_0
timestamp 1666199351
transform 1 0 72 0 -1 1650
box -1 0 297 1
<< labels >>
flabel metal1 s 940 1345 968 1373 3 FreeSans 280 180 0 0 OUT
port 1 nsew
flabel metal1 s 305 1739 462 1826 3 FreeSans 520 0 0 0 VPWR
port 2 nsew
flabel metal1 s 94 617 94 617 3 FreeSans 520 0 0 0 VGND
port 3 nsew
flabel locali s 946 109 974 137 3 FreeSans 280 270 0 0 IN1
port 4 nsew
flabel locali s 322 109 350 137 3 FreeSans 280 270 0 0 IN0
port 5 nsew
flabel locali s 636 109 664 137 3 FreeSans 280 270 0 0 IN3
port 6 nsew
flabel locali s 790 109 818 137 3 FreeSans 280 270 0 0 IN2
port 7 nsew
flabel locali s 482 109 510 137 3 FreeSans 280 270 0 0 IN4
port 8 nsew
<< properties >>
string GDS_END 43891746
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43877292
<< end >>
