magic
tech sky130B
timestamp 1666199351
<< properties >>
string GDS_END 36254
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 35930
<< end >>
