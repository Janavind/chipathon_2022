magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect 24063 16338 24705 19291
rect 26946 14917 27112 20896
<< pwell >>
rect 27181 37181 27657 37657
rect 23635 22873 28026 23379
rect 26249 22054 28026 22873
rect 16801 9534 17639 9620
rect 2294 3728 28026 4086
rect 2294 3404 3342 3728
rect 6423 3404 28026 3728
<< ndiff >>
rect 27319 37504 27519 37519
rect 27319 37334 27334 37504
rect 27504 37334 27519 37504
rect 27319 37319 27519 37334
<< ndiffc >>
rect 27334 37334 27504 37504
<< psubdiff >>
rect 27207 37619 27631 37631
rect 27207 37585 27287 37619
rect 27321 37585 27355 37619
rect 27389 37585 27423 37619
rect 27457 37585 27491 37619
rect 27525 37585 27631 37619
rect 27207 37573 27585 37585
rect 27207 37559 27265 37573
rect 27207 37525 27219 37559
rect 27253 37525 27265 37559
rect 27207 37491 27265 37525
rect 27573 37551 27585 37573
rect 27619 37551 27631 37585
rect 27207 37457 27219 37491
rect 27253 37457 27265 37491
rect 27207 37423 27265 37457
rect 27207 37389 27219 37423
rect 27253 37389 27265 37423
rect 27207 37355 27265 37389
rect 27207 37321 27219 37355
rect 27253 37321 27265 37355
rect 27207 37287 27265 37321
rect 27573 37517 27631 37551
rect 27573 37483 27585 37517
rect 27619 37483 27631 37517
rect 27573 37449 27631 37483
rect 27573 37415 27585 37449
rect 27619 37415 27631 37449
rect 27573 37381 27631 37415
rect 27573 37347 27585 37381
rect 27619 37347 27631 37381
rect 27207 37253 27219 37287
rect 27253 37265 27265 37287
rect 27573 37265 27631 37347
rect 27253 37253 27631 37265
rect 27207 37219 27347 37253
rect 27381 37219 27415 37253
rect 27449 37219 27483 37253
rect 27517 37219 27551 37253
rect 27585 37219 27631 37253
rect 27207 37207 27631 37219
rect 2320 4058 3350 4060
rect 2320 4024 2344 4058
rect 2378 4024 2415 4058
rect 2449 4024 2486 4058
rect 2520 4024 2557 4058
rect 2591 4024 2628 4058
rect 2662 4024 2698 4058
rect 2732 4024 2768 4058
rect 2802 4024 2838 4058
rect 2872 4024 2908 4058
rect 2942 4024 2978 4058
rect 3012 4024 3048 4058
rect 3082 4024 3118 4058
rect 3152 4024 3188 4058
rect 3222 4024 3258 4058
rect 3292 4026 3350 4058
rect 3384 4026 3419 4060
rect 3453 4026 3488 4060
rect 3522 4026 3557 4060
rect 3591 4026 3626 4060
rect 3660 4026 3695 4060
rect 3729 4026 3764 4060
rect 3798 4026 3833 4060
rect 3867 4026 3902 4060
rect 3936 4026 3971 4060
rect 4005 4026 4040 4060
rect 4074 4026 4109 4060
rect 4143 4026 4178 4060
rect 4212 4026 4247 4060
rect 4281 4026 4316 4060
rect 4350 4026 4385 4060
rect 4419 4026 4454 4060
rect 4488 4026 4523 4060
rect 4557 4026 4592 4060
rect 4626 4026 4661 4060
rect 4695 4026 4730 4060
rect 4764 4026 4799 4060
rect 4833 4026 4868 4060
rect 4902 4026 4937 4060
rect 4971 4026 5006 4060
rect 5040 4026 5075 4060
rect 5109 4026 5144 4060
rect 5178 4026 5213 4060
rect 5247 4026 5282 4060
rect 5316 4026 5351 4060
rect 5385 4026 5420 4060
rect 5454 4026 5489 4060
rect 5523 4026 5558 4060
rect 5592 4026 5627 4060
rect 5661 4026 5696 4060
rect 5730 4026 5765 4060
rect 5799 4026 5834 4060
rect 5868 4026 5903 4060
rect 5937 4026 5972 4060
rect 6006 4026 6041 4060
rect 3292 4024 6041 4026
rect 2320 3992 6041 4024
rect 2320 3984 3350 3992
rect 2320 3950 2344 3984
rect 2378 3950 2415 3984
rect 2449 3950 2486 3984
rect 2520 3950 2557 3984
rect 2591 3950 2628 3984
rect 2662 3950 2698 3984
rect 2732 3950 2768 3984
rect 2802 3950 2838 3984
rect 2872 3950 2908 3984
rect 2942 3950 2978 3984
rect 3012 3950 3048 3984
rect 3082 3950 3118 3984
rect 3152 3950 3188 3984
rect 3222 3950 3258 3984
rect 3292 3958 3350 3984
rect 3384 3958 3419 3992
rect 3453 3958 3488 3992
rect 3522 3958 3557 3992
rect 3591 3958 3626 3992
rect 3660 3958 3695 3992
rect 3729 3958 3764 3992
rect 3798 3958 3833 3992
rect 3867 3958 3902 3992
rect 3936 3958 3971 3992
rect 4005 3958 4040 3992
rect 4074 3958 4109 3992
rect 4143 3958 4178 3992
rect 4212 3958 4247 3992
rect 4281 3958 4316 3992
rect 4350 3958 4385 3992
rect 4419 3958 4454 3992
rect 4488 3958 4523 3992
rect 4557 3958 4592 3992
rect 4626 3958 4661 3992
rect 4695 3958 4730 3992
rect 4764 3958 4799 3992
rect 4833 3958 4868 3992
rect 4902 3958 4937 3992
rect 4971 3958 5006 3992
rect 5040 3958 5075 3992
rect 5109 3958 5144 3992
rect 5178 3958 5213 3992
rect 5247 3958 5282 3992
rect 5316 3958 5351 3992
rect 5385 3958 5420 3992
rect 5454 3958 5489 3992
rect 5523 3958 5558 3992
rect 5592 3958 5627 3992
rect 5661 3958 5696 3992
rect 5730 3958 5765 3992
rect 5799 3958 5834 3992
rect 5868 3958 5903 3992
rect 5937 3958 5972 3992
rect 6006 3958 6041 3992
rect 3292 3950 6041 3958
rect 2320 3924 6041 3950
rect 2320 3910 3350 3924
rect 2320 3876 2344 3910
rect 2378 3876 2415 3910
rect 2449 3876 2486 3910
rect 2520 3876 2557 3910
rect 2591 3876 2628 3910
rect 2662 3876 2698 3910
rect 2732 3876 2768 3910
rect 2802 3876 2838 3910
rect 2872 3876 2908 3910
rect 2942 3876 2978 3910
rect 3012 3876 3048 3910
rect 3082 3876 3118 3910
rect 3152 3876 3188 3910
rect 3222 3876 3258 3910
rect 3292 3890 3350 3910
rect 3384 3890 3419 3924
rect 3453 3890 3488 3924
rect 3522 3890 3557 3924
rect 3591 3890 3626 3924
rect 3660 3890 3695 3924
rect 3729 3890 3764 3924
rect 3798 3890 3833 3924
rect 3867 3890 3902 3924
rect 3936 3890 3971 3924
rect 4005 3890 4040 3924
rect 4074 3890 4109 3924
rect 4143 3890 4178 3924
rect 4212 3890 4247 3924
rect 4281 3890 4316 3924
rect 4350 3890 4385 3924
rect 4419 3890 4454 3924
rect 4488 3890 4523 3924
rect 4557 3890 4592 3924
rect 4626 3890 4661 3924
rect 4695 3890 4730 3924
rect 4764 3890 4799 3924
rect 4833 3890 4868 3924
rect 4902 3890 4937 3924
rect 4971 3890 5006 3924
rect 5040 3890 5075 3924
rect 5109 3890 5144 3924
rect 5178 3890 5213 3924
rect 5247 3890 5282 3924
rect 5316 3890 5351 3924
rect 5385 3890 5420 3924
rect 5454 3890 5489 3924
rect 5523 3890 5558 3924
rect 5592 3890 5627 3924
rect 5661 3890 5696 3924
rect 5730 3890 5765 3924
rect 5799 3890 5834 3924
rect 5868 3890 5903 3924
rect 5937 3890 5972 3924
rect 6006 3890 6041 3924
rect 3292 3876 6041 3890
rect 2320 3856 6041 3876
rect 2320 3836 3350 3856
rect 2320 3802 2344 3836
rect 2378 3802 2415 3836
rect 2449 3802 2486 3836
rect 2520 3802 2557 3836
rect 2591 3802 2628 3836
rect 2662 3802 2698 3836
rect 2732 3802 2768 3836
rect 2802 3802 2838 3836
rect 2872 3802 2908 3836
rect 2942 3802 2978 3836
rect 3012 3802 3048 3836
rect 3082 3802 3118 3836
rect 3152 3802 3188 3836
rect 3222 3802 3258 3836
rect 3292 3822 3350 3836
rect 3384 3822 3419 3856
rect 3453 3822 3488 3856
rect 3522 3822 3557 3856
rect 3591 3822 3626 3856
rect 3660 3822 3695 3856
rect 3729 3822 3764 3856
rect 3798 3822 3833 3856
rect 3867 3822 3902 3856
rect 3936 3822 3971 3856
rect 4005 3822 4040 3856
rect 4074 3822 4109 3856
rect 4143 3822 4178 3856
rect 4212 3822 4247 3856
rect 4281 3822 4316 3856
rect 4350 3822 4385 3856
rect 4419 3822 4454 3856
rect 4488 3822 4523 3856
rect 4557 3822 4592 3856
rect 4626 3822 4661 3856
rect 4695 3822 4730 3856
rect 4764 3822 4799 3856
rect 4833 3822 4868 3856
rect 4902 3822 4937 3856
rect 4971 3822 5006 3856
rect 5040 3822 5075 3856
rect 5109 3822 5144 3856
rect 5178 3822 5213 3856
rect 5247 3822 5282 3856
rect 5316 3822 5351 3856
rect 5385 3822 5420 3856
rect 5454 3822 5489 3856
rect 5523 3822 5558 3856
rect 5592 3822 5627 3856
rect 5661 3822 5696 3856
rect 5730 3822 5765 3856
rect 5799 3822 5834 3856
rect 5868 3822 5903 3856
rect 5937 3822 5972 3856
rect 6006 3822 6041 3856
rect 3292 3802 6041 3822
rect 2320 3788 6041 3802
rect 2320 3762 3350 3788
rect 2320 3728 2344 3762
rect 2378 3728 2415 3762
rect 2449 3728 2486 3762
rect 2520 3728 2557 3762
rect 2591 3728 2628 3762
rect 2662 3728 2698 3762
rect 2732 3728 2768 3762
rect 2802 3728 2838 3762
rect 2872 3728 2908 3762
rect 2942 3728 2978 3762
rect 3012 3728 3048 3762
rect 3082 3728 3118 3762
rect 3152 3728 3188 3762
rect 3222 3728 3258 3762
rect 3292 3754 3350 3762
rect 3384 3754 3419 3788
rect 3453 3754 3488 3788
rect 3522 3754 3557 3788
rect 3591 3754 3626 3788
rect 3660 3754 3695 3788
rect 3729 3754 3764 3788
rect 3798 3754 3833 3788
rect 3867 3754 3902 3788
rect 3936 3754 3971 3788
rect 4005 3754 4040 3788
rect 4074 3754 4109 3788
rect 4143 3754 4178 3788
rect 4212 3754 4247 3788
rect 4281 3754 4316 3788
rect 4350 3754 4385 3788
rect 4419 3754 4454 3788
rect 4488 3754 4523 3788
rect 4557 3754 4592 3788
rect 4626 3754 4661 3788
rect 4695 3754 4730 3788
rect 4764 3754 4799 3788
rect 4833 3754 4868 3788
rect 4902 3754 4937 3788
rect 4971 3754 5006 3788
rect 5040 3754 5075 3788
rect 5109 3754 5144 3788
rect 5178 3754 5213 3788
rect 5247 3754 5282 3788
rect 5316 3754 5351 3788
rect 5385 3754 5420 3788
rect 5454 3754 5489 3788
rect 5523 3754 5558 3788
rect 5592 3754 5627 3788
rect 5661 3754 5696 3788
rect 5730 3754 5765 3788
rect 5799 3754 5834 3788
rect 5868 3754 5903 3788
rect 5937 3754 5972 3788
rect 6006 3754 6041 3788
rect 6415 4058 28000 4060
rect 6415 4024 6473 4058
rect 6507 4024 6542 4058
rect 6576 4024 6611 4058
rect 6645 4024 6680 4058
rect 6714 4024 6749 4058
rect 6783 4024 6818 4058
rect 6852 4024 6887 4058
rect 6921 4024 6956 4058
rect 6990 4024 7025 4058
rect 7059 4024 7094 4058
rect 7128 4024 7163 4058
rect 7197 4024 7232 4058
rect 7266 4024 7301 4058
rect 7335 4024 7370 4058
rect 7404 4024 7439 4058
rect 7473 4024 7508 4058
rect 7542 4024 7577 4058
rect 7611 4024 7646 4058
rect 7680 4024 7715 4058
rect 7749 4024 7784 4058
rect 7818 4024 7853 4058
rect 7887 4024 7922 4058
rect 7956 4024 7991 4058
rect 8025 4024 8060 4058
rect 8094 4024 8129 4058
rect 8163 4024 8198 4058
rect 8232 4024 8267 4058
rect 8301 4024 8336 4058
rect 8370 4024 8405 4058
rect 8439 4024 8474 4058
rect 8508 4024 8543 4058
rect 8577 4024 8612 4058
rect 8646 4024 8681 4058
rect 8715 4024 8750 4058
rect 8784 4024 8819 4058
rect 8853 4024 8888 4058
rect 8922 4024 8957 4058
rect 8991 4024 9026 4058
rect 9060 4024 9095 4058
rect 9129 4024 9164 4058
rect 9198 4024 9233 4058
rect 9267 4024 9302 4058
rect 9336 4024 9371 4058
rect 9405 4024 9440 4058
rect 9474 4024 9509 4058
rect 9543 4024 9578 4058
rect 9612 4024 9647 4058
rect 9681 4024 9716 4058
rect 9750 4024 9785 4058
rect 9819 4024 9854 4058
rect 9888 4024 9922 4058
rect 9956 4024 9990 4058
rect 10024 4024 10058 4058
rect 10092 4024 10126 4058
rect 10160 4024 10194 4058
rect 10228 4024 10262 4058
rect 10296 4024 10330 4058
rect 10364 4024 10398 4058
rect 10432 4024 10466 4058
rect 10500 4024 10534 4058
rect 10568 4024 10602 4058
rect 10636 4024 10670 4058
rect 10704 4024 10738 4058
rect 10772 4024 10806 4058
rect 10840 4024 10874 4058
rect 10908 4024 10942 4058
rect 10976 4024 11010 4058
rect 11044 4024 11078 4058
rect 11112 4024 11146 4058
rect 11180 4024 11214 4058
rect 11248 4024 11282 4058
rect 11316 4024 11350 4058
rect 11384 4024 11418 4058
rect 11452 4024 11486 4058
rect 11520 4024 11554 4058
rect 11588 4024 11622 4058
rect 11656 4024 11690 4058
rect 11724 4024 11758 4058
rect 11792 4024 11826 4058
rect 11860 4024 11894 4058
rect 11928 4024 11962 4058
rect 11996 4024 12030 4058
rect 12064 4024 12098 4058
rect 12132 4024 12166 4058
rect 12200 4024 12234 4058
rect 12268 4024 12302 4058
rect 12336 4024 12370 4058
rect 12404 4024 12438 4058
rect 12472 4024 12506 4058
rect 12540 4024 12574 4058
rect 12608 4024 12642 4058
rect 12676 4024 12710 4058
rect 12744 4024 12778 4058
rect 12812 4024 12846 4058
rect 12880 4024 12914 4058
rect 12948 4024 12982 4058
rect 13016 4024 13050 4058
rect 13084 4024 13118 4058
rect 13152 4024 13186 4058
rect 13220 4024 13254 4058
rect 13288 4024 13322 4058
rect 13356 4024 13390 4058
rect 13424 4024 13458 4058
rect 13492 4024 13526 4058
rect 13560 4024 13594 4058
rect 13628 4024 13662 4058
rect 13696 4024 13730 4058
rect 13764 4024 13798 4058
rect 13832 4024 13866 4058
rect 13900 4024 13934 4058
rect 13968 4024 14002 4058
rect 14036 4024 14070 4058
rect 14104 4024 14138 4058
rect 14172 4024 14206 4058
rect 14240 4024 14274 4058
rect 14308 4024 14342 4058
rect 14376 4024 14410 4058
rect 14444 4024 14478 4058
rect 14512 4024 14546 4058
rect 14580 4024 14614 4058
rect 14648 4024 14682 4058
rect 14716 4024 14750 4058
rect 14784 4024 14818 4058
rect 14852 4024 14886 4058
rect 14920 4024 14954 4058
rect 14988 4024 15022 4058
rect 15056 4024 15090 4058
rect 15124 4024 15158 4058
rect 15192 4024 15226 4058
rect 15260 4024 15294 4058
rect 15328 4024 15362 4058
rect 15396 4024 15430 4058
rect 15464 4024 15498 4058
rect 15532 4024 15566 4058
rect 15600 4024 15634 4058
rect 15668 4024 15702 4058
rect 15736 4024 15770 4058
rect 15804 4024 15838 4058
rect 15872 4024 15906 4058
rect 15940 4024 15974 4058
rect 16008 4024 16042 4058
rect 16076 4024 16110 4058
rect 16144 4024 16178 4058
rect 16212 4024 16246 4058
rect 16280 4024 16314 4058
rect 16348 4024 16382 4058
rect 16416 4024 16450 4058
rect 16484 4024 16518 4058
rect 16552 4024 16586 4058
rect 16620 4024 16654 4058
rect 16688 4024 16722 4058
rect 16756 4024 16790 4058
rect 16824 4024 16858 4058
rect 16892 4024 16926 4058
rect 16960 4024 16994 4058
rect 17028 4024 17062 4058
rect 17096 4024 17130 4058
rect 17164 4024 17198 4058
rect 17232 4024 17266 4058
rect 17300 4024 17334 4058
rect 17368 4024 17402 4058
rect 17436 4024 17470 4058
rect 17504 4024 17538 4058
rect 17572 4024 17606 4058
rect 17640 4024 17674 4058
rect 17708 4024 17742 4058
rect 17776 4024 17810 4058
rect 17844 4024 17878 4058
rect 17912 4024 17946 4058
rect 17980 4024 18014 4058
rect 18048 4024 18082 4058
rect 18116 4024 18150 4058
rect 18184 4024 18218 4058
rect 18252 4024 18286 4058
rect 18320 4024 18354 4058
rect 18388 4024 18422 4058
rect 18456 4024 18490 4058
rect 18524 4024 18558 4058
rect 18592 4024 18626 4058
rect 18660 4024 18694 4058
rect 18728 4024 18762 4058
rect 18796 4024 18830 4058
rect 18864 4024 18898 4058
rect 18932 4024 18966 4058
rect 19000 4024 19034 4058
rect 19068 4024 19102 4058
rect 19136 4024 19170 4058
rect 19204 4024 19238 4058
rect 19272 4024 19306 4058
rect 19340 4024 19374 4058
rect 19408 4024 19442 4058
rect 19476 4024 19510 4058
rect 19544 4024 19578 4058
rect 19612 4024 19646 4058
rect 19680 4024 19714 4058
rect 19748 4024 19782 4058
rect 19816 4024 19850 4058
rect 19884 4024 19918 4058
rect 19952 4024 19986 4058
rect 20020 4024 20054 4058
rect 20088 4024 20122 4058
rect 20156 4024 20190 4058
rect 20224 4024 20258 4058
rect 20292 4024 20326 4058
rect 20360 4024 20394 4058
rect 20428 4024 20462 4058
rect 20496 4024 20530 4058
rect 20564 4024 20598 4058
rect 20632 4024 20666 4058
rect 20700 4024 20734 4058
rect 20768 4024 20802 4058
rect 20836 4024 20870 4058
rect 20904 4024 20938 4058
rect 20972 4024 21006 4058
rect 21040 4024 21074 4058
rect 21108 4024 21142 4058
rect 21176 4024 21210 4058
rect 21244 4024 21278 4058
rect 21312 4024 21346 4058
rect 21380 4024 21414 4058
rect 21448 4024 21482 4058
rect 21516 4024 21550 4058
rect 21584 4024 21618 4058
rect 21652 4024 21686 4058
rect 21720 4024 21754 4058
rect 21788 4024 21822 4058
rect 21856 4024 21890 4058
rect 21924 4024 21958 4058
rect 21992 4024 22026 4058
rect 22060 4024 22094 4058
rect 22128 4024 22162 4058
rect 22196 4024 22230 4058
rect 22264 4024 22298 4058
rect 22332 4024 22366 4058
rect 22400 4024 22434 4058
rect 22468 4024 22502 4058
rect 22536 4024 22570 4058
rect 22604 4024 22638 4058
rect 22672 4024 22706 4058
rect 22740 4024 22774 4058
rect 22808 4024 22842 4058
rect 22876 4024 22910 4058
rect 22944 4024 22978 4058
rect 23012 4024 23046 4058
rect 23080 4024 23114 4058
rect 23148 4024 23182 4058
rect 23216 4024 23250 4058
rect 23284 4024 23318 4058
rect 23352 4024 23386 4058
rect 23420 4024 23454 4058
rect 23488 4024 23522 4058
rect 23556 4024 23590 4058
rect 23624 4024 23658 4058
rect 23692 4024 23726 4058
rect 23760 4024 23794 4058
rect 23828 4024 23862 4058
rect 23896 4024 23930 4058
rect 23964 4024 23998 4058
rect 24032 4024 24066 4058
rect 24100 4024 24134 4058
rect 24168 4024 24202 4058
rect 24236 4024 24270 4058
rect 24304 4024 24338 4058
rect 24372 4024 24406 4058
rect 24440 4024 24474 4058
rect 24508 4024 24542 4058
rect 24576 4024 24610 4058
rect 24644 4024 24678 4058
rect 24712 4024 24746 4058
rect 24780 4024 24814 4058
rect 24848 4024 24882 4058
rect 24916 4024 24950 4058
rect 24984 4024 25018 4058
rect 25052 4024 25086 4058
rect 25120 4024 25154 4058
rect 25188 4024 25222 4058
rect 25256 4024 25290 4058
rect 25324 4024 25358 4058
rect 25392 4024 25426 4058
rect 25460 4024 25494 4058
rect 25528 4024 25562 4058
rect 25596 4024 25630 4058
rect 25664 4024 25698 4058
rect 25732 4024 25766 4058
rect 25800 4024 25834 4058
rect 25868 4024 25902 4058
rect 25936 4024 25970 4058
rect 26004 4024 26038 4058
rect 26072 4024 26106 4058
rect 26140 4024 26174 4058
rect 26208 4024 26242 4058
rect 26276 4024 26310 4058
rect 26344 4024 26378 4058
rect 26412 4024 26446 4058
rect 26480 4024 26514 4058
rect 26548 4024 26582 4058
rect 26616 4024 26650 4058
rect 26684 4024 26718 4058
rect 26752 4024 26786 4058
rect 26820 4024 26854 4058
rect 26888 4024 26922 4058
rect 26956 4024 26990 4058
rect 27024 4024 27058 4058
rect 27092 4024 27126 4058
rect 27160 4024 27194 4058
rect 27228 4024 27262 4058
rect 27296 4024 27330 4058
rect 27364 4024 27398 4058
rect 27432 4024 27466 4058
rect 27500 4024 27534 4058
rect 27568 4024 27602 4058
rect 27636 4024 27670 4058
rect 27704 4024 27738 4058
rect 27772 4024 27806 4058
rect 27840 4024 27874 4058
rect 27908 4024 27942 4058
rect 27976 4024 28000 4058
rect 6415 3984 28000 4024
rect 6415 3950 6473 3984
rect 6507 3950 6542 3984
rect 6576 3950 6611 3984
rect 6645 3950 6680 3984
rect 6714 3950 6749 3984
rect 6783 3950 6818 3984
rect 6852 3950 6887 3984
rect 6921 3950 6956 3984
rect 6990 3950 7025 3984
rect 7059 3950 7094 3984
rect 7128 3950 7163 3984
rect 7197 3950 7232 3984
rect 7266 3950 7301 3984
rect 7335 3950 7370 3984
rect 7404 3950 7439 3984
rect 7473 3950 7508 3984
rect 7542 3950 7577 3984
rect 7611 3950 7646 3984
rect 7680 3950 7715 3984
rect 7749 3950 7784 3984
rect 7818 3950 7853 3984
rect 7887 3950 7922 3984
rect 7956 3950 7991 3984
rect 8025 3950 8060 3984
rect 8094 3950 8129 3984
rect 8163 3950 8198 3984
rect 8232 3950 8267 3984
rect 8301 3950 8336 3984
rect 8370 3950 8405 3984
rect 8439 3950 8474 3984
rect 8508 3950 8543 3984
rect 8577 3950 8612 3984
rect 8646 3950 8681 3984
rect 8715 3950 8750 3984
rect 8784 3950 8819 3984
rect 8853 3950 8888 3984
rect 8922 3950 8957 3984
rect 8991 3950 9026 3984
rect 9060 3950 9095 3984
rect 9129 3950 9164 3984
rect 9198 3950 9233 3984
rect 9267 3950 9302 3984
rect 9336 3950 9371 3984
rect 9405 3950 9440 3984
rect 9474 3950 9509 3984
rect 9543 3950 9578 3984
rect 9612 3950 9647 3984
rect 9681 3950 9716 3984
rect 9750 3950 9785 3984
rect 9819 3950 9854 3984
rect 9888 3950 9922 3984
rect 9956 3950 9990 3984
rect 10024 3950 10058 3984
rect 10092 3950 10126 3984
rect 10160 3950 10194 3984
rect 10228 3950 10262 3984
rect 10296 3950 10330 3984
rect 10364 3950 10398 3984
rect 10432 3950 10466 3984
rect 10500 3950 10534 3984
rect 10568 3950 10602 3984
rect 10636 3950 10670 3984
rect 10704 3950 10738 3984
rect 10772 3950 10806 3984
rect 10840 3950 10874 3984
rect 10908 3950 10942 3984
rect 10976 3950 11010 3984
rect 11044 3950 11078 3984
rect 11112 3950 11146 3984
rect 11180 3950 11214 3984
rect 11248 3950 11282 3984
rect 11316 3950 11350 3984
rect 11384 3950 11418 3984
rect 11452 3950 11486 3984
rect 11520 3950 11554 3984
rect 11588 3950 11622 3984
rect 11656 3950 11690 3984
rect 11724 3950 11758 3984
rect 11792 3950 11826 3984
rect 11860 3950 11894 3984
rect 11928 3950 11962 3984
rect 11996 3950 12030 3984
rect 12064 3950 12098 3984
rect 12132 3950 12166 3984
rect 12200 3950 12234 3984
rect 12268 3950 12302 3984
rect 12336 3950 12370 3984
rect 12404 3950 12438 3984
rect 12472 3950 12506 3984
rect 12540 3950 12574 3984
rect 12608 3950 12642 3984
rect 12676 3950 12710 3984
rect 12744 3950 12778 3984
rect 12812 3950 12846 3984
rect 12880 3950 12914 3984
rect 12948 3950 12982 3984
rect 13016 3950 13050 3984
rect 13084 3950 13118 3984
rect 13152 3950 13186 3984
rect 13220 3950 13254 3984
rect 13288 3950 13322 3984
rect 13356 3950 13390 3984
rect 13424 3950 13458 3984
rect 13492 3950 13526 3984
rect 13560 3950 13594 3984
rect 13628 3950 13662 3984
rect 13696 3950 13730 3984
rect 13764 3950 13798 3984
rect 13832 3950 13866 3984
rect 13900 3950 13934 3984
rect 13968 3950 14002 3984
rect 14036 3950 14070 3984
rect 14104 3950 14138 3984
rect 14172 3950 14206 3984
rect 14240 3950 14274 3984
rect 14308 3950 14342 3984
rect 14376 3950 14410 3984
rect 14444 3950 14478 3984
rect 14512 3950 14546 3984
rect 14580 3950 14614 3984
rect 14648 3950 14682 3984
rect 14716 3950 14750 3984
rect 14784 3950 14818 3984
rect 14852 3950 14886 3984
rect 14920 3950 14954 3984
rect 14988 3950 15022 3984
rect 15056 3950 15090 3984
rect 15124 3950 15158 3984
rect 15192 3950 15226 3984
rect 15260 3950 15294 3984
rect 15328 3950 15362 3984
rect 15396 3950 15430 3984
rect 15464 3950 15498 3984
rect 15532 3950 15566 3984
rect 15600 3950 15634 3984
rect 15668 3950 15702 3984
rect 15736 3950 15770 3984
rect 15804 3950 15838 3984
rect 15872 3950 15906 3984
rect 15940 3950 15974 3984
rect 16008 3950 16042 3984
rect 16076 3950 16110 3984
rect 16144 3950 16178 3984
rect 16212 3950 16246 3984
rect 16280 3950 16314 3984
rect 16348 3950 16382 3984
rect 16416 3950 16450 3984
rect 16484 3950 16518 3984
rect 16552 3950 16586 3984
rect 16620 3950 16654 3984
rect 16688 3950 16722 3984
rect 16756 3950 16790 3984
rect 16824 3950 16858 3984
rect 16892 3950 16926 3984
rect 16960 3950 16994 3984
rect 17028 3950 17062 3984
rect 17096 3950 17130 3984
rect 17164 3950 17198 3984
rect 17232 3950 17266 3984
rect 17300 3950 17334 3984
rect 17368 3950 17402 3984
rect 17436 3950 17470 3984
rect 17504 3950 17538 3984
rect 17572 3950 17606 3984
rect 17640 3950 17674 3984
rect 17708 3950 17742 3984
rect 17776 3950 17810 3984
rect 17844 3950 17878 3984
rect 17912 3950 17946 3984
rect 17980 3950 18014 3984
rect 18048 3950 18082 3984
rect 18116 3950 18150 3984
rect 18184 3950 18218 3984
rect 18252 3950 18286 3984
rect 18320 3950 18354 3984
rect 18388 3950 18422 3984
rect 18456 3950 18490 3984
rect 18524 3950 18558 3984
rect 18592 3950 18626 3984
rect 18660 3950 18694 3984
rect 18728 3950 18762 3984
rect 18796 3950 18830 3984
rect 18864 3950 18898 3984
rect 18932 3950 18966 3984
rect 19000 3950 19034 3984
rect 19068 3950 19102 3984
rect 19136 3950 19170 3984
rect 19204 3950 19238 3984
rect 19272 3950 19306 3984
rect 19340 3950 19374 3984
rect 19408 3950 19442 3984
rect 19476 3950 19510 3984
rect 19544 3950 19578 3984
rect 19612 3950 19646 3984
rect 19680 3950 19714 3984
rect 19748 3950 19782 3984
rect 19816 3950 19850 3984
rect 19884 3950 19918 3984
rect 19952 3950 19986 3984
rect 20020 3950 20054 3984
rect 20088 3950 20122 3984
rect 20156 3950 20190 3984
rect 20224 3950 20258 3984
rect 20292 3950 20326 3984
rect 20360 3950 20394 3984
rect 20428 3950 20462 3984
rect 20496 3950 20530 3984
rect 20564 3950 20598 3984
rect 20632 3950 20666 3984
rect 20700 3950 20734 3984
rect 20768 3950 20802 3984
rect 20836 3950 20870 3984
rect 20904 3950 20938 3984
rect 20972 3950 21006 3984
rect 21040 3950 21074 3984
rect 21108 3950 21142 3984
rect 21176 3950 21210 3984
rect 21244 3950 21278 3984
rect 21312 3950 21346 3984
rect 21380 3950 21414 3984
rect 21448 3950 21482 3984
rect 21516 3950 21550 3984
rect 21584 3950 21618 3984
rect 21652 3950 21686 3984
rect 21720 3950 21754 3984
rect 21788 3950 21822 3984
rect 21856 3950 21890 3984
rect 21924 3950 21958 3984
rect 21992 3950 22026 3984
rect 22060 3950 22094 3984
rect 22128 3950 22162 3984
rect 22196 3950 22230 3984
rect 22264 3950 22298 3984
rect 22332 3950 22366 3984
rect 22400 3950 22434 3984
rect 22468 3950 22502 3984
rect 22536 3950 22570 3984
rect 22604 3950 22638 3984
rect 22672 3950 22706 3984
rect 22740 3950 22774 3984
rect 22808 3950 22842 3984
rect 22876 3950 22910 3984
rect 22944 3950 22978 3984
rect 23012 3950 23046 3984
rect 23080 3950 23114 3984
rect 23148 3950 23182 3984
rect 23216 3950 23250 3984
rect 23284 3950 23318 3984
rect 23352 3950 23386 3984
rect 23420 3950 23454 3984
rect 23488 3950 23522 3984
rect 23556 3950 23590 3984
rect 23624 3950 23658 3984
rect 23692 3950 23726 3984
rect 23760 3950 23794 3984
rect 23828 3950 23862 3984
rect 23896 3950 23930 3984
rect 23964 3950 23998 3984
rect 24032 3950 24066 3984
rect 24100 3950 24134 3984
rect 24168 3950 24202 3984
rect 24236 3950 24270 3984
rect 24304 3950 24338 3984
rect 24372 3950 24406 3984
rect 24440 3950 24474 3984
rect 24508 3950 24542 3984
rect 24576 3950 24610 3984
rect 24644 3950 24678 3984
rect 24712 3950 24746 3984
rect 24780 3950 24814 3984
rect 24848 3950 24882 3984
rect 24916 3950 24950 3984
rect 24984 3950 25018 3984
rect 25052 3950 25086 3984
rect 25120 3950 25154 3984
rect 25188 3950 25222 3984
rect 25256 3950 25290 3984
rect 25324 3950 25358 3984
rect 25392 3950 25426 3984
rect 25460 3950 25494 3984
rect 25528 3950 25562 3984
rect 25596 3950 25630 3984
rect 25664 3950 25698 3984
rect 25732 3950 25766 3984
rect 25800 3950 25834 3984
rect 25868 3950 25902 3984
rect 25936 3950 25970 3984
rect 26004 3950 26038 3984
rect 26072 3950 26106 3984
rect 26140 3950 26174 3984
rect 26208 3950 26242 3984
rect 26276 3950 26310 3984
rect 26344 3950 26378 3984
rect 26412 3950 26446 3984
rect 26480 3950 26514 3984
rect 26548 3950 26582 3984
rect 26616 3950 26650 3984
rect 26684 3950 26718 3984
rect 26752 3950 26786 3984
rect 26820 3950 26854 3984
rect 26888 3950 26922 3984
rect 26956 3950 26990 3984
rect 27024 3950 27058 3984
rect 27092 3950 27126 3984
rect 27160 3950 27194 3984
rect 27228 3950 27262 3984
rect 27296 3950 27330 3984
rect 27364 3950 27398 3984
rect 27432 3950 27466 3984
rect 27500 3950 27534 3984
rect 27568 3950 27602 3984
rect 27636 3950 27670 3984
rect 27704 3950 27738 3984
rect 27772 3950 27806 3984
rect 27840 3950 27874 3984
rect 27908 3950 27942 3984
rect 27976 3950 28000 3984
rect 6415 3910 28000 3950
rect 6415 3876 6473 3910
rect 6507 3876 6542 3910
rect 6576 3876 6611 3910
rect 6645 3876 6680 3910
rect 6714 3876 6749 3910
rect 6783 3876 6818 3910
rect 6852 3876 6887 3910
rect 6921 3876 6956 3910
rect 6990 3876 7025 3910
rect 7059 3876 7094 3910
rect 7128 3876 7163 3910
rect 7197 3876 7232 3910
rect 7266 3876 7301 3910
rect 7335 3876 7370 3910
rect 7404 3876 7439 3910
rect 7473 3876 7508 3910
rect 7542 3876 7577 3910
rect 7611 3876 7646 3910
rect 7680 3876 7715 3910
rect 7749 3876 7784 3910
rect 7818 3876 7853 3910
rect 7887 3876 7922 3910
rect 7956 3876 7991 3910
rect 8025 3876 8060 3910
rect 8094 3876 8129 3910
rect 8163 3876 8198 3910
rect 8232 3876 8267 3910
rect 8301 3876 8336 3910
rect 8370 3876 8405 3910
rect 8439 3876 8474 3910
rect 8508 3876 8543 3910
rect 8577 3876 8612 3910
rect 8646 3876 8681 3910
rect 8715 3876 8750 3910
rect 8784 3876 8819 3910
rect 8853 3876 8888 3910
rect 8922 3876 8957 3910
rect 8991 3876 9026 3910
rect 9060 3876 9095 3910
rect 9129 3876 9164 3910
rect 9198 3876 9233 3910
rect 9267 3876 9302 3910
rect 9336 3876 9371 3910
rect 9405 3876 9440 3910
rect 9474 3876 9509 3910
rect 9543 3876 9578 3910
rect 9612 3876 9647 3910
rect 9681 3876 9716 3910
rect 9750 3876 9785 3910
rect 9819 3876 9854 3910
rect 9888 3876 9922 3910
rect 9956 3876 9990 3910
rect 10024 3876 10058 3910
rect 10092 3876 10126 3910
rect 10160 3876 10194 3910
rect 10228 3876 10262 3910
rect 10296 3876 10330 3910
rect 10364 3876 10398 3910
rect 10432 3876 10466 3910
rect 10500 3876 10534 3910
rect 10568 3876 10602 3910
rect 10636 3876 10670 3910
rect 10704 3876 10738 3910
rect 10772 3876 10806 3910
rect 10840 3876 10874 3910
rect 10908 3876 10942 3910
rect 10976 3876 11010 3910
rect 11044 3876 11078 3910
rect 11112 3876 11146 3910
rect 11180 3876 11214 3910
rect 11248 3876 11282 3910
rect 11316 3876 11350 3910
rect 11384 3876 11418 3910
rect 11452 3876 11486 3910
rect 11520 3876 11554 3910
rect 11588 3876 11622 3910
rect 11656 3876 11690 3910
rect 11724 3876 11758 3910
rect 11792 3876 11826 3910
rect 11860 3876 11894 3910
rect 11928 3876 11962 3910
rect 11996 3876 12030 3910
rect 12064 3876 12098 3910
rect 12132 3876 12166 3910
rect 12200 3876 12234 3910
rect 12268 3876 12302 3910
rect 12336 3876 12370 3910
rect 12404 3876 12438 3910
rect 12472 3876 12506 3910
rect 12540 3876 12574 3910
rect 12608 3876 12642 3910
rect 12676 3876 12710 3910
rect 12744 3876 12778 3910
rect 12812 3876 12846 3910
rect 12880 3876 12914 3910
rect 12948 3876 12982 3910
rect 13016 3876 13050 3910
rect 13084 3876 13118 3910
rect 13152 3876 13186 3910
rect 13220 3876 13254 3910
rect 13288 3876 13322 3910
rect 13356 3876 13390 3910
rect 13424 3876 13458 3910
rect 13492 3876 13526 3910
rect 13560 3876 13594 3910
rect 13628 3876 13662 3910
rect 13696 3876 13730 3910
rect 13764 3876 13798 3910
rect 13832 3876 13866 3910
rect 13900 3876 13934 3910
rect 13968 3876 14002 3910
rect 14036 3876 14070 3910
rect 14104 3876 14138 3910
rect 14172 3876 14206 3910
rect 14240 3876 14274 3910
rect 14308 3876 14342 3910
rect 14376 3876 14410 3910
rect 14444 3876 14478 3910
rect 14512 3876 14546 3910
rect 14580 3876 14614 3910
rect 14648 3876 14682 3910
rect 14716 3876 14750 3910
rect 14784 3876 14818 3910
rect 14852 3876 14886 3910
rect 14920 3876 14954 3910
rect 14988 3876 15022 3910
rect 15056 3876 15090 3910
rect 15124 3876 15158 3910
rect 15192 3876 15226 3910
rect 15260 3876 15294 3910
rect 15328 3876 15362 3910
rect 15396 3876 15430 3910
rect 15464 3876 15498 3910
rect 15532 3876 15566 3910
rect 15600 3876 15634 3910
rect 15668 3876 15702 3910
rect 15736 3876 15770 3910
rect 15804 3876 15838 3910
rect 15872 3876 15906 3910
rect 15940 3876 15974 3910
rect 16008 3876 16042 3910
rect 16076 3876 16110 3910
rect 16144 3876 16178 3910
rect 16212 3876 16246 3910
rect 16280 3876 16314 3910
rect 16348 3876 16382 3910
rect 16416 3876 16450 3910
rect 16484 3876 16518 3910
rect 16552 3876 16586 3910
rect 16620 3876 16654 3910
rect 16688 3876 16722 3910
rect 16756 3876 16790 3910
rect 16824 3876 16858 3910
rect 16892 3876 16926 3910
rect 16960 3876 16994 3910
rect 17028 3876 17062 3910
rect 17096 3876 17130 3910
rect 17164 3876 17198 3910
rect 17232 3876 17266 3910
rect 17300 3876 17334 3910
rect 17368 3876 17402 3910
rect 17436 3876 17470 3910
rect 17504 3876 17538 3910
rect 17572 3876 17606 3910
rect 17640 3876 17674 3910
rect 17708 3876 17742 3910
rect 17776 3876 17810 3910
rect 17844 3876 17878 3910
rect 17912 3876 17946 3910
rect 17980 3876 18014 3910
rect 18048 3876 18082 3910
rect 18116 3876 18150 3910
rect 18184 3876 18218 3910
rect 18252 3876 18286 3910
rect 18320 3876 18354 3910
rect 18388 3876 18422 3910
rect 18456 3876 18490 3910
rect 18524 3876 18558 3910
rect 18592 3876 18626 3910
rect 18660 3876 18694 3910
rect 18728 3876 18762 3910
rect 18796 3876 18830 3910
rect 18864 3876 18898 3910
rect 18932 3876 18966 3910
rect 19000 3876 19034 3910
rect 19068 3876 19102 3910
rect 19136 3876 19170 3910
rect 19204 3876 19238 3910
rect 19272 3876 19306 3910
rect 19340 3876 19374 3910
rect 19408 3876 19442 3910
rect 19476 3876 19510 3910
rect 19544 3876 19578 3910
rect 19612 3876 19646 3910
rect 19680 3876 19714 3910
rect 19748 3876 19782 3910
rect 19816 3876 19850 3910
rect 19884 3876 19918 3910
rect 19952 3876 19986 3910
rect 20020 3876 20054 3910
rect 20088 3876 20122 3910
rect 20156 3876 20190 3910
rect 20224 3876 20258 3910
rect 20292 3876 20326 3910
rect 20360 3876 20394 3910
rect 20428 3876 20462 3910
rect 20496 3876 20530 3910
rect 20564 3876 20598 3910
rect 20632 3876 20666 3910
rect 20700 3876 20734 3910
rect 20768 3876 20802 3910
rect 20836 3876 20870 3910
rect 20904 3876 20938 3910
rect 20972 3876 21006 3910
rect 21040 3876 21074 3910
rect 21108 3876 21142 3910
rect 21176 3876 21210 3910
rect 21244 3876 21278 3910
rect 21312 3876 21346 3910
rect 21380 3876 21414 3910
rect 21448 3876 21482 3910
rect 21516 3876 21550 3910
rect 21584 3876 21618 3910
rect 21652 3876 21686 3910
rect 21720 3876 21754 3910
rect 21788 3876 21822 3910
rect 21856 3876 21890 3910
rect 21924 3876 21958 3910
rect 21992 3876 22026 3910
rect 22060 3876 22094 3910
rect 22128 3876 22162 3910
rect 22196 3876 22230 3910
rect 22264 3876 22298 3910
rect 22332 3876 22366 3910
rect 22400 3876 22434 3910
rect 22468 3876 22502 3910
rect 22536 3876 22570 3910
rect 22604 3876 22638 3910
rect 22672 3876 22706 3910
rect 22740 3876 22774 3910
rect 22808 3876 22842 3910
rect 22876 3876 22910 3910
rect 22944 3876 22978 3910
rect 23012 3876 23046 3910
rect 23080 3876 23114 3910
rect 23148 3876 23182 3910
rect 23216 3876 23250 3910
rect 23284 3876 23318 3910
rect 23352 3876 23386 3910
rect 23420 3876 23454 3910
rect 23488 3876 23522 3910
rect 23556 3876 23590 3910
rect 23624 3876 23658 3910
rect 23692 3876 23726 3910
rect 23760 3876 23794 3910
rect 23828 3876 23862 3910
rect 23896 3876 23930 3910
rect 23964 3876 23998 3910
rect 24032 3876 24066 3910
rect 24100 3876 24134 3910
rect 24168 3876 24202 3910
rect 24236 3876 24270 3910
rect 24304 3876 24338 3910
rect 24372 3876 24406 3910
rect 24440 3876 24474 3910
rect 24508 3876 24542 3910
rect 24576 3876 24610 3910
rect 24644 3876 24678 3910
rect 24712 3876 24746 3910
rect 24780 3876 24814 3910
rect 24848 3876 24882 3910
rect 24916 3876 24950 3910
rect 24984 3876 25018 3910
rect 25052 3876 25086 3910
rect 25120 3876 25154 3910
rect 25188 3876 25222 3910
rect 25256 3876 25290 3910
rect 25324 3876 25358 3910
rect 25392 3876 25426 3910
rect 25460 3876 25494 3910
rect 25528 3876 25562 3910
rect 25596 3876 25630 3910
rect 25664 3876 25698 3910
rect 25732 3876 25766 3910
rect 25800 3876 25834 3910
rect 25868 3876 25902 3910
rect 25936 3876 25970 3910
rect 26004 3876 26038 3910
rect 26072 3876 26106 3910
rect 26140 3876 26174 3910
rect 26208 3876 26242 3910
rect 26276 3876 26310 3910
rect 26344 3876 26378 3910
rect 26412 3876 26446 3910
rect 26480 3876 26514 3910
rect 26548 3876 26582 3910
rect 26616 3876 26650 3910
rect 26684 3876 26718 3910
rect 26752 3876 26786 3910
rect 26820 3876 26854 3910
rect 26888 3876 26922 3910
rect 26956 3876 26990 3910
rect 27024 3876 27058 3910
rect 27092 3876 27126 3910
rect 27160 3876 27194 3910
rect 27228 3876 27262 3910
rect 27296 3876 27330 3910
rect 27364 3876 27398 3910
rect 27432 3876 27466 3910
rect 27500 3876 27534 3910
rect 27568 3876 27602 3910
rect 27636 3876 27670 3910
rect 27704 3876 27738 3910
rect 27772 3876 27806 3910
rect 27840 3876 27874 3910
rect 27908 3876 27942 3910
rect 27976 3876 28000 3910
rect 6415 3836 28000 3876
rect 6415 3802 6473 3836
rect 6507 3802 6542 3836
rect 6576 3802 6611 3836
rect 6645 3802 6680 3836
rect 6714 3802 6749 3836
rect 6783 3802 6818 3836
rect 6852 3802 6887 3836
rect 6921 3802 6956 3836
rect 6990 3802 7025 3836
rect 7059 3802 7094 3836
rect 7128 3802 7163 3836
rect 7197 3802 7232 3836
rect 7266 3802 7301 3836
rect 7335 3802 7370 3836
rect 7404 3802 7439 3836
rect 7473 3802 7508 3836
rect 7542 3802 7577 3836
rect 7611 3802 7646 3836
rect 7680 3802 7715 3836
rect 7749 3802 7784 3836
rect 7818 3802 7853 3836
rect 7887 3802 7922 3836
rect 7956 3802 7991 3836
rect 8025 3802 8060 3836
rect 8094 3802 8129 3836
rect 8163 3802 8198 3836
rect 8232 3802 8267 3836
rect 8301 3802 8336 3836
rect 8370 3802 8405 3836
rect 8439 3802 8474 3836
rect 8508 3802 8543 3836
rect 8577 3802 8612 3836
rect 8646 3802 8681 3836
rect 8715 3802 8750 3836
rect 8784 3802 8819 3836
rect 8853 3802 8888 3836
rect 8922 3802 8957 3836
rect 8991 3802 9026 3836
rect 9060 3802 9095 3836
rect 9129 3802 9164 3836
rect 9198 3802 9233 3836
rect 9267 3802 9302 3836
rect 9336 3802 9371 3836
rect 9405 3802 9440 3836
rect 9474 3802 9509 3836
rect 9543 3802 9578 3836
rect 9612 3802 9647 3836
rect 9681 3802 9716 3836
rect 9750 3802 9785 3836
rect 9819 3802 9854 3836
rect 9888 3802 9922 3836
rect 9956 3802 9990 3836
rect 10024 3802 10058 3836
rect 10092 3802 10126 3836
rect 10160 3802 10194 3836
rect 10228 3802 10262 3836
rect 10296 3802 10330 3836
rect 10364 3802 10398 3836
rect 10432 3802 10466 3836
rect 10500 3802 10534 3836
rect 10568 3802 10602 3836
rect 10636 3802 10670 3836
rect 10704 3802 10738 3836
rect 10772 3802 10806 3836
rect 10840 3802 10874 3836
rect 10908 3802 10942 3836
rect 10976 3802 11010 3836
rect 11044 3802 11078 3836
rect 11112 3802 11146 3836
rect 11180 3802 11214 3836
rect 11248 3802 11282 3836
rect 11316 3802 11350 3836
rect 11384 3802 11418 3836
rect 11452 3802 11486 3836
rect 11520 3802 11554 3836
rect 11588 3802 11622 3836
rect 11656 3802 11690 3836
rect 11724 3802 11758 3836
rect 11792 3802 11826 3836
rect 11860 3802 11894 3836
rect 11928 3802 11962 3836
rect 11996 3802 12030 3836
rect 12064 3802 12098 3836
rect 12132 3802 12166 3836
rect 12200 3802 12234 3836
rect 12268 3802 12302 3836
rect 12336 3802 12370 3836
rect 12404 3802 12438 3836
rect 12472 3802 12506 3836
rect 12540 3802 12574 3836
rect 12608 3802 12642 3836
rect 12676 3802 12710 3836
rect 12744 3802 12778 3836
rect 12812 3802 12846 3836
rect 12880 3802 12914 3836
rect 12948 3802 12982 3836
rect 13016 3802 13050 3836
rect 13084 3802 13118 3836
rect 13152 3802 13186 3836
rect 13220 3802 13254 3836
rect 13288 3802 13322 3836
rect 13356 3802 13390 3836
rect 13424 3802 13458 3836
rect 13492 3802 13526 3836
rect 13560 3802 13594 3836
rect 13628 3802 13662 3836
rect 13696 3802 13730 3836
rect 13764 3802 13798 3836
rect 13832 3802 13866 3836
rect 13900 3802 13934 3836
rect 13968 3802 14002 3836
rect 14036 3802 14070 3836
rect 14104 3802 14138 3836
rect 14172 3802 14206 3836
rect 14240 3802 14274 3836
rect 14308 3802 14342 3836
rect 14376 3802 14410 3836
rect 14444 3802 14478 3836
rect 14512 3802 14546 3836
rect 14580 3802 14614 3836
rect 14648 3802 14682 3836
rect 14716 3802 14750 3836
rect 14784 3802 14818 3836
rect 14852 3802 14886 3836
rect 14920 3802 14954 3836
rect 14988 3802 15022 3836
rect 15056 3802 15090 3836
rect 15124 3802 15158 3836
rect 15192 3802 15226 3836
rect 15260 3802 15294 3836
rect 15328 3802 15362 3836
rect 15396 3802 15430 3836
rect 15464 3802 15498 3836
rect 15532 3802 15566 3836
rect 15600 3802 15634 3836
rect 15668 3802 15702 3836
rect 15736 3802 15770 3836
rect 15804 3802 15838 3836
rect 15872 3802 15906 3836
rect 15940 3802 15974 3836
rect 16008 3802 16042 3836
rect 16076 3802 16110 3836
rect 16144 3802 16178 3836
rect 16212 3802 16246 3836
rect 16280 3802 16314 3836
rect 16348 3802 16382 3836
rect 16416 3802 16450 3836
rect 16484 3802 16518 3836
rect 16552 3802 16586 3836
rect 16620 3802 16654 3836
rect 16688 3802 16722 3836
rect 16756 3802 16790 3836
rect 16824 3802 16858 3836
rect 16892 3802 16926 3836
rect 16960 3802 16994 3836
rect 17028 3802 17062 3836
rect 17096 3802 17130 3836
rect 17164 3802 17198 3836
rect 17232 3802 17266 3836
rect 17300 3802 17334 3836
rect 17368 3802 17402 3836
rect 17436 3802 17470 3836
rect 17504 3802 17538 3836
rect 17572 3802 17606 3836
rect 17640 3802 17674 3836
rect 17708 3802 17742 3836
rect 17776 3802 17810 3836
rect 17844 3802 17878 3836
rect 17912 3802 17946 3836
rect 17980 3802 18014 3836
rect 18048 3802 18082 3836
rect 18116 3802 18150 3836
rect 18184 3802 18218 3836
rect 18252 3802 18286 3836
rect 18320 3802 18354 3836
rect 18388 3802 18422 3836
rect 18456 3802 18490 3836
rect 18524 3802 18558 3836
rect 18592 3802 18626 3836
rect 18660 3802 18694 3836
rect 18728 3802 18762 3836
rect 18796 3802 18830 3836
rect 18864 3802 18898 3836
rect 18932 3802 18966 3836
rect 19000 3802 19034 3836
rect 19068 3802 19102 3836
rect 19136 3802 19170 3836
rect 19204 3802 19238 3836
rect 19272 3802 19306 3836
rect 19340 3802 19374 3836
rect 19408 3802 19442 3836
rect 19476 3802 19510 3836
rect 19544 3802 19578 3836
rect 19612 3802 19646 3836
rect 19680 3802 19714 3836
rect 19748 3802 19782 3836
rect 19816 3802 19850 3836
rect 19884 3802 19918 3836
rect 19952 3802 19986 3836
rect 20020 3802 20054 3836
rect 20088 3802 20122 3836
rect 20156 3802 20190 3836
rect 20224 3802 20258 3836
rect 20292 3802 20326 3836
rect 20360 3802 20394 3836
rect 20428 3802 20462 3836
rect 20496 3802 20530 3836
rect 20564 3802 20598 3836
rect 20632 3802 20666 3836
rect 20700 3802 20734 3836
rect 20768 3802 20802 3836
rect 20836 3802 20870 3836
rect 20904 3802 20938 3836
rect 20972 3802 21006 3836
rect 21040 3802 21074 3836
rect 21108 3802 21142 3836
rect 21176 3802 21210 3836
rect 21244 3802 21278 3836
rect 21312 3802 21346 3836
rect 21380 3802 21414 3836
rect 21448 3802 21482 3836
rect 21516 3802 21550 3836
rect 21584 3802 21618 3836
rect 21652 3802 21686 3836
rect 21720 3802 21754 3836
rect 21788 3802 21822 3836
rect 21856 3802 21890 3836
rect 21924 3802 21958 3836
rect 21992 3802 22026 3836
rect 22060 3802 22094 3836
rect 22128 3802 22162 3836
rect 22196 3802 22230 3836
rect 22264 3802 22298 3836
rect 22332 3802 22366 3836
rect 22400 3802 22434 3836
rect 22468 3802 22502 3836
rect 22536 3802 22570 3836
rect 22604 3802 22638 3836
rect 22672 3802 22706 3836
rect 22740 3802 22774 3836
rect 22808 3802 22842 3836
rect 22876 3802 22910 3836
rect 22944 3802 22978 3836
rect 23012 3802 23046 3836
rect 23080 3802 23114 3836
rect 23148 3802 23182 3836
rect 23216 3802 23250 3836
rect 23284 3802 23318 3836
rect 23352 3802 23386 3836
rect 23420 3802 23454 3836
rect 23488 3802 23522 3836
rect 23556 3802 23590 3836
rect 23624 3802 23658 3836
rect 23692 3802 23726 3836
rect 23760 3802 23794 3836
rect 23828 3802 23862 3836
rect 23896 3802 23930 3836
rect 23964 3802 23998 3836
rect 24032 3802 24066 3836
rect 24100 3802 24134 3836
rect 24168 3802 24202 3836
rect 24236 3802 24270 3836
rect 24304 3802 24338 3836
rect 24372 3802 24406 3836
rect 24440 3802 24474 3836
rect 24508 3802 24542 3836
rect 24576 3802 24610 3836
rect 24644 3802 24678 3836
rect 24712 3802 24746 3836
rect 24780 3802 24814 3836
rect 24848 3802 24882 3836
rect 24916 3802 24950 3836
rect 24984 3802 25018 3836
rect 25052 3802 25086 3836
rect 25120 3802 25154 3836
rect 25188 3802 25222 3836
rect 25256 3802 25290 3836
rect 25324 3802 25358 3836
rect 25392 3802 25426 3836
rect 25460 3802 25494 3836
rect 25528 3802 25562 3836
rect 25596 3802 25630 3836
rect 25664 3802 25698 3836
rect 25732 3802 25766 3836
rect 25800 3802 25834 3836
rect 25868 3802 25902 3836
rect 25936 3802 25970 3836
rect 26004 3802 26038 3836
rect 26072 3802 26106 3836
rect 26140 3802 26174 3836
rect 26208 3802 26242 3836
rect 26276 3802 26310 3836
rect 26344 3802 26378 3836
rect 26412 3802 26446 3836
rect 26480 3802 26514 3836
rect 26548 3802 26582 3836
rect 26616 3802 26650 3836
rect 26684 3802 26718 3836
rect 26752 3802 26786 3836
rect 26820 3802 26854 3836
rect 26888 3802 26922 3836
rect 26956 3802 26990 3836
rect 27024 3802 27058 3836
rect 27092 3802 27126 3836
rect 27160 3802 27194 3836
rect 27228 3802 27262 3836
rect 27296 3802 27330 3836
rect 27364 3802 27398 3836
rect 27432 3802 27466 3836
rect 27500 3802 27534 3836
rect 27568 3802 27602 3836
rect 27636 3802 27670 3836
rect 27704 3802 27738 3836
rect 27772 3802 27806 3836
rect 27840 3802 27874 3836
rect 27908 3802 27942 3836
rect 27976 3802 28000 3836
rect 6415 3762 28000 3802
rect 6415 3754 6473 3762
rect 3292 3728 3316 3754
rect 2320 3688 3316 3728
rect 2320 3654 2344 3688
rect 2378 3654 2415 3688
rect 2449 3654 2486 3688
rect 2520 3654 2557 3688
rect 2591 3654 2628 3688
rect 2662 3654 2698 3688
rect 2732 3654 2768 3688
rect 2802 3654 2838 3688
rect 2872 3654 2908 3688
rect 2942 3654 2978 3688
rect 3012 3654 3048 3688
rect 3082 3654 3118 3688
rect 3152 3654 3188 3688
rect 3222 3654 3258 3688
rect 3292 3654 3316 3688
rect 2320 3614 3316 3654
rect 2320 3580 2344 3614
rect 2378 3580 2415 3614
rect 2449 3580 2486 3614
rect 2520 3580 2557 3614
rect 2591 3580 2628 3614
rect 2662 3580 2698 3614
rect 2732 3580 2768 3614
rect 2802 3580 2838 3614
rect 2872 3580 2908 3614
rect 2942 3580 2978 3614
rect 3012 3580 3048 3614
rect 3082 3580 3118 3614
rect 3152 3580 3188 3614
rect 3222 3580 3258 3614
rect 3292 3580 3316 3614
rect 2320 3540 3316 3580
rect 2320 3506 2344 3540
rect 2378 3506 2415 3540
rect 2449 3506 2486 3540
rect 2520 3506 2557 3540
rect 2591 3506 2628 3540
rect 2662 3506 2698 3540
rect 2732 3506 2768 3540
rect 2802 3506 2838 3540
rect 2872 3506 2908 3540
rect 2942 3506 2978 3540
rect 3012 3506 3048 3540
rect 3082 3506 3118 3540
rect 3152 3506 3188 3540
rect 3222 3506 3258 3540
rect 3292 3506 3316 3540
rect 2320 3466 3316 3506
rect 2320 3432 2344 3466
rect 2378 3432 2415 3466
rect 2449 3432 2486 3466
rect 2520 3432 2557 3466
rect 2591 3432 2628 3466
rect 2662 3432 2698 3466
rect 2732 3432 2768 3466
rect 2802 3432 2838 3466
rect 2872 3432 2908 3466
rect 2942 3432 2978 3466
rect 3012 3432 3048 3466
rect 3082 3432 3118 3466
rect 3152 3432 3188 3466
rect 3222 3432 3258 3466
rect 3292 3432 3316 3466
rect 2320 3430 3316 3432
rect 6449 3728 6473 3754
rect 6507 3728 6542 3762
rect 6576 3728 6611 3762
rect 6645 3728 6680 3762
rect 6714 3728 6749 3762
rect 6783 3728 6818 3762
rect 6852 3728 6887 3762
rect 6921 3728 6956 3762
rect 6990 3728 7025 3762
rect 7059 3728 7094 3762
rect 7128 3728 7163 3762
rect 7197 3728 7232 3762
rect 7266 3728 7301 3762
rect 7335 3728 7370 3762
rect 7404 3728 7439 3762
rect 7473 3728 7508 3762
rect 7542 3728 7577 3762
rect 7611 3728 7646 3762
rect 7680 3728 7715 3762
rect 7749 3728 7784 3762
rect 7818 3728 7853 3762
rect 7887 3728 7922 3762
rect 7956 3728 7991 3762
rect 8025 3728 8060 3762
rect 8094 3728 8129 3762
rect 8163 3728 8198 3762
rect 8232 3728 8267 3762
rect 8301 3728 8336 3762
rect 8370 3728 8405 3762
rect 8439 3728 8474 3762
rect 8508 3728 8543 3762
rect 8577 3728 8612 3762
rect 8646 3728 8681 3762
rect 8715 3728 8750 3762
rect 8784 3728 8819 3762
rect 8853 3728 8888 3762
rect 8922 3728 8957 3762
rect 8991 3728 9026 3762
rect 9060 3728 9095 3762
rect 9129 3728 9164 3762
rect 9198 3728 9233 3762
rect 9267 3728 9302 3762
rect 9336 3728 9371 3762
rect 9405 3728 9440 3762
rect 9474 3728 9509 3762
rect 9543 3728 9578 3762
rect 9612 3728 9647 3762
rect 9681 3728 9716 3762
rect 9750 3728 9785 3762
rect 9819 3728 9854 3762
rect 9888 3728 9922 3762
rect 9956 3728 9990 3762
rect 10024 3728 10058 3762
rect 10092 3728 10126 3762
rect 10160 3728 10194 3762
rect 10228 3728 10262 3762
rect 10296 3728 10330 3762
rect 10364 3728 10398 3762
rect 10432 3728 10466 3762
rect 10500 3728 10534 3762
rect 10568 3728 10602 3762
rect 10636 3728 10670 3762
rect 10704 3728 10738 3762
rect 10772 3728 10806 3762
rect 10840 3728 10874 3762
rect 10908 3728 10942 3762
rect 10976 3728 11010 3762
rect 11044 3728 11078 3762
rect 11112 3728 11146 3762
rect 11180 3728 11214 3762
rect 11248 3728 11282 3762
rect 11316 3728 11350 3762
rect 11384 3728 11418 3762
rect 11452 3728 11486 3762
rect 11520 3728 11554 3762
rect 11588 3728 11622 3762
rect 11656 3728 11690 3762
rect 11724 3728 11758 3762
rect 11792 3728 11826 3762
rect 11860 3728 11894 3762
rect 11928 3728 11962 3762
rect 11996 3728 12030 3762
rect 12064 3728 12098 3762
rect 12132 3728 12166 3762
rect 12200 3728 12234 3762
rect 12268 3728 12302 3762
rect 12336 3728 12370 3762
rect 12404 3728 12438 3762
rect 12472 3728 12506 3762
rect 12540 3728 12574 3762
rect 12608 3728 12642 3762
rect 12676 3728 12710 3762
rect 12744 3728 12778 3762
rect 12812 3728 12846 3762
rect 12880 3728 12914 3762
rect 12948 3728 12982 3762
rect 13016 3728 13050 3762
rect 13084 3728 13118 3762
rect 13152 3728 13186 3762
rect 13220 3728 13254 3762
rect 13288 3728 13322 3762
rect 13356 3728 13390 3762
rect 13424 3728 13458 3762
rect 13492 3728 13526 3762
rect 13560 3728 13594 3762
rect 13628 3728 13662 3762
rect 13696 3728 13730 3762
rect 13764 3728 13798 3762
rect 13832 3728 13866 3762
rect 13900 3728 13934 3762
rect 13968 3728 14002 3762
rect 14036 3728 14070 3762
rect 14104 3728 14138 3762
rect 14172 3728 14206 3762
rect 14240 3728 14274 3762
rect 14308 3728 14342 3762
rect 14376 3728 14410 3762
rect 14444 3728 14478 3762
rect 14512 3728 14546 3762
rect 14580 3728 14614 3762
rect 14648 3728 14682 3762
rect 14716 3728 14750 3762
rect 14784 3728 14818 3762
rect 14852 3728 14886 3762
rect 14920 3728 14954 3762
rect 14988 3728 15022 3762
rect 15056 3728 15090 3762
rect 15124 3728 15158 3762
rect 15192 3728 15226 3762
rect 15260 3728 15294 3762
rect 15328 3728 15362 3762
rect 15396 3728 15430 3762
rect 15464 3728 15498 3762
rect 15532 3728 15566 3762
rect 15600 3728 15634 3762
rect 15668 3728 15702 3762
rect 15736 3728 15770 3762
rect 15804 3728 15838 3762
rect 15872 3728 15906 3762
rect 15940 3728 15974 3762
rect 16008 3728 16042 3762
rect 16076 3728 16110 3762
rect 16144 3728 16178 3762
rect 16212 3728 16246 3762
rect 16280 3728 16314 3762
rect 16348 3728 16382 3762
rect 16416 3728 16450 3762
rect 16484 3728 16518 3762
rect 16552 3728 16586 3762
rect 16620 3728 16654 3762
rect 16688 3728 16722 3762
rect 16756 3728 16790 3762
rect 16824 3728 16858 3762
rect 16892 3728 16926 3762
rect 16960 3728 16994 3762
rect 17028 3728 17062 3762
rect 17096 3728 17130 3762
rect 17164 3728 17198 3762
rect 17232 3728 17266 3762
rect 17300 3728 17334 3762
rect 17368 3728 17402 3762
rect 17436 3728 17470 3762
rect 17504 3728 17538 3762
rect 17572 3728 17606 3762
rect 17640 3728 17674 3762
rect 17708 3728 17742 3762
rect 17776 3728 17810 3762
rect 17844 3728 17878 3762
rect 17912 3728 17946 3762
rect 17980 3728 18014 3762
rect 18048 3728 18082 3762
rect 18116 3728 18150 3762
rect 18184 3728 18218 3762
rect 18252 3728 18286 3762
rect 18320 3728 18354 3762
rect 18388 3728 18422 3762
rect 18456 3728 18490 3762
rect 18524 3728 18558 3762
rect 18592 3728 18626 3762
rect 18660 3728 18694 3762
rect 18728 3728 18762 3762
rect 18796 3728 18830 3762
rect 18864 3728 18898 3762
rect 18932 3728 18966 3762
rect 19000 3728 19034 3762
rect 19068 3728 19102 3762
rect 19136 3728 19170 3762
rect 19204 3728 19238 3762
rect 19272 3728 19306 3762
rect 19340 3728 19374 3762
rect 19408 3728 19442 3762
rect 19476 3728 19510 3762
rect 19544 3728 19578 3762
rect 19612 3728 19646 3762
rect 19680 3728 19714 3762
rect 19748 3728 19782 3762
rect 19816 3728 19850 3762
rect 19884 3728 19918 3762
rect 19952 3728 19986 3762
rect 20020 3728 20054 3762
rect 20088 3728 20122 3762
rect 20156 3728 20190 3762
rect 20224 3728 20258 3762
rect 20292 3728 20326 3762
rect 20360 3728 20394 3762
rect 20428 3728 20462 3762
rect 20496 3728 20530 3762
rect 20564 3728 20598 3762
rect 20632 3728 20666 3762
rect 20700 3728 20734 3762
rect 20768 3728 20802 3762
rect 20836 3728 20870 3762
rect 20904 3728 20938 3762
rect 20972 3728 21006 3762
rect 21040 3728 21074 3762
rect 21108 3728 21142 3762
rect 21176 3728 21210 3762
rect 21244 3728 21278 3762
rect 21312 3728 21346 3762
rect 21380 3728 21414 3762
rect 21448 3728 21482 3762
rect 21516 3728 21550 3762
rect 21584 3728 21618 3762
rect 21652 3728 21686 3762
rect 21720 3728 21754 3762
rect 21788 3728 21822 3762
rect 21856 3728 21890 3762
rect 21924 3728 21958 3762
rect 21992 3728 22026 3762
rect 22060 3728 22094 3762
rect 22128 3728 22162 3762
rect 22196 3728 22230 3762
rect 22264 3728 22298 3762
rect 22332 3728 22366 3762
rect 22400 3728 22434 3762
rect 22468 3728 22502 3762
rect 22536 3728 22570 3762
rect 22604 3728 22638 3762
rect 22672 3728 22706 3762
rect 22740 3728 22774 3762
rect 22808 3728 22842 3762
rect 22876 3728 22910 3762
rect 22944 3728 22978 3762
rect 23012 3728 23046 3762
rect 23080 3728 23114 3762
rect 23148 3728 23182 3762
rect 23216 3728 23250 3762
rect 23284 3728 23318 3762
rect 23352 3728 23386 3762
rect 23420 3728 23454 3762
rect 23488 3728 23522 3762
rect 23556 3728 23590 3762
rect 23624 3728 23658 3762
rect 23692 3728 23726 3762
rect 23760 3728 23794 3762
rect 23828 3728 23862 3762
rect 23896 3728 23930 3762
rect 23964 3728 23998 3762
rect 24032 3728 24066 3762
rect 24100 3728 24134 3762
rect 24168 3728 24202 3762
rect 24236 3728 24270 3762
rect 24304 3728 24338 3762
rect 24372 3728 24406 3762
rect 24440 3728 24474 3762
rect 24508 3728 24542 3762
rect 24576 3728 24610 3762
rect 24644 3728 24678 3762
rect 24712 3728 24746 3762
rect 24780 3728 24814 3762
rect 24848 3728 24882 3762
rect 24916 3728 24950 3762
rect 24984 3728 25018 3762
rect 25052 3728 25086 3762
rect 25120 3728 25154 3762
rect 25188 3728 25222 3762
rect 25256 3728 25290 3762
rect 25324 3728 25358 3762
rect 25392 3728 25426 3762
rect 25460 3728 25494 3762
rect 25528 3728 25562 3762
rect 25596 3728 25630 3762
rect 25664 3728 25698 3762
rect 25732 3728 25766 3762
rect 25800 3728 25834 3762
rect 25868 3728 25902 3762
rect 25936 3728 25970 3762
rect 26004 3728 26038 3762
rect 26072 3728 26106 3762
rect 26140 3728 26174 3762
rect 26208 3728 26242 3762
rect 26276 3728 26310 3762
rect 26344 3728 26378 3762
rect 26412 3728 26446 3762
rect 26480 3728 26514 3762
rect 26548 3728 26582 3762
rect 26616 3728 26650 3762
rect 26684 3728 26718 3762
rect 26752 3728 26786 3762
rect 26820 3728 26854 3762
rect 26888 3728 26922 3762
rect 26956 3728 26990 3762
rect 27024 3728 27058 3762
rect 27092 3728 27126 3762
rect 27160 3728 27194 3762
rect 27228 3728 27262 3762
rect 27296 3728 27330 3762
rect 27364 3728 27398 3762
rect 27432 3728 27466 3762
rect 27500 3728 27534 3762
rect 27568 3728 27602 3762
rect 27636 3728 27670 3762
rect 27704 3728 27738 3762
rect 27772 3728 27806 3762
rect 27840 3728 27874 3762
rect 27908 3728 27942 3762
rect 27976 3728 28000 3762
rect 6449 3688 28000 3728
rect 6449 3654 6473 3688
rect 6507 3654 6542 3688
rect 6576 3654 6611 3688
rect 6645 3654 6680 3688
rect 6714 3654 6749 3688
rect 6783 3654 6818 3688
rect 6852 3654 6887 3688
rect 6921 3654 6956 3688
rect 6990 3654 7025 3688
rect 7059 3654 7094 3688
rect 7128 3654 7163 3688
rect 7197 3654 7232 3688
rect 7266 3654 7301 3688
rect 7335 3654 7370 3688
rect 7404 3654 7439 3688
rect 7473 3654 7508 3688
rect 7542 3654 7577 3688
rect 7611 3654 7646 3688
rect 7680 3654 7715 3688
rect 7749 3654 7784 3688
rect 7818 3654 7853 3688
rect 7887 3654 7922 3688
rect 7956 3654 7991 3688
rect 8025 3654 8060 3688
rect 8094 3654 8129 3688
rect 8163 3654 8198 3688
rect 8232 3654 8267 3688
rect 8301 3654 8336 3688
rect 8370 3654 8405 3688
rect 8439 3654 8474 3688
rect 8508 3654 8543 3688
rect 8577 3654 8612 3688
rect 8646 3654 8681 3688
rect 8715 3654 8750 3688
rect 8784 3654 8819 3688
rect 8853 3654 8888 3688
rect 8922 3654 8957 3688
rect 8991 3654 9026 3688
rect 9060 3654 9095 3688
rect 9129 3654 9164 3688
rect 9198 3654 9233 3688
rect 9267 3654 9302 3688
rect 9336 3654 9371 3688
rect 9405 3654 9440 3688
rect 9474 3654 9509 3688
rect 9543 3654 9578 3688
rect 9612 3654 9647 3688
rect 9681 3654 9716 3688
rect 9750 3654 9785 3688
rect 9819 3654 9854 3688
rect 9888 3654 9922 3688
rect 9956 3654 9990 3688
rect 10024 3654 10058 3688
rect 10092 3654 10126 3688
rect 10160 3654 10194 3688
rect 10228 3654 10262 3688
rect 10296 3654 10330 3688
rect 10364 3654 10398 3688
rect 10432 3654 10466 3688
rect 10500 3654 10534 3688
rect 10568 3654 10602 3688
rect 10636 3654 10670 3688
rect 10704 3654 10738 3688
rect 10772 3654 10806 3688
rect 10840 3654 10874 3688
rect 10908 3654 10942 3688
rect 10976 3654 11010 3688
rect 11044 3654 11078 3688
rect 11112 3654 11146 3688
rect 11180 3654 11214 3688
rect 11248 3654 11282 3688
rect 11316 3654 11350 3688
rect 11384 3654 11418 3688
rect 11452 3654 11486 3688
rect 11520 3654 11554 3688
rect 11588 3654 11622 3688
rect 11656 3654 11690 3688
rect 11724 3654 11758 3688
rect 11792 3654 11826 3688
rect 11860 3654 11894 3688
rect 11928 3654 11962 3688
rect 11996 3654 12030 3688
rect 12064 3654 12098 3688
rect 12132 3654 12166 3688
rect 12200 3654 12234 3688
rect 12268 3654 12302 3688
rect 12336 3654 12370 3688
rect 12404 3654 12438 3688
rect 12472 3654 12506 3688
rect 12540 3654 12574 3688
rect 12608 3654 12642 3688
rect 12676 3654 12710 3688
rect 12744 3654 12778 3688
rect 12812 3654 12846 3688
rect 12880 3654 12914 3688
rect 12948 3654 12982 3688
rect 13016 3654 13050 3688
rect 13084 3654 13118 3688
rect 13152 3654 13186 3688
rect 13220 3654 13254 3688
rect 13288 3654 13322 3688
rect 13356 3654 13390 3688
rect 13424 3654 13458 3688
rect 13492 3654 13526 3688
rect 13560 3654 13594 3688
rect 13628 3654 13662 3688
rect 13696 3654 13730 3688
rect 13764 3654 13798 3688
rect 13832 3654 13866 3688
rect 13900 3654 13934 3688
rect 13968 3654 14002 3688
rect 14036 3654 14070 3688
rect 14104 3654 14138 3688
rect 14172 3654 14206 3688
rect 14240 3654 14274 3688
rect 14308 3654 14342 3688
rect 14376 3654 14410 3688
rect 14444 3654 14478 3688
rect 14512 3654 14546 3688
rect 14580 3654 14614 3688
rect 14648 3654 14682 3688
rect 14716 3654 14750 3688
rect 14784 3654 14818 3688
rect 14852 3654 14886 3688
rect 14920 3654 14954 3688
rect 14988 3654 15022 3688
rect 15056 3654 15090 3688
rect 15124 3654 15158 3688
rect 15192 3654 15226 3688
rect 15260 3654 15294 3688
rect 15328 3654 15362 3688
rect 15396 3654 15430 3688
rect 15464 3654 15498 3688
rect 15532 3654 15566 3688
rect 15600 3654 15634 3688
rect 15668 3654 15702 3688
rect 15736 3654 15770 3688
rect 15804 3654 15838 3688
rect 15872 3654 15906 3688
rect 15940 3654 15974 3688
rect 16008 3654 16042 3688
rect 16076 3654 16110 3688
rect 16144 3654 16178 3688
rect 16212 3654 16246 3688
rect 16280 3654 16314 3688
rect 16348 3654 16382 3688
rect 16416 3654 16450 3688
rect 16484 3654 16518 3688
rect 16552 3654 16586 3688
rect 16620 3654 16654 3688
rect 16688 3654 16722 3688
rect 16756 3654 16790 3688
rect 16824 3654 16858 3688
rect 16892 3654 16926 3688
rect 16960 3654 16994 3688
rect 17028 3654 17062 3688
rect 17096 3654 17130 3688
rect 17164 3654 17198 3688
rect 17232 3654 17266 3688
rect 17300 3654 17334 3688
rect 17368 3654 17402 3688
rect 17436 3654 17470 3688
rect 17504 3654 17538 3688
rect 17572 3654 17606 3688
rect 17640 3654 17674 3688
rect 17708 3654 17742 3688
rect 17776 3654 17810 3688
rect 17844 3654 17878 3688
rect 17912 3654 17946 3688
rect 17980 3654 18014 3688
rect 18048 3654 18082 3688
rect 18116 3654 18150 3688
rect 18184 3654 18218 3688
rect 18252 3654 18286 3688
rect 18320 3654 18354 3688
rect 18388 3654 18422 3688
rect 18456 3654 18490 3688
rect 18524 3654 18558 3688
rect 18592 3654 18626 3688
rect 18660 3654 18694 3688
rect 18728 3654 18762 3688
rect 18796 3654 18830 3688
rect 18864 3654 18898 3688
rect 18932 3654 18966 3688
rect 19000 3654 19034 3688
rect 19068 3654 19102 3688
rect 19136 3654 19170 3688
rect 19204 3654 19238 3688
rect 19272 3654 19306 3688
rect 19340 3654 19374 3688
rect 19408 3654 19442 3688
rect 19476 3654 19510 3688
rect 19544 3654 19578 3688
rect 19612 3654 19646 3688
rect 19680 3654 19714 3688
rect 19748 3654 19782 3688
rect 19816 3654 19850 3688
rect 19884 3654 19918 3688
rect 19952 3654 19986 3688
rect 20020 3654 20054 3688
rect 20088 3654 20122 3688
rect 20156 3654 20190 3688
rect 20224 3654 20258 3688
rect 20292 3654 20326 3688
rect 20360 3654 20394 3688
rect 20428 3654 20462 3688
rect 20496 3654 20530 3688
rect 20564 3654 20598 3688
rect 20632 3654 20666 3688
rect 20700 3654 20734 3688
rect 20768 3654 20802 3688
rect 20836 3654 20870 3688
rect 20904 3654 20938 3688
rect 20972 3654 21006 3688
rect 21040 3654 21074 3688
rect 21108 3654 21142 3688
rect 21176 3654 21210 3688
rect 21244 3654 21278 3688
rect 21312 3654 21346 3688
rect 21380 3654 21414 3688
rect 21448 3654 21482 3688
rect 21516 3654 21550 3688
rect 21584 3654 21618 3688
rect 21652 3654 21686 3688
rect 21720 3654 21754 3688
rect 21788 3654 21822 3688
rect 21856 3654 21890 3688
rect 21924 3654 21958 3688
rect 21992 3654 22026 3688
rect 22060 3654 22094 3688
rect 22128 3654 22162 3688
rect 22196 3654 22230 3688
rect 22264 3654 22298 3688
rect 22332 3654 22366 3688
rect 22400 3654 22434 3688
rect 22468 3654 22502 3688
rect 22536 3654 22570 3688
rect 22604 3654 22638 3688
rect 22672 3654 22706 3688
rect 22740 3654 22774 3688
rect 22808 3654 22842 3688
rect 22876 3654 22910 3688
rect 22944 3654 22978 3688
rect 23012 3654 23046 3688
rect 23080 3654 23114 3688
rect 23148 3654 23182 3688
rect 23216 3654 23250 3688
rect 23284 3654 23318 3688
rect 23352 3654 23386 3688
rect 23420 3654 23454 3688
rect 23488 3654 23522 3688
rect 23556 3654 23590 3688
rect 23624 3654 23658 3688
rect 23692 3654 23726 3688
rect 23760 3654 23794 3688
rect 23828 3654 23862 3688
rect 23896 3654 23930 3688
rect 23964 3654 23998 3688
rect 24032 3654 24066 3688
rect 24100 3654 24134 3688
rect 24168 3654 24202 3688
rect 24236 3654 24270 3688
rect 24304 3654 24338 3688
rect 24372 3654 24406 3688
rect 24440 3654 24474 3688
rect 24508 3654 24542 3688
rect 24576 3654 24610 3688
rect 24644 3654 24678 3688
rect 24712 3654 24746 3688
rect 24780 3654 24814 3688
rect 24848 3654 24882 3688
rect 24916 3654 24950 3688
rect 24984 3654 25018 3688
rect 25052 3654 25086 3688
rect 25120 3654 25154 3688
rect 25188 3654 25222 3688
rect 25256 3654 25290 3688
rect 25324 3654 25358 3688
rect 25392 3654 25426 3688
rect 25460 3654 25494 3688
rect 25528 3654 25562 3688
rect 25596 3654 25630 3688
rect 25664 3654 25698 3688
rect 25732 3654 25766 3688
rect 25800 3654 25834 3688
rect 25868 3654 25902 3688
rect 25936 3654 25970 3688
rect 26004 3654 26038 3688
rect 26072 3654 26106 3688
rect 26140 3654 26174 3688
rect 26208 3654 26242 3688
rect 26276 3654 26310 3688
rect 26344 3654 26378 3688
rect 26412 3654 26446 3688
rect 26480 3654 26514 3688
rect 26548 3654 26582 3688
rect 26616 3654 26650 3688
rect 26684 3654 26718 3688
rect 26752 3654 26786 3688
rect 26820 3654 26854 3688
rect 26888 3654 26922 3688
rect 26956 3654 26990 3688
rect 27024 3654 27058 3688
rect 27092 3654 27126 3688
rect 27160 3654 27194 3688
rect 27228 3654 27262 3688
rect 27296 3654 27330 3688
rect 27364 3654 27398 3688
rect 27432 3654 27466 3688
rect 27500 3654 27534 3688
rect 27568 3654 27602 3688
rect 27636 3654 27670 3688
rect 27704 3654 27738 3688
rect 27772 3654 27806 3688
rect 27840 3654 27874 3688
rect 27908 3654 27942 3688
rect 27976 3654 28000 3688
rect 6449 3614 28000 3654
rect 6449 3580 6473 3614
rect 6507 3580 6542 3614
rect 6576 3580 6611 3614
rect 6645 3580 6680 3614
rect 6714 3580 6749 3614
rect 6783 3580 6818 3614
rect 6852 3580 6887 3614
rect 6921 3580 6956 3614
rect 6990 3580 7025 3614
rect 7059 3580 7094 3614
rect 7128 3580 7163 3614
rect 7197 3580 7232 3614
rect 7266 3580 7301 3614
rect 7335 3580 7370 3614
rect 7404 3580 7439 3614
rect 7473 3580 7508 3614
rect 7542 3580 7577 3614
rect 7611 3580 7646 3614
rect 7680 3580 7715 3614
rect 7749 3580 7784 3614
rect 7818 3580 7853 3614
rect 7887 3580 7922 3614
rect 7956 3580 7991 3614
rect 8025 3580 8060 3614
rect 8094 3580 8129 3614
rect 8163 3580 8198 3614
rect 8232 3580 8267 3614
rect 8301 3580 8336 3614
rect 8370 3580 8405 3614
rect 8439 3580 8474 3614
rect 8508 3580 8543 3614
rect 8577 3580 8612 3614
rect 8646 3580 8681 3614
rect 8715 3580 8750 3614
rect 8784 3580 8819 3614
rect 8853 3580 8888 3614
rect 8922 3580 8957 3614
rect 8991 3580 9026 3614
rect 9060 3580 9095 3614
rect 9129 3580 9164 3614
rect 9198 3580 9233 3614
rect 9267 3580 9302 3614
rect 9336 3580 9371 3614
rect 9405 3580 9440 3614
rect 9474 3580 9509 3614
rect 9543 3580 9578 3614
rect 9612 3580 9647 3614
rect 9681 3580 9716 3614
rect 9750 3580 9785 3614
rect 9819 3580 9854 3614
rect 9888 3580 9922 3614
rect 9956 3580 9990 3614
rect 10024 3580 10058 3614
rect 10092 3580 10126 3614
rect 10160 3580 10194 3614
rect 10228 3580 10262 3614
rect 10296 3580 10330 3614
rect 10364 3580 10398 3614
rect 10432 3580 10466 3614
rect 10500 3580 10534 3614
rect 10568 3580 10602 3614
rect 10636 3580 10670 3614
rect 10704 3580 10738 3614
rect 10772 3580 10806 3614
rect 10840 3580 10874 3614
rect 10908 3580 10942 3614
rect 10976 3580 11010 3614
rect 11044 3580 11078 3614
rect 11112 3580 11146 3614
rect 11180 3580 11214 3614
rect 11248 3580 11282 3614
rect 11316 3580 11350 3614
rect 11384 3580 11418 3614
rect 11452 3580 11486 3614
rect 11520 3580 11554 3614
rect 11588 3580 11622 3614
rect 11656 3580 11690 3614
rect 11724 3580 11758 3614
rect 11792 3580 11826 3614
rect 11860 3580 11894 3614
rect 11928 3580 11962 3614
rect 11996 3580 12030 3614
rect 12064 3580 12098 3614
rect 12132 3580 12166 3614
rect 12200 3580 12234 3614
rect 12268 3580 12302 3614
rect 12336 3580 12370 3614
rect 12404 3580 12438 3614
rect 12472 3580 12506 3614
rect 12540 3580 12574 3614
rect 12608 3580 12642 3614
rect 12676 3580 12710 3614
rect 12744 3580 12778 3614
rect 12812 3580 12846 3614
rect 12880 3580 12914 3614
rect 12948 3580 12982 3614
rect 13016 3580 13050 3614
rect 13084 3580 13118 3614
rect 13152 3580 13186 3614
rect 13220 3580 13254 3614
rect 13288 3580 13322 3614
rect 13356 3580 13390 3614
rect 13424 3580 13458 3614
rect 13492 3580 13526 3614
rect 13560 3580 13594 3614
rect 13628 3580 13662 3614
rect 13696 3580 13730 3614
rect 13764 3580 13798 3614
rect 13832 3580 13866 3614
rect 13900 3580 13934 3614
rect 13968 3580 14002 3614
rect 14036 3580 14070 3614
rect 14104 3580 14138 3614
rect 14172 3580 14206 3614
rect 14240 3580 14274 3614
rect 14308 3580 14342 3614
rect 14376 3580 14410 3614
rect 14444 3580 14478 3614
rect 14512 3580 14546 3614
rect 14580 3580 14614 3614
rect 14648 3580 14682 3614
rect 14716 3580 14750 3614
rect 14784 3580 14818 3614
rect 14852 3580 14886 3614
rect 14920 3580 14954 3614
rect 14988 3580 15022 3614
rect 15056 3580 15090 3614
rect 15124 3580 15158 3614
rect 15192 3580 15226 3614
rect 15260 3580 15294 3614
rect 15328 3580 15362 3614
rect 15396 3580 15430 3614
rect 15464 3580 15498 3614
rect 15532 3580 15566 3614
rect 15600 3580 15634 3614
rect 15668 3580 15702 3614
rect 15736 3580 15770 3614
rect 15804 3580 15838 3614
rect 15872 3580 15906 3614
rect 15940 3580 15974 3614
rect 16008 3580 16042 3614
rect 16076 3580 16110 3614
rect 16144 3580 16178 3614
rect 16212 3580 16246 3614
rect 16280 3580 16314 3614
rect 16348 3580 16382 3614
rect 16416 3580 16450 3614
rect 16484 3580 16518 3614
rect 16552 3580 16586 3614
rect 16620 3580 16654 3614
rect 16688 3580 16722 3614
rect 16756 3580 16790 3614
rect 16824 3580 16858 3614
rect 16892 3580 16926 3614
rect 16960 3580 16994 3614
rect 17028 3580 17062 3614
rect 17096 3580 17130 3614
rect 17164 3580 17198 3614
rect 17232 3580 17266 3614
rect 17300 3580 17334 3614
rect 17368 3580 17402 3614
rect 17436 3580 17470 3614
rect 17504 3580 17538 3614
rect 17572 3580 17606 3614
rect 17640 3580 17674 3614
rect 17708 3580 17742 3614
rect 17776 3580 17810 3614
rect 17844 3580 17878 3614
rect 17912 3580 17946 3614
rect 17980 3580 18014 3614
rect 18048 3580 18082 3614
rect 18116 3580 18150 3614
rect 18184 3580 18218 3614
rect 18252 3580 18286 3614
rect 18320 3580 18354 3614
rect 18388 3580 18422 3614
rect 18456 3580 18490 3614
rect 18524 3580 18558 3614
rect 18592 3580 18626 3614
rect 18660 3580 18694 3614
rect 18728 3580 18762 3614
rect 18796 3580 18830 3614
rect 18864 3580 18898 3614
rect 18932 3580 18966 3614
rect 19000 3580 19034 3614
rect 19068 3580 19102 3614
rect 19136 3580 19170 3614
rect 19204 3580 19238 3614
rect 19272 3580 19306 3614
rect 19340 3580 19374 3614
rect 19408 3580 19442 3614
rect 19476 3580 19510 3614
rect 19544 3580 19578 3614
rect 19612 3580 19646 3614
rect 19680 3580 19714 3614
rect 19748 3580 19782 3614
rect 19816 3580 19850 3614
rect 19884 3580 19918 3614
rect 19952 3580 19986 3614
rect 20020 3580 20054 3614
rect 20088 3580 20122 3614
rect 20156 3580 20190 3614
rect 20224 3580 20258 3614
rect 20292 3580 20326 3614
rect 20360 3580 20394 3614
rect 20428 3580 20462 3614
rect 20496 3580 20530 3614
rect 20564 3580 20598 3614
rect 20632 3580 20666 3614
rect 20700 3580 20734 3614
rect 20768 3580 20802 3614
rect 20836 3580 20870 3614
rect 20904 3580 20938 3614
rect 20972 3580 21006 3614
rect 21040 3580 21074 3614
rect 21108 3580 21142 3614
rect 21176 3580 21210 3614
rect 21244 3580 21278 3614
rect 21312 3580 21346 3614
rect 21380 3580 21414 3614
rect 21448 3580 21482 3614
rect 21516 3580 21550 3614
rect 21584 3580 21618 3614
rect 21652 3580 21686 3614
rect 21720 3580 21754 3614
rect 21788 3580 21822 3614
rect 21856 3580 21890 3614
rect 21924 3580 21958 3614
rect 21992 3580 22026 3614
rect 22060 3580 22094 3614
rect 22128 3580 22162 3614
rect 22196 3580 22230 3614
rect 22264 3580 22298 3614
rect 22332 3580 22366 3614
rect 22400 3580 22434 3614
rect 22468 3580 22502 3614
rect 22536 3580 22570 3614
rect 22604 3580 22638 3614
rect 22672 3580 22706 3614
rect 22740 3580 22774 3614
rect 22808 3580 22842 3614
rect 22876 3580 22910 3614
rect 22944 3580 22978 3614
rect 23012 3580 23046 3614
rect 23080 3580 23114 3614
rect 23148 3580 23182 3614
rect 23216 3580 23250 3614
rect 23284 3580 23318 3614
rect 23352 3580 23386 3614
rect 23420 3580 23454 3614
rect 23488 3580 23522 3614
rect 23556 3580 23590 3614
rect 23624 3580 23658 3614
rect 23692 3580 23726 3614
rect 23760 3580 23794 3614
rect 23828 3580 23862 3614
rect 23896 3580 23930 3614
rect 23964 3580 23998 3614
rect 24032 3580 24066 3614
rect 24100 3580 24134 3614
rect 24168 3580 24202 3614
rect 24236 3580 24270 3614
rect 24304 3580 24338 3614
rect 24372 3580 24406 3614
rect 24440 3580 24474 3614
rect 24508 3580 24542 3614
rect 24576 3580 24610 3614
rect 24644 3580 24678 3614
rect 24712 3580 24746 3614
rect 24780 3580 24814 3614
rect 24848 3580 24882 3614
rect 24916 3580 24950 3614
rect 24984 3580 25018 3614
rect 25052 3580 25086 3614
rect 25120 3580 25154 3614
rect 25188 3580 25222 3614
rect 25256 3580 25290 3614
rect 25324 3580 25358 3614
rect 25392 3580 25426 3614
rect 25460 3580 25494 3614
rect 25528 3580 25562 3614
rect 25596 3580 25630 3614
rect 25664 3580 25698 3614
rect 25732 3580 25766 3614
rect 25800 3580 25834 3614
rect 25868 3580 25902 3614
rect 25936 3580 25970 3614
rect 26004 3580 26038 3614
rect 26072 3580 26106 3614
rect 26140 3580 26174 3614
rect 26208 3580 26242 3614
rect 26276 3580 26310 3614
rect 26344 3580 26378 3614
rect 26412 3580 26446 3614
rect 26480 3580 26514 3614
rect 26548 3580 26582 3614
rect 26616 3580 26650 3614
rect 26684 3580 26718 3614
rect 26752 3580 26786 3614
rect 26820 3580 26854 3614
rect 26888 3580 26922 3614
rect 26956 3580 26990 3614
rect 27024 3580 27058 3614
rect 27092 3580 27126 3614
rect 27160 3580 27194 3614
rect 27228 3580 27262 3614
rect 27296 3580 27330 3614
rect 27364 3580 27398 3614
rect 27432 3580 27466 3614
rect 27500 3580 27534 3614
rect 27568 3580 27602 3614
rect 27636 3580 27670 3614
rect 27704 3580 27738 3614
rect 27772 3580 27806 3614
rect 27840 3580 27874 3614
rect 27908 3580 27942 3614
rect 27976 3580 28000 3614
rect 6449 3540 28000 3580
rect 6449 3506 6473 3540
rect 6507 3506 6542 3540
rect 6576 3506 6611 3540
rect 6645 3506 6680 3540
rect 6714 3506 6749 3540
rect 6783 3506 6818 3540
rect 6852 3506 6887 3540
rect 6921 3506 6956 3540
rect 6990 3506 7025 3540
rect 7059 3506 7094 3540
rect 7128 3506 7163 3540
rect 7197 3506 7232 3540
rect 7266 3506 7301 3540
rect 7335 3506 7370 3540
rect 7404 3506 7439 3540
rect 7473 3506 7508 3540
rect 7542 3506 7577 3540
rect 7611 3506 7646 3540
rect 7680 3506 7715 3540
rect 7749 3506 7784 3540
rect 7818 3506 7853 3540
rect 7887 3506 7922 3540
rect 7956 3506 7991 3540
rect 8025 3506 8060 3540
rect 8094 3506 8129 3540
rect 8163 3506 8198 3540
rect 8232 3506 8267 3540
rect 8301 3506 8336 3540
rect 8370 3506 8405 3540
rect 8439 3506 8474 3540
rect 8508 3506 8543 3540
rect 8577 3506 8612 3540
rect 8646 3506 8681 3540
rect 8715 3506 8750 3540
rect 8784 3506 8819 3540
rect 8853 3506 8888 3540
rect 8922 3506 8957 3540
rect 8991 3506 9026 3540
rect 9060 3506 9095 3540
rect 9129 3506 9164 3540
rect 9198 3506 9233 3540
rect 9267 3506 9302 3540
rect 9336 3506 9371 3540
rect 9405 3506 9440 3540
rect 9474 3506 9509 3540
rect 9543 3506 9578 3540
rect 9612 3506 9647 3540
rect 9681 3506 9716 3540
rect 9750 3506 9785 3540
rect 9819 3506 9854 3540
rect 9888 3506 9922 3540
rect 9956 3506 9990 3540
rect 10024 3506 10058 3540
rect 10092 3506 10126 3540
rect 10160 3506 10194 3540
rect 10228 3506 10262 3540
rect 10296 3506 10330 3540
rect 10364 3506 10398 3540
rect 10432 3506 10466 3540
rect 10500 3506 10534 3540
rect 10568 3506 10602 3540
rect 10636 3506 10670 3540
rect 10704 3506 10738 3540
rect 10772 3506 10806 3540
rect 10840 3506 10874 3540
rect 10908 3506 10942 3540
rect 10976 3506 11010 3540
rect 11044 3506 11078 3540
rect 11112 3506 11146 3540
rect 11180 3506 11214 3540
rect 11248 3506 11282 3540
rect 11316 3506 11350 3540
rect 11384 3506 11418 3540
rect 11452 3506 11486 3540
rect 11520 3506 11554 3540
rect 11588 3506 11622 3540
rect 11656 3506 11690 3540
rect 11724 3506 11758 3540
rect 11792 3506 11826 3540
rect 11860 3506 11894 3540
rect 11928 3506 11962 3540
rect 11996 3506 12030 3540
rect 12064 3506 12098 3540
rect 12132 3506 12166 3540
rect 12200 3506 12234 3540
rect 12268 3506 12302 3540
rect 12336 3506 12370 3540
rect 12404 3506 12438 3540
rect 12472 3506 12506 3540
rect 12540 3506 12574 3540
rect 12608 3506 12642 3540
rect 12676 3506 12710 3540
rect 12744 3506 12778 3540
rect 12812 3506 12846 3540
rect 12880 3506 12914 3540
rect 12948 3506 12982 3540
rect 13016 3506 13050 3540
rect 13084 3506 13118 3540
rect 13152 3506 13186 3540
rect 13220 3506 13254 3540
rect 13288 3506 13322 3540
rect 13356 3506 13390 3540
rect 13424 3506 13458 3540
rect 13492 3506 13526 3540
rect 13560 3506 13594 3540
rect 13628 3506 13662 3540
rect 13696 3506 13730 3540
rect 13764 3506 13798 3540
rect 13832 3506 13866 3540
rect 13900 3506 13934 3540
rect 13968 3506 14002 3540
rect 14036 3506 14070 3540
rect 14104 3506 14138 3540
rect 14172 3506 14206 3540
rect 14240 3506 14274 3540
rect 14308 3506 14342 3540
rect 14376 3506 14410 3540
rect 14444 3506 14478 3540
rect 14512 3506 14546 3540
rect 14580 3506 14614 3540
rect 14648 3506 14682 3540
rect 14716 3506 14750 3540
rect 14784 3506 14818 3540
rect 14852 3506 14886 3540
rect 14920 3506 14954 3540
rect 14988 3506 15022 3540
rect 15056 3506 15090 3540
rect 15124 3506 15158 3540
rect 15192 3506 15226 3540
rect 15260 3506 15294 3540
rect 15328 3506 15362 3540
rect 15396 3506 15430 3540
rect 15464 3506 15498 3540
rect 15532 3506 15566 3540
rect 15600 3506 15634 3540
rect 15668 3506 15702 3540
rect 15736 3506 15770 3540
rect 15804 3506 15838 3540
rect 15872 3506 15906 3540
rect 15940 3506 15974 3540
rect 16008 3506 16042 3540
rect 16076 3506 16110 3540
rect 16144 3506 16178 3540
rect 16212 3506 16246 3540
rect 16280 3506 16314 3540
rect 16348 3506 16382 3540
rect 16416 3506 16450 3540
rect 16484 3506 16518 3540
rect 16552 3506 16586 3540
rect 16620 3506 16654 3540
rect 16688 3506 16722 3540
rect 16756 3506 16790 3540
rect 16824 3506 16858 3540
rect 16892 3506 16926 3540
rect 16960 3506 16994 3540
rect 17028 3506 17062 3540
rect 17096 3506 17130 3540
rect 17164 3506 17198 3540
rect 17232 3506 17266 3540
rect 17300 3506 17334 3540
rect 17368 3506 17402 3540
rect 17436 3506 17470 3540
rect 17504 3506 17538 3540
rect 17572 3506 17606 3540
rect 17640 3506 17674 3540
rect 17708 3506 17742 3540
rect 17776 3506 17810 3540
rect 17844 3506 17878 3540
rect 17912 3506 17946 3540
rect 17980 3506 18014 3540
rect 18048 3506 18082 3540
rect 18116 3506 18150 3540
rect 18184 3506 18218 3540
rect 18252 3506 18286 3540
rect 18320 3506 18354 3540
rect 18388 3506 18422 3540
rect 18456 3506 18490 3540
rect 18524 3506 18558 3540
rect 18592 3506 18626 3540
rect 18660 3506 18694 3540
rect 18728 3506 18762 3540
rect 18796 3506 18830 3540
rect 18864 3506 18898 3540
rect 18932 3506 18966 3540
rect 19000 3506 19034 3540
rect 19068 3506 19102 3540
rect 19136 3506 19170 3540
rect 19204 3506 19238 3540
rect 19272 3506 19306 3540
rect 19340 3506 19374 3540
rect 19408 3506 19442 3540
rect 19476 3506 19510 3540
rect 19544 3506 19578 3540
rect 19612 3506 19646 3540
rect 19680 3506 19714 3540
rect 19748 3506 19782 3540
rect 19816 3506 19850 3540
rect 19884 3506 19918 3540
rect 19952 3506 19986 3540
rect 20020 3506 20054 3540
rect 20088 3506 20122 3540
rect 20156 3506 20190 3540
rect 20224 3506 20258 3540
rect 20292 3506 20326 3540
rect 20360 3506 20394 3540
rect 20428 3506 20462 3540
rect 20496 3506 20530 3540
rect 20564 3506 20598 3540
rect 20632 3506 20666 3540
rect 20700 3506 20734 3540
rect 20768 3506 20802 3540
rect 20836 3506 20870 3540
rect 20904 3506 20938 3540
rect 20972 3506 21006 3540
rect 21040 3506 21074 3540
rect 21108 3506 21142 3540
rect 21176 3506 21210 3540
rect 21244 3506 21278 3540
rect 21312 3506 21346 3540
rect 21380 3506 21414 3540
rect 21448 3506 21482 3540
rect 21516 3506 21550 3540
rect 21584 3506 21618 3540
rect 21652 3506 21686 3540
rect 21720 3506 21754 3540
rect 21788 3506 21822 3540
rect 21856 3506 21890 3540
rect 21924 3506 21958 3540
rect 21992 3506 22026 3540
rect 22060 3506 22094 3540
rect 22128 3506 22162 3540
rect 22196 3506 22230 3540
rect 22264 3506 22298 3540
rect 22332 3506 22366 3540
rect 22400 3506 22434 3540
rect 22468 3506 22502 3540
rect 22536 3506 22570 3540
rect 22604 3506 22638 3540
rect 22672 3506 22706 3540
rect 22740 3506 22774 3540
rect 22808 3506 22842 3540
rect 22876 3506 22910 3540
rect 22944 3506 22978 3540
rect 23012 3506 23046 3540
rect 23080 3506 23114 3540
rect 23148 3506 23182 3540
rect 23216 3506 23250 3540
rect 23284 3506 23318 3540
rect 23352 3506 23386 3540
rect 23420 3506 23454 3540
rect 23488 3506 23522 3540
rect 23556 3506 23590 3540
rect 23624 3506 23658 3540
rect 23692 3506 23726 3540
rect 23760 3506 23794 3540
rect 23828 3506 23862 3540
rect 23896 3506 23930 3540
rect 23964 3506 23998 3540
rect 24032 3506 24066 3540
rect 24100 3506 24134 3540
rect 24168 3506 24202 3540
rect 24236 3506 24270 3540
rect 24304 3506 24338 3540
rect 24372 3506 24406 3540
rect 24440 3506 24474 3540
rect 24508 3506 24542 3540
rect 24576 3506 24610 3540
rect 24644 3506 24678 3540
rect 24712 3506 24746 3540
rect 24780 3506 24814 3540
rect 24848 3506 24882 3540
rect 24916 3506 24950 3540
rect 24984 3506 25018 3540
rect 25052 3506 25086 3540
rect 25120 3506 25154 3540
rect 25188 3506 25222 3540
rect 25256 3506 25290 3540
rect 25324 3506 25358 3540
rect 25392 3506 25426 3540
rect 25460 3506 25494 3540
rect 25528 3506 25562 3540
rect 25596 3506 25630 3540
rect 25664 3506 25698 3540
rect 25732 3506 25766 3540
rect 25800 3506 25834 3540
rect 25868 3506 25902 3540
rect 25936 3506 25970 3540
rect 26004 3506 26038 3540
rect 26072 3506 26106 3540
rect 26140 3506 26174 3540
rect 26208 3506 26242 3540
rect 26276 3506 26310 3540
rect 26344 3506 26378 3540
rect 26412 3506 26446 3540
rect 26480 3506 26514 3540
rect 26548 3506 26582 3540
rect 26616 3506 26650 3540
rect 26684 3506 26718 3540
rect 26752 3506 26786 3540
rect 26820 3506 26854 3540
rect 26888 3506 26922 3540
rect 26956 3506 26990 3540
rect 27024 3506 27058 3540
rect 27092 3506 27126 3540
rect 27160 3506 27194 3540
rect 27228 3506 27262 3540
rect 27296 3506 27330 3540
rect 27364 3506 27398 3540
rect 27432 3506 27466 3540
rect 27500 3506 27534 3540
rect 27568 3506 27602 3540
rect 27636 3506 27670 3540
rect 27704 3506 27738 3540
rect 27772 3506 27806 3540
rect 27840 3506 27874 3540
rect 27908 3506 27942 3540
rect 27976 3506 28000 3540
rect 6449 3466 28000 3506
rect 6449 3432 6473 3466
rect 6507 3432 6542 3466
rect 6576 3432 6611 3466
rect 6645 3432 6680 3466
rect 6714 3432 6749 3466
rect 6783 3432 6818 3466
rect 6852 3432 6887 3466
rect 6921 3432 6956 3466
rect 6990 3432 7025 3466
rect 7059 3432 7094 3466
rect 7128 3432 7163 3466
rect 7197 3432 7232 3466
rect 7266 3432 7301 3466
rect 7335 3432 7370 3466
rect 7404 3432 7439 3466
rect 7473 3432 7508 3466
rect 7542 3432 7577 3466
rect 7611 3432 7646 3466
rect 7680 3432 7715 3466
rect 7749 3432 7784 3466
rect 7818 3432 7853 3466
rect 7887 3432 7922 3466
rect 7956 3432 7991 3466
rect 8025 3432 8060 3466
rect 8094 3432 8129 3466
rect 8163 3432 8198 3466
rect 8232 3432 8267 3466
rect 8301 3432 8336 3466
rect 8370 3432 8405 3466
rect 8439 3432 8474 3466
rect 8508 3432 8543 3466
rect 8577 3432 8612 3466
rect 8646 3432 8681 3466
rect 8715 3432 8750 3466
rect 8784 3432 8819 3466
rect 8853 3432 8888 3466
rect 8922 3432 8957 3466
rect 8991 3432 9026 3466
rect 9060 3432 9095 3466
rect 9129 3432 9164 3466
rect 9198 3432 9233 3466
rect 9267 3432 9302 3466
rect 9336 3432 9371 3466
rect 9405 3432 9440 3466
rect 9474 3432 9509 3466
rect 9543 3432 9578 3466
rect 9612 3432 9647 3466
rect 9681 3432 9716 3466
rect 9750 3432 9785 3466
rect 9819 3432 9854 3466
rect 9888 3432 9922 3466
rect 9956 3432 9990 3466
rect 10024 3432 10058 3466
rect 10092 3432 10126 3466
rect 10160 3432 10194 3466
rect 10228 3432 10262 3466
rect 10296 3432 10330 3466
rect 10364 3432 10398 3466
rect 10432 3432 10466 3466
rect 10500 3432 10534 3466
rect 10568 3432 10602 3466
rect 10636 3432 10670 3466
rect 10704 3432 10738 3466
rect 10772 3432 10806 3466
rect 10840 3432 10874 3466
rect 10908 3432 10942 3466
rect 10976 3432 11010 3466
rect 11044 3432 11078 3466
rect 11112 3432 11146 3466
rect 11180 3432 11214 3466
rect 11248 3432 11282 3466
rect 11316 3432 11350 3466
rect 11384 3432 11418 3466
rect 11452 3432 11486 3466
rect 11520 3432 11554 3466
rect 11588 3432 11622 3466
rect 11656 3432 11690 3466
rect 11724 3432 11758 3466
rect 11792 3432 11826 3466
rect 11860 3432 11894 3466
rect 11928 3432 11962 3466
rect 11996 3432 12030 3466
rect 12064 3432 12098 3466
rect 12132 3432 12166 3466
rect 12200 3432 12234 3466
rect 12268 3432 12302 3466
rect 12336 3432 12370 3466
rect 12404 3432 12438 3466
rect 12472 3432 12506 3466
rect 12540 3432 12574 3466
rect 12608 3432 12642 3466
rect 12676 3432 12710 3466
rect 12744 3432 12778 3466
rect 12812 3432 12846 3466
rect 12880 3432 12914 3466
rect 12948 3432 12982 3466
rect 13016 3432 13050 3466
rect 13084 3432 13118 3466
rect 13152 3432 13186 3466
rect 13220 3432 13254 3466
rect 13288 3432 13322 3466
rect 13356 3432 13390 3466
rect 13424 3432 13458 3466
rect 13492 3432 13526 3466
rect 13560 3432 13594 3466
rect 13628 3432 13662 3466
rect 13696 3432 13730 3466
rect 13764 3432 13798 3466
rect 13832 3432 13866 3466
rect 13900 3432 13934 3466
rect 13968 3432 14002 3466
rect 14036 3432 14070 3466
rect 14104 3432 14138 3466
rect 14172 3432 14206 3466
rect 14240 3432 14274 3466
rect 14308 3432 14342 3466
rect 14376 3432 14410 3466
rect 14444 3432 14478 3466
rect 14512 3432 14546 3466
rect 14580 3432 14614 3466
rect 14648 3432 14682 3466
rect 14716 3432 14750 3466
rect 14784 3432 14818 3466
rect 14852 3432 14886 3466
rect 14920 3432 14954 3466
rect 14988 3432 15022 3466
rect 15056 3432 15090 3466
rect 15124 3432 15158 3466
rect 15192 3432 15226 3466
rect 15260 3432 15294 3466
rect 15328 3432 15362 3466
rect 15396 3432 15430 3466
rect 15464 3432 15498 3466
rect 15532 3432 15566 3466
rect 15600 3432 15634 3466
rect 15668 3432 15702 3466
rect 15736 3432 15770 3466
rect 15804 3432 15838 3466
rect 15872 3432 15906 3466
rect 15940 3432 15974 3466
rect 16008 3432 16042 3466
rect 16076 3432 16110 3466
rect 16144 3432 16178 3466
rect 16212 3432 16246 3466
rect 16280 3432 16314 3466
rect 16348 3432 16382 3466
rect 16416 3432 16450 3466
rect 16484 3432 16518 3466
rect 16552 3432 16586 3466
rect 16620 3432 16654 3466
rect 16688 3432 16722 3466
rect 16756 3432 16790 3466
rect 16824 3432 16858 3466
rect 16892 3432 16926 3466
rect 16960 3432 16994 3466
rect 17028 3432 17062 3466
rect 17096 3432 17130 3466
rect 17164 3432 17198 3466
rect 17232 3432 17266 3466
rect 17300 3432 17334 3466
rect 17368 3432 17402 3466
rect 17436 3432 17470 3466
rect 17504 3432 17538 3466
rect 17572 3432 17606 3466
rect 17640 3432 17674 3466
rect 17708 3432 17742 3466
rect 17776 3432 17810 3466
rect 17844 3432 17878 3466
rect 17912 3432 17946 3466
rect 17980 3432 18014 3466
rect 18048 3432 18082 3466
rect 18116 3432 18150 3466
rect 18184 3432 18218 3466
rect 18252 3432 18286 3466
rect 18320 3432 18354 3466
rect 18388 3432 18422 3466
rect 18456 3432 18490 3466
rect 18524 3432 18558 3466
rect 18592 3432 18626 3466
rect 18660 3432 18694 3466
rect 18728 3432 18762 3466
rect 18796 3432 18830 3466
rect 18864 3432 18898 3466
rect 18932 3432 18966 3466
rect 19000 3432 19034 3466
rect 19068 3432 19102 3466
rect 19136 3432 19170 3466
rect 19204 3432 19238 3466
rect 19272 3432 19306 3466
rect 19340 3432 19374 3466
rect 19408 3432 19442 3466
rect 19476 3432 19510 3466
rect 19544 3432 19578 3466
rect 19612 3432 19646 3466
rect 19680 3432 19714 3466
rect 19748 3432 19782 3466
rect 19816 3432 19850 3466
rect 19884 3432 19918 3466
rect 19952 3432 19986 3466
rect 20020 3432 20054 3466
rect 20088 3432 20122 3466
rect 20156 3432 20190 3466
rect 20224 3432 20258 3466
rect 20292 3432 20326 3466
rect 20360 3432 20394 3466
rect 20428 3432 20462 3466
rect 20496 3432 20530 3466
rect 20564 3432 20598 3466
rect 20632 3432 20666 3466
rect 20700 3432 20734 3466
rect 20768 3432 20802 3466
rect 20836 3432 20870 3466
rect 20904 3432 20938 3466
rect 20972 3432 21006 3466
rect 21040 3432 21074 3466
rect 21108 3432 21142 3466
rect 21176 3432 21210 3466
rect 21244 3432 21278 3466
rect 21312 3432 21346 3466
rect 21380 3432 21414 3466
rect 21448 3432 21482 3466
rect 21516 3432 21550 3466
rect 21584 3432 21618 3466
rect 21652 3432 21686 3466
rect 21720 3432 21754 3466
rect 21788 3432 21822 3466
rect 21856 3432 21890 3466
rect 21924 3432 21958 3466
rect 21992 3432 22026 3466
rect 22060 3432 22094 3466
rect 22128 3432 22162 3466
rect 22196 3432 22230 3466
rect 22264 3432 22298 3466
rect 22332 3432 22366 3466
rect 22400 3432 22434 3466
rect 22468 3432 22502 3466
rect 22536 3432 22570 3466
rect 22604 3432 22638 3466
rect 22672 3432 22706 3466
rect 22740 3432 22774 3466
rect 22808 3432 22842 3466
rect 22876 3432 22910 3466
rect 22944 3432 22978 3466
rect 23012 3432 23046 3466
rect 23080 3432 23114 3466
rect 23148 3432 23182 3466
rect 23216 3432 23250 3466
rect 23284 3432 23318 3466
rect 23352 3432 23386 3466
rect 23420 3432 23454 3466
rect 23488 3432 23522 3466
rect 23556 3432 23590 3466
rect 23624 3432 23658 3466
rect 23692 3432 23726 3466
rect 23760 3432 23794 3466
rect 23828 3432 23862 3466
rect 23896 3432 23930 3466
rect 23964 3432 23998 3466
rect 24032 3432 24066 3466
rect 24100 3432 24134 3466
rect 24168 3432 24202 3466
rect 24236 3432 24270 3466
rect 24304 3432 24338 3466
rect 24372 3432 24406 3466
rect 24440 3432 24474 3466
rect 24508 3432 24542 3466
rect 24576 3432 24610 3466
rect 24644 3432 24678 3466
rect 24712 3432 24746 3466
rect 24780 3432 24814 3466
rect 24848 3432 24882 3466
rect 24916 3432 24950 3466
rect 24984 3432 25018 3466
rect 25052 3432 25086 3466
rect 25120 3432 25154 3466
rect 25188 3432 25222 3466
rect 25256 3432 25290 3466
rect 25324 3432 25358 3466
rect 25392 3432 25426 3466
rect 25460 3432 25494 3466
rect 25528 3432 25562 3466
rect 25596 3432 25630 3466
rect 25664 3432 25698 3466
rect 25732 3432 25766 3466
rect 25800 3432 25834 3466
rect 25868 3432 25902 3466
rect 25936 3432 25970 3466
rect 26004 3432 26038 3466
rect 26072 3432 26106 3466
rect 26140 3432 26174 3466
rect 26208 3432 26242 3466
rect 26276 3432 26310 3466
rect 26344 3432 26378 3466
rect 26412 3432 26446 3466
rect 26480 3432 26514 3466
rect 26548 3432 26582 3466
rect 26616 3432 26650 3466
rect 26684 3432 26718 3466
rect 26752 3432 26786 3466
rect 26820 3432 26854 3466
rect 26888 3432 26922 3466
rect 26956 3432 26990 3466
rect 27024 3432 27058 3466
rect 27092 3432 27126 3466
rect 27160 3432 27194 3466
rect 27228 3432 27262 3466
rect 27296 3432 27330 3466
rect 27364 3432 27398 3466
rect 27432 3432 27466 3466
rect 27500 3432 27534 3466
rect 27568 3432 27602 3466
rect 27636 3432 27670 3466
rect 27704 3432 27738 3466
rect 27772 3432 27806 3466
rect 27840 3432 27874 3466
rect 27908 3432 27942 3466
rect 27976 3432 28000 3466
rect 6449 3430 28000 3432
<< mvpsubdiff >>
rect 23687 23319 23747 23353
rect 23781 23319 23816 23353
rect 23850 23319 23885 23353
rect 23919 23319 23954 23353
rect 23988 23319 24023 23353
rect 24057 23319 24092 23353
rect 24126 23319 24161 23353
rect 24195 23319 24230 23353
rect 24264 23319 24299 23353
rect 24333 23319 24368 23353
rect 24402 23319 24437 23353
rect 24471 23319 24506 23353
rect 24540 23319 24575 23353
rect 24609 23319 24644 23353
rect 24678 23319 24713 23353
rect 24747 23319 24782 23353
rect 24816 23319 24851 23353
rect 24885 23319 24920 23353
rect 24954 23319 24989 23353
rect 25023 23319 25058 23353
rect 25092 23319 25127 23353
rect 25161 23319 25196 23353
rect 25230 23319 25265 23353
rect 25299 23319 25334 23353
rect 25368 23319 25403 23353
rect 25437 23319 25472 23353
rect 25506 23319 25541 23353
rect 25575 23319 25610 23353
rect 25644 23319 25679 23353
rect 25713 23319 25748 23353
rect 25782 23319 25817 23353
rect 25851 23319 25886 23353
rect 25920 23319 25955 23353
rect 25989 23319 26024 23353
rect 26058 23319 26093 23353
rect 26127 23319 26162 23353
rect 26196 23319 26231 23353
rect 26265 23319 26300 23353
rect 26334 23319 26368 23353
rect 26402 23319 26436 23353
rect 26470 23319 26504 23353
rect 26538 23319 26572 23353
rect 26606 23319 26640 23353
rect 26674 23319 26708 23353
rect 26742 23319 26776 23353
rect 26810 23319 26844 23353
rect 26878 23319 26912 23353
rect 26946 23319 26980 23353
rect 27014 23319 27048 23353
rect 27082 23319 27116 23353
rect 27150 23319 27184 23353
rect 27218 23319 27252 23353
rect 27286 23319 27320 23353
rect 27354 23319 27388 23353
rect 27422 23319 27456 23353
rect 27490 23319 27524 23353
rect 27558 23319 27592 23353
rect 27626 23319 27660 23353
rect 27694 23319 27728 23353
rect 27762 23319 27796 23353
rect 27830 23319 27864 23353
rect 27898 23319 27932 23353
rect 27966 23319 28000 23353
rect 23687 23283 28000 23319
rect 23687 23249 23747 23283
rect 23781 23249 23816 23283
rect 23850 23249 23885 23283
rect 23919 23249 23954 23283
rect 23988 23249 24023 23283
rect 24057 23249 24092 23283
rect 24126 23249 24161 23283
rect 24195 23249 24230 23283
rect 24264 23249 24299 23283
rect 24333 23249 24368 23283
rect 24402 23249 24437 23283
rect 24471 23249 24506 23283
rect 24540 23249 24575 23283
rect 24609 23249 24644 23283
rect 24678 23249 24713 23283
rect 24747 23249 24782 23283
rect 24816 23249 24851 23283
rect 24885 23249 24920 23283
rect 24954 23249 24989 23283
rect 25023 23249 25058 23283
rect 25092 23249 25127 23283
rect 25161 23249 25196 23283
rect 25230 23249 25265 23283
rect 25299 23249 25334 23283
rect 25368 23249 25403 23283
rect 25437 23249 25472 23283
rect 25506 23249 25541 23283
rect 25575 23249 25610 23283
rect 25644 23249 25679 23283
rect 25713 23249 25748 23283
rect 25782 23249 25817 23283
rect 25851 23249 25886 23283
rect 25920 23249 25955 23283
rect 25989 23249 26024 23283
rect 26058 23249 26093 23283
rect 26127 23249 26162 23283
rect 26196 23249 26231 23283
rect 26265 23249 26300 23283
rect 26334 23249 26368 23283
rect 26402 23249 26436 23283
rect 26470 23249 26504 23283
rect 26538 23249 26572 23283
rect 26606 23249 26640 23283
rect 26674 23249 26708 23283
rect 26742 23249 26776 23283
rect 26810 23249 26844 23283
rect 26878 23249 26912 23283
rect 26946 23249 26980 23283
rect 27014 23249 27048 23283
rect 27082 23249 27116 23283
rect 27150 23249 27184 23283
rect 27218 23249 27252 23283
rect 27286 23249 27320 23283
rect 27354 23249 27388 23283
rect 27422 23249 27456 23283
rect 27490 23249 27524 23283
rect 27558 23249 27592 23283
rect 27626 23249 27660 23283
rect 27694 23249 27728 23283
rect 27762 23249 27796 23283
rect 27830 23249 27864 23283
rect 27898 23249 27932 23283
rect 27966 23249 28000 23283
rect 23687 23213 28000 23249
rect 23687 23179 23747 23213
rect 23781 23179 23816 23213
rect 23850 23179 23885 23213
rect 23919 23179 23954 23213
rect 23988 23179 24023 23213
rect 24057 23179 24092 23213
rect 24126 23179 24161 23213
rect 24195 23179 24230 23213
rect 24264 23179 24299 23213
rect 24333 23179 24368 23213
rect 24402 23179 24437 23213
rect 24471 23179 24506 23213
rect 24540 23179 24575 23213
rect 24609 23179 24644 23213
rect 24678 23179 24713 23213
rect 24747 23179 24782 23213
rect 24816 23179 24851 23213
rect 24885 23179 24920 23213
rect 24954 23179 24989 23213
rect 25023 23179 25058 23213
rect 25092 23179 25127 23213
rect 25161 23179 25196 23213
rect 25230 23179 25265 23213
rect 25299 23179 25334 23213
rect 25368 23179 25403 23213
rect 25437 23179 25472 23213
rect 25506 23179 25541 23213
rect 25575 23179 25610 23213
rect 25644 23179 25679 23213
rect 25713 23179 25748 23213
rect 25782 23179 25817 23213
rect 25851 23179 25886 23213
rect 25920 23179 25955 23213
rect 25989 23179 26024 23213
rect 26058 23179 26093 23213
rect 26127 23179 26162 23213
rect 26196 23179 26231 23213
rect 26265 23179 26300 23213
rect 26334 23179 26368 23213
rect 26402 23179 26436 23213
rect 26470 23179 26504 23213
rect 26538 23179 26572 23213
rect 26606 23179 26640 23213
rect 26674 23179 26708 23213
rect 26742 23179 26776 23213
rect 26810 23179 26844 23213
rect 26878 23179 26912 23213
rect 26946 23179 26980 23213
rect 27014 23179 27048 23213
rect 27082 23179 27116 23213
rect 27150 23179 27184 23213
rect 27218 23179 27252 23213
rect 27286 23179 27320 23213
rect 27354 23179 27388 23213
rect 27422 23179 27456 23213
rect 27490 23179 27524 23213
rect 27558 23179 27592 23213
rect 27626 23179 27660 23213
rect 27694 23179 27728 23213
rect 27762 23179 27796 23213
rect 27830 23179 27864 23213
rect 27898 23179 27932 23213
rect 27966 23179 28000 23213
rect 23687 23143 28000 23179
rect 23687 23109 23747 23143
rect 23781 23109 23816 23143
rect 23850 23109 23885 23143
rect 23919 23109 23954 23143
rect 23988 23109 24023 23143
rect 24057 23109 24092 23143
rect 24126 23109 24161 23143
rect 24195 23109 24230 23143
rect 24264 23109 24299 23143
rect 24333 23109 24368 23143
rect 24402 23109 24437 23143
rect 24471 23109 24506 23143
rect 24540 23109 24575 23143
rect 24609 23109 24644 23143
rect 24678 23109 24713 23143
rect 24747 23109 24782 23143
rect 24816 23109 24851 23143
rect 24885 23109 24920 23143
rect 24954 23109 24989 23143
rect 25023 23109 25058 23143
rect 25092 23109 25127 23143
rect 25161 23109 25196 23143
rect 25230 23109 25265 23143
rect 25299 23109 25334 23143
rect 25368 23109 25403 23143
rect 25437 23109 25472 23143
rect 25506 23109 25541 23143
rect 25575 23109 25610 23143
rect 25644 23109 25679 23143
rect 25713 23109 25748 23143
rect 25782 23109 25817 23143
rect 25851 23109 25886 23143
rect 25920 23109 25955 23143
rect 25989 23109 26024 23143
rect 26058 23109 26093 23143
rect 26127 23109 26162 23143
rect 26196 23109 26231 23143
rect 26265 23109 26300 23143
rect 26334 23109 26368 23143
rect 26402 23109 26436 23143
rect 26470 23109 26504 23143
rect 26538 23109 26572 23143
rect 26606 23109 26640 23143
rect 26674 23109 26708 23143
rect 26742 23109 26776 23143
rect 26810 23109 26844 23143
rect 26878 23109 26912 23143
rect 26946 23109 26980 23143
rect 27014 23109 27048 23143
rect 27082 23109 27116 23143
rect 27150 23109 27184 23143
rect 27218 23109 27252 23143
rect 27286 23109 27320 23143
rect 27354 23109 27388 23143
rect 27422 23109 27456 23143
rect 27490 23109 27524 23143
rect 27558 23109 27592 23143
rect 27626 23109 27660 23143
rect 27694 23109 27728 23143
rect 27762 23109 27796 23143
rect 27830 23109 27864 23143
rect 27898 23109 27932 23143
rect 27966 23109 28000 23143
rect 23687 23073 28000 23109
rect 23687 23039 23747 23073
rect 23781 23039 23816 23073
rect 23850 23039 23885 23073
rect 23919 23039 23954 23073
rect 23988 23039 24023 23073
rect 24057 23039 24092 23073
rect 24126 23039 24161 23073
rect 24195 23039 24230 23073
rect 24264 23039 24299 23073
rect 24333 23039 24368 23073
rect 24402 23039 24437 23073
rect 24471 23039 24506 23073
rect 24540 23039 24575 23073
rect 24609 23039 24644 23073
rect 24678 23039 24713 23073
rect 24747 23039 24782 23073
rect 24816 23039 24851 23073
rect 24885 23039 24920 23073
rect 24954 23039 24989 23073
rect 25023 23039 25058 23073
rect 25092 23039 25127 23073
rect 25161 23039 25196 23073
rect 25230 23039 25265 23073
rect 25299 23039 25334 23073
rect 25368 23039 25403 23073
rect 25437 23039 25472 23073
rect 25506 23039 25541 23073
rect 25575 23039 25610 23073
rect 25644 23039 25679 23073
rect 25713 23039 25748 23073
rect 25782 23039 25817 23073
rect 25851 23039 25886 23073
rect 25920 23039 25955 23073
rect 25989 23039 26024 23073
rect 26058 23039 26093 23073
rect 26127 23039 26162 23073
rect 26196 23039 26231 23073
rect 26265 23039 26300 23073
rect 26334 23039 26368 23073
rect 26402 23039 26436 23073
rect 26470 23039 26504 23073
rect 26538 23039 26572 23073
rect 26606 23039 26640 23073
rect 26674 23039 26708 23073
rect 26742 23039 26776 23073
rect 26810 23039 26844 23073
rect 26878 23039 26912 23073
rect 26946 23039 26980 23073
rect 27014 23039 27048 23073
rect 27082 23039 27116 23073
rect 27150 23039 27184 23073
rect 27218 23039 27252 23073
rect 27286 23039 27320 23073
rect 27354 23039 27388 23073
rect 27422 23039 27456 23073
rect 27490 23039 27524 23073
rect 27558 23039 27592 23073
rect 27626 23039 27660 23073
rect 27694 23039 27728 23073
rect 27762 23039 27796 23073
rect 27830 23039 27864 23073
rect 27898 23039 27932 23073
rect 27966 23039 28000 23073
rect 23687 23003 28000 23039
rect 23687 22969 23747 23003
rect 23781 22969 23816 23003
rect 23850 22969 23885 23003
rect 23919 22969 23954 23003
rect 23988 22969 24023 23003
rect 24057 22969 24092 23003
rect 24126 22969 24161 23003
rect 24195 22969 24230 23003
rect 24264 22969 24299 23003
rect 24333 22969 24368 23003
rect 24402 22969 24437 23003
rect 24471 22969 24506 23003
rect 24540 22969 24575 23003
rect 24609 22969 24644 23003
rect 24678 22969 24713 23003
rect 24747 22969 24782 23003
rect 24816 22969 24851 23003
rect 24885 22969 24920 23003
rect 24954 22969 24989 23003
rect 25023 22969 25058 23003
rect 25092 22969 25127 23003
rect 25161 22969 25196 23003
rect 25230 22969 25265 23003
rect 25299 22969 25334 23003
rect 25368 22969 25403 23003
rect 25437 22969 25472 23003
rect 25506 22969 25541 23003
rect 25575 22969 25610 23003
rect 25644 22969 25679 23003
rect 25713 22969 25748 23003
rect 25782 22969 25817 23003
rect 25851 22969 25886 23003
rect 25920 22969 25955 23003
rect 25989 22969 26024 23003
rect 26058 22969 26093 23003
rect 26127 22969 26162 23003
rect 26196 22969 26231 23003
rect 26265 22969 26300 23003
rect 26334 22969 26368 23003
rect 26402 22969 26436 23003
rect 26470 22969 26504 23003
rect 26538 22969 26572 23003
rect 26606 22969 26640 23003
rect 26674 22969 26708 23003
rect 26742 22969 26776 23003
rect 26810 22969 26844 23003
rect 26878 22969 26912 23003
rect 26946 22969 26980 23003
rect 27014 22969 27048 23003
rect 27082 22969 27116 23003
rect 27150 22969 27184 23003
rect 27218 22969 27252 23003
rect 27286 22969 27320 23003
rect 27354 22969 27388 23003
rect 27422 22969 27456 23003
rect 27490 22969 27524 23003
rect 27558 22969 27592 23003
rect 27626 22969 27660 23003
rect 27694 22969 27728 23003
rect 27762 22969 27796 23003
rect 27830 22969 27864 23003
rect 27898 22969 27932 23003
rect 27966 22969 28000 23003
rect 23687 22933 28000 22969
rect 23687 22899 23747 22933
rect 23781 22899 23816 22933
rect 23850 22899 23885 22933
rect 23919 22899 23954 22933
rect 23988 22899 24023 22933
rect 24057 22899 24092 22933
rect 24126 22899 24161 22933
rect 24195 22899 24230 22933
rect 24264 22899 24299 22933
rect 24333 22899 24368 22933
rect 24402 22899 24437 22933
rect 24471 22899 24506 22933
rect 24540 22899 24575 22933
rect 24609 22899 24644 22933
rect 24678 22899 24713 22933
rect 24747 22899 24782 22933
rect 24816 22899 24851 22933
rect 24885 22899 24920 22933
rect 24954 22899 24989 22933
rect 25023 22899 25058 22933
rect 25092 22899 25127 22933
rect 25161 22899 25196 22933
rect 25230 22899 25265 22933
rect 25299 22899 25334 22933
rect 25368 22899 25403 22933
rect 25437 22899 25472 22933
rect 25506 22899 25541 22933
rect 25575 22899 25610 22933
rect 25644 22899 25679 22933
rect 25713 22899 25748 22933
rect 25782 22899 25817 22933
rect 25851 22899 25886 22933
rect 25920 22899 25955 22933
rect 25989 22899 26024 22933
rect 26058 22899 26093 22933
rect 26127 22899 26162 22933
rect 26196 22899 26231 22933
rect 26265 22899 26300 22933
rect 26334 22899 26368 22933
rect 26402 22899 26436 22933
rect 26470 22899 26504 22933
rect 26538 22899 26572 22933
rect 26606 22899 26640 22933
rect 26674 22899 26708 22933
rect 26742 22899 26776 22933
rect 26810 22899 26844 22933
rect 26878 22899 26912 22933
rect 26946 22899 26980 22933
rect 27014 22899 27048 22933
rect 27082 22899 27116 22933
rect 27150 22899 27184 22933
rect 27218 22899 27252 22933
rect 27286 22899 27320 22933
rect 27354 22899 27388 22933
rect 27422 22899 27456 22933
rect 27490 22899 27524 22933
rect 27558 22899 27592 22933
rect 27626 22899 27660 22933
rect 27694 22899 27728 22933
rect 27762 22899 27796 22933
rect 27830 22899 27864 22933
rect 27898 22899 27932 22933
rect 27966 22899 28000 22933
rect 26275 22856 28000 22899
rect 26275 22822 26309 22856
rect 26343 22822 26380 22856
rect 26414 22822 26451 22856
rect 26485 22822 26522 22856
rect 26556 22822 26593 22856
rect 26627 22822 26664 22856
rect 26698 22822 26735 22856
rect 26769 22822 26806 22856
rect 26840 22822 26877 22856
rect 26911 22822 26948 22856
rect 26982 22822 27019 22856
rect 27053 22822 27090 22856
rect 27124 22822 27161 22856
rect 27195 22822 27232 22856
rect 27266 22822 27302 22856
rect 27336 22822 27372 22856
rect 27406 22822 27442 22856
rect 27476 22822 27512 22856
rect 27546 22822 27582 22856
rect 27616 22822 27652 22856
rect 27686 22822 27722 22856
rect 27756 22822 27792 22856
rect 27826 22822 27862 22856
rect 27896 22822 27932 22856
rect 27966 22822 28000 22856
rect 26275 22782 28000 22822
rect 26275 22748 26309 22782
rect 26343 22748 26380 22782
rect 26414 22748 26451 22782
rect 26485 22748 26522 22782
rect 26556 22748 26593 22782
rect 26627 22748 26664 22782
rect 26698 22748 26735 22782
rect 26769 22748 26806 22782
rect 26840 22748 26877 22782
rect 26911 22748 26948 22782
rect 26982 22748 27019 22782
rect 27053 22748 27090 22782
rect 27124 22748 27161 22782
rect 27195 22748 27232 22782
rect 27266 22748 27302 22782
rect 27336 22748 27372 22782
rect 27406 22748 27442 22782
rect 27476 22748 27512 22782
rect 27546 22748 27582 22782
rect 27616 22748 27652 22782
rect 27686 22748 27722 22782
rect 27756 22748 27792 22782
rect 27826 22748 27862 22782
rect 27896 22748 27932 22782
rect 27966 22748 28000 22782
rect 26275 22708 28000 22748
rect 26275 22674 26309 22708
rect 26343 22674 26380 22708
rect 26414 22674 26451 22708
rect 26485 22674 26522 22708
rect 26556 22674 26593 22708
rect 26627 22674 26664 22708
rect 26698 22674 26735 22708
rect 26769 22674 26806 22708
rect 26840 22674 26877 22708
rect 26911 22674 26948 22708
rect 26982 22674 27019 22708
rect 27053 22674 27090 22708
rect 27124 22674 27161 22708
rect 27195 22674 27232 22708
rect 27266 22674 27302 22708
rect 27336 22674 27372 22708
rect 27406 22674 27442 22708
rect 27476 22674 27512 22708
rect 27546 22674 27582 22708
rect 27616 22674 27652 22708
rect 27686 22674 27722 22708
rect 27756 22674 27792 22708
rect 27826 22674 27862 22708
rect 27896 22674 27932 22708
rect 27966 22674 28000 22708
rect 26275 22634 28000 22674
rect 26275 22600 26309 22634
rect 26343 22600 26380 22634
rect 26414 22600 26451 22634
rect 26485 22600 26522 22634
rect 26556 22600 26593 22634
rect 26627 22600 26664 22634
rect 26698 22600 26735 22634
rect 26769 22600 26806 22634
rect 26840 22600 26877 22634
rect 26911 22600 26948 22634
rect 26982 22600 27019 22634
rect 27053 22600 27090 22634
rect 27124 22600 27161 22634
rect 27195 22600 27232 22634
rect 27266 22600 27302 22634
rect 27336 22600 27372 22634
rect 27406 22600 27442 22634
rect 27476 22600 27512 22634
rect 27546 22600 27582 22634
rect 27616 22600 27652 22634
rect 27686 22600 27722 22634
rect 27756 22600 27792 22634
rect 27826 22600 27862 22634
rect 27896 22600 27932 22634
rect 27966 22600 28000 22634
rect 26275 22560 28000 22600
rect 26275 22526 26309 22560
rect 26343 22526 26380 22560
rect 26414 22526 26451 22560
rect 26485 22526 26522 22560
rect 26556 22526 26593 22560
rect 26627 22526 26664 22560
rect 26698 22526 26735 22560
rect 26769 22526 26806 22560
rect 26840 22526 26877 22560
rect 26911 22526 26948 22560
rect 26982 22526 27019 22560
rect 27053 22526 27090 22560
rect 27124 22526 27161 22560
rect 27195 22526 27232 22560
rect 27266 22526 27302 22560
rect 27336 22526 27372 22560
rect 27406 22526 27442 22560
rect 27476 22526 27512 22560
rect 27546 22526 27582 22560
rect 27616 22526 27652 22560
rect 27686 22526 27722 22560
rect 27756 22526 27792 22560
rect 27826 22526 27862 22560
rect 27896 22526 27932 22560
rect 27966 22526 28000 22560
rect 26275 22486 28000 22526
rect 26275 22452 26309 22486
rect 26343 22452 26380 22486
rect 26414 22452 26451 22486
rect 26485 22452 26522 22486
rect 26556 22452 26593 22486
rect 26627 22452 26664 22486
rect 26698 22452 26735 22486
rect 26769 22452 26806 22486
rect 26840 22452 26877 22486
rect 26911 22452 26948 22486
rect 26982 22452 27019 22486
rect 27053 22452 27090 22486
rect 27124 22452 27161 22486
rect 27195 22452 27232 22486
rect 27266 22452 27302 22486
rect 27336 22452 27372 22486
rect 27406 22452 27442 22486
rect 27476 22452 27512 22486
rect 27546 22452 27582 22486
rect 27616 22452 27652 22486
rect 27686 22452 27722 22486
rect 27756 22452 27792 22486
rect 27826 22452 27862 22486
rect 27896 22452 27932 22486
rect 27966 22452 28000 22486
rect 26275 22412 28000 22452
rect 26275 22378 26309 22412
rect 26343 22378 26380 22412
rect 26414 22378 26451 22412
rect 26485 22378 26522 22412
rect 26556 22378 26593 22412
rect 26627 22378 26664 22412
rect 26698 22378 26735 22412
rect 26769 22378 26806 22412
rect 26840 22378 26877 22412
rect 26911 22378 26948 22412
rect 26982 22378 27019 22412
rect 27053 22378 27090 22412
rect 27124 22378 27161 22412
rect 27195 22378 27232 22412
rect 27266 22378 27302 22412
rect 27336 22378 27372 22412
rect 27406 22378 27442 22412
rect 27476 22378 27512 22412
rect 27546 22378 27582 22412
rect 27616 22378 27652 22412
rect 27686 22378 27722 22412
rect 27756 22378 27792 22412
rect 27826 22378 27862 22412
rect 27896 22378 27932 22412
rect 27966 22378 28000 22412
rect 26275 22338 28000 22378
rect 26275 22304 26309 22338
rect 26343 22304 26380 22338
rect 26414 22304 26451 22338
rect 26485 22304 26522 22338
rect 26556 22304 26593 22338
rect 26627 22304 26664 22338
rect 26698 22304 26735 22338
rect 26769 22304 26806 22338
rect 26840 22304 26877 22338
rect 26911 22304 26948 22338
rect 26982 22304 27019 22338
rect 27053 22304 27090 22338
rect 27124 22304 27161 22338
rect 27195 22304 27232 22338
rect 27266 22304 27302 22338
rect 27336 22304 27372 22338
rect 27406 22304 27442 22338
rect 27476 22304 27512 22338
rect 27546 22304 27582 22338
rect 27616 22304 27652 22338
rect 27686 22304 27722 22338
rect 27756 22304 27792 22338
rect 27826 22304 27862 22338
rect 27896 22304 27932 22338
rect 27966 22304 28000 22338
rect 26275 22264 28000 22304
rect 26275 22230 26309 22264
rect 26343 22230 26380 22264
rect 26414 22230 26451 22264
rect 26485 22230 26522 22264
rect 26556 22230 26593 22264
rect 26627 22230 26664 22264
rect 26698 22230 26735 22264
rect 26769 22230 26806 22264
rect 26840 22230 26877 22264
rect 26911 22230 26948 22264
rect 26982 22230 27019 22264
rect 27053 22230 27090 22264
rect 27124 22230 27161 22264
rect 27195 22230 27232 22264
rect 27266 22230 27302 22264
rect 27336 22230 27372 22264
rect 27406 22230 27442 22264
rect 27476 22230 27512 22264
rect 27546 22230 27582 22264
rect 27616 22230 27652 22264
rect 27686 22230 27722 22264
rect 27756 22230 27792 22264
rect 27826 22230 27862 22264
rect 27896 22230 27932 22264
rect 27966 22230 28000 22264
rect 26275 22190 28000 22230
rect 26275 22156 26309 22190
rect 26343 22156 26380 22190
rect 26414 22156 26451 22190
rect 26485 22156 26522 22190
rect 26556 22156 26593 22190
rect 26627 22156 26664 22190
rect 26698 22156 26735 22190
rect 26769 22156 26806 22190
rect 26840 22156 26877 22190
rect 26911 22156 26948 22190
rect 26982 22156 27019 22190
rect 27053 22156 27090 22190
rect 27124 22156 27161 22190
rect 27195 22156 27232 22190
rect 27266 22156 27302 22190
rect 27336 22156 27372 22190
rect 27406 22156 27442 22190
rect 27476 22156 27512 22190
rect 27546 22156 27582 22190
rect 27616 22156 27652 22190
rect 27686 22156 27722 22190
rect 27756 22156 27792 22190
rect 27826 22156 27862 22190
rect 27896 22156 27932 22190
rect 27966 22156 28000 22190
rect 26275 22116 28000 22156
rect 26275 22082 26309 22116
rect 26343 22082 26380 22116
rect 26414 22082 26451 22116
rect 26485 22082 26522 22116
rect 26556 22082 26593 22116
rect 26627 22082 26664 22116
rect 26698 22082 26735 22116
rect 26769 22082 26806 22116
rect 26840 22082 26877 22116
rect 26911 22082 26948 22116
rect 26982 22082 27019 22116
rect 27053 22082 27090 22116
rect 27124 22082 27161 22116
rect 27195 22082 27232 22116
rect 27266 22082 27302 22116
rect 27336 22082 27372 22116
rect 27406 22082 27442 22116
rect 27476 22082 27512 22116
rect 27546 22082 27582 22116
rect 27616 22082 27652 22116
rect 27686 22082 27722 22116
rect 27756 22082 27792 22116
rect 27826 22082 27862 22116
rect 27896 22082 27932 22116
rect 27966 22082 28000 22116
rect 26275 22080 28000 22082
rect 16853 9560 16903 9594
rect 16937 9560 16976 9594
rect 17010 9560 17049 9594
rect 17083 9560 17122 9594
rect 17156 9560 17195 9594
rect 17229 9560 17267 9594
rect 17301 9560 17339 9594
rect 17373 9560 17411 9594
rect 17445 9560 17483 9594
rect 17517 9560 17555 9594
rect 17589 9560 17613 9594
<< mvnsubdiff >>
rect 26978 20796 27172 20956
rect 26978 20762 27012 20796
rect 27046 20762 27172 20796
rect 26978 20728 27172 20762
rect 26978 20694 27012 20728
rect 27046 20694 27172 20728
rect 26978 20660 27172 20694
rect 26978 20626 27012 20660
rect 27046 20626 27172 20660
rect 26978 20592 27172 20626
rect 26978 20558 27012 20592
rect 27046 20558 27172 20592
rect 26978 20524 27172 20558
rect 26978 20490 27012 20524
rect 27046 20490 27172 20524
rect 26978 20456 27172 20490
rect 26978 20422 27012 20456
rect 27046 20422 27172 20456
rect 26978 20388 27172 20422
rect 26978 20354 27012 20388
rect 27046 20354 27172 20388
rect 26978 20320 27172 20354
rect 26978 20286 27012 20320
rect 27046 20286 27172 20320
rect 26978 20252 27172 20286
rect 26978 20218 27012 20252
rect 27046 20218 27172 20252
rect 26978 20184 27172 20218
rect 26978 20150 27012 20184
rect 27046 20150 27172 20184
rect 26978 20116 27172 20150
rect 26978 20082 27012 20116
rect 27046 20082 27172 20116
rect 26978 20048 27172 20082
rect 26978 20014 27012 20048
rect 27046 20014 27172 20048
rect 26978 19980 27172 20014
rect 26978 19946 27012 19980
rect 27046 19946 27172 19980
rect 26978 19912 27172 19946
rect 26978 19878 27012 19912
rect 27046 19878 27172 19912
rect 26978 19844 27172 19878
rect 26978 19810 27012 19844
rect 27046 19810 27172 19844
rect 26978 19776 27172 19810
rect 26978 19742 27012 19776
rect 27046 19742 27172 19776
rect 26978 19708 27172 19742
rect 26978 19674 27012 19708
rect 27046 19674 27172 19708
rect 26978 19640 27172 19674
rect 26978 19606 27012 19640
rect 27046 19606 27172 19640
rect 26978 19572 27172 19606
rect 26978 19538 27012 19572
rect 27046 19538 27172 19572
rect 26978 19504 27172 19538
rect 26978 19470 27012 19504
rect 27046 19470 27172 19504
rect 26978 19436 27172 19470
rect 26978 19402 27012 19436
rect 27046 19402 27172 19436
rect 26978 19368 27172 19402
rect 26978 19334 27012 19368
rect 27046 19334 27172 19368
rect 26978 19300 27172 19334
rect 26978 19266 27012 19300
rect 27046 19266 27172 19300
rect 26978 19232 27172 19266
rect 24129 19201 24639 19225
rect 24129 17704 24639 17739
rect 24163 17670 24197 17704
rect 24231 17670 24265 17704
rect 24299 17670 24333 17704
rect 24367 17670 24401 17704
rect 24435 17670 24469 17704
rect 24503 17670 24537 17704
rect 24571 17670 24605 17704
rect 24129 17635 24639 17670
rect 24163 17601 24197 17635
rect 24231 17601 24265 17635
rect 24299 17601 24333 17635
rect 24367 17601 24401 17635
rect 24435 17601 24469 17635
rect 24503 17601 24537 17635
rect 24571 17601 24605 17635
rect 24129 17566 24639 17601
rect 24163 17532 24197 17566
rect 24231 17532 24265 17566
rect 24299 17532 24333 17566
rect 24367 17532 24401 17566
rect 24435 17532 24469 17566
rect 24503 17532 24537 17566
rect 24571 17532 24605 17566
rect 24129 17497 24639 17532
rect 24163 17463 24197 17497
rect 24231 17463 24265 17497
rect 24299 17463 24333 17497
rect 24367 17463 24401 17497
rect 24435 17463 24469 17497
rect 24503 17463 24537 17497
rect 24571 17463 24605 17497
rect 24129 17428 24639 17463
rect 24163 17394 24197 17428
rect 24231 17394 24265 17428
rect 24299 17394 24333 17428
rect 24367 17394 24401 17428
rect 24435 17394 24469 17428
rect 24503 17394 24537 17428
rect 24571 17394 24605 17428
rect 24129 17359 24639 17394
rect 24163 17325 24197 17359
rect 24231 17325 24265 17359
rect 24299 17325 24333 17359
rect 24367 17325 24401 17359
rect 24435 17325 24469 17359
rect 24503 17325 24537 17359
rect 24571 17325 24605 17359
rect 24129 17290 24639 17325
rect 24163 17256 24197 17290
rect 24231 17256 24265 17290
rect 24299 17256 24333 17290
rect 24367 17256 24401 17290
rect 24435 17256 24469 17290
rect 24503 17256 24537 17290
rect 24571 17256 24605 17290
rect 24129 17221 24639 17256
rect 24163 17187 24197 17221
rect 24231 17187 24265 17221
rect 24299 17187 24333 17221
rect 24367 17187 24401 17221
rect 24435 17187 24469 17221
rect 24503 17187 24537 17221
rect 24571 17187 24605 17221
rect 24129 17152 24639 17187
rect 24163 17118 24197 17152
rect 24231 17118 24265 17152
rect 24299 17118 24333 17152
rect 24367 17118 24401 17152
rect 24435 17118 24469 17152
rect 24503 17118 24537 17152
rect 24571 17118 24605 17152
rect 24129 17083 24639 17118
rect 24163 17049 24197 17083
rect 24231 17049 24265 17083
rect 24299 17049 24333 17083
rect 24367 17049 24401 17083
rect 24435 17049 24469 17083
rect 24503 17049 24537 17083
rect 24571 17049 24605 17083
rect 24129 17014 24639 17049
rect 24163 16980 24197 17014
rect 24231 16980 24265 17014
rect 24299 16980 24333 17014
rect 24367 16980 24401 17014
rect 24435 16980 24469 17014
rect 24503 16980 24537 17014
rect 24571 16980 24605 17014
rect 24129 16945 24639 16980
rect 24163 16911 24197 16945
rect 24231 16911 24265 16945
rect 24299 16911 24333 16945
rect 24367 16911 24401 16945
rect 24435 16911 24469 16945
rect 24503 16911 24537 16945
rect 24571 16911 24605 16945
rect 24129 16876 24639 16911
rect 24163 16842 24197 16876
rect 24231 16842 24265 16876
rect 24299 16842 24333 16876
rect 24367 16842 24401 16876
rect 24435 16842 24469 16876
rect 24503 16842 24537 16876
rect 24571 16842 24605 16876
rect 24129 16807 24639 16842
rect 24163 16773 24197 16807
rect 24231 16773 24265 16807
rect 24299 16773 24333 16807
rect 24367 16773 24401 16807
rect 24435 16773 24469 16807
rect 24503 16773 24537 16807
rect 24571 16773 24605 16807
rect 24129 16738 24639 16773
rect 24163 16704 24197 16738
rect 24231 16704 24265 16738
rect 24299 16704 24333 16738
rect 24367 16704 24401 16738
rect 24435 16704 24469 16738
rect 24503 16704 24537 16738
rect 24571 16704 24605 16738
rect 24129 16669 24639 16704
rect 24163 16635 24197 16669
rect 24231 16635 24265 16669
rect 24299 16635 24333 16669
rect 24367 16635 24401 16669
rect 24435 16635 24469 16669
rect 24503 16635 24537 16669
rect 24571 16635 24605 16669
rect 24129 16600 24639 16635
rect 24163 16566 24197 16600
rect 24231 16566 24265 16600
rect 24299 16566 24333 16600
rect 24367 16566 24401 16600
rect 24435 16566 24469 16600
rect 24503 16566 24537 16600
rect 24571 16566 24605 16600
rect 24129 16531 24639 16566
rect 24163 16497 24197 16531
rect 24231 16497 24265 16531
rect 24299 16497 24333 16531
rect 24367 16497 24401 16531
rect 24435 16497 24469 16531
rect 24503 16497 24537 16531
rect 24571 16497 24605 16531
rect 24129 16462 24639 16497
rect 24163 16428 24197 16462
rect 24231 16428 24265 16462
rect 24299 16428 24333 16462
rect 24367 16428 24401 16462
rect 24435 16428 24469 16462
rect 24503 16428 24537 16462
rect 24571 16428 24605 16462
rect 24129 16404 24639 16428
rect 24145 16338 24639 16404
rect 26978 19198 27012 19232
rect 27046 19198 27172 19232
rect 26978 19164 27172 19198
rect 26978 19130 27012 19164
rect 27046 19130 27172 19164
rect 26978 19096 27172 19130
rect 26978 19062 27012 19096
rect 27046 19062 27172 19096
rect 26978 19028 27172 19062
rect 26978 18994 27012 19028
rect 27046 18994 27172 19028
rect 26978 18960 27172 18994
rect 26978 18926 27012 18960
rect 27046 18926 27172 18960
rect 26978 18892 27172 18926
rect 26978 18858 27012 18892
rect 27046 18858 27172 18892
rect 26978 18824 27172 18858
rect 26978 18790 27012 18824
rect 27046 18790 27172 18824
rect 26978 18756 27172 18790
rect 26978 18722 27012 18756
rect 27046 18722 27172 18756
rect 26978 18688 27172 18722
rect 26978 18654 27012 18688
rect 27046 18654 27172 18688
rect 26978 18620 27172 18654
rect 26978 18586 27012 18620
rect 27046 18586 27172 18620
rect 26978 18552 27172 18586
rect 26978 18518 27012 18552
rect 27046 18518 27172 18552
rect 26978 18484 27172 18518
rect 26978 18450 27012 18484
rect 27046 18450 27172 18484
rect 26978 18416 27172 18450
rect 26978 18382 27012 18416
rect 27046 18382 27172 18416
rect 26978 18348 27172 18382
rect 26978 18314 27012 18348
rect 27046 18314 27172 18348
rect 26978 18280 27172 18314
rect 26978 18246 27012 18280
rect 27046 18246 27172 18280
rect 26978 18212 27172 18246
rect 26978 18178 27012 18212
rect 27046 18178 27172 18212
rect 26978 18144 27172 18178
rect 26978 18110 27012 18144
rect 27046 18110 27172 18144
rect 26978 18076 27172 18110
rect 26978 18042 27012 18076
rect 27046 18042 27172 18076
rect 26978 18008 27172 18042
rect 26978 17974 27012 18008
rect 27046 17974 27172 18008
rect 26978 17940 27172 17974
rect 26978 17906 27012 17940
rect 27046 17906 27172 17940
rect 26978 17872 27172 17906
rect 26978 17838 27012 17872
rect 27046 17838 27172 17872
rect 26978 17804 27172 17838
rect 26978 17770 27012 17804
rect 27046 17770 27172 17804
rect 26978 17736 27172 17770
rect 26978 17702 27012 17736
rect 27046 17702 27172 17736
rect 26978 17668 27172 17702
rect 26978 17634 27012 17668
rect 27046 17634 27172 17668
rect 26978 17600 27172 17634
rect 26978 17566 27012 17600
rect 27046 17566 27172 17600
rect 26978 17532 27172 17566
rect 26978 17498 27012 17532
rect 27046 17498 27172 17532
rect 26978 17464 27172 17498
rect 26978 17430 27012 17464
rect 27046 17430 27172 17464
rect 26978 17396 27172 17430
rect 26978 17362 27012 17396
rect 27046 17362 27172 17396
rect 26978 17328 27172 17362
rect 26978 17294 27012 17328
rect 27046 17294 27172 17328
rect 26978 17259 27172 17294
rect 26978 17225 27012 17259
rect 27046 17225 27172 17259
rect 26978 17190 27172 17225
rect 26978 17156 27012 17190
rect 27046 17156 27172 17190
rect 26978 17121 27172 17156
rect 26978 17087 27012 17121
rect 27046 17087 27172 17121
rect 26978 17052 27172 17087
rect 26978 17018 27012 17052
rect 27046 17018 27172 17052
rect 26978 16983 27172 17018
rect 26978 16949 27012 16983
rect 27046 16949 27172 16983
rect 26978 16914 27172 16949
rect 26978 16880 27012 16914
rect 27046 16880 27172 16914
rect 26978 16845 27172 16880
rect 26978 16811 27012 16845
rect 27046 16811 27172 16845
rect 26978 16776 27172 16811
rect 26978 16742 27012 16776
rect 27046 16742 27172 16776
rect 26978 16707 27172 16742
rect 26978 16673 27012 16707
rect 27046 16673 27172 16707
rect 26978 16638 27172 16673
rect 26978 16604 27012 16638
rect 27046 16604 27172 16638
rect 26978 16569 27172 16604
rect 26978 16535 27012 16569
rect 27046 16535 27172 16569
rect 26978 16500 27172 16535
rect 26978 16466 27012 16500
rect 27046 16466 27172 16500
rect 26978 16431 27172 16466
rect 26978 16397 27012 16431
rect 27046 16397 27172 16431
rect 26978 16362 27172 16397
rect 26978 16328 27012 16362
rect 27046 16328 27172 16362
rect 26978 16293 27172 16328
rect 26978 16259 27012 16293
rect 27046 16259 27172 16293
rect 26978 16224 27172 16259
rect 26978 16190 27012 16224
rect 27046 16190 27172 16224
rect 26978 16155 27172 16190
rect 26978 16121 27012 16155
rect 27046 16121 27172 16155
rect 26978 16086 27172 16121
rect 26978 16052 27012 16086
rect 27046 16052 27172 16086
rect 26978 16017 27172 16052
rect 26978 15983 27012 16017
rect 27046 15983 27172 16017
rect 26978 15948 27172 15983
rect 26978 15914 27012 15948
rect 27046 15914 27172 15948
rect 26978 15879 27172 15914
rect 26978 15845 27012 15879
rect 27046 15845 27172 15879
rect 26978 15810 27172 15845
rect 26978 15776 27012 15810
rect 27046 15776 27172 15810
rect 26978 15741 27172 15776
rect 26978 15707 27012 15741
rect 27046 15707 27172 15741
rect 26978 15672 27172 15707
rect 26978 15638 27012 15672
rect 27046 15638 27172 15672
rect 26978 15603 27172 15638
rect 26978 15569 27012 15603
rect 27046 15569 27172 15603
rect 26978 15534 27172 15569
rect 26978 15500 27012 15534
rect 27046 15500 27172 15534
rect 26978 15465 27172 15500
rect 26978 15431 27012 15465
rect 27046 15431 27172 15465
rect 26978 15396 27172 15431
rect 26978 15362 27012 15396
rect 27046 15362 27172 15396
rect 26978 15327 27172 15362
rect 26978 15293 27012 15327
rect 27046 15293 27172 15327
rect 26978 15258 27172 15293
rect 26978 15224 27012 15258
rect 27046 15224 27172 15258
rect 26978 15189 27172 15224
rect 26978 15155 27012 15189
rect 27046 15155 27172 15189
rect 26978 15120 27172 15155
rect 26978 15086 27012 15120
rect 27046 15086 27172 15120
rect 26978 15051 27172 15086
rect 26978 15017 27012 15051
rect 27046 15017 27172 15051
rect 26978 14857 27172 15017
<< psubdiffcont >>
rect 27287 37585 27321 37619
rect 27355 37585 27389 37619
rect 27423 37585 27457 37619
rect 27491 37585 27525 37619
rect 27219 37525 27253 37559
rect 27585 37551 27619 37585
rect 27219 37457 27253 37491
rect 27219 37389 27253 37423
rect 27219 37321 27253 37355
rect 27585 37483 27619 37517
rect 27585 37415 27619 37449
rect 27585 37347 27619 37381
rect 27219 37253 27253 37287
rect 27347 37219 27381 37253
rect 27415 37219 27449 37253
rect 27483 37219 27517 37253
rect 27551 37219 27585 37253
rect 2344 4024 2378 4058
rect 2415 4024 2449 4058
rect 2486 4024 2520 4058
rect 2557 4024 2591 4058
rect 2628 4024 2662 4058
rect 2698 4024 2732 4058
rect 2768 4024 2802 4058
rect 2838 4024 2872 4058
rect 2908 4024 2942 4058
rect 2978 4024 3012 4058
rect 3048 4024 3082 4058
rect 3118 4024 3152 4058
rect 3188 4024 3222 4058
rect 3258 4024 3292 4058
rect 3350 4026 3384 4060
rect 3419 4026 3453 4060
rect 3488 4026 3522 4060
rect 3557 4026 3591 4060
rect 3626 4026 3660 4060
rect 3695 4026 3729 4060
rect 3764 4026 3798 4060
rect 3833 4026 3867 4060
rect 3902 4026 3936 4060
rect 3971 4026 4005 4060
rect 4040 4026 4074 4060
rect 4109 4026 4143 4060
rect 4178 4026 4212 4060
rect 4247 4026 4281 4060
rect 4316 4026 4350 4060
rect 4385 4026 4419 4060
rect 4454 4026 4488 4060
rect 4523 4026 4557 4060
rect 4592 4026 4626 4060
rect 4661 4026 4695 4060
rect 4730 4026 4764 4060
rect 4799 4026 4833 4060
rect 4868 4026 4902 4060
rect 4937 4026 4971 4060
rect 5006 4026 5040 4060
rect 5075 4026 5109 4060
rect 5144 4026 5178 4060
rect 5213 4026 5247 4060
rect 5282 4026 5316 4060
rect 5351 4026 5385 4060
rect 5420 4026 5454 4060
rect 5489 4026 5523 4060
rect 5558 4026 5592 4060
rect 5627 4026 5661 4060
rect 5696 4026 5730 4060
rect 5765 4026 5799 4060
rect 5834 4026 5868 4060
rect 5903 4026 5937 4060
rect 5972 4026 6006 4060
rect 2344 3950 2378 3984
rect 2415 3950 2449 3984
rect 2486 3950 2520 3984
rect 2557 3950 2591 3984
rect 2628 3950 2662 3984
rect 2698 3950 2732 3984
rect 2768 3950 2802 3984
rect 2838 3950 2872 3984
rect 2908 3950 2942 3984
rect 2978 3950 3012 3984
rect 3048 3950 3082 3984
rect 3118 3950 3152 3984
rect 3188 3950 3222 3984
rect 3258 3950 3292 3984
rect 3350 3958 3384 3992
rect 3419 3958 3453 3992
rect 3488 3958 3522 3992
rect 3557 3958 3591 3992
rect 3626 3958 3660 3992
rect 3695 3958 3729 3992
rect 3764 3958 3798 3992
rect 3833 3958 3867 3992
rect 3902 3958 3936 3992
rect 3971 3958 4005 3992
rect 4040 3958 4074 3992
rect 4109 3958 4143 3992
rect 4178 3958 4212 3992
rect 4247 3958 4281 3992
rect 4316 3958 4350 3992
rect 4385 3958 4419 3992
rect 4454 3958 4488 3992
rect 4523 3958 4557 3992
rect 4592 3958 4626 3992
rect 4661 3958 4695 3992
rect 4730 3958 4764 3992
rect 4799 3958 4833 3992
rect 4868 3958 4902 3992
rect 4937 3958 4971 3992
rect 5006 3958 5040 3992
rect 5075 3958 5109 3992
rect 5144 3958 5178 3992
rect 5213 3958 5247 3992
rect 5282 3958 5316 3992
rect 5351 3958 5385 3992
rect 5420 3958 5454 3992
rect 5489 3958 5523 3992
rect 5558 3958 5592 3992
rect 5627 3958 5661 3992
rect 5696 3958 5730 3992
rect 5765 3958 5799 3992
rect 5834 3958 5868 3992
rect 5903 3958 5937 3992
rect 5972 3958 6006 3992
rect 2344 3876 2378 3910
rect 2415 3876 2449 3910
rect 2486 3876 2520 3910
rect 2557 3876 2591 3910
rect 2628 3876 2662 3910
rect 2698 3876 2732 3910
rect 2768 3876 2802 3910
rect 2838 3876 2872 3910
rect 2908 3876 2942 3910
rect 2978 3876 3012 3910
rect 3048 3876 3082 3910
rect 3118 3876 3152 3910
rect 3188 3876 3222 3910
rect 3258 3876 3292 3910
rect 3350 3890 3384 3924
rect 3419 3890 3453 3924
rect 3488 3890 3522 3924
rect 3557 3890 3591 3924
rect 3626 3890 3660 3924
rect 3695 3890 3729 3924
rect 3764 3890 3798 3924
rect 3833 3890 3867 3924
rect 3902 3890 3936 3924
rect 3971 3890 4005 3924
rect 4040 3890 4074 3924
rect 4109 3890 4143 3924
rect 4178 3890 4212 3924
rect 4247 3890 4281 3924
rect 4316 3890 4350 3924
rect 4385 3890 4419 3924
rect 4454 3890 4488 3924
rect 4523 3890 4557 3924
rect 4592 3890 4626 3924
rect 4661 3890 4695 3924
rect 4730 3890 4764 3924
rect 4799 3890 4833 3924
rect 4868 3890 4902 3924
rect 4937 3890 4971 3924
rect 5006 3890 5040 3924
rect 5075 3890 5109 3924
rect 5144 3890 5178 3924
rect 5213 3890 5247 3924
rect 5282 3890 5316 3924
rect 5351 3890 5385 3924
rect 5420 3890 5454 3924
rect 5489 3890 5523 3924
rect 5558 3890 5592 3924
rect 5627 3890 5661 3924
rect 5696 3890 5730 3924
rect 5765 3890 5799 3924
rect 5834 3890 5868 3924
rect 5903 3890 5937 3924
rect 5972 3890 6006 3924
rect 2344 3802 2378 3836
rect 2415 3802 2449 3836
rect 2486 3802 2520 3836
rect 2557 3802 2591 3836
rect 2628 3802 2662 3836
rect 2698 3802 2732 3836
rect 2768 3802 2802 3836
rect 2838 3802 2872 3836
rect 2908 3802 2942 3836
rect 2978 3802 3012 3836
rect 3048 3802 3082 3836
rect 3118 3802 3152 3836
rect 3188 3802 3222 3836
rect 3258 3802 3292 3836
rect 3350 3822 3384 3856
rect 3419 3822 3453 3856
rect 3488 3822 3522 3856
rect 3557 3822 3591 3856
rect 3626 3822 3660 3856
rect 3695 3822 3729 3856
rect 3764 3822 3798 3856
rect 3833 3822 3867 3856
rect 3902 3822 3936 3856
rect 3971 3822 4005 3856
rect 4040 3822 4074 3856
rect 4109 3822 4143 3856
rect 4178 3822 4212 3856
rect 4247 3822 4281 3856
rect 4316 3822 4350 3856
rect 4385 3822 4419 3856
rect 4454 3822 4488 3856
rect 4523 3822 4557 3856
rect 4592 3822 4626 3856
rect 4661 3822 4695 3856
rect 4730 3822 4764 3856
rect 4799 3822 4833 3856
rect 4868 3822 4902 3856
rect 4937 3822 4971 3856
rect 5006 3822 5040 3856
rect 5075 3822 5109 3856
rect 5144 3822 5178 3856
rect 5213 3822 5247 3856
rect 5282 3822 5316 3856
rect 5351 3822 5385 3856
rect 5420 3822 5454 3856
rect 5489 3822 5523 3856
rect 5558 3822 5592 3856
rect 5627 3822 5661 3856
rect 5696 3822 5730 3856
rect 5765 3822 5799 3856
rect 5834 3822 5868 3856
rect 5903 3822 5937 3856
rect 5972 3822 6006 3856
rect 2344 3728 2378 3762
rect 2415 3728 2449 3762
rect 2486 3728 2520 3762
rect 2557 3728 2591 3762
rect 2628 3728 2662 3762
rect 2698 3728 2732 3762
rect 2768 3728 2802 3762
rect 2838 3728 2872 3762
rect 2908 3728 2942 3762
rect 2978 3728 3012 3762
rect 3048 3728 3082 3762
rect 3118 3728 3152 3762
rect 3188 3728 3222 3762
rect 3258 3728 3292 3762
rect 3350 3754 3384 3788
rect 3419 3754 3453 3788
rect 3488 3754 3522 3788
rect 3557 3754 3591 3788
rect 3626 3754 3660 3788
rect 3695 3754 3729 3788
rect 3764 3754 3798 3788
rect 3833 3754 3867 3788
rect 3902 3754 3936 3788
rect 3971 3754 4005 3788
rect 4040 3754 4074 3788
rect 4109 3754 4143 3788
rect 4178 3754 4212 3788
rect 4247 3754 4281 3788
rect 4316 3754 4350 3788
rect 4385 3754 4419 3788
rect 4454 3754 4488 3788
rect 4523 3754 4557 3788
rect 4592 3754 4626 3788
rect 4661 3754 4695 3788
rect 4730 3754 4764 3788
rect 4799 3754 4833 3788
rect 4868 3754 4902 3788
rect 4937 3754 4971 3788
rect 5006 3754 5040 3788
rect 5075 3754 5109 3788
rect 5144 3754 5178 3788
rect 5213 3754 5247 3788
rect 5282 3754 5316 3788
rect 5351 3754 5385 3788
rect 5420 3754 5454 3788
rect 5489 3754 5523 3788
rect 5558 3754 5592 3788
rect 5627 3754 5661 3788
rect 5696 3754 5730 3788
rect 5765 3754 5799 3788
rect 5834 3754 5868 3788
rect 5903 3754 5937 3788
rect 5972 3754 6006 3788
rect 6041 3754 6415 4060
rect 6473 4024 6507 4058
rect 6542 4024 6576 4058
rect 6611 4024 6645 4058
rect 6680 4024 6714 4058
rect 6749 4024 6783 4058
rect 6818 4024 6852 4058
rect 6887 4024 6921 4058
rect 6956 4024 6990 4058
rect 7025 4024 7059 4058
rect 7094 4024 7128 4058
rect 7163 4024 7197 4058
rect 7232 4024 7266 4058
rect 7301 4024 7335 4058
rect 7370 4024 7404 4058
rect 7439 4024 7473 4058
rect 7508 4024 7542 4058
rect 7577 4024 7611 4058
rect 7646 4024 7680 4058
rect 7715 4024 7749 4058
rect 7784 4024 7818 4058
rect 7853 4024 7887 4058
rect 7922 4024 7956 4058
rect 7991 4024 8025 4058
rect 8060 4024 8094 4058
rect 8129 4024 8163 4058
rect 8198 4024 8232 4058
rect 8267 4024 8301 4058
rect 8336 4024 8370 4058
rect 8405 4024 8439 4058
rect 8474 4024 8508 4058
rect 8543 4024 8577 4058
rect 8612 4024 8646 4058
rect 8681 4024 8715 4058
rect 8750 4024 8784 4058
rect 8819 4024 8853 4058
rect 8888 4024 8922 4058
rect 8957 4024 8991 4058
rect 9026 4024 9060 4058
rect 9095 4024 9129 4058
rect 9164 4024 9198 4058
rect 9233 4024 9267 4058
rect 9302 4024 9336 4058
rect 9371 4024 9405 4058
rect 9440 4024 9474 4058
rect 9509 4024 9543 4058
rect 9578 4024 9612 4058
rect 9647 4024 9681 4058
rect 9716 4024 9750 4058
rect 9785 4024 9819 4058
rect 9854 4024 9888 4058
rect 9922 4024 9956 4058
rect 9990 4024 10024 4058
rect 10058 4024 10092 4058
rect 10126 4024 10160 4058
rect 10194 4024 10228 4058
rect 10262 4024 10296 4058
rect 10330 4024 10364 4058
rect 10398 4024 10432 4058
rect 10466 4024 10500 4058
rect 10534 4024 10568 4058
rect 10602 4024 10636 4058
rect 10670 4024 10704 4058
rect 10738 4024 10772 4058
rect 10806 4024 10840 4058
rect 10874 4024 10908 4058
rect 10942 4024 10976 4058
rect 11010 4024 11044 4058
rect 11078 4024 11112 4058
rect 11146 4024 11180 4058
rect 11214 4024 11248 4058
rect 11282 4024 11316 4058
rect 11350 4024 11384 4058
rect 11418 4024 11452 4058
rect 11486 4024 11520 4058
rect 11554 4024 11588 4058
rect 11622 4024 11656 4058
rect 11690 4024 11724 4058
rect 11758 4024 11792 4058
rect 11826 4024 11860 4058
rect 11894 4024 11928 4058
rect 11962 4024 11996 4058
rect 12030 4024 12064 4058
rect 12098 4024 12132 4058
rect 12166 4024 12200 4058
rect 12234 4024 12268 4058
rect 12302 4024 12336 4058
rect 12370 4024 12404 4058
rect 12438 4024 12472 4058
rect 12506 4024 12540 4058
rect 12574 4024 12608 4058
rect 12642 4024 12676 4058
rect 12710 4024 12744 4058
rect 12778 4024 12812 4058
rect 12846 4024 12880 4058
rect 12914 4024 12948 4058
rect 12982 4024 13016 4058
rect 13050 4024 13084 4058
rect 13118 4024 13152 4058
rect 13186 4024 13220 4058
rect 13254 4024 13288 4058
rect 13322 4024 13356 4058
rect 13390 4024 13424 4058
rect 13458 4024 13492 4058
rect 13526 4024 13560 4058
rect 13594 4024 13628 4058
rect 13662 4024 13696 4058
rect 13730 4024 13764 4058
rect 13798 4024 13832 4058
rect 13866 4024 13900 4058
rect 13934 4024 13968 4058
rect 14002 4024 14036 4058
rect 14070 4024 14104 4058
rect 14138 4024 14172 4058
rect 14206 4024 14240 4058
rect 14274 4024 14308 4058
rect 14342 4024 14376 4058
rect 14410 4024 14444 4058
rect 14478 4024 14512 4058
rect 14546 4024 14580 4058
rect 14614 4024 14648 4058
rect 14682 4024 14716 4058
rect 14750 4024 14784 4058
rect 14818 4024 14852 4058
rect 14886 4024 14920 4058
rect 14954 4024 14988 4058
rect 15022 4024 15056 4058
rect 15090 4024 15124 4058
rect 15158 4024 15192 4058
rect 15226 4024 15260 4058
rect 15294 4024 15328 4058
rect 15362 4024 15396 4058
rect 15430 4024 15464 4058
rect 15498 4024 15532 4058
rect 15566 4024 15600 4058
rect 15634 4024 15668 4058
rect 15702 4024 15736 4058
rect 15770 4024 15804 4058
rect 15838 4024 15872 4058
rect 15906 4024 15940 4058
rect 15974 4024 16008 4058
rect 16042 4024 16076 4058
rect 16110 4024 16144 4058
rect 16178 4024 16212 4058
rect 16246 4024 16280 4058
rect 16314 4024 16348 4058
rect 16382 4024 16416 4058
rect 16450 4024 16484 4058
rect 16518 4024 16552 4058
rect 16586 4024 16620 4058
rect 16654 4024 16688 4058
rect 16722 4024 16756 4058
rect 16790 4024 16824 4058
rect 16858 4024 16892 4058
rect 16926 4024 16960 4058
rect 16994 4024 17028 4058
rect 17062 4024 17096 4058
rect 17130 4024 17164 4058
rect 17198 4024 17232 4058
rect 17266 4024 17300 4058
rect 17334 4024 17368 4058
rect 17402 4024 17436 4058
rect 17470 4024 17504 4058
rect 17538 4024 17572 4058
rect 17606 4024 17640 4058
rect 17674 4024 17708 4058
rect 17742 4024 17776 4058
rect 17810 4024 17844 4058
rect 17878 4024 17912 4058
rect 17946 4024 17980 4058
rect 18014 4024 18048 4058
rect 18082 4024 18116 4058
rect 18150 4024 18184 4058
rect 18218 4024 18252 4058
rect 18286 4024 18320 4058
rect 18354 4024 18388 4058
rect 18422 4024 18456 4058
rect 18490 4024 18524 4058
rect 18558 4024 18592 4058
rect 18626 4024 18660 4058
rect 18694 4024 18728 4058
rect 18762 4024 18796 4058
rect 18830 4024 18864 4058
rect 18898 4024 18932 4058
rect 18966 4024 19000 4058
rect 19034 4024 19068 4058
rect 19102 4024 19136 4058
rect 19170 4024 19204 4058
rect 19238 4024 19272 4058
rect 19306 4024 19340 4058
rect 19374 4024 19408 4058
rect 19442 4024 19476 4058
rect 19510 4024 19544 4058
rect 19578 4024 19612 4058
rect 19646 4024 19680 4058
rect 19714 4024 19748 4058
rect 19782 4024 19816 4058
rect 19850 4024 19884 4058
rect 19918 4024 19952 4058
rect 19986 4024 20020 4058
rect 20054 4024 20088 4058
rect 20122 4024 20156 4058
rect 20190 4024 20224 4058
rect 20258 4024 20292 4058
rect 20326 4024 20360 4058
rect 20394 4024 20428 4058
rect 20462 4024 20496 4058
rect 20530 4024 20564 4058
rect 20598 4024 20632 4058
rect 20666 4024 20700 4058
rect 20734 4024 20768 4058
rect 20802 4024 20836 4058
rect 20870 4024 20904 4058
rect 20938 4024 20972 4058
rect 21006 4024 21040 4058
rect 21074 4024 21108 4058
rect 21142 4024 21176 4058
rect 21210 4024 21244 4058
rect 21278 4024 21312 4058
rect 21346 4024 21380 4058
rect 21414 4024 21448 4058
rect 21482 4024 21516 4058
rect 21550 4024 21584 4058
rect 21618 4024 21652 4058
rect 21686 4024 21720 4058
rect 21754 4024 21788 4058
rect 21822 4024 21856 4058
rect 21890 4024 21924 4058
rect 21958 4024 21992 4058
rect 22026 4024 22060 4058
rect 22094 4024 22128 4058
rect 22162 4024 22196 4058
rect 22230 4024 22264 4058
rect 22298 4024 22332 4058
rect 22366 4024 22400 4058
rect 22434 4024 22468 4058
rect 22502 4024 22536 4058
rect 22570 4024 22604 4058
rect 22638 4024 22672 4058
rect 22706 4024 22740 4058
rect 22774 4024 22808 4058
rect 22842 4024 22876 4058
rect 22910 4024 22944 4058
rect 22978 4024 23012 4058
rect 23046 4024 23080 4058
rect 23114 4024 23148 4058
rect 23182 4024 23216 4058
rect 23250 4024 23284 4058
rect 23318 4024 23352 4058
rect 23386 4024 23420 4058
rect 23454 4024 23488 4058
rect 23522 4024 23556 4058
rect 23590 4024 23624 4058
rect 23658 4024 23692 4058
rect 23726 4024 23760 4058
rect 23794 4024 23828 4058
rect 23862 4024 23896 4058
rect 23930 4024 23964 4058
rect 23998 4024 24032 4058
rect 24066 4024 24100 4058
rect 24134 4024 24168 4058
rect 24202 4024 24236 4058
rect 24270 4024 24304 4058
rect 24338 4024 24372 4058
rect 24406 4024 24440 4058
rect 24474 4024 24508 4058
rect 24542 4024 24576 4058
rect 24610 4024 24644 4058
rect 24678 4024 24712 4058
rect 24746 4024 24780 4058
rect 24814 4024 24848 4058
rect 24882 4024 24916 4058
rect 24950 4024 24984 4058
rect 25018 4024 25052 4058
rect 25086 4024 25120 4058
rect 25154 4024 25188 4058
rect 25222 4024 25256 4058
rect 25290 4024 25324 4058
rect 25358 4024 25392 4058
rect 25426 4024 25460 4058
rect 25494 4024 25528 4058
rect 25562 4024 25596 4058
rect 25630 4024 25664 4058
rect 25698 4024 25732 4058
rect 25766 4024 25800 4058
rect 25834 4024 25868 4058
rect 25902 4024 25936 4058
rect 25970 4024 26004 4058
rect 26038 4024 26072 4058
rect 26106 4024 26140 4058
rect 26174 4024 26208 4058
rect 26242 4024 26276 4058
rect 26310 4024 26344 4058
rect 26378 4024 26412 4058
rect 26446 4024 26480 4058
rect 26514 4024 26548 4058
rect 26582 4024 26616 4058
rect 26650 4024 26684 4058
rect 26718 4024 26752 4058
rect 26786 4024 26820 4058
rect 26854 4024 26888 4058
rect 26922 4024 26956 4058
rect 26990 4024 27024 4058
rect 27058 4024 27092 4058
rect 27126 4024 27160 4058
rect 27194 4024 27228 4058
rect 27262 4024 27296 4058
rect 27330 4024 27364 4058
rect 27398 4024 27432 4058
rect 27466 4024 27500 4058
rect 27534 4024 27568 4058
rect 27602 4024 27636 4058
rect 27670 4024 27704 4058
rect 27738 4024 27772 4058
rect 27806 4024 27840 4058
rect 27874 4024 27908 4058
rect 27942 4024 27976 4058
rect 6473 3950 6507 3984
rect 6542 3950 6576 3984
rect 6611 3950 6645 3984
rect 6680 3950 6714 3984
rect 6749 3950 6783 3984
rect 6818 3950 6852 3984
rect 6887 3950 6921 3984
rect 6956 3950 6990 3984
rect 7025 3950 7059 3984
rect 7094 3950 7128 3984
rect 7163 3950 7197 3984
rect 7232 3950 7266 3984
rect 7301 3950 7335 3984
rect 7370 3950 7404 3984
rect 7439 3950 7473 3984
rect 7508 3950 7542 3984
rect 7577 3950 7611 3984
rect 7646 3950 7680 3984
rect 7715 3950 7749 3984
rect 7784 3950 7818 3984
rect 7853 3950 7887 3984
rect 7922 3950 7956 3984
rect 7991 3950 8025 3984
rect 8060 3950 8094 3984
rect 8129 3950 8163 3984
rect 8198 3950 8232 3984
rect 8267 3950 8301 3984
rect 8336 3950 8370 3984
rect 8405 3950 8439 3984
rect 8474 3950 8508 3984
rect 8543 3950 8577 3984
rect 8612 3950 8646 3984
rect 8681 3950 8715 3984
rect 8750 3950 8784 3984
rect 8819 3950 8853 3984
rect 8888 3950 8922 3984
rect 8957 3950 8991 3984
rect 9026 3950 9060 3984
rect 9095 3950 9129 3984
rect 9164 3950 9198 3984
rect 9233 3950 9267 3984
rect 9302 3950 9336 3984
rect 9371 3950 9405 3984
rect 9440 3950 9474 3984
rect 9509 3950 9543 3984
rect 9578 3950 9612 3984
rect 9647 3950 9681 3984
rect 9716 3950 9750 3984
rect 9785 3950 9819 3984
rect 9854 3950 9888 3984
rect 9922 3950 9956 3984
rect 9990 3950 10024 3984
rect 10058 3950 10092 3984
rect 10126 3950 10160 3984
rect 10194 3950 10228 3984
rect 10262 3950 10296 3984
rect 10330 3950 10364 3984
rect 10398 3950 10432 3984
rect 10466 3950 10500 3984
rect 10534 3950 10568 3984
rect 10602 3950 10636 3984
rect 10670 3950 10704 3984
rect 10738 3950 10772 3984
rect 10806 3950 10840 3984
rect 10874 3950 10908 3984
rect 10942 3950 10976 3984
rect 11010 3950 11044 3984
rect 11078 3950 11112 3984
rect 11146 3950 11180 3984
rect 11214 3950 11248 3984
rect 11282 3950 11316 3984
rect 11350 3950 11384 3984
rect 11418 3950 11452 3984
rect 11486 3950 11520 3984
rect 11554 3950 11588 3984
rect 11622 3950 11656 3984
rect 11690 3950 11724 3984
rect 11758 3950 11792 3984
rect 11826 3950 11860 3984
rect 11894 3950 11928 3984
rect 11962 3950 11996 3984
rect 12030 3950 12064 3984
rect 12098 3950 12132 3984
rect 12166 3950 12200 3984
rect 12234 3950 12268 3984
rect 12302 3950 12336 3984
rect 12370 3950 12404 3984
rect 12438 3950 12472 3984
rect 12506 3950 12540 3984
rect 12574 3950 12608 3984
rect 12642 3950 12676 3984
rect 12710 3950 12744 3984
rect 12778 3950 12812 3984
rect 12846 3950 12880 3984
rect 12914 3950 12948 3984
rect 12982 3950 13016 3984
rect 13050 3950 13084 3984
rect 13118 3950 13152 3984
rect 13186 3950 13220 3984
rect 13254 3950 13288 3984
rect 13322 3950 13356 3984
rect 13390 3950 13424 3984
rect 13458 3950 13492 3984
rect 13526 3950 13560 3984
rect 13594 3950 13628 3984
rect 13662 3950 13696 3984
rect 13730 3950 13764 3984
rect 13798 3950 13832 3984
rect 13866 3950 13900 3984
rect 13934 3950 13968 3984
rect 14002 3950 14036 3984
rect 14070 3950 14104 3984
rect 14138 3950 14172 3984
rect 14206 3950 14240 3984
rect 14274 3950 14308 3984
rect 14342 3950 14376 3984
rect 14410 3950 14444 3984
rect 14478 3950 14512 3984
rect 14546 3950 14580 3984
rect 14614 3950 14648 3984
rect 14682 3950 14716 3984
rect 14750 3950 14784 3984
rect 14818 3950 14852 3984
rect 14886 3950 14920 3984
rect 14954 3950 14988 3984
rect 15022 3950 15056 3984
rect 15090 3950 15124 3984
rect 15158 3950 15192 3984
rect 15226 3950 15260 3984
rect 15294 3950 15328 3984
rect 15362 3950 15396 3984
rect 15430 3950 15464 3984
rect 15498 3950 15532 3984
rect 15566 3950 15600 3984
rect 15634 3950 15668 3984
rect 15702 3950 15736 3984
rect 15770 3950 15804 3984
rect 15838 3950 15872 3984
rect 15906 3950 15940 3984
rect 15974 3950 16008 3984
rect 16042 3950 16076 3984
rect 16110 3950 16144 3984
rect 16178 3950 16212 3984
rect 16246 3950 16280 3984
rect 16314 3950 16348 3984
rect 16382 3950 16416 3984
rect 16450 3950 16484 3984
rect 16518 3950 16552 3984
rect 16586 3950 16620 3984
rect 16654 3950 16688 3984
rect 16722 3950 16756 3984
rect 16790 3950 16824 3984
rect 16858 3950 16892 3984
rect 16926 3950 16960 3984
rect 16994 3950 17028 3984
rect 17062 3950 17096 3984
rect 17130 3950 17164 3984
rect 17198 3950 17232 3984
rect 17266 3950 17300 3984
rect 17334 3950 17368 3984
rect 17402 3950 17436 3984
rect 17470 3950 17504 3984
rect 17538 3950 17572 3984
rect 17606 3950 17640 3984
rect 17674 3950 17708 3984
rect 17742 3950 17776 3984
rect 17810 3950 17844 3984
rect 17878 3950 17912 3984
rect 17946 3950 17980 3984
rect 18014 3950 18048 3984
rect 18082 3950 18116 3984
rect 18150 3950 18184 3984
rect 18218 3950 18252 3984
rect 18286 3950 18320 3984
rect 18354 3950 18388 3984
rect 18422 3950 18456 3984
rect 18490 3950 18524 3984
rect 18558 3950 18592 3984
rect 18626 3950 18660 3984
rect 18694 3950 18728 3984
rect 18762 3950 18796 3984
rect 18830 3950 18864 3984
rect 18898 3950 18932 3984
rect 18966 3950 19000 3984
rect 19034 3950 19068 3984
rect 19102 3950 19136 3984
rect 19170 3950 19204 3984
rect 19238 3950 19272 3984
rect 19306 3950 19340 3984
rect 19374 3950 19408 3984
rect 19442 3950 19476 3984
rect 19510 3950 19544 3984
rect 19578 3950 19612 3984
rect 19646 3950 19680 3984
rect 19714 3950 19748 3984
rect 19782 3950 19816 3984
rect 19850 3950 19884 3984
rect 19918 3950 19952 3984
rect 19986 3950 20020 3984
rect 20054 3950 20088 3984
rect 20122 3950 20156 3984
rect 20190 3950 20224 3984
rect 20258 3950 20292 3984
rect 20326 3950 20360 3984
rect 20394 3950 20428 3984
rect 20462 3950 20496 3984
rect 20530 3950 20564 3984
rect 20598 3950 20632 3984
rect 20666 3950 20700 3984
rect 20734 3950 20768 3984
rect 20802 3950 20836 3984
rect 20870 3950 20904 3984
rect 20938 3950 20972 3984
rect 21006 3950 21040 3984
rect 21074 3950 21108 3984
rect 21142 3950 21176 3984
rect 21210 3950 21244 3984
rect 21278 3950 21312 3984
rect 21346 3950 21380 3984
rect 21414 3950 21448 3984
rect 21482 3950 21516 3984
rect 21550 3950 21584 3984
rect 21618 3950 21652 3984
rect 21686 3950 21720 3984
rect 21754 3950 21788 3984
rect 21822 3950 21856 3984
rect 21890 3950 21924 3984
rect 21958 3950 21992 3984
rect 22026 3950 22060 3984
rect 22094 3950 22128 3984
rect 22162 3950 22196 3984
rect 22230 3950 22264 3984
rect 22298 3950 22332 3984
rect 22366 3950 22400 3984
rect 22434 3950 22468 3984
rect 22502 3950 22536 3984
rect 22570 3950 22604 3984
rect 22638 3950 22672 3984
rect 22706 3950 22740 3984
rect 22774 3950 22808 3984
rect 22842 3950 22876 3984
rect 22910 3950 22944 3984
rect 22978 3950 23012 3984
rect 23046 3950 23080 3984
rect 23114 3950 23148 3984
rect 23182 3950 23216 3984
rect 23250 3950 23284 3984
rect 23318 3950 23352 3984
rect 23386 3950 23420 3984
rect 23454 3950 23488 3984
rect 23522 3950 23556 3984
rect 23590 3950 23624 3984
rect 23658 3950 23692 3984
rect 23726 3950 23760 3984
rect 23794 3950 23828 3984
rect 23862 3950 23896 3984
rect 23930 3950 23964 3984
rect 23998 3950 24032 3984
rect 24066 3950 24100 3984
rect 24134 3950 24168 3984
rect 24202 3950 24236 3984
rect 24270 3950 24304 3984
rect 24338 3950 24372 3984
rect 24406 3950 24440 3984
rect 24474 3950 24508 3984
rect 24542 3950 24576 3984
rect 24610 3950 24644 3984
rect 24678 3950 24712 3984
rect 24746 3950 24780 3984
rect 24814 3950 24848 3984
rect 24882 3950 24916 3984
rect 24950 3950 24984 3984
rect 25018 3950 25052 3984
rect 25086 3950 25120 3984
rect 25154 3950 25188 3984
rect 25222 3950 25256 3984
rect 25290 3950 25324 3984
rect 25358 3950 25392 3984
rect 25426 3950 25460 3984
rect 25494 3950 25528 3984
rect 25562 3950 25596 3984
rect 25630 3950 25664 3984
rect 25698 3950 25732 3984
rect 25766 3950 25800 3984
rect 25834 3950 25868 3984
rect 25902 3950 25936 3984
rect 25970 3950 26004 3984
rect 26038 3950 26072 3984
rect 26106 3950 26140 3984
rect 26174 3950 26208 3984
rect 26242 3950 26276 3984
rect 26310 3950 26344 3984
rect 26378 3950 26412 3984
rect 26446 3950 26480 3984
rect 26514 3950 26548 3984
rect 26582 3950 26616 3984
rect 26650 3950 26684 3984
rect 26718 3950 26752 3984
rect 26786 3950 26820 3984
rect 26854 3950 26888 3984
rect 26922 3950 26956 3984
rect 26990 3950 27024 3984
rect 27058 3950 27092 3984
rect 27126 3950 27160 3984
rect 27194 3950 27228 3984
rect 27262 3950 27296 3984
rect 27330 3950 27364 3984
rect 27398 3950 27432 3984
rect 27466 3950 27500 3984
rect 27534 3950 27568 3984
rect 27602 3950 27636 3984
rect 27670 3950 27704 3984
rect 27738 3950 27772 3984
rect 27806 3950 27840 3984
rect 27874 3950 27908 3984
rect 27942 3950 27976 3984
rect 6473 3876 6507 3910
rect 6542 3876 6576 3910
rect 6611 3876 6645 3910
rect 6680 3876 6714 3910
rect 6749 3876 6783 3910
rect 6818 3876 6852 3910
rect 6887 3876 6921 3910
rect 6956 3876 6990 3910
rect 7025 3876 7059 3910
rect 7094 3876 7128 3910
rect 7163 3876 7197 3910
rect 7232 3876 7266 3910
rect 7301 3876 7335 3910
rect 7370 3876 7404 3910
rect 7439 3876 7473 3910
rect 7508 3876 7542 3910
rect 7577 3876 7611 3910
rect 7646 3876 7680 3910
rect 7715 3876 7749 3910
rect 7784 3876 7818 3910
rect 7853 3876 7887 3910
rect 7922 3876 7956 3910
rect 7991 3876 8025 3910
rect 8060 3876 8094 3910
rect 8129 3876 8163 3910
rect 8198 3876 8232 3910
rect 8267 3876 8301 3910
rect 8336 3876 8370 3910
rect 8405 3876 8439 3910
rect 8474 3876 8508 3910
rect 8543 3876 8577 3910
rect 8612 3876 8646 3910
rect 8681 3876 8715 3910
rect 8750 3876 8784 3910
rect 8819 3876 8853 3910
rect 8888 3876 8922 3910
rect 8957 3876 8991 3910
rect 9026 3876 9060 3910
rect 9095 3876 9129 3910
rect 9164 3876 9198 3910
rect 9233 3876 9267 3910
rect 9302 3876 9336 3910
rect 9371 3876 9405 3910
rect 9440 3876 9474 3910
rect 9509 3876 9543 3910
rect 9578 3876 9612 3910
rect 9647 3876 9681 3910
rect 9716 3876 9750 3910
rect 9785 3876 9819 3910
rect 9854 3876 9888 3910
rect 9922 3876 9956 3910
rect 9990 3876 10024 3910
rect 10058 3876 10092 3910
rect 10126 3876 10160 3910
rect 10194 3876 10228 3910
rect 10262 3876 10296 3910
rect 10330 3876 10364 3910
rect 10398 3876 10432 3910
rect 10466 3876 10500 3910
rect 10534 3876 10568 3910
rect 10602 3876 10636 3910
rect 10670 3876 10704 3910
rect 10738 3876 10772 3910
rect 10806 3876 10840 3910
rect 10874 3876 10908 3910
rect 10942 3876 10976 3910
rect 11010 3876 11044 3910
rect 11078 3876 11112 3910
rect 11146 3876 11180 3910
rect 11214 3876 11248 3910
rect 11282 3876 11316 3910
rect 11350 3876 11384 3910
rect 11418 3876 11452 3910
rect 11486 3876 11520 3910
rect 11554 3876 11588 3910
rect 11622 3876 11656 3910
rect 11690 3876 11724 3910
rect 11758 3876 11792 3910
rect 11826 3876 11860 3910
rect 11894 3876 11928 3910
rect 11962 3876 11996 3910
rect 12030 3876 12064 3910
rect 12098 3876 12132 3910
rect 12166 3876 12200 3910
rect 12234 3876 12268 3910
rect 12302 3876 12336 3910
rect 12370 3876 12404 3910
rect 12438 3876 12472 3910
rect 12506 3876 12540 3910
rect 12574 3876 12608 3910
rect 12642 3876 12676 3910
rect 12710 3876 12744 3910
rect 12778 3876 12812 3910
rect 12846 3876 12880 3910
rect 12914 3876 12948 3910
rect 12982 3876 13016 3910
rect 13050 3876 13084 3910
rect 13118 3876 13152 3910
rect 13186 3876 13220 3910
rect 13254 3876 13288 3910
rect 13322 3876 13356 3910
rect 13390 3876 13424 3910
rect 13458 3876 13492 3910
rect 13526 3876 13560 3910
rect 13594 3876 13628 3910
rect 13662 3876 13696 3910
rect 13730 3876 13764 3910
rect 13798 3876 13832 3910
rect 13866 3876 13900 3910
rect 13934 3876 13968 3910
rect 14002 3876 14036 3910
rect 14070 3876 14104 3910
rect 14138 3876 14172 3910
rect 14206 3876 14240 3910
rect 14274 3876 14308 3910
rect 14342 3876 14376 3910
rect 14410 3876 14444 3910
rect 14478 3876 14512 3910
rect 14546 3876 14580 3910
rect 14614 3876 14648 3910
rect 14682 3876 14716 3910
rect 14750 3876 14784 3910
rect 14818 3876 14852 3910
rect 14886 3876 14920 3910
rect 14954 3876 14988 3910
rect 15022 3876 15056 3910
rect 15090 3876 15124 3910
rect 15158 3876 15192 3910
rect 15226 3876 15260 3910
rect 15294 3876 15328 3910
rect 15362 3876 15396 3910
rect 15430 3876 15464 3910
rect 15498 3876 15532 3910
rect 15566 3876 15600 3910
rect 15634 3876 15668 3910
rect 15702 3876 15736 3910
rect 15770 3876 15804 3910
rect 15838 3876 15872 3910
rect 15906 3876 15940 3910
rect 15974 3876 16008 3910
rect 16042 3876 16076 3910
rect 16110 3876 16144 3910
rect 16178 3876 16212 3910
rect 16246 3876 16280 3910
rect 16314 3876 16348 3910
rect 16382 3876 16416 3910
rect 16450 3876 16484 3910
rect 16518 3876 16552 3910
rect 16586 3876 16620 3910
rect 16654 3876 16688 3910
rect 16722 3876 16756 3910
rect 16790 3876 16824 3910
rect 16858 3876 16892 3910
rect 16926 3876 16960 3910
rect 16994 3876 17028 3910
rect 17062 3876 17096 3910
rect 17130 3876 17164 3910
rect 17198 3876 17232 3910
rect 17266 3876 17300 3910
rect 17334 3876 17368 3910
rect 17402 3876 17436 3910
rect 17470 3876 17504 3910
rect 17538 3876 17572 3910
rect 17606 3876 17640 3910
rect 17674 3876 17708 3910
rect 17742 3876 17776 3910
rect 17810 3876 17844 3910
rect 17878 3876 17912 3910
rect 17946 3876 17980 3910
rect 18014 3876 18048 3910
rect 18082 3876 18116 3910
rect 18150 3876 18184 3910
rect 18218 3876 18252 3910
rect 18286 3876 18320 3910
rect 18354 3876 18388 3910
rect 18422 3876 18456 3910
rect 18490 3876 18524 3910
rect 18558 3876 18592 3910
rect 18626 3876 18660 3910
rect 18694 3876 18728 3910
rect 18762 3876 18796 3910
rect 18830 3876 18864 3910
rect 18898 3876 18932 3910
rect 18966 3876 19000 3910
rect 19034 3876 19068 3910
rect 19102 3876 19136 3910
rect 19170 3876 19204 3910
rect 19238 3876 19272 3910
rect 19306 3876 19340 3910
rect 19374 3876 19408 3910
rect 19442 3876 19476 3910
rect 19510 3876 19544 3910
rect 19578 3876 19612 3910
rect 19646 3876 19680 3910
rect 19714 3876 19748 3910
rect 19782 3876 19816 3910
rect 19850 3876 19884 3910
rect 19918 3876 19952 3910
rect 19986 3876 20020 3910
rect 20054 3876 20088 3910
rect 20122 3876 20156 3910
rect 20190 3876 20224 3910
rect 20258 3876 20292 3910
rect 20326 3876 20360 3910
rect 20394 3876 20428 3910
rect 20462 3876 20496 3910
rect 20530 3876 20564 3910
rect 20598 3876 20632 3910
rect 20666 3876 20700 3910
rect 20734 3876 20768 3910
rect 20802 3876 20836 3910
rect 20870 3876 20904 3910
rect 20938 3876 20972 3910
rect 21006 3876 21040 3910
rect 21074 3876 21108 3910
rect 21142 3876 21176 3910
rect 21210 3876 21244 3910
rect 21278 3876 21312 3910
rect 21346 3876 21380 3910
rect 21414 3876 21448 3910
rect 21482 3876 21516 3910
rect 21550 3876 21584 3910
rect 21618 3876 21652 3910
rect 21686 3876 21720 3910
rect 21754 3876 21788 3910
rect 21822 3876 21856 3910
rect 21890 3876 21924 3910
rect 21958 3876 21992 3910
rect 22026 3876 22060 3910
rect 22094 3876 22128 3910
rect 22162 3876 22196 3910
rect 22230 3876 22264 3910
rect 22298 3876 22332 3910
rect 22366 3876 22400 3910
rect 22434 3876 22468 3910
rect 22502 3876 22536 3910
rect 22570 3876 22604 3910
rect 22638 3876 22672 3910
rect 22706 3876 22740 3910
rect 22774 3876 22808 3910
rect 22842 3876 22876 3910
rect 22910 3876 22944 3910
rect 22978 3876 23012 3910
rect 23046 3876 23080 3910
rect 23114 3876 23148 3910
rect 23182 3876 23216 3910
rect 23250 3876 23284 3910
rect 23318 3876 23352 3910
rect 23386 3876 23420 3910
rect 23454 3876 23488 3910
rect 23522 3876 23556 3910
rect 23590 3876 23624 3910
rect 23658 3876 23692 3910
rect 23726 3876 23760 3910
rect 23794 3876 23828 3910
rect 23862 3876 23896 3910
rect 23930 3876 23964 3910
rect 23998 3876 24032 3910
rect 24066 3876 24100 3910
rect 24134 3876 24168 3910
rect 24202 3876 24236 3910
rect 24270 3876 24304 3910
rect 24338 3876 24372 3910
rect 24406 3876 24440 3910
rect 24474 3876 24508 3910
rect 24542 3876 24576 3910
rect 24610 3876 24644 3910
rect 24678 3876 24712 3910
rect 24746 3876 24780 3910
rect 24814 3876 24848 3910
rect 24882 3876 24916 3910
rect 24950 3876 24984 3910
rect 25018 3876 25052 3910
rect 25086 3876 25120 3910
rect 25154 3876 25188 3910
rect 25222 3876 25256 3910
rect 25290 3876 25324 3910
rect 25358 3876 25392 3910
rect 25426 3876 25460 3910
rect 25494 3876 25528 3910
rect 25562 3876 25596 3910
rect 25630 3876 25664 3910
rect 25698 3876 25732 3910
rect 25766 3876 25800 3910
rect 25834 3876 25868 3910
rect 25902 3876 25936 3910
rect 25970 3876 26004 3910
rect 26038 3876 26072 3910
rect 26106 3876 26140 3910
rect 26174 3876 26208 3910
rect 26242 3876 26276 3910
rect 26310 3876 26344 3910
rect 26378 3876 26412 3910
rect 26446 3876 26480 3910
rect 26514 3876 26548 3910
rect 26582 3876 26616 3910
rect 26650 3876 26684 3910
rect 26718 3876 26752 3910
rect 26786 3876 26820 3910
rect 26854 3876 26888 3910
rect 26922 3876 26956 3910
rect 26990 3876 27024 3910
rect 27058 3876 27092 3910
rect 27126 3876 27160 3910
rect 27194 3876 27228 3910
rect 27262 3876 27296 3910
rect 27330 3876 27364 3910
rect 27398 3876 27432 3910
rect 27466 3876 27500 3910
rect 27534 3876 27568 3910
rect 27602 3876 27636 3910
rect 27670 3876 27704 3910
rect 27738 3876 27772 3910
rect 27806 3876 27840 3910
rect 27874 3876 27908 3910
rect 27942 3876 27976 3910
rect 6473 3802 6507 3836
rect 6542 3802 6576 3836
rect 6611 3802 6645 3836
rect 6680 3802 6714 3836
rect 6749 3802 6783 3836
rect 6818 3802 6852 3836
rect 6887 3802 6921 3836
rect 6956 3802 6990 3836
rect 7025 3802 7059 3836
rect 7094 3802 7128 3836
rect 7163 3802 7197 3836
rect 7232 3802 7266 3836
rect 7301 3802 7335 3836
rect 7370 3802 7404 3836
rect 7439 3802 7473 3836
rect 7508 3802 7542 3836
rect 7577 3802 7611 3836
rect 7646 3802 7680 3836
rect 7715 3802 7749 3836
rect 7784 3802 7818 3836
rect 7853 3802 7887 3836
rect 7922 3802 7956 3836
rect 7991 3802 8025 3836
rect 8060 3802 8094 3836
rect 8129 3802 8163 3836
rect 8198 3802 8232 3836
rect 8267 3802 8301 3836
rect 8336 3802 8370 3836
rect 8405 3802 8439 3836
rect 8474 3802 8508 3836
rect 8543 3802 8577 3836
rect 8612 3802 8646 3836
rect 8681 3802 8715 3836
rect 8750 3802 8784 3836
rect 8819 3802 8853 3836
rect 8888 3802 8922 3836
rect 8957 3802 8991 3836
rect 9026 3802 9060 3836
rect 9095 3802 9129 3836
rect 9164 3802 9198 3836
rect 9233 3802 9267 3836
rect 9302 3802 9336 3836
rect 9371 3802 9405 3836
rect 9440 3802 9474 3836
rect 9509 3802 9543 3836
rect 9578 3802 9612 3836
rect 9647 3802 9681 3836
rect 9716 3802 9750 3836
rect 9785 3802 9819 3836
rect 9854 3802 9888 3836
rect 9922 3802 9956 3836
rect 9990 3802 10024 3836
rect 10058 3802 10092 3836
rect 10126 3802 10160 3836
rect 10194 3802 10228 3836
rect 10262 3802 10296 3836
rect 10330 3802 10364 3836
rect 10398 3802 10432 3836
rect 10466 3802 10500 3836
rect 10534 3802 10568 3836
rect 10602 3802 10636 3836
rect 10670 3802 10704 3836
rect 10738 3802 10772 3836
rect 10806 3802 10840 3836
rect 10874 3802 10908 3836
rect 10942 3802 10976 3836
rect 11010 3802 11044 3836
rect 11078 3802 11112 3836
rect 11146 3802 11180 3836
rect 11214 3802 11248 3836
rect 11282 3802 11316 3836
rect 11350 3802 11384 3836
rect 11418 3802 11452 3836
rect 11486 3802 11520 3836
rect 11554 3802 11588 3836
rect 11622 3802 11656 3836
rect 11690 3802 11724 3836
rect 11758 3802 11792 3836
rect 11826 3802 11860 3836
rect 11894 3802 11928 3836
rect 11962 3802 11996 3836
rect 12030 3802 12064 3836
rect 12098 3802 12132 3836
rect 12166 3802 12200 3836
rect 12234 3802 12268 3836
rect 12302 3802 12336 3836
rect 12370 3802 12404 3836
rect 12438 3802 12472 3836
rect 12506 3802 12540 3836
rect 12574 3802 12608 3836
rect 12642 3802 12676 3836
rect 12710 3802 12744 3836
rect 12778 3802 12812 3836
rect 12846 3802 12880 3836
rect 12914 3802 12948 3836
rect 12982 3802 13016 3836
rect 13050 3802 13084 3836
rect 13118 3802 13152 3836
rect 13186 3802 13220 3836
rect 13254 3802 13288 3836
rect 13322 3802 13356 3836
rect 13390 3802 13424 3836
rect 13458 3802 13492 3836
rect 13526 3802 13560 3836
rect 13594 3802 13628 3836
rect 13662 3802 13696 3836
rect 13730 3802 13764 3836
rect 13798 3802 13832 3836
rect 13866 3802 13900 3836
rect 13934 3802 13968 3836
rect 14002 3802 14036 3836
rect 14070 3802 14104 3836
rect 14138 3802 14172 3836
rect 14206 3802 14240 3836
rect 14274 3802 14308 3836
rect 14342 3802 14376 3836
rect 14410 3802 14444 3836
rect 14478 3802 14512 3836
rect 14546 3802 14580 3836
rect 14614 3802 14648 3836
rect 14682 3802 14716 3836
rect 14750 3802 14784 3836
rect 14818 3802 14852 3836
rect 14886 3802 14920 3836
rect 14954 3802 14988 3836
rect 15022 3802 15056 3836
rect 15090 3802 15124 3836
rect 15158 3802 15192 3836
rect 15226 3802 15260 3836
rect 15294 3802 15328 3836
rect 15362 3802 15396 3836
rect 15430 3802 15464 3836
rect 15498 3802 15532 3836
rect 15566 3802 15600 3836
rect 15634 3802 15668 3836
rect 15702 3802 15736 3836
rect 15770 3802 15804 3836
rect 15838 3802 15872 3836
rect 15906 3802 15940 3836
rect 15974 3802 16008 3836
rect 16042 3802 16076 3836
rect 16110 3802 16144 3836
rect 16178 3802 16212 3836
rect 16246 3802 16280 3836
rect 16314 3802 16348 3836
rect 16382 3802 16416 3836
rect 16450 3802 16484 3836
rect 16518 3802 16552 3836
rect 16586 3802 16620 3836
rect 16654 3802 16688 3836
rect 16722 3802 16756 3836
rect 16790 3802 16824 3836
rect 16858 3802 16892 3836
rect 16926 3802 16960 3836
rect 16994 3802 17028 3836
rect 17062 3802 17096 3836
rect 17130 3802 17164 3836
rect 17198 3802 17232 3836
rect 17266 3802 17300 3836
rect 17334 3802 17368 3836
rect 17402 3802 17436 3836
rect 17470 3802 17504 3836
rect 17538 3802 17572 3836
rect 17606 3802 17640 3836
rect 17674 3802 17708 3836
rect 17742 3802 17776 3836
rect 17810 3802 17844 3836
rect 17878 3802 17912 3836
rect 17946 3802 17980 3836
rect 18014 3802 18048 3836
rect 18082 3802 18116 3836
rect 18150 3802 18184 3836
rect 18218 3802 18252 3836
rect 18286 3802 18320 3836
rect 18354 3802 18388 3836
rect 18422 3802 18456 3836
rect 18490 3802 18524 3836
rect 18558 3802 18592 3836
rect 18626 3802 18660 3836
rect 18694 3802 18728 3836
rect 18762 3802 18796 3836
rect 18830 3802 18864 3836
rect 18898 3802 18932 3836
rect 18966 3802 19000 3836
rect 19034 3802 19068 3836
rect 19102 3802 19136 3836
rect 19170 3802 19204 3836
rect 19238 3802 19272 3836
rect 19306 3802 19340 3836
rect 19374 3802 19408 3836
rect 19442 3802 19476 3836
rect 19510 3802 19544 3836
rect 19578 3802 19612 3836
rect 19646 3802 19680 3836
rect 19714 3802 19748 3836
rect 19782 3802 19816 3836
rect 19850 3802 19884 3836
rect 19918 3802 19952 3836
rect 19986 3802 20020 3836
rect 20054 3802 20088 3836
rect 20122 3802 20156 3836
rect 20190 3802 20224 3836
rect 20258 3802 20292 3836
rect 20326 3802 20360 3836
rect 20394 3802 20428 3836
rect 20462 3802 20496 3836
rect 20530 3802 20564 3836
rect 20598 3802 20632 3836
rect 20666 3802 20700 3836
rect 20734 3802 20768 3836
rect 20802 3802 20836 3836
rect 20870 3802 20904 3836
rect 20938 3802 20972 3836
rect 21006 3802 21040 3836
rect 21074 3802 21108 3836
rect 21142 3802 21176 3836
rect 21210 3802 21244 3836
rect 21278 3802 21312 3836
rect 21346 3802 21380 3836
rect 21414 3802 21448 3836
rect 21482 3802 21516 3836
rect 21550 3802 21584 3836
rect 21618 3802 21652 3836
rect 21686 3802 21720 3836
rect 21754 3802 21788 3836
rect 21822 3802 21856 3836
rect 21890 3802 21924 3836
rect 21958 3802 21992 3836
rect 22026 3802 22060 3836
rect 22094 3802 22128 3836
rect 22162 3802 22196 3836
rect 22230 3802 22264 3836
rect 22298 3802 22332 3836
rect 22366 3802 22400 3836
rect 22434 3802 22468 3836
rect 22502 3802 22536 3836
rect 22570 3802 22604 3836
rect 22638 3802 22672 3836
rect 22706 3802 22740 3836
rect 22774 3802 22808 3836
rect 22842 3802 22876 3836
rect 22910 3802 22944 3836
rect 22978 3802 23012 3836
rect 23046 3802 23080 3836
rect 23114 3802 23148 3836
rect 23182 3802 23216 3836
rect 23250 3802 23284 3836
rect 23318 3802 23352 3836
rect 23386 3802 23420 3836
rect 23454 3802 23488 3836
rect 23522 3802 23556 3836
rect 23590 3802 23624 3836
rect 23658 3802 23692 3836
rect 23726 3802 23760 3836
rect 23794 3802 23828 3836
rect 23862 3802 23896 3836
rect 23930 3802 23964 3836
rect 23998 3802 24032 3836
rect 24066 3802 24100 3836
rect 24134 3802 24168 3836
rect 24202 3802 24236 3836
rect 24270 3802 24304 3836
rect 24338 3802 24372 3836
rect 24406 3802 24440 3836
rect 24474 3802 24508 3836
rect 24542 3802 24576 3836
rect 24610 3802 24644 3836
rect 24678 3802 24712 3836
rect 24746 3802 24780 3836
rect 24814 3802 24848 3836
rect 24882 3802 24916 3836
rect 24950 3802 24984 3836
rect 25018 3802 25052 3836
rect 25086 3802 25120 3836
rect 25154 3802 25188 3836
rect 25222 3802 25256 3836
rect 25290 3802 25324 3836
rect 25358 3802 25392 3836
rect 25426 3802 25460 3836
rect 25494 3802 25528 3836
rect 25562 3802 25596 3836
rect 25630 3802 25664 3836
rect 25698 3802 25732 3836
rect 25766 3802 25800 3836
rect 25834 3802 25868 3836
rect 25902 3802 25936 3836
rect 25970 3802 26004 3836
rect 26038 3802 26072 3836
rect 26106 3802 26140 3836
rect 26174 3802 26208 3836
rect 26242 3802 26276 3836
rect 26310 3802 26344 3836
rect 26378 3802 26412 3836
rect 26446 3802 26480 3836
rect 26514 3802 26548 3836
rect 26582 3802 26616 3836
rect 26650 3802 26684 3836
rect 26718 3802 26752 3836
rect 26786 3802 26820 3836
rect 26854 3802 26888 3836
rect 26922 3802 26956 3836
rect 26990 3802 27024 3836
rect 27058 3802 27092 3836
rect 27126 3802 27160 3836
rect 27194 3802 27228 3836
rect 27262 3802 27296 3836
rect 27330 3802 27364 3836
rect 27398 3802 27432 3836
rect 27466 3802 27500 3836
rect 27534 3802 27568 3836
rect 27602 3802 27636 3836
rect 27670 3802 27704 3836
rect 27738 3802 27772 3836
rect 27806 3802 27840 3836
rect 27874 3802 27908 3836
rect 27942 3802 27976 3836
rect 2344 3654 2378 3688
rect 2415 3654 2449 3688
rect 2486 3654 2520 3688
rect 2557 3654 2591 3688
rect 2628 3654 2662 3688
rect 2698 3654 2732 3688
rect 2768 3654 2802 3688
rect 2838 3654 2872 3688
rect 2908 3654 2942 3688
rect 2978 3654 3012 3688
rect 3048 3654 3082 3688
rect 3118 3654 3152 3688
rect 3188 3654 3222 3688
rect 3258 3654 3292 3688
rect 2344 3580 2378 3614
rect 2415 3580 2449 3614
rect 2486 3580 2520 3614
rect 2557 3580 2591 3614
rect 2628 3580 2662 3614
rect 2698 3580 2732 3614
rect 2768 3580 2802 3614
rect 2838 3580 2872 3614
rect 2908 3580 2942 3614
rect 2978 3580 3012 3614
rect 3048 3580 3082 3614
rect 3118 3580 3152 3614
rect 3188 3580 3222 3614
rect 3258 3580 3292 3614
rect 2344 3506 2378 3540
rect 2415 3506 2449 3540
rect 2486 3506 2520 3540
rect 2557 3506 2591 3540
rect 2628 3506 2662 3540
rect 2698 3506 2732 3540
rect 2768 3506 2802 3540
rect 2838 3506 2872 3540
rect 2908 3506 2942 3540
rect 2978 3506 3012 3540
rect 3048 3506 3082 3540
rect 3118 3506 3152 3540
rect 3188 3506 3222 3540
rect 3258 3506 3292 3540
rect 2344 3432 2378 3466
rect 2415 3432 2449 3466
rect 2486 3432 2520 3466
rect 2557 3432 2591 3466
rect 2628 3432 2662 3466
rect 2698 3432 2732 3466
rect 2768 3432 2802 3466
rect 2838 3432 2872 3466
rect 2908 3432 2942 3466
rect 2978 3432 3012 3466
rect 3048 3432 3082 3466
rect 3118 3432 3152 3466
rect 3188 3432 3222 3466
rect 3258 3432 3292 3466
rect 6473 3728 6507 3762
rect 6542 3728 6576 3762
rect 6611 3728 6645 3762
rect 6680 3728 6714 3762
rect 6749 3728 6783 3762
rect 6818 3728 6852 3762
rect 6887 3728 6921 3762
rect 6956 3728 6990 3762
rect 7025 3728 7059 3762
rect 7094 3728 7128 3762
rect 7163 3728 7197 3762
rect 7232 3728 7266 3762
rect 7301 3728 7335 3762
rect 7370 3728 7404 3762
rect 7439 3728 7473 3762
rect 7508 3728 7542 3762
rect 7577 3728 7611 3762
rect 7646 3728 7680 3762
rect 7715 3728 7749 3762
rect 7784 3728 7818 3762
rect 7853 3728 7887 3762
rect 7922 3728 7956 3762
rect 7991 3728 8025 3762
rect 8060 3728 8094 3762
rect 8129 3728 8163 3762
rect 8198 3728 8232 3762
rect 8267 3728 8301 3762
rect 8336 3728 8370 3762
rect 8405 3728 8439 3762
rect 8474 3728 8508 3762
rect 8543 3728 8577 3762
rect 8612 3728 8646 3762
rect 8681 3728 8715 3762
rect 8750 3728 8784 3762
rect 8819 3728 8853 3762
rect 8888 3728 8922 3762
rect 8957 3728 8991 3762
rect 9026 3728 9060 3762
rect 9095 3728 9129 3762
rect 9164 3728 9198 3762
rect 9233 3728 9267 3762
rect 9302 3728 9336 3762
rect 9371 3728 9405 3762
rect 9440 3728 9474 3762
rect 9509 3728 9543 3762
rect 9578 3728 9612 3762
rect 9647 3728 9681 3762
rect 9716 3728 9750 3762
rect 9785 3728 9819 3762
rect 9854 3728 9888 3762
rect 9922 3728 9956 3762
rect 9990 3728 10024 3762
rect 10058 3728 10092 3762
rect 10126 3728 10160 3762
rect 10194 3728 10228 3762
rect 10262 3728 10296 3762
rect 10330 3728 10364 3762
rect 10398 3728 10432 3762
rect 10466 3728 10500 3762
rect 10534 3728 10568 3762
rect 10602 3728 10636 3762
rect 10670 3728 10704 3762
rect 10738 3728 10772 3762
rect 10806 3728 10840 3762
rect 10874 3728 10908 3762
rect 10942 3728 10976 3762
rect 11010 3728 11044 3762
rect 11078 3728 11112 3762
rect 11146 3728 11180 3762
rect 11214 3728 11248 3762
rect 11282 3728 11316 3762
rect 11350 3728 11384 3762
rect 11418 3728 11452 3762
rect 11486 3728 11520 3762
rect 11554 3728 11588 3762
rect 11622 3728 11656 3762
rect 11690 3728 11724 3762
rect 11758 3728 11792 3762
rect 11826 3728 11860 3762
rect 11894 3728 11928 3762
rect 11962 3728 11996 3762
rect 12030 3728 12064 3762
rect 12098 3728 12132 3762
rect 12166 3728 12200 3762
rect 12234 3728 12268 3762
rect 12302 3728 12336 3762
rect 12370 3728 12404 3762
rect 12438 3728 12472 3762
rect 12506 3728 12540 3762
rect 12574 3728 12608 3762
rect 12642 3728 12676 3762
rect 12710 3728 12744 3762
rect 12778 3728 12812 3762
rect 12846 3728 12880 3762
rect 12914 3728 12948 3762
rect 12982 3728 13016 3762
rect 13050 3728 13084 3762
rect 13118 3728 13152 3762
rect 13186 3728 13220 3762
rect 13254 3728 13288 3762
rect 13322 3728 13356 3762
rect 13390 3728 13424 3762
rect 13458 3728 13492 3762
rect 13526 3728 13560 3762
rect 13594 3728 13628 3762
rect 13662 3728 13696 3762
rect 13730 3728 13764 3762
rect 13798 3728 13832 3762
rect 13866 3728 13900 3762
rect 13934 3728 13968 3762
rect 14002 3728 14036 3762
rect 14070 3728 14104 3762
rect 14138 3728 14172 3762
rect 14206 3728 14240 3762
rect 14274 3728 14308 3762
rect 14342 3728 14376 3762
rect 14410 3728 14444 3762
rect 14478 3728 14512 3762
rect 14546 3728 14580 3762
rect 14614 3728 14648 3762
rect 14682 3728 14716 3762
rect 14750 3728 14784 3762
rect 14818 3728 14852 3762
rect 14886 3728 14920 3762
rect 14954 3728 14988 3762
rect 15022 3728 15056 3762
rect 15090 3728 15124 3762
rect 15158 3728 15192 3762
rect 15226 3728 15260 3762
rect 15294 3728 15328 3762
rect 15362 3728 15396 3762
rect 15430 3728 15464 3762
rect 15498 3728 15532 3762
rect 15566 3728 15600 3762
rect 15634 3728 15668 3762
rect 15702 3728 15736 3762
rect 15770 3728 15804 3762
rect 15838 3728 15872 3762
rect 15906 3728 15940 3762
rect 15974 3728 16008 3762
rect 16042 3728 16076 3762
rect 16110 3728 16144 3762
rect 16178 3728 16212 3762
rect 16246 3728 16280 3762
rect 16314 3728 16348 3762
rect 16382 3728 16416 3762
rect 16450 3728 16484 3762
rect 16518 3728 16552 3762
rect 16586 3728 16620 3762
rect 16654 3728 16688 3762
rect 16722 3728 16756 3762
rect 16790 3728 16824 3762
rect 16858 3728 16892 3762
rect 16926 3728 16960 3762
rect 16994 3728 17028 3762
rect 17062 3728 17096 3762
rect 17130 3728 17164 3762
rect 17198 3728 17232 3762
rect 17266 3728 17300 3762
rect 17334 3728 17368 3762
rect 17402 3728 17436 3762
rect 17470 3728 17504 3762
rect 17538 3728 17572 3762
rect 17606 3728 17640 3762
rect 17674 3728 17708 3762
rect 17742 3728 17776 3762
rect 17810 3728 17844 3762
rect 17878 3728 17912 3762
rect 17946 3728 17980 3762
rect 18014 3728 18048 3762
rect 18082 3728 18116 3762
rect 18150 3728 18184 3762
rect 18218 3728 18252 3762
rect 18286 3728 18320 3762
rect 18354 3728 18388 3762
rect 18422 3728 18456 3762
rect 18490 3728 18524 3762
rect 18558 3728 18592 3762
rect 18626 3728 18660 3762
rect 18694 3728 18728 3762
rect 18762 3728 18796 3762
rect 18830 3728 18864 3762
rect 18898 3728 18932 3762
rect 18966 3728 19000 3762
rect 19034 3728 19068 3762
rect 19102 3728 19136 3762
rect 19170 3728 19204 3762
rect 19238 3728 19272 3762
rect 19306 3728 19340 3762
rect 19374 3728 19408 3762
rect 19442 3728 19476 3762
rect 19510 3728 19544 3762
rect 19578 3728 19612 3762
rect 19646 3728 19680 3762
rect 19714 3728 19748 3762
rect 19782 3728 19816 3762
rect 19850 3728 19884 3762
rect 19918 3728 19952 3762
rect 19986 3728 20020 3762
rect 20054 3728 20088 3762
rect 20122 3728 20156 3762
rect 20190 3728 20224 3762
rect 20258 3728 20292 3762
rect 20326 3728 20360 3762
rect 20394 3728 20428 3762
rect 20462 3728 20496 3762
rect 20530 3728 20564 3762
rect 20598 3728 20632 3762
rect 20666 3728 20700 3762
rect 20734 3728 20768 3762
rect 20802 3728 20836 3762
rect 20870 3728 20904 3762
rect 20938 3728 20972 3762
rect 21006 3728 21040 3762
rect 21074 3728 21108 3762
rect 21142 3728 21176 3762
rect 21210 3728 21244 3762
rect 21278 3728 21312 3762
rect 21346 3728 21380 3762
rect 21414 3728 21448 3762
rect 21482 3728 21516 3762
rect 21550 3728 21584 3762
rect 21618 3728 21652 3762
rect 21686 3728 21720 3762
rect 21754 3728 21788 3762
rect 21822 3728 21856 3762
rect 21890 3728 21924 3762
rect 21958 3728 21992 3762
rect 22026 3728 22060 3762
rect 22094 3728 22128 3762
rect 22162 3728 22196 3762
rect 22230 3728 22264 3762
rect 22298 3728 22332 3762
rect 22366 3728 22400 3762
rect 22434 3728 22468 3762
rect 22502 3728 22536 3762
rect 22570 3728 22604 3762
rect 22638 3728 22672 3762
rect 22706 3728 22740 3762
rect 22774 3728 22808 3762
rect 22842 3728 22876 3762
rect 22910 3728 22944 3762
rect 22978 3728 23012 3762
rect 23046 3728 23080 3762
rect 23114 3728 23148 3762
rect 23182 3728 23216 3762
rect 23250 3728 23284 3762
rect 23318 3728 23352 3762
rect 23386 3728 23420 3762
rect 23454 3728 23488 3762
rect 23522 3728 23556 3762
rect 23590 3728 23624 3762
rect 23658 3728 23692 3762
rect 23726 3728 23760 3762
rect 23794 3728 23828 3762
rect 23862 3728 23896 3762
rect 23930 3728 23964 3762
rect 23998 3728 24032 3762
rect 24066 3728 24100 3762
rect 24134 3728 24168 3762
rect 24202 3728 24236 3762
rect 24270 3728 24304 3762
rect 24338 3728 24372 3762
rect 24406 3728 24440 3762
rect 24474 3728 24508 3762
rect 24542 3728 24576 3762
rect 24610 3728 24644 3762
rect 24678 3728 24712 3762
rect 24746 3728 24780 3762
rect 24814 3728 24848 3762
rect 24882 3728 24916 3762
rect 24950 3728 24984 3762
rect 25018 3728 25052 3762
rect 25086 3728 25120 3762
rect 25154 3728 25188 3762
rect 25222 3728 25256 3762
rect 25290 3728 25324 3762
rect 25358 3728 25392 3762
rect 25426 3728 25460 3762
rect 25494 3728 25528 3762
rect 25562 3728 25596 3762
rect 25630 3728 25664 3762
rect 25698 3728 25732 3762
rect 25766 3728 25800 3762
rect 25834 3728 25868 3762
rect 25902 3728 25936 3762
rect 25970 3728 26004 3762
rect 26038 3728 26072 3762
rect 26106 3728 26140 3762
rect 26174 3728 26208 3762
rect 26242 3728 26276 3762
rect 26310 3728 26344 3762
rect 26378 3728 26412 3762
rect 26446 3728 26480 3762
rect 26514 3728 26548 3762
rect 26582 3728 26616 3762
rect 26650 3728 26684 3762
rect 26718 3728 26752 3762
rect 26786 3728 26820 3762
rect 26854 3728 26888 3762
rect 26922 3728 26956 3762
rect 26990 3728 27024 3762
rect 27058 3728 27092 3762
rect 27126 3728 27160 3762
rect 27194 3728 27228 3762
rect 27262 3728 27296 3762
rect 27330 3728 27364 3762
rect 27398 3728 27432 3762
rect 27466 3728 27500 3762
rect 27534 3728 27568 3762
rect 27602 3728 27636 3762
rect 27670 3728 27704 3762
rect 27738 3728 27772 3762
rect 27806 3728 27840 3762
rect 27874 3728 27908 3762
rect 27942 3728 27976 3762
rect 6473 3654 6507 3688
rect 6542 3654 6576 3688
rect 6611 3654 6645 3688
rect 6680 3654 6714 3688
rect 6749 3654 6783 3688
rect 6818 3654 6852 3688
rect 6887 3654 6921 3688
rect 6956 3654 6990 3688
rect 7025 3654 7059 3688
rect 7094 3654 7128 3688
rect 7163 3654 7197 3688
rect 7232 3654 7266 3688
rect 7301 3654 7335 3688
rect 7370 3654 7404 3688
rect 7439 3654 7473 3688
rect 7508 3654 7542 3688
rect 7577 3654 7611 3688
rect 7646 3654 7680 3688
rect 7715 3654 7749 3688
rect 7784 3654 7818 3688
rect 7853 3654 7887 3688
rect 7922 3654 7956 3688
rect 7991 3654 8025 3688
rect 8060 3654 8094 3688
rect 8129 3654 8163 3688
rect 8198 3654 8232 3688
rect 8267 3654 8301 3688
rect 8336 3654 8370 3688
rect 8405 3654 8439 3688
rect 8474 3654 8508 3688
rect 8543 3654 8577 3688
rect 8612 3654 8646 3688
rect 8681 3654 8715 3688
rect 8750 3654 8784 3688
rect 8819 3654 8853 3688
rect 8888 3654 8922 3688
rect 8957 3654 8991 3688
rect 9026 3654 9060 3688
rect 9095 3654 9129 3688
rect 9164 3654 9198 3688
rect 9233 3654 9267 3688
rect 9302 3654 9336 3688
rect 9371 3654 9405 3688
rect 9440 3654 9474 3688
rect 9509 3654 9543 3688
rect 9578 3654 9612 3688
rect 9647 3654 9681 3688
rect 9716 3654 9750 3688
rect 9785 3654 9819 3688
rect 9854 3654 9888 3688
rect 9922 3654 9956 3688
rect 9990 3654 10024 3688
rect 10058 3654 10092 3688
rect 10126 3654 10160 3688
rect 10194 3654 10228 3688
rect 10262 3654 10296 3688
rect 10330 3654 10364 3688
rect 10398 3654 10432 3688
rect 10466 3654 10500 3688
rect 10534 3654 10568 3688
rect 10602 3654 10636 3688
rect 10670 3654 10704 3688
rect 10738 3654 10772 3688
rect 10806 3654 10840 3688
rect 10874 3654 10908 3688
rect 10942 3654 10976 3688
rect 11010 3654 11044 3688
rect 11078 3654 11112 3688
rect 11146 3654 11180 3688
rect 11214 3654 11248 3688
rect 11282 3654 11316 3688
rect 11350 3654 11384 3688
rect 11418 3654 11452 3688
rect 11486 3654 11520 3688
rect 11554 3654 11588 3688
rect 11622 3654 11656 3688
rect 11690 3654 11724 3688
rect 11758 3654 11792 3688
rect 11826 3654 11860 3688
rect 11894 3654 11928 3688
rect 11962 3654 11996 3688
rect 12030 3654 12064 3688
rect 12098 3654 12132 3688
rect 12166 3654 12200 3688
rect 12234 3654 12268 3688
rect 12302 3654 12336 3688
rect 12370 3654 12404 3688
rect 12438 3654 12472 3688
rect 12506 3654 12540 3688
rect 12574 3654 12608 3688
rect 12642 3654 12676 3688
rect 12710 3654 12744 3688
rect 12778 3654 12812 3688
rect 12846 3654 12880 3688
rect 12914 3654 12948 3688
rect 12982 3654 13016 3688
rect 13050 3654 13084 3688
rect 13118 3654 13152 3688
rect 13186 3654 13220 3688
rect 13254 3654 13288 3688
rect 13322 3654 13356 3688
rect 13390 3654 13424 3688
rect 13458 3654 13492 3688
rect 13526 3654 13560 3688
rect 13594 3654 13628 3688
rect 13662 3654 13696 3688
rect 13730 3654 13764 3688
rect 13798 3654 13832 3688
rect 13866 3654 13900 3688
rect 13934 3654 13968 3688
rect 14002 3654 14036 3688
rect 14070 3654 14104 3688
rect 14138 3654 14172 3688
rect 14206 3654 14240 3688
rect 14274 3654 14308 3688
rect 14342 3654 14376 3688
rect 14410 3654 14444 3688
rect 14478 3654 14512 3688
rect 14546 3654 14580 3688
rect 14614 3654 14648 3688
rect 14682 3654 14716 3688
rect 14750 3654 14784 3688
rect 14818 3654 14852 3688
rect 14886 3654 14920 3688
rect 14954 3654 14988 3688
rect 15022 3654 15056 3688
rect 15090 3654 15124 3688
rect 15158 3654 15192 3688
rect 15226 3654 15260 3688
rect 15294 3654 15328 3688
rect 15362 3654 15396 3688
rect 15430 3654 15464 3688
rect 15498 3654 15532 3688
rect 15566 3654 15600 3688
rect 15634 3654 15668 3688
rect 15702 3654 15736 3688
rect 15770 3654 15804 3688
rect 15838 3654 15872 3688
rect 15906 3654 15940 3688
rect 15974 3654 16008 3688
rect 16042 3654 16076 3688
rect 16110 3654 16144 3688
rect 16178 3654 16212 3688
rect 16246 3654 16280 3688
rect 16314 3654 16348 3688
rect 16382 3654 16416 3688
rect 16450 3654 16484 3688
rect 16518 3654 16552 3688
rect 16586 3654 16620 3688
rect 16654 3654 16688 3688
rect 16722 3654 16756 3688
rect 16790 3654 16824 3688
rect 16858 3654 16892 3688
rect 16926 3654 16960 3688
rect 16994 3654 17028 3688
rect 17062 3654 17096 3688
rect 17130 3654 17164 3688
rect 17198 3654 17232 3688
rect 17266 3654 17300 3688
rect 17334 3654 17368 3688
rect 17402 3654 17436 3688
rect 17470 3654 17504 3688
rect 17538 3654 17572 3688
rect 17606 3654 17640 3688
rect 17674 3654 17708 3688
rect 17742 3654 17776 3688
rect 17810 3654 17844 3688
rect 17878 3654 17912 3688
rect 17946 3654 17980 3688
rect 18014 3654 18048 3688
rect 18082 3654 18116 3688
rect 18150 3654 18184 3688
rect 18218 3654 18252 3688
rect 18286 3654 18320 3688
rect 18354 3654 18388 3688
rect 18422 3654 18456 3688
rect 18490 3654 18524 3688
rect 18558 3654 18592 3688
rect 18626 3654 18660 3688
rect 18694 3654 18728 3688
rect 18762 3654 18796 3688
rect 18830 3654 18864 3688
rect 18898 3654 18932 3688
rect 18966 3654 19000 3688
rect 19034 3654 19068 3688
rect 19102 3654 19136 3688
rect 19170 3654 19204 3688
rect 19238 3654 19272 3688
rect 19306 3654 19340 3688
rect 19374 3654 19408 3688
rect 19442 3654 19476 3688
rect 19510 3654 19544 3688
rect 19578 3654 19612 3688
rect 19646 3654 19680 3688
rect 19714 3654 19748 3688
rect 19782 3654 19816 3688
rect 19850 3654 19884 3688
rect 19918 3654 19952 3688
rect 19986 3654 20020 3688
rect 20054 3654 20088 3688
rect 20122 3654 20156 3688
rect 20190 3654 20224 3688
rect 20258 3654 20292 3688
rect 20326 3654 20360 3688
rect 20394 3654 20428 3688
rect 20462 3654 20496 3688
rect 20530 3654 20564 3688
rect 20598 3654 20632 3688
rect 20666 3654 20700 3688
rect 20734 3654 20768 3688
rect 20802 3654 20836 3688
rect 20870 3654 20904 3688
rect 20938 3654 20972 3688
rect 21006 3654 21040 3688
rect 21074 3654 21108 3688
rect 21142 3654 21176 3688
rect 21210 3654 21244 3688
rect 21278 3654 21312 3688
rect 21346 3654 21380 3688
rect 21414 3654 21448 3688
rect 21482 3654 21516 3688
rect 21550 3654 21584 3688
rect 21618 3654 21652 3688
rect 21686 3654 21720 3688
rect 21754 3654 21788 3688
rect 21822 3654 21856 3688
rect 21890 3654 21924 3688
rect 21958 3654 21992 3688
rect 22026 3654 22060 3688
rect 22094 3654 22128 3688
rect 22162 3654 22196 3688
rect 22230 3654 22264 3688
rect 22298 3654 22332 3688
rect 22366 3654 22400 3688
rect 22434 3654 22468 3688
rect 22502 3654 22536 3688
rect 22570 3654 22604 3688
rect 22638 3654 22672 3688
rect 22706 3654 22740 3688
rect 22774 3654 22808 3688
rect 22842 3654 22876 3688
rect 22910 3654 22944 3688
rect 22978 3654 23012 3688
rect 23046 3654 23080 3688
rect 23114 3654 23148 3688
rect 23182 3654 23216 3688
rect 23250 3654 23284 3688
rect 23318 3654 23352 3688
rect 23386 3654 23420 3688
rect 23454 3654 23488 3688
rect 23522 3654 23556 3688
rect 23590 3654 23624 3688
rect 23658 3654 23692 3688
rect 23726 3654 23760 3688
rect 23794 3654 23828 3688
rect 23862 3654 23896 3688
rect 23930 3654 23964 3688
rect 23998 3654 24032 3688
rect 24066 3654 24100 3688
rect 24134 3654 24168 3688
rect 24202 3654 24236 3688
rect 24270 3654 24304 3688
rect 24338 3654 24372 3688
rect 24406 3654 24440 3688
rect 24474 3654 24508 3688
rect 24542 3654 24576 3688
rect 24610 3654 24644 3688
rect 24678 3654 24712 3688
rect 24746 3654 24780 3688
rect 24814 3654 24848 3688
rect 24882 3654 24916 3688
rect 24950 3654 24984 3688
rect 25018 3654 25052 3688
rect 25086 3654 25120 3688
rect 25154 3654 25188 3688
rect 25222 3654 25256 3688
rect 25290 3654 25324 3688
rect 25358 3654 25392 3688
rect 25426 3654 25460 3688
rect 25494 3654 25528 3688
rect 25562 3654 25596 3688
rect 25630 3654 25664 3688
rect 25698 3654 25732 3688
rect 25766 3654 25800 3688
rect 25834 3654 25868 3688
rect 25902 3654 25936 3688
rect 25970 3654 26004 3688
rect 26038 3654 26072 3688
rect 26106 3654 26140 3688
rect 26174 3654 26208 3688
rect 26242 3654 26276 3688
rect 26310 3654 26344 3688
rect 26378 3654 26412 3688
rect 26446 3654 26480 3688
rect 26514 3654 26548 3688
rect 26582 3654 26616 3688
rect 26650 3654 26684 3688
rect 26718 3654 26752 3688
rect 26786 3654 26820 3688
rect 26854 3654 26888 3688
rect 26922 3654 26956 3688
rect 26990 3654 27024 3688
rect 27058 3654 27092 3688
rect 27126 3654 27160 3688
rect 27194 3654 27228 3688
rect 27262 3654 27296 3688
rect 27330 3654 27364 3688
rect 27398 3654 27432 3688
rect 27466 3654 27500 3688
rect 27534 3654 27568 3688
rect 27602 3654 27636 3688
rect 27670 3654 27704 3688
rect 27738 3654 27772 3688
rect 27806 3654 27840 3688
rect 27874 3654 27908 3688
rect 27942 3654 27976 3688
rect 6473 3580 6507 3614
rect 6542 3580 6576 3614
rect 6611 3580 6645 3614
rect 6680 3580 6714 3614
rect 6749 3580 6783 3614
rect 6818 3580 6852 3614
rect 6887 3580 6921 3614
rect 6956 3580 6990 3614
rect 7025 3580 7059 3614
rect 7094 3580 7128 3614
rect 7163 3580 7197 3614
rect 7232 3580 7266 3614
rect 7301 3580 7335 3614
rect 7370 3580 7404 3614
rect 7439 3580 7473 3614
rect 7508 3580 7542 3614
rect 7577 3580 7611 3614
rect 7646 3580 7680 3614
rect 7715 3580 7749 3614
rect 7784 3580 7818 3614
rect 7853 3580 7887 3614
rect 7922 3580 7956 3614
rect 7991 3580 8025 3614
rect 8060 3580 8094 3614
rect 8129 3580 8163 3614
rect 8198 3580 8232 3614
rect 8267 3580 8301 3614
rect 8336 3580 8370 3614
rect 8405 3580 8439 3614
rect 8474 3580 8508 3614
rect 8543 3580 8577 3614
rect 8612 3580 8646 3614
rect 8681 3580 8715 3614
rect 8750 3580 8784 3614
rect 8819 3580 8853 3614
rect 8888 3580 8922 3614
rect 8957 3580 8991 3614
rect 9026 3580 9060 3614
rect 9095 3580 9129 3614
rect 9164 3580 9198 3614
rect 9233 3580 9267 3614
rect 9302 3580 9336 3614
rect 9371 3580 9405 3614
rect 9440 3580 9474 3614
rect 9509 3580 9543 3614
rect 9578 3580 9612 3614
rect 9647 3580 9681 3614
rect 9716 3580 9750 3614
rect 9785 3580 9819 3614
rect 9854 3580 9888 3614
rect 9922 3580 9956 3614
rect 9990 3580 10024 3614
rect 10058 3580 10092 3614
rect 10126 3580 10160 3614
rect 10194 3580 10228 3614
rect 10262 3580 10296 3614
rect 10330 3580 10364 3614
rect 10398 3580 10432 3614
rect 10466 3580 10500 3614
rect 10534 3580 10568 3614
rect 10602 3580 10636 3614
rect 10670 3580 10704 3614
rect 10738 3580 10772 3614
rect 10806 3580 10840 3614
rect 10874 3580 10908 3614
rect 10942 3580 10976 3614
rect 11010 3580 11044 3614
rect 11078 3580 11112 3614
rect 11146 3580 11180 3614
rect 11214 3580 11248 3614
rect 11282 3580 11316 3614
rect 11350 3580 11384 3614
rect 11418 3580 11452 3614
rect 11486 3580 11520 3614
rect 11554 3580 11588 3614
rect 11622 3580 11656 3614
rect 11690 3580 11724 3614
rect 11758 3580 11792 3614
rect 11826 3580 11860 3614
rect 11894 3580 11928 3614
rect 11962 3580 11996 3614
rect 12030 3580 12064 3614
rect 12098 3580 12132 3614
rect 12166 3580 12200 3614
rect 12234 3580 12268 3614
rect 12302 3580 12336 3614
rect 12370 3580 12404 3614
rect 12438 3580 12472 3614
rect 12506 3580 12540 3614
rect 12574 3580 12608 3614
rect 12642 3580 12676 3614
rect 12710 3580 12744 3614
rect 12778 3580 12812 3614
rect 12846 3580 12880 3614
rect 12914 3580 12948 3614
rect 12982 3580 13016 3614
rect 13050 3580 13084 3614
rect 13118 3580 13152 3614
rect 13186 3580 13220 3614
rect 13254 3580 13288 3614
rect 13322 3580 13356 3614
rect 13390 3580 13424 3614
rect 13458 3580 13492 3614
rect 13526 3580 13560 3614
rect 13594 3580 13628 3614
rect 13662 3580 13696 3614
rect 13730 3580 13764 3614
rect 13798 3580 13832 3614
rect 13866 3580 13900 3614
rect 13934 3580 13968 3614
rect 14002 3580 14036 3614
rect 14070 3580 14104 3614
rect 14138 3580 14172 3614
rect 14206 3580 14240 3614
rect 14274 3580 14308 3614
rect 14342 3580 14376 3614
rect 14410 3580 14444 3614
rect 14478 3580 14512 3614
rect 14546 3580 14580 3614
rect 14614 3580 14648 3614
rect 14682 3580 14716 3614
rect 14750 3580 14784 3614
rect 14818 3580 14852 3614
rect 14886 3580 14920 3614
rect 14954 3580 14988 3614
rect 15022 3580 15056 3614
rect 15090 3580 15124 3614
rect 15158 3580 15192 3614
rect 15226 3580 15260 3614
rect 15294 3580 15328 3614
rect 15362 3580 15396 3614
rect 15430 3580 15464 3614
rect 15498 3580 15532 3614
rect 15566 3580 15600 3614
rect 15634 3580 15668 3614
rect 15702 3580 15736 3614
rect 15770 3580 15804 3614
rect 15838 3580 15872 3614
rect 15906 3580 15940 3614
rect 15974 3580 16008 3614
rect 16042 3580 16076 3614
rect 16110 3580 16144 3614
rect 16178 3580 16212 3614
rect 16246 3580 16280 3614
rect 16314 3580 16348 3614
rect 16382 3580 16416 3614
rect 16450 3580 16484 3614
rect 16518 3580 16552 3614
rect 16586 3580 16620 3614
rect 16654 3580 16688 3614
rect 16722 3580 16756 3614
rect 16790 3580 16824 3614
rect 16858 3580 16892 3614
rect 16926 3580 16960 3614
rect 16994 3580 17028 3614
rect 17062 3580 17096 3614
rect 17130 3580 17164 3614
rect 17198 3580 17232 3614
rect 17266 3580 17300 3614
rect 17334 3580 17368 3614
rect 17402 3580 17436 3614
rect 17470 3580 17504 3614
rect 17538 3580 17572 3614
rect 17606 3580 17640 3614
rect 17674 3580 17708 3614
rect 17742 3580 17776 3614
rect 17810 3580 17844 3614
rect 17878 3580 17912 3614
rect 17946 3580 17980 3614
rect 18014 3580 18048 3614
rect 18082 3580 18116 3614
rect 18150 3580 18184 3614
rect 18218 3580 18252 3614
rect 18286 3580 18320 3614
rect 18354 3580 18388 3614
rect 18422 3580 18456 3614
rect 18490 3580 18524 3614
rect 18558 3580 18592 3614
rect 18626 3580 18660 3614
rect 18694 3580 18728 3614
rect 18762 3580 18796 3614
rect 18830 3580 18864 3614
rect 18898 3580 18932 3614
rect 18966 3580 19000 3614
rect 19034 3580 19068 3614
rect 19102 3580 19136 3614
rect 19170 3580 19204 3614
rect 19238 3580 19272 3614
rect 19306 3580 19340 3614
rect 19374 3580 19408 3614
rect 19442 3580 19476 3614
rect 19510 3580 19544 3614
rect 19578 3580 19612 3614
rect 19646 3580 19680 3614
rect 19714 3580 19748 3614
rect 19782 3580 19816 3614
rect 19850 3580 19884 3614
rect 19918 3580 19952 3614
rect 19986 3580 20020 3614
rect 20054 3580 20088 3614
rect 20122 3580 20156 3614
rect 20190 3580 20224 3614
rect 20258 3580 20292 3614
rect 20326 3580 20360 3614
rect 20394 3580 20428 3614
rect 20462 3580 20496 3614
rect 20530 3580 20564 3614
rect 20598 3580 20632 3614
rect 20666 3580 20700 3614
rect 20734 3580 20768 3614
rect 20802 3580 20836 3614
rect 20870 3580 20904 3614
rect 20938 3580 20972 3614
rect 21006 3580 21040 3614
rect 21074 3580 21108 3614
rect 21142 3580 21176 3614
rect 21210 3580 21244 3614
rect 21278 3580 21312 3614
rect 21346 3580 21380 3614
rect 21414 3580 21448 3614
rect 21482 3580 21516 3614
rect 21550 3580 21584 3614
rect 21618 3580 21652 3614
rect 21686 3580 21720 3614
rect 21754 3580 21788 3614
rect 21822 3580 21856 3614
rect 21890 3580 21924 3614
rect 21958 3580 21992 3614
rect 22026 3580 22060 3614
rect 22094 3580 22128 3614
rect 22162 3580 22196 3614
rect 22230 3580 22264 3614
rect 22298 3580 22332 3614
rect 22366 3580 22400 3614
rect 22434 3580 22468 3614
rect 22502 3580 22536 3614
rect 22570 3580 22604 3614
rect 22638 3580 22672 3614
rect 22706 3580 22740 3614
rect 22774 3580 22808 3614
rect 22842 3580 22876 3614
rect 22910 3580 22944 3614
rect 22978 3580 23012 3614
rect 23046 3580 23080 3614
rect 23114 3580 23148 3614
rect 23182 3580 23216 3614
rect 23250 3580 23284 3614
rect 23318 3580 23352 3614
rect 23386 3580 23420 3614
rect 23454 3580 23488 3614
rect 23522 3580 23556 3614
rect 23590 3580 23624 3614
rect 23658 3580 23692 3614
rect 23726 3580 23760 3614
rect 23794 3580 23828 3614
rect 23862 3580 23896 3614
rect 23930 3580 23964 3614
rect 23998 3580 24032 3614
rect 24066 3580 24100 3614
rect 24134 3580 24168 3614
rect 24202 3580 24236 3614
rect 24270 3580 24304 3614
rect 24338 3580 24372 3614
rect 24406 3580 24440 3614
rect 24474 3580 24508 3614
rect 24542 3580 24576 3614
rect 24610 3580 24644 3614
rect 24678 3580 24712 3614
rect 24746 3580 24780 3614
rect 24814 3580 24848 3614
rect 24882 3580 24916 3614
rect 24950 3580 24984 3614
rect 25018 3580 25052 3614
rect 25086 3580 25120 3614
rect 25154 3580 25188 3614
rect 25222 3580 25256 3614
rect 25290 3580 25324 3614
rect 25358 3580 25392 3614
rect 25426 3580 25460 3614
rect 25494 3580 25528 3614
rect 25562 3580 25596 3614
rect 25630 3580 25664 3614
rect 25698 3580 25732 3614
rect 25766 3580 25800 3614
rect 25834 3580 25868 3614
rect 25902 3580 25936 3614
rect 25970 3580 26004 3614
rect 26038 3580 26072 3614
rect 26106 3580 26140 3614
rect 26174 3580 26208 3614
rect 26242 3580 26276 3614
rect 26310 3580 26344 3614
rect 26378 3580 26412 3614
rect 26446 3580 26480 3614
rect 26514 3580 26548 3614
rect 26582 3580 26616 3614
rect 26650 3580 26684 3614
rect 26718 3580 26752 3614
rect 26786 3580 26820 3614
rect 26854 3580 26888 3614
rect 26922 3580 26956 3614
rect 26990 3580 27024 3614
rect 27058 3580 27092 3614
rect 27126 3580 27160 3614
rect 27194 3580 27228 3614
rect 27262 3580 27296 3614
rect 27330 3580 27364 3614
rect 27398 3580 27432 3614
rect 27466 3580 27500 3614
rect 27534 3580 27568 3614
rect 27602 3580 27636 3614
rect 27670 3580 27704 3614
rect 27738 3580 27772 3614
rect 27806 3580 27840 3614
rect 27874 3580 27908 3614
rect 27942 3580 27976 3614
rect 6473 3506 6507 3540
rect 6542 3506 6576 3540
rect 6611 3506 6645 3540
rect 6680 3506 6714 3540
rect 6749 3506 6783 3540
rect 6818 3506 6852 3540
rect 6887 3506 6921 3540
rect 6956 3506 6990 3540
rect 7025 3506 7059 3540
rect 7094 3506 7128 3540
rect 7163 3506 7197 3540
rect 7232 3506 7266 3540
rect 7301 3506 7335 3540
rect 7370 3506 7404 3540
rect 7439 3506 7473 3540
rect 7508 3506 7542 3540
rect 7577 3506 7611 3540
rect 7646 3506 7680 3540
rect 7715 3506 7749 3540
rect 7784 3506 7818 3540
rect 7853 3506 7887 3540
rect 7922 3506 7956 3540
rect 7991 3506 8025 3540
rect 8060 3506 8094 3540
rect 8129 3506 8163 3540
rect 8198 3506 8232 3540
rect 8267 3506 8301 3540
rect 8336 3506 8370 3540
rect 8405 3506 8439 3540
rect 8474 3506 8508 3540
rect 8543 3506 8577 3540
rect 8612 3506 8646 3540
rect 8681 3506 8715 3540
rect 8750 3506 8784 3540
rect 8819 3506 8853 3540
rect 8888 3506 8922 3540
rect 8957 3506 8991 3540
rect 9026 3506 9060 3540
rect 9095 3506 9129 3540
rect 9164 3506 9198 3540
rect 9233 3506 9267 3540
rect 9302 3506 9336 3540
rect 9371 3506 9405 3540
rect 9440 3506 9474 3540
rect 9509 3506 9543 3540
rect 9578 3506 9612 3540
rect 9647 3506 9681 3540
rect 9716 3506 9750 3540
rect 9785 3506 9819 3540
rect 9854 3506 9888 3540
rect 9922 3506 9956 3540
rect 9990 3506 10024 3540
rect 10058 3506 10092 3540
rect 10126 3506 10160 3540
rect 10194 3506 10228 3540
rect 10262 3506 10296 3540
rect 10330 3506 10364 3540
rect 10398 3506 10432 3540
rect 10466 3506 10500 3540
rect 10534 3506 10568 3540
rect 10602 3506 10636 3540
rect 10670 3506 10704 3540
rect 10738 3506 10772 3540
rect 10806 3506 10840 3540
rect 10874 3506 10908 3540
rect 10942 3506 10976 3540
rect 11010 3506 11044 3540
rect 11078 3506 11112 3540
rect 11146 3506 11180 3540
rect 11214 3506 11248 3540
rect 11282 3506 11316 3540
rect 11350 3506 11384 3540
rect 11418 3506 11452 3540
rect 11486 3506 11520 3540
rect 11554 3506 11588 3540
rect 11622 3506 11656 3540
rect 11690 3506 11724 3540
rect 11758 3506 11792 3540
rect 11826 3506 11860 3540
rect 11894 3506 11928 3540
rect 11962 3506 11996 3540
rect 12030 3506 12064 3540
rect 12098 3506 12132 3540
rect 12166 3506 12200 3540
rect 12234 3506 12268 3540
rect 12302 3506 12336 3540
rect 12370 3506 12404 3540
rect 12438 3506 12472 3540
rect 12506 3506 12540 3540
rect 12574 3506 12608 3540
rect 12642 3506 12676 3540
rect 12710 3506 12744 3540
rect 12778 3506 12812 3540
rect 12846 3506 12880 3540
rect 12914 3506 12948 3540
rect 12982 3506 13016 3540
rect 13050 3506 13084 3540
rect 13118 3506 13152 3540
rect 13186 3506 13220 3540
rect 13254 3506 13288 3540
rect 13322 3506 13356 3540
rect 13390 3506 13424 3540
rect 13458 3506 13492 3540
rect 13526 3506 13560 3540
rect 13594 3506 13628 3540
rect 13662 3506 13696 3540
rect 13730 3506 13764 3540
rect 13798 3506 13832 3540
rect 13866 3506 13900 3540
rect 13934 3506 13968 3540
rect 14002 3506 14036 3540
rect 14070 3506 14104 3540
rect 14138 3506 14172 3540
rect 14206 3506 14240 3540
rect 14274 3506 14308 3540
rect 14342 3506 14376 3540
rect 14410 3506 14444 3540
rect 14478 3506 14512 3540
rect 14546 3506 14580 3540
rect 14614 3506 14648 3540
rect 14682 3506 14716 3540
rect 14750 3506 14784 3540
rect 14818 3506 14852 3540
rect 14886 3506 14920 3540
rect 14954 3506 14988 3540
rect 15022 3506 15056 3540
rect 15090 3506 15124 3540
rect 15158 3506 15192 3540
rect 15226 3506 15260 3540
rect 15294 3506 15328 3540
rect 15362 3506 15396 3540
rect 15430 3506 15464 3540
rect 15498 3506 15532 3540
rect 15566 3506 15600 3540
rect 15634 3506 15668 3540
rect 15702 3506 15736 3540
rect 15770 3506 15804 3540
rect 15838 3506 15872 3540
rect 15906 3506 15940 3540
rect 15974 3506 16008 3540
rect 16042 3506 16076 3540
rect 16110 3506 16144 3540
rect 16178 3506 16212 3540
rect 16246 3506 16280 3540
rect 16314 3506 16348 3540
rect 16382 3506 16416 3540
rect 16450 3506 16484 3540
rect 16518 3506 16552 3540
rect 16586 3506 16620 3540
rect 16654 3506 16688 3540
rect 16722 3506 16756 3540
rect 16790 3506 16824 3540
rect 16858 3506 16892 3540
rect 16926 3506 16960 3540
rect 16994 3506 17028 3540
rect 17062 3506 17096 3540
rect 17130 3506 17164 3540
rect 17198 3506 17232 3540
rect 17266 3506 17300 3540
rect 17334 3506 17368 3540
rect 17402 3506 17436 3540
rect 17470 3506 17504 3540
rect 17538 3506 17572 3540
rect 17606 3506 17640 3540
rect 17674 3506 17708 3540
rect 17742 3506 17776 3540
rect 17810 3506 17844 3540
rect 17878 3506 17912 3540
rect 17946 3506 17980 3540
rect 18014 3506 18048 3540
rect 18082 3506 18116 3540
rect 18150 3506 18184 3540
rect 18218 3506 18252 3540
rect 18286 3506 18320 3540
rect 18354 3506 18388 3540
rect 18422 3506 18456 3540
rect 18490 3506 18524 3540
rect 18558 3506 18592 3540
rect 18626 3506 18660 3540
rect 18694 3506 18728 3540
rect 18762 3506 18796 3540
rect 18830 3506 18864 3540
rect 18898 3506 18932 3540
rect 18966 3506 19000 3540
rect 19034 3506 19068 3540
rect 19102 3506 19136 3540
rect 19170 3506 19204 3540
rect 19238 3506 19272 3540
rect 19306 3506 19340 3540
rect 19374 3506 19408 3540
rect 19442 3506 19476 3540
rect 19510 3506 19544 3540
rect 19578 3506 19612 3540
rect 19646 3506 19680 3540
rect 19714 3506 19748 3540
rect 19782 3506 19816 3540
rect 19850 3506 19884 3540
rect 19918 3506 19952 3540
rect 19986 3506 20020 3540
rect 20054 3506 20088 3540
rect 20122 3506 20156 3540
rect 20190 3506 20224 3540
rect 20258 3506 20292 3540
rect 20326 3506 20360 3540
rect 20394 3506 20428 3540
rect 20462 3506 20496 3540
rect 20530 3506 20564 3540
rect 20598 3506 20632 3540
rect 20666 3506 20700 3540
rect 20734 3506 20768 3540
rect 20802 3506 20836 3540
rect 20870 3506 20904 3540
rect 20938 3506 20972 3540
rect 21006 3506 21040 3540
rect 21074 3506 21108 3540
rect 21142 3506 21176 3540
rect 21210 3506 21244 3540
rect 21278 3506 21312 3540
rect 21346 3506 21380 3540
rect 21414 3506 21448 3540
rect 21482 3506 21516 3540
rect 21550 3506 21584 3540
rect 21618 3506 21652 3540
rect 21686 3506 21720 3540
rect 21754 3506 21788 3540
rect 21822 3506 21856 3540
rect 21890 3506 21924 3540
rect 21958 3506 21992 3540
rect 22026 3506 22060 3540
rect 22094 3506 22128 3540
rect 22162 3506 22196 3540
rect 22230 3506 22264 3540
rect 22298 3506 22332 3540
rect 22366 3506 22400 3540
rect 22434 3506 22468 3540
rect 22502 3506 22536 3540
rect 22570 3506 22604 3540
rect 22638 3506 22672 3540
rect 22706 3506 22740 3540
rect 22774 3506 22808 3540
rect 22842 3506 22876 3540
rect 22910 3506 22944 3540
rect 22978 3506 23012 3540
rect 23046 3506 23080 3540
rect 23114 3506 23148 3540
rect 23182 3506 23216 3540
rect 23250 3506 23284 3540
rect 23318 3506 23352 3540
rect 23386 3506 23420 3540
rect 23454 3506 23488 3540
rect 23522 3506 23556 3540
rect 23590 3506 23624 3540
rect 23658 3506 23692 3540
rect 23726 3506 23760 3540
rect 23794 3506 23828 3540
rect 23862 3506 23896 3540
rect 23930 3506 23964 3540
rect 23998 3506 24032 3540
rect 24066 3506 24100 3540
rect 24134 3506 24168 3540
rect 24202 3506 24236 3540
rect 24270 3506 24304 3540
rect 24338 3506 24372 3540
rect 24406 3506 24440 3540
rect 24474 3506 24508 3540
rect 24542 3506 24576 3540
rect 24610 3506 24644 3540
rect 24678 3506 24712 3540
rect 24746 3506 24780 3540
rect 24814 3506 24848 3540
rect 24882 3506 24916 3540
rect 24950 3506 24984 3540
rect 25018 3506 25052 3540
rect 25086 3506 25120 3540
rect 25154 3506 25188 3540
rect 25222 3506 25256 3540
rect 25290 3506 25324 3540
rect 25358 3506 25392 3540
rect 25426 3506 25460 3540
rect 25494 3506 25528 3540
rect 25562 3506 25596 3540
rect 25630 3506 25664 3540
rect 25698 3506 25732 3540
rect 25766 3506 25800 3540
rect 25834 3506 25868 3540
rect 25902 3506 25936 3540
rect 25970 3506 26004 3540
rect 26038 3506 26072 3540
rect 26106 3506 26140 3540
rect 26174 3506 26208 3540
rect 26242 3506 26276 3540
rect 26310 3506 26344 3540
rect 26378 3506 26412 3540
rect 26446 3506 26480 3540
rect 26514 3506 26548 3540
rect 26582 3506 26616 3540
rect 26650 3506 26684 3540
rect 26718 3506 26752 3540
rect 26786 3506 26820 3540
rect 26854 3506 26888 3540
rect 26922 3506 26956 3540
rect 26990 3506 27024 3540
rect 27058 3506 27092 3540
rect 27126 3506 27160 3540
rect 27194 3506 27228 3540
rect 27262 3506 27296 3540
rect 27330 3506 27364 3540
rect 27398 3506 27432 3540
rect 27466 3506 27500 3540
rect 27534 3506 27568 3540
rect 27602 3506 27636 3540
rect 27670 3506 27704 3540
rect 27738 3506 27772 3540
rect 27806 3506 27840 3540
rect 27874 3506 27908 3540
rect 27942 3506 27976 3540
rect 6473 3432 6507 3466
rect 6542 3432 6576 3466
rect 6611 3432 6645 3466
rect 6680 3432 6714 3466
rect 6749 3432 6783 3466
rect 6818 3432 6852 3466
rect 6887 3432 6921 3466
rect 6956 3432 6990 3466
rect 7025 3432 7059 3466
rect 7094 3432 7128 3466
rect 7163 3432 7197 3466
rect 7232 3432 7266 3466
rect 7301 3432 7335 3466
rect 7370 3432 7404 3466
rect 7439 3432 7473 3466
rect 7508 3432 7542 3466
rect 7577 3432 7611 3466
rect 7646 3432 7680 3466
rect 7715 3432 7749 3466
rect 7784 3432 7818 3466
rect 7853 3432 7887 3466
rect 7922 3432 7956 3466
rect 7991 3432 8025 3466
rect 8060 3432 8094 3466
rect 8129 3432 8163 3466
rect 8198 3432 8232 3466
rect 8267 3432 8301 3466
rect 8336 3432 8370 3466
rect 8405 3432 8439 3466
rect 8474 3432 8508 3466
rect 8543 3432 8577 3466
rect 8612 3432 8646 3466
rect 8681 3432 8715 3466
rect 8750 3432 8784 3466
rect 8819 3432 8853 3466
rect 8888 3432 8922 3466
rect 8957 3432 8991 3466
rect 9026 3432 9060 3466
rect 9095 3432 9129 3466
rect 9164 3432 9198 3466
rect 9233 3432 9267 3466
rect 9302 3432 9336 3466
rect 9371 3432 9405 3466
rect 9440 3432 9474 3466
rect 9509 3432 9543 3466
rect 9578 3432 9612 3466
rect 9647 3432 9681 3466
rect 9716 3432 9750 3466
rect 9785 3432 9819 3466
rect 9854 3432 9888 3466
rect 9922 3432 9956 3466
rect 9990 3432 10024 3466
rect 10058 3432 10092 3466
rect 10126 3432 10160 3466
rect 10194 3432 10228 3466
rect 10262 3432 10296 3466
rect 10330 3432 10364 3466
rect 10398 3432 10432 3466
rect 10466 3432 10500 3466
rect 10534 3432 10568 3466
rect 10602 3432 10636 3466
rect 10670 3432 10704 3466
rect 10738 3432 10772 3466
rect 10806 3432 10840 3466
rect 10874 3432 10908 3466
rect 10942 3432 10976 3466
rect 11010 3432 11044 3466
rect 11078 3432 11112 3466
rect 11146 3432 11180 3466
rect 11214 3432 11248 3466
rect 11282 3432 11316 3466
rect 11350 3432 11384 3466
rect 11418 3432 11452 3466
rect 11486 3432 11520 3466
rect 11554 3432 11588 3466
rect 11622 3432 11656 3466
rect 11690 3432 11724 3466
rect 11758 3432 11792 3466
rect 11826 3432 11860 3466
rect 11894 3432 11928 3466
rect 11962 3432 11996 3466
rect 12030 3432 12064 3466
rect 12098 3432 12132 3466
rect 12166 3432 12200 3466
rect 12234 3432 12268 3466
rect 12302 3432 12336 3466
rect 12370 3432 12404 3466
rect 12438 3432 12472 3466
rect 12506 3432 12540 3466
rect 12574 3432 12608 3466
rect 12642 3432 12676 3466
rect 12710 3432 12744 3466
rect 12778 3432 12812 3466
rect 12846 3432 12880 3466
rect 12914 3432 12948 3466
rect 12982 3432 13016 3466
rect 13050 3432 13084 3466
rect 13118 3432 13152 3466
rect 13186 3432 13220 3466
rect 13254 3432 13288 3466
rect 13322 3432 13356 3466
rect 13390 3432 13424 3466
rect 13458 3432 13492 3466
rect 13526 3432 13560 3466
rect 13594 3432 13628 3466
rect 13662 3432 13696 3466
rect 13730 3432 13764 3466
rect 13798 3432 13832 3466
rect 13866 3432 13900 3466
rect 13934 3432 13968 3466
rect 14002 3432 14036 3466
rect 14070 3432 14104 3466
rect 14138 3432 14172 3466
rect 14206 3432 14240 3466
rect 14274 3432 14308 3466
rect 14342 3432 14376 3466
rect 14410 3432 14444 3466
rect 14478 3432 14512 3466
rect 14546 3432 14580 3466
rect 14614 3432 14648 3466
rect 14682 3432 14716 3466
rect 14750 3432 14784 3466
rect 14818 3432 14852 3466
rect 14886 3432 14920 3466
rect 14954 3432 14988 3466
rect 15022 3432 15056 3466
rect 15090 3432 15124 3466
rect 15158 3432 15192 3466
rect 15226 3432 15260 3466
rect 15294 3432 15328 3466
rect 15362 3432 15396 3466
rect 15430 3432 15464 3466
rect 15498 3432 15532 3466
rect 15566 3432 15600 3466
rect 15634 3432 15668 3466
rect 15702 3432 15736 3466
rect 15770 3432 15804 3466
rect 15838 3432 15872 3466
rect 15906 3432 15940 3466
rect 15974 3432 16008 3466
rect 16042 3432 16076 3466
rect 16110 3432 16144 3466
rect 16178 3432 16212 3466
rect 16246 3432 16280 3466
rect 16314 3432 16348 3466
rect 16382 3432 16416 3466
rect 16450 3432 16484 3466
rect 16518 3432 16552 3466
rect 16586 3432 16620 3466
rect 16654 3432 16688 3466
rect 16722 3432 16756 3466
rect 16790 3432 16824 3466
rect 16858 3432 16892 3466
rect 16926 3432 16960 3466
rect 16994 3432 17028 3466
rect 17062 3432 17096 3466
rect 17130 3432 17164 3466
rect 17198 3432 17232 3466
rect 17266 3432 17300 3466
rect 17334 3432 17368 3466
rect 17402 3432 17436 3466
rect 17470 3432 17504 3466
rect 17538 3432 17572 3466
rect 17606 3432 17640 3466
rect 17674 3432 17708 3466
rect 17742 3432 17776 3466
rect 17810 3432 17844 3466
rect 17878 3432 17912 3466
rect 17946 3432 17980 3466
rect 18014 3432 18048 3466
rect 18082 3432 18116 3466
rect 18150 3432 18184 3466
rect 18218 3432 18252 3466
rect 18286 3432 18320 3466
rect 18354 3432 18388 3466
rect 18422 3432 18456 3466
rect 18490 3432 18524 3466
rect 18558 3432 18592 3466
rect 18626 3432 18660 3466
rect 18694 3432 18728 3466
rect 18762 3432 18796 3466
rect 18830 3432 18864 3466
rect 18898 3432 18932 3466
rect 18966 3432 19000 3466
rect 19034 3432 19068 3466
rect 19102 3432 19136 3466
rect 19170 3432 19204 3466
rect 19238 3432 19272 3466
rect 19306 3432 19340 3466
rect 19374 3432 19408 3466
rect 19442 3432 19476 3466
rect 19510 3432 19544 3466
rect 19578 3432 19612 3466
rect 19646 3432 19680 3466
rect 19714 3432 19748 3466
rect 19782 3432 19816 3466
rect 19850 3432 19884 3466
rect 19918 3432 19952 3466
rect 19986 3432 20020 3466
rect 20054 3432 20088 3466
rect 20122 3432 20156 3466
rect 20190 3432 20224 3466
rect 20258 3432 20292 3466
rect 20326 3432 20360 3466
rect 20394 3432 20428 3466
rect 20462 3432 20496 3466
rect 20530 3432 20564 3466
rect 20598 3432 20632 3466
rect 20666 3432 20700 3466
rect 20734 3432 20768 3466
rect 20802 3432 20836 3466
rect 20870 3432 20904 3466
rect 20938 3432 20972 3466
rect 21006 3432 21040 3466
rect 21074 3432 21108 3466
rect 21142 3432 21176 3466
rect 21210 3432 21244 3466
rect 21278 3432 21312 3466
rect 21346 3432 21380 3466
rect 21414 3432 21448 3466
rect 21482 3432 21516 3466
rect 21550 3432 21584 3466
rect 21618 3432 21652 3466
rect 21686 3432 21720 3466
rect 21754 3432 21788 3466
rect 21822 3432 21856 3466
rect 21890 3432 21924 3466
rect 21958 3432 21992 3466
rect 22026 3432 22060 3466
rect 22094 3432 22128 3466
rect 22162 3432 22196 3466
rect 22230 3432 22264 3466
rect 22298 3432 22332 3466
rect 22366 3432 22400 3466
rect 22434 3432 22468 3466
rect 22502 3432 22536 3466
rect 22570 3432 22604 3466
rect 22638 3432 22672 3466
rect 22706 3432 22740 3466
rect 22774 3432 22808 3466
rect 22842 3432 22876 3466
rect 22910 3432 22944 3466
rect 22978 3432 23012 3466
rect 23046 3432 23080 3466
rect 23114 3432 23148 3466
rect 23182 3432 23216 3466
rect 23250 3432 23284 3466
rect 23318 3432 23352 3466
rect 23386 3432 23420 3466
rect 23454 3432 23488 3466
rect 23522 3432 23556 3466
rect 23590 3432 23624 3466
rect 23658 3432 23692 3466
rect 23726 3432 23760 3466
rect 23794 3432 23828 3466
rect 23862 3432 23896 3466
rect 23930 3432 23964 3466
rect 23998 3432 24032 3466
rect 24066 3432 24100 3466
rect 24134 3432 24168 3466
rect 24202 3432 24236 3466
rect 24270 3432 24304 3466
rect 24338 3432 24372 3466
rect 24406 3432 24440 3466
rect 24474 3432 24508 3466
rect 24542 3432 24576 3466
rect 24610 3432 24644 3466
rect 24678 3432 24712 3466
rect 24746 3432 24780 3466
rect 24814 3432 24848 3466
rect 24882 3432 24916 3466
rect 24950 3432 24984 3466
rect 25018 3432 25052 3466
rect 25086 3432 25120 3466
rect 25154 3432 25188 3466
rect 25222 3432 25256 3466
rect 25290 3432 25324 3466
rect 25358 3432 25392 3466
rect 25426 3432 25460 3466
rect 25494 3432 25528 3466
rect 25562 3432 25596 3466
rect 25630 3432 25664 3466
rect 25698 3432 25732 3466
rect 25766 3432 25800 3466
rect 25834 3432 25868 3466
rect 25902 3432 25936 3466
rect 25970 3432 26004 3466
rect 26038 3432 26072 3466
rect 26106 3432 26140 3466
rect 26174 3432 26208 3466
rect 26242 3432 26276 3466
rect 26310 3432 26344 3466
rect 26378 3432 26412 3466
rect 26446 3432 26480 3466
rect 26514 3432 26548 3466
rect 26582 3432 26616 3466
rect 26650 3432 26684 3466
rect 26718 3432 26752 3466
rect 26786 3432 26820 3466
rect 26854 3432 26888 3466
rect 26922 3432 26956 3466
rect 26990 3432 27024 3466
rect 27058 3432 27092 3466
rect 27126 3432 27160 3466
rect 27194 3432 27228 3466
rect 27262 3432 27296 3466
rect 27330 3432 27364 3466
rect 27398 3432 27432 3466
rect 27466 3432 27500 3466
rect 27534 3432 27568 3466
rect 27602 3432 27636 3466
rect 27670 3432 27704 3466
rect 27738 3432 27772 3466
rect 27806 3432 27840 3466
rect 27874 3432 27908 3466
rect 27942 3432 27976 3466
<< mvpsubdiffcont >>
rect 23747 23319 23781 23353
rect 23816 23319 23850 23353
rect 23885 23319 23919 23353
rect 23954 23319 23988 23353
rect 24023 23319 24057 23353
rect 24092 23319 24126 23353
rect 24161 23319 24195 23353
rect 24230 23319 24264 23353
rect 24299 23319 24333 23353
rect 24368 23319 24402 23353
rect 24437 23319 24471 23353
rect 24506 23319 24540 23353
rect 24575 23319 24609 23353
rect 24644 23319 24678 23353
rect 24713 23319 24747 23353
rect 24782 23319 24816 23353
rect 24851 23319 24885 23353
rect 24920 23319 24954 23353
rect 24989 23319 25023 23353
rect 25058 23319 25092 23353
rect 25127 23319 25161 23353
rect 25196 23319 25230 23353
rect 25265 23319 25299 23353
rect 25334 23319 25368 23353
rect 25403 23319 25437 23353
rect 25472 23319 25506 23353
rect 25541 23319 25575 23353
rect 25610 23319 25644 23353
rect 25679 23319 25713 23353
rect 25748 23319 25782 23353
rect 25817 23319 25851 23353
rect 25886 23319 25920 23353
rect 25955 23319 25989 23353
rect 26024 23319 26058 23353
rect 26093 23319 26127 23353
rect 26162 23319 26196 23353
rect 26231 23319 26265 23353
rect 26300 23319 26334 23353
rect 26368 23319 26402 23353
rect 26436 23319 26470 23353
rect 26504 23319 26538 23353
rect 26572 23319 26606 23353
rect 26640 23319 26674 23353
rect 26708 23319 26742 23353
rect 26776 23319 26810 23353
rect 26844 23319 26878 23353
rect 26912 23319 26946 23353
rect 26980 23319 27014 23353
rect 27048 23319 27082 23353
rect 27116 23319 27150 23353
rect 27184 23319 27218 23353
rect 27252 23319 27286 23353
rect 27320 23319 27354 23353
rect 27388 23319 27422 23353
rect 27456 23319 27490 23353
rect 27524 23319 27558 23353
rect 27592 23319 27626 23353
rect 27660 23319 27694 23353
rect 27728 23319 27762 23353
rect 27796 23319 27830 23353
rect 27864 23319 27898 23353
rect 27932 23319 27966 23353
rect 23747 23249 23781 23283
rect 23816 23249 23850 23283
rect 23885 23249 23919 23283
rect 23954 23249 23988 23283
rect 24023 23249 24057 23283
rect 24092 23249 24126 23283
rect 24161 23249 24195 23283
rect 24230 23249 24264 23283
rect 24299 23249 24333 23283
rect 24368 23249 24402 23283
rect 24437 23249 24471 23283
rect 24506 23249 24540 23283
rect 24575 23249 24609 23283
rect 24644 23249 24678 23283
rect 24713 23249 24747 23283
rect 24782 23249 24816 23283
rect 24851 23249 24885 23283
rect 24920 23249 24954 23283
rect 24989 23249 25023 23283
rect 25058 23249 25092 23283
rect 25127 23249 25161 23283
rect 25196 23249 25230 23283
rect 25265 23249 25299 23283
rect 25334 23249 25368 23283
rect 25403 23249 25437 23283
rect 25472 23249 25506 23283
rect 25541 23249 25575 23283
rect 25610 23249 25644 23283
rect 25679 23249 25713 23283
rect 25748 23249 25782 23283
rect 25817 23249 25851 23283
rect 25886 23249 25920 23283
rect 25955 23249 25989 23283
rect 26024 23249 26058 23283
rect 26093 23249 26127 23283
rect 26162 23249 26196 23283
rect 26231 23249 26265 23283
rect 26300 23249 26334 23283
rect 26368 23249 26402 23283
rect 26436 23249 26470 23283
rect 26504 23249 26538 23283
rect 26572 23249 26606 23283
rect 26640 23249 26674 23283
rect 26708 23249 26742 23283
rect 26776 23249 26810 23283
rect 26844 23249 26878 23283
rect 26912 23249 26946 23283
rect 26980 23249 27014 23283
rect 27048 23249 27082 23283
rect 27116 23249 27150 23283
rect 27184 23249 27218 23283
rect 27252 23249 27286 23283
rect 27320 23249 27354 23283
rect 27388 23249 27422 23283
rect 27456 23249 27490 23283
rect 27524 23249 27558 23283
rect 27592 23249 27626 23283
rect 27660 23249 27694 23283
rect 27728 23249 27762 23283
rect 27796 23249 27830 23283
rect 27864 23249 27898 23283
rect 27932 23249 27966 23283
rect 23747 23179 23781 23213
rect 23816 23179 23850 23213
rect 23885 23179 23919 23213
rect 23954 23179 23988 23213
rect 24023 23179 24057 23213
rect 24092 23179 24126 23213
rect 24161 23179 24195 23213
rect 24230 23179 24264 23213
rect 24299 23179 24333 23213
rect 24368 23179 24402 23213
rect 24437 23179 24471 23213
rect 24506 23179 24540 23213
rect 24575 23179 24609 23213
rect 24644 23179 24678 23213
rect 24713 23179 24747 23213
rect 24782 23179 24816 23213
rect 24851 23179 24885 23213
rect 24920 23179 24954 23213
rect 24989 23179 25023 23213
rect 25058 23179 25092 23213
rect 25127 23179 25161 23213
rect 25196 23179 25230 23213
rect 25265 23179 25299 23213
rect 25334 23179 25368 23213
rect 25403 23179 25437 23213
rect 25472 23179 25506 23213
rect 25541 23179 25575 23213
rect 25610 23179 25644 23213
rect 25679 23179 25713 23213
rect 25748 23179 25782 23213
rect 25817 23179 25851 23213
rect 25886 23179 25920 23213
rect 25955 23179 25989 23213
rect 26024 23179 26058 23213
rect 26093 23179 26127 23213
rect 26162 23179 26196 23213
rect 26231 23179 26265 23213
rect 26300 23179 26334 23213
rect 26368 23179 26402 23213
rect 26436 23179 26470 23213
rect 26504 23179 26538 23213
rect 26572 23179 26606 23213
rect 26640 23179 26674 23213
rect 26708 23179 26742 23213
rect 26776 23179 26810 23213
rect 26844 23179 26878 23213
rect 26912 23179 26946 23213
rect 26980 23179 27014 23213
rect 27048 23179 27082 23213
rect 27116 23179 27150 23213
rect 27184 23179 27218 23213
rect 27252 23179 27286 23213
rect 27320 23179 27354 23213
rect 27388 23179 27422 23213
rect 27456 23179 27490 23213
rect 27524 23179 27558 23213
rect 27592 23179 27626 23213
rect 27660 23179 27694 23213
rect 27728 23179 27762 23213
rect 27796 23179 27830 23213
rect 27864 23179 27898 23213
rect 27932 23179 27966 23213
rect 23747 23109 23781 23143
rect 23816 23109 23850 23143
rect 23885 23109 23919 23143
rect 23954 23109 23988 23143
rect 24023 23109 24057 23143
rect 24092 23109 24126 23143
rect 24161 23109 24195 23143
rect 24230 23109 24264 23143
rect 24299 23109 24333 23143
rect 24368 23109 24402 23143
rect 24437 23109 24471 23143
rect 24506 23109 24540 23143
rect 24575 23109 24609 23143
rect 24644 23109 24678 23143
rect 24713 23109 24747 23143
rect 24782 23109 24816 23143
rect 24851 23109 24885 23143
rect 24920 23109 24954 23143
rect 24989 23109 25023 23143
rect 25058 23109 25092 23143
rect 25127 23109 25161 23143
rect 25196 23109 25230 23143
rect 25265 23109 25299 23143
rect 25334 23109 25368 23143
rect 25403 23109 25437 23143
rect 25472 23109 25506 23143
rect 25541 23109 25575 23143
rect 25610 23109 25644 23143
rect 25679 23109 25713 23143
rect 25748 23109 25782 23143
rect 25817 23109 25851 23143
rect 25886 23109 25920 23143
rect 25955 23109 25989 23143
rect 26024 23109 26058 23143
rect 26093 23109 26127 23143
rect 26162 23109 26196 23143
rect 26231 23109 26265 23143
rect 26300 23109 26334 23143
rect 26368 23109 26402 23143
rect 26436 23109 26470 23143
rect 26504 23109 26538 23143
rect 26572 23109 26606 23143
rect 26640 23109 26674 23143
rect 26708 23109 26742 23143
rect 26776 23109 26810 23143
rect 26844 23109 26878 23143
rect 26912 23109 26946 23143
rect 26980 23109 27014 23143
rect 27048 23109 27082 23143
rect 27116 23109 27150 23143
rect 27184 23109 27218 23143
rect 27252 23109 27286 23143
rect 27320 23109 27354 23143
rect 27388 23109 27422 23143
rect 27456 23109 27490 23143
rect 27524 23109 27558 23143
rect 27592 23109 27626 23143
rect 27660 23109 27694 23143
rect 27728 23109 27762 23143
rect 27796 23109 27830 23143
rect 27864 23109 27898 23143
rect 27932 23109 27966 23143
rect 23747 23039 23781 23073
rect 23816 23039 23850 23073
rect 23885 23039 23919 23073
rect 23954 23039 23988 23073
rect 24023 23039 24057 23073
rect 24092 23039 24126 23073
rect 24161 23039 24195 23073
rect 24230 23039 24264 23073
rect 24299 23039 24333 23073
rect 24368 23039 24402 23073
rect 24437 23039 24471 23073
rect 24506 23039 24540 23073
rect 24575 23039 24609 23073
rect 24644 23039 24678 23073
rect 24713 23039 24747 23073
rect 24782 23039 24816 23073
rect 24851 23039 24885 23073
rect 24920 23039 24954 23073
rect 24989 23039 25023 23073
rect 25058 23039 25092 23073
rect 25127 23039 25161 23073
rect 25196 23039 25230 23073
rect 25265 23039 25299 23073
rect 25334 23039 25368 23073
rect 25403 23039 25437 23073
rect 25472 23039 25506 23073
rect 25541 23039 25575 23073
rect 25610 23039 25644 23073
rect 25679 23039 25713 23073
rect 25748 23039 25782 23073
rect 25817 23039 25851 23073
rect 25886 23039 25920 23073
rect 25955 23039 25989 23073
rect 26024 23039 26058 23073
rect 26093 23039 26127 23073
rect 26162 23039 26196 23073
rect 26231 23039 26265 23073
rect 26300 23039 26334 23073
rect 26368 23039 26402 23073
rect 26436 23039 26470 23073
rect 26504 23039 26538 23073
rect 26572 23039 26606 23073
rect 26640 23039 26674 23073
rect 26708 23039 26742 23073
rect 26776 23039 26810 23073
rect 26844 23039 26878 23073
rect 26912 23039 26946 23073
rect 26980 23039 27014 23073
rect 27048 23039 27082 23073
rect 27116 23039 27150 23073
rect 27184 23039 27218 23073
rect 27252 23039 27286 23073
rect 27320 23039 27354 23073
rect 27388 23039 27422 23073
rect 27456 23039 27490 23073
rect 27524 23039 27558 23073
rect 27592 23039 27626 23073
rect 27660 23039 27694 23073
rect 27728 23039 27762 23073
rect 27796 23039 27830 23073
rect 27864 23039 27898 23073
rect 27932 23039 27966 23073
rect 23747 22969 23781 23003
rect 23816 22969 23850 23003
rect 23885 22969 23919 23003
rect 23954 22969 23988 23003
rect 24023 22969 24057 23003
rect 24092 22969 24126 23003
rect 24161 22969 24195 23003
rect 24230 22969 24264 23003
rect 24299 22969 24333 23003
rect 24368 22969 24402 23003
rect 24437 22969 24471 23003
rect 24506 22969 24540 23003
rect 24575 22969 24609 23003
rect 24644 22969 24678 23003
rect 24713 22969 24747 23003
rect 24782 22969 24816 23003
rect 24851 22969 24885 23003
rect 24920 22969 24954 23003
rect 24989 22969 25023 23003
rect 25058 22969 25092 23003
rect 25127 22969 25161 23003
rect 25196 22969 25230 23003
rect 25265 22969 25299 23003
rect 25334 22969 25368 23003
rect 25403 22969 25437 23003
rect 25472 22969 25506 23003
rect 25541 22969 25575 23003
rect 25610 22969 25644 23003
rect 25679 22969 25713 23003
rect 25748 22969 25782 23003
rect 25817 22969 25851 23003
rect 25886 22969 25920 23003
rect 25955 22969 25989 23003
rect 26024 22969 26058 23003
rect 26093 22969 26127 23003
rect 26162 22969 26196 23003
rect 26231 22969 26265 23003
rect 26300 22969 26334 23003
rect 26368 22969 26402 23003
rect 26436 22969 26470 23003
rect 26504 22969 26538 23003
rect 26572 22969 26606 23003
rect 26640 22969 26674 23003
rect 26708 22969 26742 23003
rect 26776 22969 26810 23003
rect 26844 22969 26878 23003
rect 26912 22969 26946 23003
rect 26980 22969 27014 23003
rect 27048 22969 27082 23003
rect 27116 22969 27150 23003
rect 27184 22969 27218 23003
rect 27252 22969 27286 23003
rect 27320 22969 27354 23003
rect 27388 22969 27422 23003
rect 27456 22969 27490 23003
rect 27524 22969 27558 23003
rect 27592 22969 27626 23003
rect 27660 22969 27694 23003
rect 27728 22969 27762 23003
rect 27796 22969 27830 23003
rect 27864 22969 27898 23003
rect 27932 22969 27966 23003
rect 23747 22899 23781 22933
rect 23816 22899 23850 22933
rect 23885 22899 23919 22933
rect 23954 22899 23988 22933
rect 24023 22899 24057 22933
rect 24092 22899 24126 22933
rect 24161 22899 24195 22933
rect 24230 22899 24264 22933
rect 24299 22899 24333 22933
rect 24368 22899 24402 22933
rect 24437 22899 24471 22933
rect 24506 22899 24540 22933
rect 24575 22899 24609 22933
rect 24644 22899 24678 22933
rect 24713 22899 24747 22933
rect 24782 22899 24816 22933
rect 24851 22899 24885 22933
rect 24920 22899 24954 22933
rect 24989 22899 25023 22933
rect 25058 22899 25092 22933
rect 25127 22899 25161 22933
rect 25196 22899 25230 22933
rect 25265 22899 25299 22933
rect 25334 22899 25368 22933
rect 25403 22899 25437 22933
rect 25472 22899 25506 22933
rect 25541 22899 25575 22933
rect 25610 22899 25644 22933
rect 25679 22899 25713 22933
rect 25748 22899 25782 22933
rect 25817 22899 25851 22933
rect 25886 22899 25920 22933
rect 25955 22899 25989 22933
rect 26024 22899 26058 22933
rect 26093 22899 26127 22933
rect 26162 22899 26196 22933
rect 26231 22899 26265 22933
rect 26300 22899 26334 22933
rect 26368 22899 26402 22933
rect 26436 22899 26470 22933
rect 26504 22899 26538 22933
rect 26572 22899 26606 22933
rect 26640 22899 26674 22933
rect 26708 22899 26742 22933
rect 26776 22899 26810 22933
rect 26844 22899 26878 22933
rect 26912 22899 26946 22933
rect 26980 22899 27014 22933
rect 27048 22899 27082 22933
rect 27116 22899 27150 22933
rect 27184 22899 27218 22933
rect 27252 22899 27286 22933
rect 27320 22899 27354 22933
rect 27388 22899 27422 22933
rect 27456 22899 27490 22933
rect 27524 22899 27558 22933
rect 27592 22899 27626 22933
rect 27660 22899 27694 22933
rect 27728 22899 27762 22933
rect 27796 22899 27830 22933
rect 27864 22899 27898 22933
rect 27932 22899 27966 22933
rect 26309 22822 26343 22856
rect 26380 22822 26414 22856
rect 26451 22822 26485 22856
rect 26522 22822 26556 22856
rect 26593 22822 26627 22856
rect 26664 22822 26698 22856
rect 26735 22822 26769 22856
rect 26806 22822 26840 22856
rect 26877 22822 26911 22856
rect 26948 22822 26982 22856
rect 27019 22822 27053 22856
rect 27090 22822 27124 22856
rect 27161 22822 27195 22856
rect 27232 22822 27266 22856
rect 27302 22822 27336 22856
rect 27372 22822 27406 22856
rect 27442 22822 27476 22856
rect 27512 22822 27546 22856
rect 27582 22822 27616 22856
rect 27652 22822 27686 22856
rect 27722 22822 27756 22856
rect 27792 22822 27826 22856
rect 27862 22822 27896 22856
rect 27932 22822 27966 22856
rect 26309 22748 26343 22782
rect 26380 22748 26414 22782
rect 26451 22748 26485 22782
rect 26522 22748 26556 22782
rect 26593 22748 26627 22782
rect 26664 22748 26698 22782
rect 26735 22748 26769 22782
rect 26806 22748 26840 22782
rect 26877 22748 26911 22782
rect 26948 22748 26982 22782
rect 27019 22748 27053 22782
rect 27090 22748 27124 22782
rect 27161 22748 27195 22782
rect 27232 22748 27266 22782
rect 27302 22748 27336 22782
rect 27372 22748 27406 22782
rect 27442 22748 27476 22782
rect 27512 22748 27546 22782
rect 27582 22748 27616 22782
rect 27652 22748 27686 22782
rect 27722 22748 27756 22782
rect 27792 22748 27826 22782
rect 27862 22748 27896 22782
rect 27932 22748 27966 22782
rect 26309 22674 26343 22708
rect 26380 22674 26414 22708
rect 26451 22674 26485 22708
rect 26522 22674 26556 22708
rect 26593 22674 26627 22708
rect 26664 22674 26698 22708
rect 26735 22674 26769 22708
rect 26806 22674 26840 22708
rect 26877 22674 26911 22708
rect 26948 22674 26982 22708
rect 27019 22674 27053 22708
rect 27090 22674 27124 22708
rect 27161 22674 27195 22708
rect 27232 22674 27266 22708
rect 27302 22674 27336 22708
rect 27372 22674 27406 22708
rect 27442 22674 27476 22708
rect 27512 22674 27546 22708
rect 27582 22674 27616 22708
rect 27652 22674 27686 22708
rect 27722 22674 27756 22708
rect 27792 22674 27826 22708
rect 27862 22674 27896 22708
rect 27932 22674 27966 22708
rect 26309 22600 26343 22634
rect 26380 22600 26414 22634
rect 26451 22600 26485 22634
rect 26522 22600 26556 22634
rect 26593 22600 26627 22634
rect 26664 22600 26698 22634
rect 26735 22600 26769 22634
rect 26806 22600 26840 22634
rect 26877 22600 26911 22634
rect 26948 22600 26982 22634
rect 27019 22600 27053 22634
rect 27090 22600 27124 22634
rect 27161 22600 27195 22634
rect 27232 22600 27266 22634
rect 27302 22600 27336 22634
rect 27372 22600 27406 22634
rect 27442 22600 27476 22634
rect 27512 22600 27546 22634
rect 27582 22600 27616 22634
rect 27652 22600 27686 22634
rect 27722 22600 27756 22634
rect 27792 22600 27826 22634
rect 27862 22600 27896 22634
rect 27932 22600 27966 22634
rect 26309 22526 26343 22560
rect 26380 22526 26414 22560
rect 26451 22526 26485 22560
rect 26522 22526 26556 22560
rect 26593 22526 26627 22560
rect 26664 22526 26698 22560
rect 26735 22526 26769 22560
rect 26806 22526 26840 22560
rect 26877 22526 26911 22560
rect 26948 22526 26982 22560
rect 27019 22526 27053 22560
rect 27090 22526 27124 22560
rect 27161 22526 27195 22560
rect 27232 22526 27266 22560
rect 27302 22526 27336 22560
rect 27372 22526 27406 22560
rect 27442 22526 27476 22560
rect 27512 22526 27546 22560
rect 27582 22526 27616 22560
rect 27652 22526 27686 22560
rect 27722 22526 27756 22560
rect 27792 22526 27826 22560
rect 27862 22526 27896 22560
rect 27932 22526 27966 22560
rect 26309 22452 26343 22486
rect 26380 22452 26414 22486
rect 26451 22452 26485 22486
rect 26522 22452 26556 22486
rect 26593 22452 26627 22486
rect 26664 22452 26698 22486
rect 26735 22452 26769 22486
rect 26806 22452 26840 22486
rect 26877 22452 26911 22486
rect 26948 22452 26982 22486
rect 27019 22452 27053 22486
rect 27090 22452 27124 22486
rect 27161 22452 27195 22486
rect 27232 22452 27266 22486
rect 27302 22452 27336 22486
rect 27372 22452 27406 22486
rect 27442 22452 27476 22486
rect 27512 22452 27546 22486
rect 27582 22452 27616 22486
rect 27652 22452 27686 22486
rect 27722 22452 27756 22486
rect 27792 22452 27826 22486
rect 27862 22452 27896 22486
rect 27932 22452 27966 22486
rect 26309 22378 26343 22412
rect 26380 22378 26414 22412
rect 26451 22378 26485 22412
rect 26522 22378 26556 22412
rect 26593 22378 26627 22412
rect 26664 22378 26698 22412
rect 26735 22378 26769 22412
rect 26806 22378 26840 22412
rect 26877 22378 26911 22412
rect 26948 22378 26982 22412
rect 27019 22378 27053 22412
rect 27090 22378 27124 22412
rect 27161 22378 27195 22412
rect 27232 22378 27266 22412
rect 27302 22378 27336 22412
rect 27372 22378 27406 22412
rect 27442 22378 27476 22412
rect 27512 22378 27546 22412
rect 27582 22378 27616 22412
rect 27652 22378 27686 22412
rect 27722 22378 27756 22412
rect 27792 22378 27826 22412
rect 27862 22378 27896 22412
rect 27932 22378 27966 22412
rect 26309 22304 26343 22338
rect 26380 22304 26414 22338
rect 26451 22304 26485 22338
rect 26522 22304 26556 22338
rect 26593 22304 26627 22338
rect 26664 22304 26698 22338
rect 26735 22304 26769 22338
rect 26806 22304 26840 22338
rect 26877 22304 26911 22338
rect 26948 22304 26982 22338
rect 27019 22304 27053 22338
rect 27090 22304 27124 22338
rect 27161 22304 27195 22338
rect 27232 22304 27266 22338
rect 27302 22304 27336 22338
rect 27372 22304 27406 22338
rect 27442 22304 27476 22338
rect 27512 22304 27546 22338
rect 27582 22304 27616 22338
rect 27652 22304 27686 22338
rect 27722 22304 27756 22338
rect 27792 22304 27826 22338
rect 27862 22304 27896 22338
rect 27932 22304 27966 22338
rect 26309 22230 26343 22264
rect 26380 22230 26414 22264
rect 26451 22230 26485 22264
rect 26522 22230 26556 22264
rect 26593 22230 26627 22264
rect 26664 22230 26698 22264
rect 26735 22230 26769 22264
rect 26806 22230 26840 22264
rect 26877 22230 26911 22264
rect 26948 22230 26982 22264
rect 27019 22230 27053 22264
rect 27090 22230 27124 22264
rect 27161 22230 27195 22264
rect 27232 22230 27266 22264
rect 27302 22230 27336 22264
rect 27372 22230 27406 22264
rect 27442 22230 27476 22264
rect 27512 22230 27546 22264
rect 27582 22230 27616 22264
rect 27652 22230 27686 22264
rect 27722 22230 27756 22264
rect 27792 22230 27826 22264
rect 27862 22230 27896 22264
rect 27932 22230 27966 22264
rect 26309 22156 26343 22190
rect 26380 22156 26414 22190
rect 26451 22156 26485 22190
rect 26522 22156 26556 22190
rect 26593 22156 26627 22190
rect 26664 22156 26698 22190
rect 26735 22156 26769 22190
rect 26806 22156 26840 22190
rect 26877 22156 26911 22190
rect 26948 22156 26982 22190
rect 27019 22156 27053 22190
rect 27090 22156 27124 22190
rect 27161 22156 27195 22190
rect 27232 22156 27266 22190
rect 27302 22156 27336 22190
rect 27372 22156 27406 22190
rect 27442 22156 27476 22190
rect 27512 22156 27546 22190
rect 27582 22156 27616 22190
rect 27652 22156 27686 22190
rect 27722 22156 27756 22190
rect 27792 22156 27826 22190
rect 27862 22156 27896 22190
rect 27932 22156 27966 22190
rect 26309 22082 26343 22116
rect 26380 22082 26414 22116
rect 26451 22082 26485 22116
rect 26522 22082 26556 22116
rect 26593 22082 26627 22116
rect 26664 22082 26698 22116
rect 26735 22082 26769 22116
rect 26806 22082 26840 22116
rect 26877 22082 26911 22116
rect 26948 22082 26982 22116
rect 27019 22082 27053 22116
rect 27090 22082 27124 22116
rect 27161 22082 27195 22116
rect 27232 22082 27266 22116
rect 27302 22082 27336 22116
rect 27372 22082 27406 22116
rect 27442 22082 27476 22116
rect 27512 22082 27546 22116
rect 27582 22082 27616 22116
rect 27652 22082 27686 22116
rect 27722 22082 27756 22116
rect 27792 22082 27826 22116
rect 27862 22082 27896 22116
rect 27932 22082 27966 22116
rect 16903 9560 16937 9594
rect 16976 9560 17010 9594
rect 17049 9560 17083 9594
rect 17122 9560 17156 9594
rect 17195 9560 17229 9594
rect 17267 9560 17301 9594
rect 17339 9560 17373 9594
rect 17411 9560 17445 9594
rect 17483 9560 17517 9594
rect 17555 9560 17589 9594
<< mvnsubdiffcont >>
rect 27012 20762 27046 20796
rect 27012 20694 27046 20728
rect 27012 20626 27046 20660
rect 27012 20558 27046 20592
rect 27012 20490 27046 20524
rect 27012 20422 27046 20456
rect 27012 20354 27046 20388
rect 27012 20286 27046 20320
rect 27012 20218 27046 20252
rect 27012 20150 27046 20184
rect 27012 20082 27046 20116
rect 27012 20014 27046 20048
rect 27012 19946 27046 19980
rect 27012 19878 27046 19912
rect 27012 19810 27046 19844
rect 27012 19742 27046 19776
rect 27012 19674 27046 19708
rect 27012 19606 27046 19640
rect 27012 19538 27046 19572
rect 27012 19470 27046 19504
rect 27012 19402 27046 19436
rect 27012 19334 27046 19368
rect 27012 19266 27046 19300
rect 24129 17739 24639 19201
rect 24129 17670 24163 17704
rect 24197 17670 24231 17704
rect 24265 17670 24299 17704
rect 24333 17670 24367 17704
rect 24401 17670 24435 17704
rect 24469 17670 24503 17704
rect 24537 17670 24571 17704
rect 24605 17670 24639 17704
rect 24129 17601 24163 17635
rect 24197 17601 24231 17635
rect 24265 17601 24299 17635
rect 24333 17601 24367 17635
rect 24401 17601 24435 17635
rect 24469 17601 24503 17635
rect 24537 17601 24571 17635
rect 24605 17601 24639 17635
rect 24129 17532 24163 17566
rect 24197 17532 24231 17566
rect 24265 17532 24299 17566
rect 24333 17532 24367 17566
rect 24401 17532 24435 17566
rect 24469 17532 24503 17566
rect 24537 17532 24571 17566
rect 24605 17532 24639 17566
rect 24129 17463 24163 17497
rect 24197 17463 24231 17497
rect 24265 17463 24299 17497
rect 24333 17463 24367 17497
rect 24401 17463 24435 17497
rect 24469 17463 24503 17497
rect 24537 17463 24571 17497
rect 24605 17463 24639 17497
rect 24129 17394 24163 17428
rect 24197 17394 24231 17428
rect 24265 17394 24299 17428
rect 24333 17394 24367 17428
rect 24401 17394 24435 17428
rect 24469 17394 24503 17428
rect 24537 17394 24571 17428
rect 24605 17394 24639 17428
rect 24129 17325 24163 17359
rect 24197 17325 24231 17359
rect 24265 17325 24299 17359
rect 24333 17325 24367 17359
rect 24401 17325 24435 17359
rect 24469 17325 24503 17359
rect 24537 17325 24571 17359
rect 24605 17325 24639 17359
rect 24129 17256 24163 17290
rect 24197 17256 24231 17290
rect 24265 17256 24299 17290
rect 24333 17256 24367 17290
rect 24401 17256 24435 17290
rect 24469 17256 24503 17290
rect 24537 17256 24571 17290
rect 24605 17256 24639 17290
rect 24129 17187 24163 17221
rect 24197 17187 24231 17221
rect 24265 17187 24299 17221
rect 24333 17187 24367 17221
rect 24401 17187 24435 17221
rect 24469 17187 24503 17221
rect 24537 17187 24571 17221
rect 24605 17187 24639 17221
rect 24129 17118 24163 17152
rect 24197 17118 24231 17152
rect 24265 17118 24299 17152
rect 24333 17118 24367 17152
rect 24401 17118 24435 17152
rect 24469 17118 24503 17152
rect 24537 17118 24571 17152
rect 24605 17118 24639 17152
rect 24129 17049 24163 17083
rect 24197 17049 24231 17083
rect 24265 17049 24299 17083
rect 24333 17049 24367 17083
rect 24401 17049 24435 17083
rect 24469 17049 24503 17083
rect 24537 17049 24571 17083
rect 24605 17049 24639 17083
rect 24129 16980 24163 17014
rect 24197 16980 24231 17014
rect 24265 16980 24299 17014
rect 24333 16980 24367 17014
rect 24401 16980 24435 17014
rect 24469 16980 24503 17014
rect 24537 16980 24571 17014
rect 24605 16980 24639 17014
rect 24129 16911 24163 16945
rect 24197 16911 24231 16945
rect 24265 16911 24299 16945
rect 24333 16911 24367 16945
rect 24401 16911 24435 16945
rect 24469 16911 24503 16945
rect 24537 16911 24571 16945
rect 24605 16911 24639 16945
rect 24129 16842 24163 16876
rect 24197 16842 24231 16876
rect 24265 16842 24299 16876
rect 24333 16842 24367 16876
rect 24401 16842 24435 16876
rect 24469 16842 24503 16876
rect 24537 16842 24571 16876
rect 24605 16842 24639 16876
rect 24129 16773 24163 16807
rect 24197 16773 24231 16807
rect 24265 16773 24299 16807
rect 24333 16773 24367 16807
rect 24401 16773 24435 16807
rect 24469 16773 24503 16807
rect 24537 16773 24571 16807
rect 24605 16773 24639 16807
rect 24129 16704 24163 16738
rect 24197 16704 24231 16738
rect 24265 16704 24299 16738
rect 24333 16704 24367 16738
rect 24401 16704 24435 16738
rect 24469 16704 24503 16738
rect 24537 16704 24571 16738
rect 24605 16704 24639 16738
rect 24129 16635 24163 16669
rect 24197 16635 24231 16669
rect 24265 16635 24299 16669
rect 24333 16635 24367 16669
rect 24401 16635 24435 16669
rect 24469 16635 24503 16669
rect 24537 16635 24571 16669
rect 24605 16635 24639 16669
rect 24129 16566 24163 16600
rect 24197 16566 24231 16600
rect 24265 16566 24299 16600
rect 24333 16566 24367 16600
rect 24401 16566 24435 16600
rect 24469 16566 24503 16600
rect 24537 16566 24571 16600
rect 24605 16566 24639 16600
rect 24129 16497 24163 16531
rect 24197 16497 24231 16531
rect 24265 16497 24299 16531
rect 24333 16497 24367 16531
rect 24401 16497 24435 16531
rect 24469 16497 24503 16531
rect 24537 16497 24571 16531
rect 24605 16497 24639 16531
rect 24129 16428 24163 16462
rect 24197 16428 24231 16462
rect 24265 16428 24299 16462
rect 24333 16428 24367 16462
rect 24401 16428 24435 16462
rect 24469 16428 24503 16462
rect 24537 16428 24571 16462
rect 24605 16428 24639 16462
rect 27012 19198 27046 19232
rect 27012 19130 27046 19164
rect 27012 19062 27046 19096
rect 27012 18994 27046 19028
rect 27012 18926 27046 18960
rect 27012 18858 27046 18892
rect 27012 18790 27046 18824
rect 27012 18722 27046 18756
rect 27012 18654 27046 18688
rect 27012 18586 27046 18620
rect 27012 18518 27046 18552
rect 27012 18450 27046 18484
rect 27012 18382 27046 18416
rect 27012 18314 27046 18348
rect 27012 18246 27046 18280
rect 27012 18178 27046 18212
rect 27012 18110 27046 18144
rect 27012 18042 27046 18076
rect 27012 17974 27046 18008
rect 27012 17906 27046 17940
rect 27012 17838 27046 17872
rect 27012 17770 27046 17804
rect 27012 17702 27046 17736
rect 27012 17634 27046 17668
rect 27012 17566 27046 17600
rect 27012 17498 27046 17532
rect 27012 17430 27046 17464
rect 27012 17362 27046 17396
rect 27012 17294 27046 17328
rect 27012 17225 27046 17259
rect 27012 17156 27046 17190
rect 27012 17087 27046 17121
rect 27012 17018 27046 17052
rect 27012 16949 27046 16983
rect 27012 16880 27046 16914
rect 27012 16811 27046 16845
rect 27012 16742 27046 16776
rect 27012 16673 27046 16707
rect 27012 16604 27046 16638
rect 27012 16535 27046 16569
rect 27012 16466 27046 16500
rect 27012 16397 27046 16431
rect 27012 16328 27046 16362
rect 27012 16259 27046 16293
rect 27012 16190 27046 16224
rect 27012 16121 27046 16155
rect 27012 16052 27046 16086
rect 27012 15983 27046 16017
rect 27012 15914 27046 15948
rect 27012 15845 27046 15879
rect 27012 15776 27046 15810
rect 27012 15707 27046 15741
rect 27012 15638 27046 15672
rect 27012 15569 27046 15603
rect 27012 15500 27046 15534
rect 27012 15431 27046 15465
rect 27012 15362 27046 15396
rect 27012 15293 27046 15327
rect 27012 15224 27046 15258
rect 27012 15155 27046 15189
rect 27012 15086 27046 15120
rect 27012 15017 27046 15051
<< poly >>
rect 2246 33392 2646 33408
rect 2750 33392 3150 33408
rect 24970 10923 25266 11010
rect 24970 10906 25090 10923
rect 25146 10906 25266 10923
rect 25322 10923 25618 11010
rect 25322 10906 25442 10923
rect 25498 10906 25618 10923
<< locali >>
rect 27213 37619 27625 37620
rect 27213 37600 27287 37619
rect 27321 37614 27355 37619
rect 27389 37614 27423 37619
rect 27457 37614 27491 37619
rect 27525 37614 27625 37619
rect 27213 37566 27219 37600
rect 27253 37585 27287 37600
rect 27326 37585 27355 37614
rect 27399 37585 27423 37614
rect 27473 37585 27491 37614
rect 27547 37585 27625 37614
rect 27253 37580 27292 37585
rect 27326 37580 27365 37585
rect 27399 37580 27439 37585
rect 27473 37580 27513 37585
rect 27547 37580 27585 37585
rect 27253 37574 27585 37580
rect 27253 37566 27259 37574
rect 27213 37559 27259 37566
rect 27213 37525 27219 37559
rect 27253 37525 27259 37559
rect 27213 37514 27259 37525
rect 27579 37551 27585 37574
rect 27619 37551 27625 37585
rect 27579 37542 27625 37551
rect 27219 37491 27253 37514
rect 2097 37421 2166 37467
rect 27219 37423 27253 37457
rect 2097 37402 2143 37421
rect 27219 37379 27253 37389
rect 27334 37504 27504 37520
rect 27213 37355 27259 37379
rect 27213 37299 27219 37355
rect 27253 37299 27259 37355
rect 27334 37318 27504 37334
rect 27579 37483 27585 37542
rect 27619 37483 27625 37542
rect 27579 37470 27625 37483
rect 27579 37415 27585 37470
rect 27619 37415 27625 37470
rect 27579 37398 27625 37415
rect 27579 37347 27585 37398
rect 27619 37347 27625 37398
rect 27579 37325 27625 37347
rect 27213 37287 27259 37299
rect 27213 37253 27219 37287
rect 27253 37259 27259 37287
rect 27579 37291 27585 37325
rect 27619 37291 27625 37325
rect 27579 37259 27625 37291
rect 27253 37253 27625 37259
rect 27213 37219 27291 37253
rect 27325 37219 27347 37253
rect 27399 37219 27415 37253
rect 27473 37219 27483 37253
rect 27546 37219 27551 37253
rect 27585 37219 27625 37253
rect 27213 37213 27625 37219
rect 2244 34506 2256 34540
rect 2290 34506 2333 34540
rect 2367 34506 2410 34540
rect 2444 34506 2487 34540
rect 2521 34506 2564 34540
rect 2598 34506 2641 34540
rect 2675 34506 2718 34540
rect 2752 34506 2795 34540
rect 2829 34506 2872 34540
rect 2906 34506 2949 34540
rect 2983 34506 3026 34540
rect 3060 34506 3103 34540
rect 3137 34506 3152 34540
rect 2244 34468 3152 34506
rect 2244 34434 2256 34468
rect 2290 34434 2333 34468
rect 2367 34434 2410 34468
rect 2444 34434 2487 34468
rect 2521 34434 2564 34468
rect 2598 34434 2641 34468
rect 2675 34434 2718 34468
rect 2752 34434 2795 34468
rect 2829 34434 2872 34468
rect 2906 34434 2949 34468
rect 2983 34434 3026 34468
rect 3060 34434 3103 34468
rect 3137 34434 3152 34468
rect 2244 34396 3152 34434
rect 2244 34362 2256 34396
rect 2290 34362 2333 34396
rect 2367 34362 2410 34396
rect 2444 34362 2487 34396
rect 2521 34362 2564 34396
rect 2598 34362 2641 34396
rect 2675 34362 2718 34396
rect 2752 34362 2795 34396
rect 2829 34362 2872 34396
rect 2906 34362 2949 34396
rect 2983 34362 3026 34396
rect 3060 34362 3103 34396
rect 3137 34362 3152 34396
rect 2244 34132 3152 34362
rect 23661 23319 23747 23353
rect 23781 23319 23816 23353
rect 23850 23319 23885 23353
rect 23919 23319 23954 23353
rect 23988 23319 24023 23353
rect 24057 23319 24092 23353
rect 24126 23319 24161 23353
rect 24195 23319 24230 23353
rect 24264 23319 24299 23353
rect 24333 23319 24368 23353
rect 24402 23319 24437 23353
rect 24471 23319 24506 23353
rect 24540 23319 24575 23353
rect 24609 23319 24644 23353
rect 24678 23319 24713 23353
rect 24747 23319 24782 23353
rect 24816 23319 24851 23353
rect 24885 23319 24920 23353
rect 24954 23319 24989 23353
rect 25023 23319 25058 23353
rect 25092 23319 25127 23353
rect 25161 23319 25196 23353
rect 25230 23319 25265 23353
rect 25299 23319 25334 23353
rect 25368 23319 25403 23353
rect 25437 23319 25472 23353
rect 25506 23319 25541 23353
rect 25575 23319 25610 23353
rect 25644 23319 25679 23353
rect 25713 23319 25748 23353
rect 25782 23319 25817 23353
rect 25851 23319 25886 23353
rect 25920 23319 25955 23353
rect 25989 23319 26024 23353
rect 26058 23319 26093 23353
rect 26127 23319 26162 23353
rect 26196 23319 26231 23353
rect 26265 23319 26300 23353
rect 26334 23319 26368 23353
rect 26402 23319 26436 23353
rect 26470 23319 26504 23353
rect 26538 23319 26572 23353
rect 26606 23319 26640 23353
rect 26674 23319 26708 23353
rect 26742 23319 26776 23353
rect 26810 23319 26844 23353
rect 26878 23319 26912 23353
rect 26946 23319 26980 23353
rect 27014 23319 27048 23353
rect 27082 23319 27116 23353
rect 27150 23319 27184 23353
rect 27218 23319 27252 23353
rect 27286 23319 27320 23353
rect 27354 23319 27388 23353
rect 27422 23319 27456 23353
rect 27490 23319 27524 23353
rect 27558 23319 27592 23353
rect 27626 23319 27660 23353
rect 27694 23319 27728 23353
rect 27762 23319 27796 23353
rect 27830 23319 27864 23353
rect 27898 23319 27932 23353
rect 27966 23319 28029 23353
rect 23661 23284 28029 23319
rect 23661 23283 23806 23284
rect 23840 23283 23879 23284
rect 23913 23283 23952 23284
rect 23986 23283 24025 23284
rect 24059 23283 24098 23284
rect 24132 23283 24171 23284
rect 24205 23283 24244 23284
rect 24278 23283 24317 23284
rect 24351 23283 24390 23284
rect 24424 23283 24462 23284
rect 24496 23283 24534 23284
rect 24568 23283 24606 23284
rect 24640 23283 24678 23284
rect 23661 23249 23747 23283
rect 23781 23250 23806 23283
rect 23850 23250 23879 23283
rect 23919 23250 23952 23283
rect 23781 23249 23816 23250
rect 23850 23249 23885 23250
rect 23919 23249 23954 23250
rect 23988 23249 24023 23283
rect 24059 23250 24092 23283
rect 24132 23250 24161 23283
rect 24205 23250 24230 23283
rect 24278 23250 24299 23283
rect 24351 23250 24368 23283
rect 24424 23250 24437 23283
rect 24496 23250 24506 23283
rect 24568 23250 24575 23283
rect 24640 23250 24644 23283
rect 24057 23249 24092 23250
rect 24126 23249 24161 23250
rect 24195 23249 24230 23250
rect 24264 23249 24299 23250
rect 24333 23249 24368 23250
rect 24402 23249 24437 23250
rect 24471 23249 24506 23250
rect 24540 23249 24575 23250
rect 24609 23249 24644 23250
rect 24712 23283 24750 23284
rect 24784 23283 24822 23284
rect 24856 23283 24894 23284
rect 24928 23283 24966 23284
rect 25000 23283 25038 23284
rect 25072 23283 25110 23284
rect 25144 23283 25182 23284
rect 25216 23283 25254 23284
rect 25288 23283 25326 23284
rect 25360 23283 25398 23284
rect 25432 23283 25470 23284
rect 25504 23283 25542 23284
rect 25576 23283 25614 23284
rect 25648 23283 25686 23284
rect 25720 23283 25758 23284
rect 25792 23283 25830 23284
rect 25864 23283 25902 23284
rect 25936 23283 25974 23284
rect 26008 23283 26046 23284
rect 26080 23283 26118 23284
rect 26152 23283 26190 23284
rect 26224 23283 26262 23284
rect 26296 23283 26334 23284
rect 24712 23250 24713 23283
rect 24678 23249 24713 23250
rect 24747 23250 24750 23283
rect 24816 23250 24822 23283
rect 24885 23250 24894 23283
rect 24954 23250 24966 23283
rect 25023 23250 25038 23283
rect 25092 23250 25110 23283
rect 25161 23250 25182 23283
rect 25230 23250 25254 23283
rect 25299 23250 25326 23283
rect 25368 23250 25398 23283
rect 25437 23250 25470 23283
rect 24747 23249 24782 23250
rect 24816 23249 24851 23250
rect 24885 23249 24920 23250
rect 24954 23249 24989 23250
rect 25023 23249 25058 23250
rect 25092 23249 25127 23250
rect 25161 23249 25196 23250
rect 25230 23249 25265 23250
rect 25299 23249 25334 23250
rect 25368 23249 25403 23250
rect 25437 23249 25472 23250
rect 25506 23249 25541 23283
rect 25576 23250 25610 23283
rect 25648 23250 25679 23283
rect 25720 23250 25748 23283
rect 25792 23250 25817 23283
rect 25864 23250 25886 23283
rect 25936 23250 25955 23283
rect 26008 23250 26024 23283
rect 26080 23250 26093 23283
rect 26152 23250 26162 23283
rect 26224 23250 26231 23283
rect 26296 23250 26300 23283
rect 25575 23249 25610 23250
rect 25644 23249 25679 23250
rect 25713 23249 25748 23250
rect 25782 23249 25817 23250
rect 25851 23249 25886 23250
rect 25920 23249 25955 23250
rect 25989 23249 26024 23250
rect 26058 23249 26093 23250
rect 26127 23249 26162 23250
rect 26196 23249 26231 23250
rect 26265 23249 26300 23250
rect 26368 23283 26406 23284
rect 26440 23283 26478 23284
rect 26512 23283 26550 23284
rect 26584 23283 26622 23284
rect 26656 23283 26694 23284
rect 26728 23283 26766 23284
rect 26800 23283 26838 23284
rect 26872 23283 26910 23284
rect 26944 23283 26982 23284
rect 27016 23283 27054 23284
rect 27088 23283 27126 23284
rect 27160 23283 27198 23284
rect 27232 23283 27270 23284
rect 27304 23283 27342 23284
rect 27376 23283 27414 23284
rect 27448 23283 27486 23284
rect 27520 23283 27558 23284
rect 26334 23249 26368 23250
rect 26402 23250 26406 23283
rect 26470 23250 26478 23283
rect 26538 23250 26550 23283
rect 26606 23250 26622 23283
rect 26674 23250 26694 23283
rect 26742 23250 26766 23283
rect 26810 23250 26838 23283
rect 26878 23250 26910 23283
rect 26402 23249 26436 23250
rect 26470 23249 26504 23250
rect 26538 23249 26572 23250
rect 26606 23249 26640 23250
rect 26674 23249 26708 23250
rect 26742 23249 26776 23250
rect 26810 23249 26844 23250
rect 26878 23249 26912 23250
rect 26946 23249 26980 23283
rect 27016 23250 27048 23283
rect 27088 23250 27116 23283
rect 27160 23250 27184 23283
rect 27232 23250 27252 23283
rect 27304 23250 27320 23283
rect 27376 23250 27388 23283
rect 27448 23250 27456 23283
rect 27520 23250 27524 23283
rect 27014 23249 27048 23250
rect 27082 23249 27116 23250
rect 27150 23249 27184 23250
rect 27218 23249 27252 23250
rect 27286 23249 27320 23250
rect 27354 23249 27388 23250
rect 27422 23249 27456 23250
rect 27490 23249 27524 23250
rect 27592 23283 27630 23284
rect 27664 23283 27702 23284
rect 27736 23283 27774 23284
rect 27808 23283 27846 23284
rect 27880 23283 27918 23284
rect 27952 23283 28029 23284
rect 27558 23249 27592 23250
rect 27626 23250 27630 23283
rect 27694 23250 27702 23283
rect 27762 23250 27774 23283
rect 27830 23250 27846 23283
rect 27898 23250 27918 23283
rect 27626 23249 27660 23250
rect 27694 23249 27728 23250
rect 27762 23249 27796 23250
rect 27830 23249 27864 23250
rect 27898 23249 27932 23250
rect 27966 23249 28029 23283
rect 23661 23213 28029 23249
rect 23661 23179 23747 23213
rect 23781 23198 23816 23213
rect 23850 23198 23885 23213
rect 23919 23198 23954 23213
rect 23781 23179 23806 23198
rect 23850 23179 23879 23198
rect 23919 23179 23952 23198
rect 23988 23179 24023 23213
rect 24057 23198 24092 23213
rect 24126 23198 24161 23213
rect 24195 23198 24230 23213
rect 24264 23198 24299 23213
rect 24333 23198 24368 23213
rect 24402 23198 24437 23213
rect 24471 23198 24506 23213
rect 24540 23198 24575 23213
rect 24609 23198 24644 23213
rect 24059 23179 24092 23198
rect 24132 23179 24161 23198
rect 24205 23179 24230 23198
rect 24278 23179 24299 23198
rect 24351 23179 24368 23198
rect 24424 23179 24437 23198
rect 24496 23179 24506 23198
rect 24568 23179 24575 23198
rect 24640 23179 24644 23198
rect 24678 23198 24713 23213
rect 23661 23164 23806 23179
rect 23840 23164 23879 23179
rect 23913 23164 23952 23179
rect 23986 23164 24025 23179
rect 24059 23164 24098 23179
rect 24132 23164 24171 23179
rect 24205 23164 24244 23179
rect 24278 23164 24317 23179
rect 24351 23164 24390 23179
rect 24424 23164 24462 23179
rect 24496 23164 24534 23179
rect 24568 23164 24606 23179
rect 24640 23164 24678 23179
rect 24712 23179 24713 23198
rect 24747 23198 24782 23213
rect 24816 23198 24851 23213
rect 24885 23198 24920 23213
rect 24954 23198 24989 23213
rect 25023 23198 25058 23213
rect 25092 23198 25127 23213
rect 25161 23198 25196 23213
rect 25230 23198 25265 23213
rect 25299 23198 25334 23213
rect 25368 23198 25403 23213
rect 25437 23198 25472 23213
rect 24747 23179 24750 23198
rect 24816 23179 24822 23198
rect 24885 23179 24894 23198
rect 24954 23179 24966 23198
rect 25023 23179 25038 23198
rect 25092 23179 25110 23198
rect 25161 23179 25182 23198
rect 25230 23179 25254 23198
rect 25299 23179 25326 23198
rect 25368 23179 25398 23198
rect 25437 23179 25470 23198
rect 25506 23179 25541 23213
rect 25575 23198 25610 23213
rect 25644 23198 25679 23213
rect 25713 23198 25748 23213
rect 25782 23198 25817 23213
rect 25851 23198 25886 23213
rect 25920 23198 25955 23213
rect 25989 23198 26024 23213
rect 26058 23198 26093 23213
rect 26127 23198 26162 23213
rect 26196 23198 26231 23213
rect 26265 23198 26300 23213
rect 25576 23179 25610 23198
rect 25648 23179 25679 23198
rect 25720 23179 25748 23198
rect 25792 23179 25817 23198
rect 25864 23179 25886 23198
rect 25936 23179 25955 23198
rect 26008 23179 26024 23198
rect 26080 23179 26093 23198
rect 26152 23179 26162 23198
rect 26224 23179 26231 23198
rect 26296 23179 26300 23198
rect 26334 23198 26368 23213
rect 24712 23164 24750 23179
rect 24784 23164 24822 23179
rect 24856 23164 24894 23179
rect 24928 23164 24966 23179
rect 25000 23164 25038 23179
rect 25072 23164 25110 23179
rect 25144 23164 25182 23179
rect 25216 23164 25254 23179
rect 25288 23164 25326 23179
rect 25360 23164 25398 23179
rect 25432 23164 25470 23179
rect 25504 23164 25542 23179
rect 25576 23164 25614 23179
rect 25648 23164 25686 23179
rect 25720 23164 25758 23179
rect 25792 23164 25830 23179
rect 25864 23164 25902 23179
rect 25936 23164 25974 23179
rect 26008 23164 26046 23179
rect 26080 23164 26118 23179
rect 26152 23164 26190 23179
rect 26224 23164 26262 23179
rect 26296 23164 26334 23179
rect 26402 23198 26436 23213
rect 26470 23198 26504 23213
rect 26538 23198 26572 23213
rect 26606 23198 26640 23213
rect 26674 23198 26708 23213
rect 26742 23198 26776 23213
rect 26810 23198 26844 23213
rect 26878 23198 26912 23213
rect 26402 23179 26406 23198
rect 26470 23179 26478 23198
rect 26538 23179 26550 23198
rect 26606 23179 26622 23198
rect 26674 23179 26694 23198
rect 26742 23179 26766 23198
rect 26810 23179 26838 23198
rect 26878 23179 26910 23198
rect 26946 23179 26980 23213
rect 27014 23198 27048 23213
rect 27082 23198 27116 23213
rect 27150 23198 27184 23213
rect 27218 23198 27252 23213
rect 27286 23198 27320 23213
rect 27354 23198 27388 23213
rect 27422 23198 27456 23213
rect 27490 23198 27524 23213
rect 27016 23179 27048 23198
rect 27088 23179 27116 23198
rect 27160 23179 27184 23198
rect 27232 23179 27252 23198
rect 27304 23179 27320 23198
rect 27376 23179 27388 23198
rect 27448 23179 27456 23198
rect 27520 23179 27524 23198
rect 27558 23198 27592 23213
rect 26368 23164 26406 23179
rect 26440 23164 26478 23179
rect 26512 23164 26550 23179
rect 26584 23164 26622 23179
rect 26656 23164 26694 23179
rect 26728 23164 26766 23179
rect 26800 23164 26838 23179
rect 26872 23164 26910 23179
rect 26944 23164 26982 23179
rect 27016 23164 27054 23179
rect 27088 23164 27126 23179
rect 27160 23164 27198 23179
rect 27232 23164 27270 23179
rect 27304 23164 27342 23179
rect 27376 23164 27414 23179
rect 27448 23164 27486 23179
rect 27520 23164 27558 23179
rect 27626 23198 27660 23213
rect 27694 23198 27728 23213
rect 27762 23198 27796 23213
rect 27830 23198 27864 23213
rect 27898 23198 27932 23213
rect 27626 23179 27630 23198
rect 27694 23179 27702 23198
rect 27762 23179 27774 23198
rect 27830 23179 27846 23198
rect 27898 23179 27918 23198
rect 27966 23179 28029 23213
rect 27592 23164 27630 23179
rect 27664 23164 27702 23179
rect 27736 23164 27774 23179
rect 27808 23164 27846 23179
rect 27880 23164 27918 23179
rect 27952 23164 28029 23179
rect 23661 23143 28029 23164
rect 23661 23109 23747 23143
rect 23781 23112 23816 23143
rect 23850 23112 23885 23143
rect 23919 23112 23954 23143
rect 23781 23109 23806 23112
rect 23850 23109 23879 23112
rect 23919 23109 23952 23112
rect 23988 23109 24023 23143
rect 24057 23112 24092 23143
rect 24126 23112 24161 23143
rect 24195 23112 24230 23143
rect 24264 23112 24299 23143
rect 24333 23112 24368 23143
rect 24402 23112 24437 23143
rect 24471 23112 24506 23143
rect 24540 23112 24575 23143
rect 24609 23112 24644 23143
rect 24059 23109 24092 23112
rect 24132 23109 24161 23112
rect 24205 23109 24230 23112
rect 24278 23109 24299 23112
rect 24351 23109 24368 23112
rect 24424 23109 24437 23112
rect 24496 23109 24506 23112
rect 24568 23109 24575 23112
rect 24640 23109 24644 23112
rect 24678 23112 24713 23143
rect 23661 23078 23806 23109
rect 23840 23078 23879 23109
rect 23913 23078 23952 23109
rect 23986 23078 24025 23109
rect 24059 23078 24098 23109
rect 24132 23078 24171 23109
rect 24205 23078 24244 23109
rect 24278 23078 24317 23109
rect 24351 23078 24390 23109
rect 24424 23078 24462 23109
rect 24496 23078 24534 23109
rect 24568 23078 24606 23109
rect 24640 23078 24678 23109
rect 24712 23109 24713 23112
rect 24747 23112 24782 23143
rect 24816 23112 24851 23143
rect 24885 23112 24920 23143
rect 24954 23112 24989 23143
rect 25023 23112 25058 23143
rect 25092 23112 25127 23143
rect 25161 23112 25196 23143
rect 25230 23112 25265 23143
rect 25299 23112 25334 23143
rect 25368 23112 25403 23143
rect 25437 23112 25472 23143
rect 24747 23109 24750 23112
rect 24816 23109 24822 23112
rect 24885 23109 24894 23112
rect 24954 23109 24966 23112
rect 25023 23109 25038 23112
rect 25092 23109 25110 23112
rect 25161 23109 25182 23112
rect 25230 23109 25254 23112
rect 25299 23109 25326 23112
rect 25368 23109 25398 23112
rect 25437 23109 25470 23112
rect 25506 23109 25541 23143
rect 25575 23112 25610 23143
rect 25644 23112 25679 23143
rect 25713 23112 25748 23143
rect 25782 23112 25817 23143
rect 25851 23112 25886 23143
rect 25920 23112 25955 23143
rect 25989 23112 26024 23143
rect 26058 23112 26093 23143
rect 26127 23112 26162 23143
rect 26196 23112 26231 23143
rect 26265 23112 26300 23143
rect 25576 23109 25610 23112
rect 25648 23109 25679 23112
rect 25720 23109 25748 23112
rect 25792 23109 25817 23112
rect 25864 23109 25886 23112
rect 25936 23109 25955 23112
rect 26008 23109 26024 23112
rect 26080 23109 26093 23112
rect 26152 23109 26162 23112
rect 26224 23109 26231 23112
rect 26296 23109 26300 23112
rect 26334 23112 26368 23143
rect 24712 23078 24750 23109
rect 24784 23078 24822 23109
rect 24856 23078 24894 23109
rect 24928 23078 24966 23109
rect 25000 23078 25038 23109
rect 25072 23078 25110 23109
rect 25144 23078 25182 23109
rect 25216 23078 25254 23109
rect 25288 23078 25326 23109
rect 25360 23078 25398 23109
rect 25432 23078 25470 23109
rect 25504 23078 25542 23109
rect 25576 23078 25614 23109
rect 25648 23078 25686 23109
rect 25720 23078 25758 23109
rect 25792 23078 25830 23109
rect 25864 23078 25902 23109
rect 25936 23078 25974 23109
rect 26008 23078 26046 23109
rect 26080 23078 26118 23109
rect 26152 23078 26190 23109
rect 26224 23078 26262 23109
rect 26296 23078 26334 23109
rect 26402 23112 26436 23143
rect 26470 23112 26504 23143
rect 26538 23112 26572 23143
rect 26606 23112 26640 23143
rect 26674 23112 26708 23143
rect 26742 23112 26776 23143
rect 26810 23112 26844 23143
rect 26878 23112 26912 23143
rect 26402 23109 26406 23112
rect 26470 23109 26478 23112
rect 26538 23109 26550 23112
rect 26606 23109 26622 23112
rect 26674 23109 26694 23112
rect 26742 23109 26766 23112
rect 26810 23109 26838 23112
rect 26878 23109 26910 23112
rect 26946 23109 26980 23143
rect 27014 23112 27048 23143
rect 27082 23112 27116 23143
rect 27150 23112 27184 23143
rect 27218 23112 27252 23143
rect 27286 23112 27320 23143
rect 27354 23112 27388 23143
rect 27422 23112 27456 23143
rect 27490 23112 27524 23143
rect 27016 23109 27048 23112
rect 27088 23109 27116 23112
rect 27160 23109 27184 23112
rect 27232 23109 27252 23112
rect 27304 23109 27320 23112
rect 27376 23109 27388 23112
rect 27448 23109 27456 23112
rect 27520 23109 27524 23112
rect 27558 23112 27592 23143
rect 26368 23078 26406 23109
rect 26440 23078 26478 23109
rect 26512 23078 26550 23109
rect 26584 23078 26622 23109
rect 26656 23078 26694 23109
rect 26728 23078 26766 23109
rect 26800 23078 26838 23109
rect 26872 23078 26910 23109
rect 26944 23078 26982 23109
rect 27016 23078 27054 23109
rect 27088 23078 27126 23109
rect 27160 23078 27198 23109
rect 27232 23078 27270 23109
rect 27304 23078 27342 23109
rect 27376 23078 27414 23109
rect 27448 23078 27486 23109
rect 27520 23078 27558 23109
rect 27626 23112 27660 23143
rect 27694 23112 27728 23143
rect 27762 23112 27796 23143
rect 27830 23112 27864 23143
rect 27898 23112 27932 23143
rect 27626 23109 27630 23112
rect 27694 23109 27702 23112
rect 27762 23109 27774 23112
rect 27830 23109 27846 23112
rect 27898 23109 27918 23112
rect 27966 23109 28029 23143
rect 27592 23078 27630 23109
rect 27664 23078 27702 23109
rect 27736 23078 27774 23109
rect 27808 23078 27846 23109
rect 27880 23078 27918 23109
rect 27952 23078 28029 23109
rect 23661 23073 28029 23078
rect 23661 23039 23747 23073
rect 23781 23039 23816 23073
rect 23850 23039 23885 23073
rect 23919 23039 23954 23073
rect 23988 23039 24023 23073
rect 24057 23039 24092 23073
rect 24126 23039 24161 23073
rect 24195 23039 24230 23073
rect 24264 23039 24299 23073
rect 24333 23039 24368 23073
rect 24402 23039 24437 23073
rect 24471 23039 24506 23073
rect 24540 23039 24575 23073
rect 24609 23039 24644 23073
rect 24678 23039 24713 23073
rect 24747 23039 24782 23073
rect 24816 23039 24851 23073
rect 24885 23039 24920 23073
rect 24954 23039 24989 23073
rect 25023 23039 25058 23073
rect 25092 23039 25127 23073
rect 25161 23039 25196 23073
rect 25230 23039 25265 23073
rect 25299 23039 25334 23073
rect 25368 23039 25403 23073
rect 25437 23039 25472 23073
rect 25506 23039 25541 23073
rect 25575 23039 25610 23073
rect 25644 23039 25679 23073
rect 25713 23039 25748 23073
rect 25782 23039 25817 23073
rect 25851 23039 25886 23073
rect 25920 23039 25955 23073
rect 25989 23039 26024 23073
rect 26058 23039 26093 23073
rect 26127 23039 26162 23073
rect 26196 23039 26231 23073
rect 26265 23039 26300 23073
rect 26334 23039 26368 23073
rect 26402 23039 26436 23073
rect 26470 23039 26504 23073
rect 26538 23039 26572 23073
rect 26606 23039 26640 23073
rect 26674 23039 26708 23073
rect 26742 23039 26776 23073
rect 26810 23039 26844 23073
rect 26878 23039 26912 23073
rect 26946 23039 26980 23073
rect 27014 23039 27048 23073
rect 27082 23039 27116 23073
rect 27150 23039 27184 23073
rect 27218 23039 27252 23073
rect 27286 23039 27320 23073
rect 27354 23039 27388 23073
rect 27422 23039 27456 23073
rect 27490 23039 27524 23073
rect 27558 23039 27592 23073
rect 27626 23039 27660 23073
rect 27694 23039 27728 23073
rect 27762 23039 27796 23073
rect 27830 23039 27864 23073
rect 27898 23039 27932 23073
rect 27966 23039 28029 23073
rect 23661 23026 28029 23039
rect 23661 23003 23806 23026
rect 23840 23003 23879 23026
rect 23913 23003 23952 23026
rect 23986 23003 24025 23026
rect 24059 23003 24098 23026
rect 24132 23003 24171 23026
rect 24205 23003 24244 23026
rect 24278 23003 24317 23026
rect 24351 23003 24390 23026
rect 24424 23003 24462 23026
rect 24496 23003 24534 23026
rect 24568 23003 24606 23026
rect 24640 23003 24678 23026
rect 23661 22969 23747 23003
rect 23781 22992 23806 23003
rect 23850 22992 23879 23003
rect 23919 22992 23952 23003
rect 23781 22969 23816 22992
rect 23850 22969 23885 22992
rect 23919 22969 23954 22992
rect 23988 22969 24023 23003
rect 24059 22992 24092 23003
rect 24132 22992 24161 23003
rect 24205 22992 24230 23003
rect 24278 22992 24299 23003
rect 24351 22992 24368 23003
rect 24424 22992 24437 23003
rect 24496 22992 24506 23003
rect 24568 22992 24575 23003
rect 24640 22992 24644 23003
rect 24057 22969 24092 22992
rect 24126 22969 24161 22992
rect 24195 22969 24230 22992
rect 24264 22969 24299 22992
rect 24333 22969 24368 22992
rect 24402 22969 24437 22992
rect 24471 22969 24506 22992
rect 24540 22969 24575 22992
rect 24609 22969 24644 22992
rect 24712 23003 24750 23026
rect 24784 23003 24822 23026
rect 24856 23003 24894 23026
rect 24928 23003 24966 23026
rect 25000 23003 25038 23026
rect 25072 23003 25110 23026
rect 25144 23003 25182 23026
rect 25216 23003 25254 23026
rect 25288 23003 25326 23026
rect 25360 23003 25398 23026
rect 25432 23003 25470 23026
rect 25504 23003 25542 23026
rect 25576 23003 25614 23026
rect 25648 23003 25686 23026
rect 25720 23003 25758 23026
rect 25792 23003 25830 23026
rect 25864 23003 25902 23026
rect 25936 23003 25974 23026
rect 26008 23003 26046 23026
rect 26080 23003 26118 23026
rect 26152 23003 26190 23026
rect 26224 23003 26262 23026
rect 26296 23003 26334 23026
rect 24712 22992 24713 23003
rect 24678 22969 24713 22992
rect 24747 22992 24750 23003
rect 24816 22992 24822 23003
rect 24885 22992 24894 23003
rect 24954 22992 24966 23003
rect 25023 22992 25038 23003
rect 25092 22992 25110 23003
rect 25161 22992 25182 23003
rect 25230 22992 25254 23003
rect 25299 22992 25326 23003
rect 25368 22992 25398 23003
rect 25437 22992 25470 23003
rect 24747 22969 24782 22992
rect 24816 22969 24851 22992
rect 24885 22969 24920 22992
rect 24954 22969 24989 22992
rect 25023 22969 25058 22992
rect 25092 22969 25127 22992
rect 25161 22969 25196 22992
rect 25230 22969 25265 22992
rect 25299 22969 25334 22992
rect 25368 22969 25403 22992
rect 25437 22969 25472 22992
rect 25506 22969 25541 23003
rect 25576 22992 25610 23003
rect 25648 22992 25679 23003
rect 25720 22992 25748 23003
rect 25792 22992 25817 23003
rect 25864 22992 25886 23003
rect 25936 22992 25955 23003
rect 26008 22992 26024 23003
rect 26080 22992 26093 23003
rect 26152 22992 26162 23003
rect 26224 22992 26231 23003
rect 26296 22992 26300 23003
rect 25575 22969 25610 22992
rect 25644 22969 25679 22992
rect 25713 22969 25748 22992
rect 25782 22969 25817 22992
rect 25851 22969 25886 22992
rect 25920 22969 25955 22992
rect 25989 22969 26024 22992
rect 26058 22969 26093 22992
rect 26127 22969 26162 22992
rect 26196 22969 26231 22992
rect 26265 22969 26300 22992
rect 26368 23003 26406 23026
rect 26440 23003 26478 23026
rect 26512 23003 26550 23026
rect 26584 23003 26622 23026
rect 26656 23003 26694 23026
rect 26728 23003 26766 23026
rect 26800 23003 26838 23026
rect 26872 23003 26910 23026
rect 26944 23003 26982 23026
rect 27016 23003 27054 23026
rect 27088 23003 27126 23026
rect 27160 23003 27198 23026
rect 27232 23003 27270 23026
rect 27304 23003 27342 23026
rect 27376 23003 27414 23026
rect 27448 23003 27486 23026
rect 27520 23003 27558 23026
rect 26334 22969 26368 22992
rect 26402 22992 26406 23003
rect 26470 22992 26478 23003
rect 26538 22992 26550 23003
rect 26606 22992 26622 23003
rect 26674 22992 26694 23003
rect 26742 22992 26766 23003
rect 26810 22992 26838 23003
rect 26878 22992 26910 23003
rect 26402 22969 26436 22992
rect 26470 22969 26504 22992
rect 26538 22969 26572 22992
rect 26606 22969 26640 22992
rect 26674 22969 26708 22992
rect 26742 22969 26776 22992
rect 26810 22969 26844 22992
rect 26878 22969 26912 22992
rect 26946 22969 26980 23003
rect 27016 22992 27048 23003
rect 27088 22992 27116 23003
rect 27160 22992 27184 23003
rect 27232 22992 27252 23003
rect 27304 22992 27320 23003
rect 27376 22992 27388 23003
rect 27448 22992 27456 23003
rect 27520 22992 27524 23003
rect 27014 22969 27048 22992
rect 27082 22969 27116 22992
rect 27150 22969 27184 22992
rect 27218 22969 27252 22992
rect 27286 22969 27320 22992
rect 27354 22969 27388 22992
rect 27422 22969 27456 22992
rect 27490 22969 27524 22992
rect 27592 23003 27630 23026
rect 27664 23003 27702 23026
rect 27736 23003 27774 23026
rect 27808 23003 27846 23026
rect 27880 23003 27918 23026
rect 27952 23003 28029 23026
rect 27558 22969 27592 22992
rect 27626 22992 27630 23003
rect 27694 22992 27702 23003
rect 27762 22992 27774 23003
rect 27830 22992 27846 23003
rect 27898 22992 27918 23003
rect 27626 22969 27660 22992
rect 27694 22969 27728 22992
rect 27762 22969 27796 22992
rect 27830 22969 27864 22992
rect 27898 22969 27932 22992
rect 27966 22969 28029 23003
rect 23661 22933 28029 22969
rect 23661 22899 23747 22933
rect 23781 22899 23816 22933
rect 23850 22899 23885 22933
rect 23919 22899 23954 22933
rect 23988 22899 24023 22933
rect 24057 22899 24092 22933
rect 24126 22899 24161 22933
rect 24195 22899 24230 22933
rect 24264 22899 24299 22933
rect 24333 22899 24368 22933
rect 24402 22899 24437 22933
rect 24471 22899 24506 22933
rect 24540 22899 24575 22933
rect 24609 22899 24644 22933
rect 24678 22899 24713 22933
rect 24747 22899 24782 22933
rect 24816 22899 24851 22933
rect 24885 22899 24920 22933
rect 24954 22899 24989 22933
rect 25023 22899 25058 22933
rect 25092 22899 25127 22933
rect 25161 22899 25196 22933
rect 25230 22899 25265 22933
rect 25299 22899 25334 22933
rect 25368 22899 25403 22933
rect 25437 22899 25472 22933
rect 25506 22899 25541 22933
rect 25575 22899 25610 22933
rect 25644 22899 25679 22933
rect 25713 22899 25748 22933
rect 25782 22899 25817 22933
rect 25851 22899 25886 22933
rect 25920 22899 25955 22933
rect 25989 22899 26024 22933
rect 26058 22899 26093 22933
rect 26127 22899 26162 22933
rect 26196 22899 26231 22933
rect 26265 22899 26300 22933
rect 26334 22899 26368 22933
rect 26402 22899 26436 22933
rect 26470 22899 26504 22933
rect 26538 22899 26572 22933
rect 26606 22899 26640 22933
rect 26674 22899 26708 22933
rect 26742 22899 26776 22933
rect 26810 22899 26844 22933
rect 26878 22899 26912 22933
rect 26946 22899 26980 22933
rect 27014 22899 27048 22933
rect 27082 22899 27116 22933
rect 27150 22899 27184 22933
rect 27218 22899 27252 22933
rect 27286 22899 27320 22933
rect 27354 22899 27388 22933
rect 27422 22899 27456 22933
rect 27490 22899 27524 22933
rect 27558 22899 27592 22933
rect 27626 22899 27660 22933
rect 27694 22899 27728 22933
rect 27762 22899 27796 22933
rect 27830 22899 27864 22933
rect 27898 22899 27932 22933
rect 27966 22899 28029 22933
rect 26275 22890 28029 22899
rect 26275 22856 26434 22890
rect 26468 22856 26509 22890
rect 26543 22856 26584 22890
rect 26618 22856 26659 22890
rect 26693 22856 26734 22890
rect 26768 22856 26808 22890
rect 26842 22856 26882 22890
rect 26916 22856 26956 22890
rect 26990 22856 27030 22890
rect 27064 22856 27104 22890
rect 27138 22856 27178 22890
rect 27212 22856 27252 22890
rect 27286 22856 27326 22890
rect 27360 22856 27400 22890
rect 27434 22856 27474 22890
rect 27508 22856 27548 22890
rect 27582 22856 27622 22890
rect 27656 22856 27696 22890
rect 27730 22856 27770 22890
rect 27804 22856 27844 22890
rect 27878 22856 27918 22890
rect 27952 22856 28029 22890
rect 26275 22822 26309 22856
rect 26343 22822 26380 22856
rect 26414 22822 26451 22856
rect 26485 22822 26522 22856
rect 26556 22822 26593 22856
rect 26627 22822 26664 22856
rect 26698 22822 26735 22856
rect 26769 22822 26806 22856
rect 26840 22822 26877 22856
rect 26911 22822 26948 22856
rect 26982 22822 27019 22856
rect 27053 22822 27090 22856
rect 27124 22822 27161 22856
rect 27195 22822 27232 22856
rect 27266 22822 27302 22856
rect 27336 22822 27372 22856
rect 27406 22822 27442 22856
rect 27476 22822 27512 22856
rect 27546 22822 27582 22856
rect 27616 22822 27652 22856
rect 27686 22822 27722 22856
rect 27756 22822 27792 22856
rect 27826 22822 27862 22856
rect 27896 22822 27932 22856
rect 27966 22822 28029 22856
rect 26275 22818 28029 22822
rect 26275 22784 26434 22818
rect 26468 22784 26509 22818
rect 26543 22784 26584 22818
rect 26618 22784 26659 22818
rect 26693 22784 26734 22818
rect 26768 22784 26808 22818
rect 26842 22784 26882 22818
rect 26916 22784 26956 22818
rect 26990 22784 27030 22818
rect 27064 22784 27104 22818
rect 27138 22784 27178 22818
rect 27212 22784 27252 22818
rect 27286 22784 27326 22818
rect 27360 22784 27400 22818
rect 27434 22784 27474 22818
rect 27508 22784 27548 22818
rect 27582 22784 27622 22818
rect 27656 22784 27696 22818
rect 27730 22784 27770 22818
rect 27804 22784 27844 22818
rect 27878 22784 27918 22818
rect 27952 22784 28029 22818
rect 26275 22782 28029 22784
rect 26275 22748 26309 22782
rect 26343 22748 26380 22782
rect 26414 22748 26451 22782
rect 26485 22748 26522 22782
rect 26556 22748 26593 22782
rect 26627 22748 26664 22782
rect 26698 22748 26735 22782
rect 26769 22748 26806 22782
rect 26840 22748 26877 22782
rect 26911 22748 26948 22782
rect 26982 22748 27019 22782
rect 27053 22748 27090 22782
rect 27124 22748 27161 22782
rect 27195 22748 27232 22782
rect 27266 22748 27302 22782
rect 27336 22748 27372 22782
rect 27406 22748 27442 22782
rect 27476 22748 27512 22782
rect 27546 22748 27582 22782
rect 27616 22748 27652 22782
rect 27686 22748 27722 22782
rect 27756 22748 27792 22782
rect 27826 22748 27862 22782
rect 27896 22748 27932 22782
rect 27966 22748 28029 22782
rect 26275 22746 28029 22748
rect 26275 22712 26434 22746
rect 26468 22712 26509 22746
rect 26543 22712 26584 22746
rect 26618 22712 26659 22746
rect 26693 22712 26734 22746
rect 26768 22712 26808 22746
rect 26842 22712 26882 22746
rect 26916 22712 26956 22746
rect 26990 22712 27030 22746
rect 27064 22712 27104 22746
rect 27138 22712 27178 22746
rect 27212 22712 27252 22746
rect 27286 22712 27326 22746
rect 27360 22712 27400 22746
rect 27434 22712 27474 22746
rect 27508 22712 27548 22746
rect 27582 22712 27622 22746
rect 27656 22712 27696 22746
rect 27730 22712 27770 22746
rect 27804 22712 27844 22746
rect 27878 22712 27918 22746
rect 27952 22712 28029 22746
rect 26275 22708 28029 22712
rect 26275 22674 26309 22708
rect 26343 22674 26380 22708
rect 26414 22674 26451 22708
rect 26485 22674 26522 22708
rect 26556 22674 26593 22708
rect 26627 22674 26664 22708
rect 26698 22674 26735 22708
rect 26769 22674 26806 22708
rect 26840 22674 26877 22708
rect 26911 22674 26948 22708
rect 26982 22674 27019 22708
rect 27053 22674 27090 22708
rect 27124 22674 27161 22708
rect 27195 22674 27232 22708
rect 27266 22674 27302 22708
rect 27336 22674 27372 22708
rect 27406 22674 27442 22708
rect 27476 22674 27512 22708
rect 27546 22674 27582 22708
rect 27616 22674 27652 22708
rect 27686 22674 27722 22708
rect 27756 22674 27792 22708
rect 27826 22674 27862 22708
rect 27896 22674 27932 22708
rect 27966 22674 28029 22708
rect 26275 22640 26434 22674
rect 26468 22640 26509 22674
rect 26543 22640 26584 22674
rect 26618 22640 26659 22674
rect 26693 22640 26734 22674
rect 26768 22640 26808 22674
rect 26842 22640 26882 22674
rect 26916 22640 26956 22674
rect 26990 22640 27030 22674
rect 27064 22640 27104 22674
rect 27138 22640 27178 22674
rect 27212 22640 27252 22674
rect 27286 22640 27326 22674
rect 27360 22640 27400 22674
rect 27434 22640 27474 22674
rect 27508 22640 27548 22674
rect 27582 22640 27622 22674
rect 27656 22640 27696 22674
rect 27730 22640 27770 22674
rect 27804 22640 27844 22674
rect 27878 22640 27918 22674
rect 27952 22640 28029 22674
rect 26275 22634 28029 22640
rect 26275 22600 26309 22634
rect 26343 22600 26380 22634
rect 26414 22602 26451 22634
rect 26485 22602 26522 22634
rect 26556 22602 26593 22634
rect 26627 22602 26664 22634
rect 26698 22602 26735 22634
rect 26414 22600 26434 22602
rect 26485 22600 26509 22602
rect 26556 22600 26584 22602
rect 26627 22600 26659 22602
rect 26698 22600 26734 22602
rect 26769 22600 26806 22634
rect 26840 22602 26877 22634
rect 26911 22602 26948 22634
rect 26982 22602 27019 22634
rect 27053 22602 27090 22634
rect 27124 22602 27161 22634
rect 27195 22602 27232 22634
rect 27266 22602 27302 22634
rect 27336 22602 27372 22634
rect 27406 22602 27442 22634
rect 27476 22602 27512 22634
rect 26842 22600 26877 22602
rect 26916 22600 26948 22602
rect 26990 22600 27019 22602
rect 27064 22600 27090 22602
rect 27138 22600 27161 22602
rect 27212 22600 27232 22602
rect 27286 22600 27302 22602
rect 27360 22600 27372 22602
rect 27434 22600 27442 22602
rect 27508 22600 27512 22602
rect 27546 22602 27582 22634
rect 27546 22600 27548 22602
rect 26275 22568 26434 22600
rect 26468 22568 26509 22600
rect 26543 22568 26584 22600
rect 26618 22568 26659 22600
rect 26693 22568 26734 22600
rect 26768 22568 26808 22600
rect 26842 22568 26882 22600
rect 26916 22568 26956 22600
rect 26990 22568 27030 22600
rect 27064 22568 27104 22600
rect 27138 22568 27178 22600
rect 27212 22568 27252 22600
rect 27286 22568 27326 22600
rect 27360 22568 27400 22600
rect 27434 22568 27474 22600
rect 27508 22568 27548 22600
rect 27616 22602 27652 22634
rect 27686 22602 27722 22634
rect 27756 22602 27792 22634
rect 27826 22602 27862 22634
rect 27896 22602 27932 22634
rect 27616 22600 27622 22602
rect 27686 22600 27696 22602
rect 27756 22600 27770 22602
rect 27826 22600 27844 22602
rect 27896 22600 27918 22602
rect 27966 22600 28029 22634
rect 27582 22568 27622 22600
rect 27656 22568 27696 22600
rect 27730 22568 27770 22600
rect 27804 22568 27844 22600
rect 27878 22568 27918 22600
rect 27952 22568 28029 22600
rect 26275 22560 28029 22568
rect 26275 22526 26309 22560
rect 26343 22526 26380 22560
rect 26414 22530 26451 22560
rect 26485 22530 26522 22560
rect 26556 22530 26593 22560
rect 26627 22530 26664 22560
rect 26698 22530 26735 22560
rect 26414 22526 26434 22530
rect 26485 22526 26509 22530
rect 26556 22526 26584 22530
rect 26627 22526 26659 22530
rect 26698 22526 26734 22530
rect 26769 22526 26806 22560
rect 26840 22530 26877 22560
rect 26911 22530 26948 22560
rect 26982 22530 27019 22560
rect 27053 22530 27090 22560
rect 27124 22530 27161 22560
rect 27195 22530 27232 22560
rect 27266 22530 27302 22560
rect 27336 22530 27372 22560
rect 27406 22530 27442 22560
rect 27476 22530 27512 22560
rect 26842 22526 26877 22530
rect 26916 22526 26948 22530
rect 26990 22526 27019 22530
rect 27064 22526 27090 22530
rect 27138 22526 27161 22530
rect 27212 22526 27232 22530
rect 27286 22526 27302 22530
rect 27360 22526 27372 22530
rect 27434 22526 27442 22530
rect 27508 22526 27512 22530
rect 27546 22530 27582 22560
rect 27546 22526 27548 22530
rect 26275 22496 26434 22526
rect 26468 22496 26509 22526
rect 26543 22496 26584 22526
rect 26618 22496 26659 22526
rect 26693 22496 26734 22526
rect 26768 22496 26808 22526
rect 26842 22496 26882 22526
rect 26916 22496 26956 22526
rect 26990 22496 27030 22526
rect 27064 22496 27104 22526
rect 27138 22496 27178 22526
rect 27212 22496 27252 22526
rect 27286 22496 27326 22526
rect 27360 22496 27400 22526
rect 27434 22496 27474 22526
rect 27508 22496 27548 22526
rect 27616 22530 27652 22560
rect 27686 22530 27722 22560
rect 27756 22530 27792 22560
rect 27826 22530 27862 22560
rect 27896 22530 27932 22560
rect 27616 22526 27622 22530
rect 27686 22526 27696 22530
rect 27756 22526 27770 22530
rect 27826 22526 27844 22530
rect 27896 22526 27918 22530
rect 27966 22526 28029 22560
rect 27582 22496 27622 22526
rect 27656 22496 27696 22526
rect 27730 22496 27770 22526
rect 27804 22496 27844 22526
rect 27878 22496 27918 22526
rect 27952 22496 28029 22526
rect 26275 22486 28029 22496
rect 26275 22452 26309 22486
rect 26343 22452 26380 22486
rect 26414 22458 26451 22486
rect 26485 22458 26522 22486
rect 26556 22458 26593 22486
rect 26627 22458 26664 22486
rect 26698 22458 26735 22486
rect 26414 22452 26434 22458
rect 26485 22452 26509 22458
rect 26556 22452 26584 22458
rect 26627 22452 26659 22458
rect 26698 22452 26734 22458
rect 26769 22452 26806 22486
rect 26840 22458 26877 22486
rect 26911 22458 26948 22486
rect 26982 22458 27019 22486
rect 27053 22458 27090 22486
rect 27124 22458 27161 22486
rect 27195 22458 27232 22486
rect 27266 22458 27302 22486
rect 27336 22458 27372 22486
rect 27406 22458 27442 22486
rect 27476 22458 27512 22486
rect 26842 22452 26877 22458
rect 26916 22452 26948 22458
rect 26990 22452 27019 22458
rect 27064 22452 27090 22458
rect 27138 22452 27161 22458
rect 27212 22452 27232 22458
rect 27286 22452 27302 22458
rect 27360 22452 27372 22458
rect 27434 22452 27442 22458
rect 27508 22452 27512 22458
rect 27546 22458 27582 22486
rect 27546 22452 27548 22458
rect 26275 22424 26434 22452
rect 26468 22424 26509 22452
rect 26543 22424 26584 22452
rect 26618 22424 26659 22452
rect 26693 22424 26734 22452
rect 26768 22424 26808 22452
rect 26842 22424 26882 22452
rect 26916 22424 26956 22452
rect 26990 22424 27030 22452
rect 27064 22424 27104 22452
rect 27138 22424 27178 22452
rect 27212 22424 27252 22452
rect 27286 22424 27326 22452
rect 27360 22424 27400 22452
rect 27434 22424 27474 22452
rect 27508 22424 27548 22452
rect 27616 22458 27652 22486
rect 27686 22458 27722 22486
rect 27756 22458 27792 22486
rect 27826 22458 27862 22486
rect 27896 22458 27932 22486
rect 27616 22452 27622 22458
rect 27686 22452 27696 22458
rect 27756 22452 27770 22458
rect 27826 22452 27844 22458
rect 27896 22452 27918 22458
rect 27966 22452 28029 22486
rect 27582 22424 27622 22452
rect 27656 22424 27696 22452
rect 27730 22424 27770 22452
rect 27804 22424 27844 22452
rect 27878 22424 27918 22452
rect 27952 22424 28029 22452
rect 26275 22412 28029 22424
rect 26275 22378 26309 22412
rect 26343 22378 26380 22412
rect 26414 22386 26451 22412
rect 26485 22386 26522 22412
rect 26556 22386 26593 22412
rect 26627 22386 26664 22412
rect 26698 22386 26735 22412
rect 26414 22378 26434 22386
rect 26485 22378 26509 22386
rect 26556 22378 26584 22386
rect 26627 22378 26659 22386
rect 26698 22378 26734 22386
rect 26769 22378 26806 22412
rect 26840 22386 26877 22412
rect 26911 22386 26948 22412
rect 26982 22386 27019 22412
rect 27053 22386 27090 22412
rect 27124 22386 27161 22412
rect 27195 22386 27232 22412
rect 27266 22386 27302 22412
rect 27336 22386 27372 22412
rect 27406 22386 27442 22412
rect 27476 22386 27512 22412
rect 26842 22378 26877 22386
rect 26916 22378 26948 22386
rect 26990 22378 27019 22386
rect 27064 22378 27090 22386
rect 27138 22378 27161 22386
rect 27212 22378 27232 22386
rect 27286 22378 27302 22386
rect 27360 22378 27372 22386
rect 27434 22378 27442 22386
rect 27508 22378 27512 22386
rect 27546 22386 27582 22412
rect 27546 22378 27548 22386
rect 26275 22352 26434 22378
rect 26468 22352 26509 22378
rect 26543 22352 26584 22378
rect 26618 22352 26659 22378
rect 26693 22352 26734 22378
rect 26768 22352 26808 22378
rect 26842 22352 26882 22378
rect 26916 22352 26956 22378
rect 26990 22352 27030 22378
rect 27064 22352 27104 22378
rect 27138 22352 27178 22378
rect 27212 22352 27252 22378
rect 27286 22352 27326 22378
rect 27360 22352 27400 22378
rect 27434 22352 27474 22378
rect 27508 22352 27548 22378
rect 27616 22386 27652 22412
rect 27686 22386 27722 22412
rect 27756 22386 27792 22412
rect 27826 22386 27862 22412
rect 27896 22386 27932 22412
rect 27616 22378 27622 22386
rect 27686 22378 27696 22386
rect 27756 22378 27770 22386
rect 27826 22378 27844 22386
rect 27896 22378 27918 22386
rect 27966 22378 28029 22412
rect 27582 22352 27622 22378
rect 27656 22352 27696 22378
rect 27730 22352 27770 22378
rect 27804 22352 27844 22378
rect 27878 22352 27918 22378
rect 27952 22352 28029 22378
rect 26275 22338 28029 22352
rect 26275 22304 26309 22338
rect 26343 22304 26380 22338
rect 26414 22314 26451 22338
rect 26485 22314 26522 22338
rect 26556 22314 26593 22338
rect 26627 22314 26664 22338
rect 26698 22314 26735 22338
rect 26414 22304 26434 22314
rect 26485 22304 26509 22314
rect 26556 22304 26584 22314
rect 26627 22304 26659 22314
rect 26698 22304 26734 22314
rect 26769 22304 26806 22338
rect 26840 22314 26877 22338
rect 26911 22314 26948 22338
rect 26982 22314 27019 22338
rect 27053 22314 27090 22338
rect 27124 22314 27161 22338
rect 27195 22314 27232 22338
rect 27266 22314 27302 22338
rect 27336 22314 27372 22338
rect 27406 22314 27442 22338
rect 27476 22314 27512 22338
rect 26842 22304 26877 22314
rect 26916 22304 26948 22314
rect 26990 22304 27019 22314
rect 27064 22304 27090 22314
rect 27138 22304 27161 22314
rect 27212 22304 27232 22314
rect 27286 22304 27302 22314
rect 27360 22304 27372 22314
rect 27434 22304 27442 22314
rect 27508 22304 27512 22314
rect 27546 22314 27582 22338
rect 27546 22304 27548 22314
rect 26275 22280 26434 22304
rect 26468 22280 26509 22304
rect 26543 22280 26584 22304
rect 26618 22280 26659 22304
rect 26693 22280 26734 22304
rect 26768 22280 26808 22304
rect 26842 22280 26882 22304
rect 26916 22280 26956 22304
rect 26990 22280 27030 22304
rect 27064 22280 27104 22304
rect 27138 22280 27178 22304
rect 27212 22280 27252 22304
rect 27286 22280 27326 22304
rect 27360 22280 27400 22304
rect 27434 22280 27474 22304
rect 27508 22280 27548 22304
rect 27616 22314 27652 22338
rect 27686 22314 27722 22338
rect 27756 22314 27792 22338
rect 27826 22314 27862 22338
rect 27896 22314 27932 22338
rect 27616 22304 27622 22314
rect 27686 22304 27696 22314
rect 27756 22304 27770 22314
rect 27826 22304 27844 22314
rect 27896 22304 27918 22314
rect 27966 22304 28029 22338
rect 27582 22280 27622 22304
rect 27656 22280 27696 22304
rect 27730 22280 27770 22304
rect 27804 22280 27844 22304
rect 27878 22280 27918 22304
rect 27952 22280 28029 22304
rect 26275 22264 28029 22280
rect 26275 22230 26309 22264
rect 26343 22230 26380 22264
rect 26414 22242 26451 22264
rect 26485 22242 26522 22264
rect 26556 22242 26593 22264
rect 26627 22242 26664 22264
rect 26698 22242 26735 22264
rect 26414 22230 26434 22242
rect 26485 22230 26509 22242
rect 26556 22230 26584 22242
rect 26627 22230 26659 22242
rect 26698 22230 26734 22242
rect 26769 22230 26806 22264
rect 26840 22242 26877 22264
rect 26911 22242 26948 22264
rect 26982 22242 27019 22264
rect 27053 22242 27090 22264
rect 27124 22242 27161 22264
rect 27195 22242 27232 22264
rect 27266 22242 27302 22264
rect 27336 22242 27372 22264
rect 27406 22242 27442 22264
rect 27476 22242 27512 22264
rect 26842 22230 26877 22242
rect 26916 22230 26948 22242
rect 26990 22230 27019 22242
rect 27064 22230 27090 22242
rect 27138 22230 27161 22242
rect 27212 22230 27232 22242
rect 27286 22230 27302 22242
rect 27360 22230 27372 22242
rect 27434 22230 27442 22242
rect 27508 22230 27512 22242
rect 27546 22242 27582 22264
rect 27546 22230 27548 22242
rect 26275 22208 26434 22230
rect 26468 22208 26509 22230
rect 26543 22208 26584 22230
rect 26618 22208 26659 22230
rect 26693 22208 26734 22230
rect 26768 22208 26808 22230
rect 26842 22208 26882 22230
rect 26916 22208 26956 22230
rect 26990 22208 27030 22230
rect 27064 22208 27104 22230
rect 27138 22208 27178 22230
rect 27212 22208 27252 22230
rect 27286 22208 27326 22230
rect 27360 22208 27400 22230
rect 27434 22208 27474 22230
rect 27508 22208 27548 22230
rect 27616 22242 27652 22264
rect 27686 22242 27722 22264
rect 27756 22242 27792 22264
rect 27826 22242 27862 22264
rect 27896 22242 27932 22264
rect 27616 22230 27622 22242
rect 27686 22230 27696 22242
rect 27756 22230 27770 22242
rect 27826 22230 27844 22242
rect 27896 22230 27918 22242
rect 27966 22230 28029 22264
rect 27582 22208 27622 22230
rect 27656 22208 27696 22230
rect 27730 22208 27770 22230
rect 27804 22208 27844 22230
rect 27878 22208 27918 22230
rect 27952 22208 28029 22230
rect 26275 22190 28029 22208
rect 26275 22156 26309 22190
rect 26343 22156 26380 22190
rect 26414 22170 26451 22190
rect 26485 22170 26522 22190
rect 26556 22170 26593 22190
rect 26627 22170 26664 22190
rect 26698 22170 26735 22190
rect 26414 22156 26434 22170
rect 26485 22156 26509 22170
rect 26556 22156 26584 22170
rect 26627 22156 26659 22170
rect 26698 22156 26734 22170
rect 26769 22156 26806 22190
rect 26840 22170 26877 22190
rect 26911 22170 26948 22190
rect 26982 22170 27019 22190
rect 27053 22170 27090 22190
rect 27124 22170 27161 22190
rect 27195 22170 27232 22190
rect 27266 22170 27302 22190
rect 27336 22170 27372 22190
rect 27406 22170 27442 22190
rect 27476 22170 27512 22190
rect 26842 22156 26877 22170
rect 26916 22156 26948 22170
rect 26990 22156 27019 22170
rect 27064 22156 27090 22170
rect 27138 22156 27161 22170
rect 27212 22156 27232 22170
rect 27286 22156 27302 22170
rect 27360 22156 27372 22170
rect 27434 22156 27442 22170
rect 27508 22156 27512 22170
rect 27546 22170 27582 22190
rect 27546 22156 27548 22170
rect 26275 22136 26434 22156
rect 26468 22136 26509 22156
rect 26543 22136 26584 22156
rect 26618 22136 26659 22156
rect 26693 22136 26734 22156
rect 26768 22136 26808 22156
rect 26842 22136 26882 22156
rect 26916 22136 26956 22156
rect 26990 22136 27030 22156
rect 27064 22136 27104 22156
rect 27138 22136 27178 22156
rect 27212 22136 27252 22156
rect 27286 22136 27326 22156
rect 27360 22136 27400 22156
rect 27434 22136 27474 22156
rect 27508 22136 27548 22156
rect 27616 22170 27652 22190
rect 27686 22170 27722 22190
rect 27756 22170 27792 22190
rect 27826 22170 27862 22190
rect 27896 22170 27932 22190
rect 27616 22156 27622 22170
rect 27686 22156 27696 22170
rect 27756 22156 27770 22170
rect 27826 22156 27844 22170
rect 27896 22156 27918 22170
rect 27966 22156 28029 22190
rect 27582 22136 27622 22156
rect 27656 22136 27696 22156
rect 27730 22136 27770 22156
rect 27804 22136 27844 22156
rect 27878 22136 27918 22156
rect 27952 22136 28029 22156
rect 26275 22116 28029 22136
rect 26275 22082 26309 22116
rect 26343 22082 26380 22116
rect 26414 22082 26451 22116
rect 26485 22082 26522 22116
rect 26556 22082 26593 22116
rect 26627 22082 26664 22116
rect 26698 22082 26735 22116
rect 26769 22082 26806 22116
rect 26840 22082 26877 22116
rect 26911 22082 26948 22116
rect 26982 22082 27019 22116
rect 27053 22082 27090 22116
rect 27124 22082 27161 22116
rect 27195 22082 27232 22116
rect 27266 22082 27302 22116
rect 27336 22082 27372 22116
rect 27406 22082 27442 22116
rect 27476 22082 27512 22116
rect 27546 22082 27582 22116
rect 27616 22082 27652 22116
rect 27686 22082 27722 22116
rect 27756 22082 27792 22116
rect 27826 22082 27862 22116
rect 27896 22082 27932 22116
rect 27966 22082 28029 22116
rect 26275 22080 28029 22082
rect 27028 20830 27113 20846
rect 27012 20796 27113 20830
rect 27046 20762 27113 20796
rect 27012 20728 27113 20762
rect 27046 20694 27113 20728
rect 27012 20660 27113 20694
rect 27046 20626 27113 20660
rect 27012 20592 27113 20626
rect 27046 20558 27113 20592
rect 27012 20524 27113 20558
rect 27046 20490 27113 20524
rect 27012 20456 27113 20490
rect 27046 20422 27113 20456
rect 27012 20388 27113 20422
rect 27046 20354 27113 20388
rect 27012 20320 27113 20354
rect 27046 20286 27113 20320
rect 27012 20252 27113 20286
rect 27046 20218 27113 20252
rect 27012 20184 27113 20218
rect 27046 20150 27113 20184
rect 27012 20116 27113 20150
rect 27046 20082 27113 20116
rect 27012 20048 27113 20082
rect 27046 20014 27113 20048
rect 27012 19980 27113 20014
rect 27046 19946 27113 19980
rect 27012 19912 27113 19946
rect 27046 19878 27113 19912
rect 27012 19844 27113 19878
rect 27046 19810 27113 19844
rect 27012 19776 27113 19810
rect 27046 19742 27113 19776
rect 27012 19708 27113 19742
rect 27046 19674 27113 19708
rect 27012 19640 27113 19674
rect 27046 19606 27113 19640
rect 27012 19572 27113 19606
rect 27046 19538 27113 19572
rect 27012 19504 27113 19538
rect 27046 19470 27113 19504
rect 27012 19436 27113 19470
rect 27046 19402 27113 19436
rect 27012 19368 27113 19402
rect 27046 19334 27113 19368
rect 27012 19300 27113 19334
rect 27046 19266 27113 19300
rect 27012 19232 27113 19266
rect 24129 19201 24639 19225
rect 24129 17704 24639 17739
rect 24163 17670 24197 17704
rect 24231 17670 24265 17704
rect 24299 17670 24333 17704
rect 24367 17670 24401 17704
rect 24435 17670 24469 17704
rect 24503 17670 24537 17704
rect 24571 17670 24605 17704
rect 24129 17635 24639 17670
rect 24163 17601 24197 17635
rect 24231 17601 24265 17635
rect 24299 17601 24333 17635
rect 24367 17601 24401 17635
rect 24435 17601 24469 17635
rect 24503 17601 24537 17635
rect 24571 17601 24605 17635
rect 24129 17566 24639 17601
rect 24163 17532 24197 17566
rect 24231 17532 24265 17566
rect 24299 17532 24333 17566
rect 24367 17532 24401 17566
rect 24435 17532 24469 17566
rect 24503 17532 24537 17566
rect 24571 17532 24605 17566
rect 24129 17497 24639 17532
rect 24163 17463 24197 17497
rect 24231 17463 24265 17497
rect 24299 17463 24333 17497
rect 24367 17463 24401 17497
rect 24435 17463 24469 17497
rect 24503 17463 24537 17497
rect 24571 17463 24605 17497
rect 24129 17428 24639 17463
rect 24163 17394 24197 17428
rect 24231 17394 24265 17428
rect 24299 17394 24333 17428
rect 24367 17394 24401 17428
rect 24435 17394 24469 17428
rect 24503 17394 24537 17428
rect 24571 17394 24605 17428
rect 24129 17359 24639 17394
rect 24163 17325 24197 17359
rect 24231 17325 24265 17359
rect 24299 17325 24333 17359
rect 24367 17325 24401 17359
rect 24435 17325 24469 17359
rect 24503 17325 24537 17359
rect 24571 17325 24605 17359
rect 24129 17290 24639 17325
rect 24163 17256 24197 17290
rect 24231 17256 24265 17290
rect 24299 17256 24333 17290
rect 24367 17256 24401 17290
rect 24435 17256 24469 17290
rect 24503 17256 24537 17290
rect 24571 17256 24605 17290
rect 24129 17221 24639 17256
rect 24163 17187 24197 17221
rect 24231 17187 24265 17221
rect 24299 17187 24333 17221
rect 24367 17187 24401 17221
rect 24435 17187 24469 17221
rect 24503 17187 24537 17221
rect 24571 17187 24605 17221
rect 24129 17152 24639 17187
rect 24163 17118 24197 17152
rect 24231 17118 24265 17152
rect 24299 17118 24333 17152
rect 24367 17118 24401 17152
rect 24435 17118 24469 17152
rect 24503 17118 24537 17152
rect 24571 17118 24605 17152
rect 24129 17083 24639 17118
rect 24163 17049 24197 17083
rect 24231 17049 24265 17083
rect 24299 17049 24333 17083
rect 24367 17049 24401 17083
rect 24435 17049 24469 17083
rect 24503 17049 24537 17083
rect 24571 17049 24605 17083
rect 24129 17014 24639 17049
rect 24163 16980 24197 17014
rect 24231 16980 24265 17014
rect 24299 16980 24333 17014
rect 24367 16980 24401 17014
rect 24435 16980 24469 17014
rect 24503 16980 24537 17014
rect 24571 16980 24605 17014
rect 24129 16945 24639 16980
rect 24163 16911 24197 16945
rect 24231 16911 24265 16945
rect 24299 16911 24333 16945
rect 24367 16911 24401 16945
rect 24435 16911 24469 16945
rect 24503 16911 24537 16945
rect 24571 16911 24605 16945
rect 24129 16876 24639 16911
rect 24163 16842 24197 16876
rect 24231 16842 24265 16876
rect 24299 16842 24333 16876
rect 24367 16842 24401 16876
rect 24435 16842 24469 16876
rect 24503 16842 24537 16876
rect 24571 16842 24605 16876
rect 24129 16807 24639 16842
rect 24163 16773 24197 16807
rect 24231 16773 24265 16807
rect 24299 16773 24333 16807
rect 24367 16773 24401 16807
rect 24435 16773 24469 16807
rect 24503 16773 24537 16807
rect 24571 16773 24605 16807
rect 24129 16738 24639 16773
rect 24163 16704 24197 16738
rect 24231 16704 24265 16738
rect 24299 16704 24333 16738
rect 24367 16704 24401 16738
rect 24435 16704 24469 16738
rect 24503 16704 24537 16738
rect 24571 16704 24605 16738
rect 24129 16669 24639 16704
rect 24163 16635 24197 16669
rect 24231 16635 24265 16669
rect 24299 16635 24333 16669
rect 24367 16635 24401 16669
rect 24435 16635 24469 16669
rect 24503 16635 24537 16669
rect 24571 16635 24605 16669
rect 24129 16600 24639 16635
rect 24163 16566 24197 16600
rect 24231 16566 24265 16600
rect 24299 16566 24333 16600
rect 24367 16566 24401 16600
rect 24435 16566 24469 16600
rect 24503 16566 24537 16600
rect 24571 16566 24605 16600
rect 24129 16531 24639 16566
rect 24163 16497 24197 16531
rect 24231 16497 24265 16531
rect 24299 16497 24333 16531
rect 24367 16497 24401 16531
rect 24435 16497 24469 16531
rect 24503 16497 24537 16531
rect 24571 16497 24605 16531
rect 24129 16462 24639 16497
rect 24163 16428 24197 16462
rect 24231 16428 24265 16462
rect 24299 16428 24333 16462
rect 24367 16428 24401 16462
rect 24435 16428 24469 16462
rect 24503 16428 24537 16462
rect 24571 16428 24605 16462
rect 24129 16404 24639 16428
rect 24145 16338 24639 16404
rect 27046 19198 27113 19232
rect 27012 19164 27113 19198
rect 27046 19130 27113 19164
rect 27012 19096 27113 19130
rect 27046 19062 27113 19096
rect 27012 19028 27113 19062
rect 27046 18994 27113 19028
rect 27012 18960 27113 18994
rect 27046 18926 27113 18960
rect 27012 18892 27113 18926
rect 27046 18858 27113 18892
rect 27012 18824 27113 18858
rect 27046 18790 27113 18824
rect 27012 18756 27113 18790
rect 27046 18722 27113 18756
rect 27012 18688 27113 18722
rect 27046 18654 27113 18688
rect 27012 18620 27113 18654
rect 27046 18586 27113 18620
rect 27012 18552 27113 18586
rect 27046 18518 27113 18552
rect 27012 18484 27113 18518
rect 27046 18450 27113 18484
rect 27012 18416 27113 18450
rect 27046 18382 27113 18416
rect 27012 18348 27113 18382
rect 27046 18314 27113 18348
rect 27012 18280 27113 18314
rect 27046 18246 27113 18280
rect 27012 18212 27113 18246
rect 27046 18178 27113 18212
rect 27012 18144 27113 18178
rect 27046 18110 27113 18144
rect 27012 18076 27113 18110
rect 27046 18042 27113 18076
rect 27012 18008 27113 18042
rect 27046 17974 27113 18008
rect 27012 17940 27113 17974
rect 27046 17906 27113 17940
rect 27012 17872 27113 17906
rect 27046 17838 27113 17872
rect 27012 17804 27113 17838
rect 27046 17770 27113 17804
rect 27012 17736 27113 17770
rect 27046 17702 27113 17736
rect 27012 17668 27113 17702
rect 27046 17634 27113 17668
rect 27012 17600 27113 17634
rect 27046 17566 27113 17600
rect 27012 17532 27113 17566
rect 27046 17498 27113 17532
rect 27012 17464 27113 17498
rect 27046 17430 27113 17464
rect 27012 17396 27113 17430
rect 27046 17362 27113 17396
rect 27012 17328 27113 17362
rect 27046 17294 27113 17328
rect 27012 17259 27113 17294
rect 27046 17225 27113 17259
rect 27012 17190 27113 17225
rect 27046 17156 27113 17190
rect 27012 17121 27113 17156
rect 27046 17087 27113 17121
rect 27012 17052 27113 17087
rect 27046 17018 27113 17052
rect 27012 16983 27113 17018
rect 27046 16949 27113 16983
rect 27012 16914 27113 16949
rect 27046 16880 27113 16914
rect 27012 16845 27113 16880
rect 27046 16811 27113 16845
rect 27012 16776 27113 16811
rect 27046 16742 27113 16776
rect 27012 16707 27113 16742
rect 27046 16673 27113 16707
rect 27012 16638 27113 16673
rect 27046 16604 27113 16638
rect 27012 16569 27113 16604
rect 27046 16535 27113 16569
rect 27012 16500 27113 16535
rect 27046 16466 27113 16500
rect 27012 16431 27113 16466
rect 27046 16397 27113 16431
rect 27012 16362 27113 16397
rect 27046 16328 27113 16362
rect 27012 16293 27113 16328
rect 27046 16259 27113 16293
rect 27012 16224 27113 16259
rect 27046 16190 27113 16224
rect 27012 16155 27113 16190
rect 27046 16121 27113 16155
rect 27012 16086 27113 16121
rect 27046 16052 27113 16086
rect 27012 16017 27113 16052
rect 27046 15983 27113 16017
rect 27012 15948 27113 15983
rect 27046 15914 27113 15948
rect 27012 15879 27113 15914
rect 27046 15845 27113 15879
rect 27012 15810 27113 15845
rect 27046 15776 27113 15810
rect 27012 15741 27113 15776
rect 27046 15707 27113 15741
rect 27012 15672 27113 15707
rect 27046 15638 27113 15672
rect 27012 15603 27113 15638
rect 27046 15569 27113 15603
rect 27012 15534 27113 15569
rect 27046 15500 27113 15534
rect 27012 15465 27113 15500
rect 27046 15431 27113 15465
rect 27012 15396 27113 15431
rect 27046 15362 27113 15396
rect 27012 15327 27113 15362
rect 27046 15293 27113 15327
rect 27012 15258 27113 15293
rect 27046 15224 27113 15258
rect 27012 15189 27113 15224
rect 27046 15155 27113 15189
rect 27012 15120 27113 15155
rect 27046 15086 27113 15120
rect 27012 15051 27113 15086
rect 27046 15017 27113 15051
rect 27012 14983 27113 15017
rect 27028 14978 27113 14983
rect 13900 11875 13964 11993
rect 25925 11489 26329 11785
rect 16827 9560 16903 9594
rect 16937 9560 16976 9594
rect 17010 9560 17049 9594
rect 17083 9560 17122 9594
rect 17156 9560 17195 9594
rect 17229 9560 17267 9594
rect 17301 9560 17339 9594
rect 17373 9560 17411 9594
rect 17445 9560 17483 9594
rect 17517 9560 17555 9594
rect 17589 9560 17613 9594
rect 2320 4060 4514 4151
rect 2320 4058 3350 4060
rect 2320 4024 2344 4058
rect 2378 4024 2415 4058
rect 2449 4024 2486 4058
rect 2520 4024 2557 4058
rect 2591 4024 2628 4058
rect 2662 4024 2698 4058
rect 2732 4024 2768 4058
rect 2802 4024 2838 4058
rect 2872 4024 2908 4058
rect 2942 4024 2978 4058
rect 3012 4024 3048 4058
rect 3082 4024 3118 4058
rect 3152 4024 3188 4058
rect 3222 4024 3258 4058
rect 3292 4026 3350 4058
rect 3384 4026 3419 4060
rect 3453 4026 3488 4060
rect 3522 4026 3557 4060
rect 3591 4026 3626 4060
rect 3660 4026 3695 4060
rect 3729 4026 3764 4060
rect 3798 4026 3833 4060
rect 3867 4026 3902 4060
rect 3936 4026 3971 4060
rect 4005 4026 4040 4060
rect 4074 4026 4109 4060
rect 4143 4026 4178 4060
rect 4212 4026 4247 4060
rect 4281 4026 4316 4060
rect 4350 4026 4385 4060
rect 4419 4026 4454 4060
rect 4488 4026 4523 4060
rect 4557 4026 4592 4060
rect 4626 4026 4661 4060
rect 4695 4026 4730 4060
rect 4764 4026 4799 4060
rect 4833 4026 4868 4060
rect 4902 4026 4937 4060
rect 4971 4026 5006 4060
rect 5040 4026 5075 4060
rect 5109 4026 5144 4060
rect 5178 4026 5213 4060
rect 5247 4026 5282 4060
rect 5316 4026 5351 4060
rect 5385 4026 5420 4060
rect 5454 4026 5489 4060
rect 5523 4026 5558 4060
rect 5592 4026 5627 4060
rect 5661 4026 5696 4060
rect 5730 4026 5765 4060
rect 5799 4026 5834 4060
rect 5868 4026 5903 4060
rect 5937 4026 5972 4060
rect 6006 4026 6041 4060
rect 3292 4024 6041 4026
rect 2320 3992 6041 4024
rect 2320 3984 3350 3992
rect 2320 3950 2344 3984
rect 2378 3950 2415 3984
rect 2449 3950 2486 3984
rect 2520 3950 2557 3984
rect 2591 3950 2628 3984
rect 2662 3950 2698 3984
rect 2732 3950 2768 3984
rect 2802 3950 2838 3984
rect 2872 3950 2908 3984
rect 2942 3950 2978 3984
rect 3012 3950 3048 3984
rect 3082 3950 3118 3984
rect 3152 3950 3188 3984
rect 3222 3950 3258 3984
rect 3292 3958 3350 3984
rect 3384 3958 3419 3992
rect 3453 3958 3488 3992
rect 3522 3958 3557 3992
rect 3591 3958 3626 3992
rect 3660 3958 3695 3992
rect 3729 3958 3764 3992
rect 3798 3958 3833 3992
rect 3867 3958 3902 3992
rect 3936 3958 3971 3992
rect 4005 3958 4040 3992
rect 4074 3958 4109 3992
rect 4143 3958 4178 3992
rect 4212 3958 4247 3992
rect 4281 3958 4316 3992
rect 4350 3958 4385 3992
rect 4419 3958 4454 3992
rect 4488 3958 4523 3992
rect 4557 3958 4592 3992
rect 4626 3958 4661 3992
rect 4695 3958 4730 3992
rect 4764 3958 4799 3992
rect 4833 3958 4868 3992
rect 4902 3958 4937 3992
rect 4971 3958 5006 3992
rect 5040 3958 5075 3992
rect 5109 3958 5144 3992
rect 5178 3958 5213 3992
rect 5247 3958 5282 3992
rect 5316 3958 5351 3992
rect 5385 3958 5420 3992
rect 5454 3958 5489 3992
rect 5523 3958 5558 3992
rect 5592 3958 5627 3992
rect 5661 3958 5696 3992
rect 5730 3958 5765 3992
rect 5799 3958 5834 3992
rect 5868 3958 5903 3992
rect 5937 3958 5972 3992
rect 6006 3958 6041 3992
rect 3292 3950 6041 3958
rect 2320 3924 6041 3950
rect 2320 3910 3350 3924
rect 2320 3876 2344 3910
rect 2378 3876 2415 3910
rect 2449 3876 2486 3910
rect 2520 3876 2557 3910
rect 2591 3876 2628 3910
rect 2662 3876 2698 3910
rect 2732 3876 2768 3910
rect 2802 3876 2838 3910
rect 2872 3876 2908 3910
rect 2942 3876 2978 3910
rect 3012 3876 3048 3910
rect 3082 3876 3118 3910
rect 3152 3876 3188 3910
rect 3222 3876 3258 3910
rect 3292 3890 3350 3910
rect 3384 3890 3419 3924
rect 3453 3890 3488 3924
rect 3522 3890 3557 3924
rect 3591 3890 3626 3924
rect 3660 3890 3695 3924
rect 3729 3890 3764 3924
rect 3798 3890 3833 3924
rect 3867 3890 3902 3924
rect 3936 3890 3971 3924
rect 4005 3890 4040 3924
rect 4074 3890 4109 3924
rect 4143 3890 4178 3924
rect 4212 3890 4247 3924
rect 4281 3890 4316 3924
rect 4350 3890 4385 3924
rect 4419 3890 4454 3924
rect 4488 3890 4523 3924
rect 4557 3890 4592 3924
rect 4626 3890 4661 3924
rect 4695 3890 4730 3924
rect 4764 3890 4799 3924
rect 4833 3890 4868 3924
rect 4902 3890 4937 3924
rect 4971 3890 5006 3924
rect 5040 3890 5075 3924
rect 5109 3890 5144 3924
rect 5178 3890 5213 3924
rect 5247 3890 5282 3924
rect 5316 3890 5351 3924
rect 5385 3890 5420 3924
rect 5454 3890 5489 3924
rect 5523 3890 5558 3924
rect 5592 3890 5627 3924
rect 5661 3890 5696 3924
rect 5730 3890 5765 3924
rect 5799 3890 5834 3924
rect 5868 3890 5903 3924
rect 5937 3890 5972 3924
rect 6006 3890 6041 3924
rect 3292 3876 6041 3890
rect 2320 3856 6041 3876
rect 2320 3836 3350 3856
rect 2320 3802 2344 3836
rect 2378 3802 2415 3836
rect 2449 3802 2486 3836
rect 2520 3802 2557 3836
rect 2591 3802 2628 3836
rect 2662 3802 2698 3836
rect 2732 3802 2768 3836
rect 2802 3831 2838 3836
rect 2802 3802 2832 3831
rect 2872 3802 2908 3836
rect 2942 3831 2978 3836
rect 3012 3831 3048 3836
rect 3082 3831 3118 3836
rect 2949 3802 2978 3831
rect 3032 3802 3048 3831
rect 3115 3802 3118 3831
rect 3152 3831 3188 3836
rect 3152 3802 3164 3831
rect 3222 3802 3258 3836
rect 3292 3822 3350 3836
rect 3384 3822 3419 3856
rect 3453 3822 3488 3856
rect 3522 3822 3557 3856
rect 3591 3822 3626 3856
rect 3660 3822 3695 3856
rect 3729 3822 3764 3856
rect 3798 3822 3833 3856
rect 3867 3822 3902 3856
rect 3936 3822 3971 3856
rect 4005 3822 4040 3856
rect 4074 3822 4109 3856
rect 4143 3822 4178 3856
rect 4212 3822 4247 3856
rect 4281 3822 4316 3856
rect 4350 3822 4385 3856
rect 4419 3822 4454 3856
rect 4488 3822 4523 3856
rect 4557 3822 4592 3856
rect 4626 3822 4661 3856
rect 4695 3822 4730 3856
rect 4764 3822 4799 3856
rect 4833 3822 4868 3856
rect 4902 3822 4937 3856
rect 4971 3822 5006 3856
rect 5040 3822 5075 3856
rect 5109 3822 5144 3856
rect 5178 3822 5213 3856
rect 5247 3822 5282 3856
rect 5316 3822 5351 3856
rect 5385 3822 5420 3856
rect 5454 3822 5489 3856
rect 5523 3822 5558 3856
rect 5592 3822 5627 3856
rect 5661 3822 5696 3856
rect 5730 3822 5765 3856
rect 5799 3822 5834 3856
rect 5868 3822 5903 3856
rect 5937 3822 5972 3856
rect 6006 3822 6041 3856
rect 3292 3802 6041 3822
rect 2320 3797 2832 3802
rect 2866 3797 2915 3802
rect 2949 3797 2998 3802
rect 3032 3797 3081 3802
rect 3115 3797 3164 3802
rect 3198 3797 6041 3802
rect 2320 3788 6041 3797
rect 2320 3779 3350 3788
rect 2320 3762 2532 3779
rect 2566 3762 2624 3779
rect 2658 3762 2716 3779
rect 2750 3762 3350 3779
rect 2320 3728 2344 3762
rect 2378 3728 2415 3762
rect 2449 3728 2486 3762
rect 2520 3745 2532 3762
rect 2591 3745 2624 3762
rect 2520 3728 2557 3745
rect 2591 3728 2628 3745
rect 2662 3728 2698 3762
rect 2750 3745 2768 3762
rect 2732 3728 2768 3745
rect 2802 3728 2838 3762
rect 2872 3728 2908 3762
rect 2942 3728 2978 3762
rect 3012 3728 3048 3762
rect 3082 3728 3118 3762
rect 3152 3728 3188 3762
rect 3222 3728 3258 3762
rect 3292 3754 3350 3762
rect 3384 3754 3419 3788
rect 3453 3754 3488 3788
rect 3522 3754 3557 3788
rect 3591 3754 3626 3788
rect 3660 3754 3695 3788
rect 3729 3754 3764 3788
rect 3798 3754 3833 3788
rect 3867 3754 3902 3788
rect 3936 3754 3971 3788
rect 4005 3754 4040 3788
rect 4074 3754 4109 3788
rect 4143 3754 4178 3788
rect 4212 3754 4247 3788
rect 4281 3754 4316 3788
rect 4350 3754 4385 3788
rect 4419 3754 4454 3788
rect 4488 3754 4523 3788
rect 4557 3754 4592 3788
rect 4626 3754 4661 3788
rect 4695 3754 4730 3788
rect 4764 3754 4799 3788
rect 4833 3754 4868 3788
rect 4902 3754 4937 3788
rect 4971 3754 5006 3788
rect 5040 3754 5075 3788
rect 5109 3754 5144 3788
rect 5178 3754 5213 3788
rect 5247 3754 5282 3788
rect 5316 3754 5351 3788
rect 5385 3754 5420 3788
rect 5454 3754 5489 3788
rect 5523 3754 5558 3788
rect 5592 3754 5627 3788
rect 5661 3754 5696 3788
rect 5730 3754 5765 3788
rect 5799 3754 5834 3788
rect 5868 3754 5903 3788
rect 5937 3754 5972 3788
rect 6006 3754 6041 3788
rect 6415 4058 28000 4060
rect 6415 4024 6473 4058
rect 6507 4024 6542 4058
rect 6576 4024 6611 4058
rect 6645 4024 6680 4058
rect 6714 4024 6749 4058
rect 6783 4024 6818 4058
rect 6852 4024 6887 4058
rect 6921 4024 6956 4058
rect 6990 4024 7025 4058
rect 7059 4024 7094 4058
rect 7128 4024 7163 4058
rect 7197 4024 7232 4058
rect 7266 4024 7301 4058
rect 7335 4024 7370 4058
rect 7404 4024 7439 4058
rect 7473 4024 7508 4058
rect 7542 4024 7577 4058
rect 7611 4024 7646 4058
rect 7680 4024 7715 4058
rect 7749 4024 7784 4058
rect 7818 4024 7853 4058
rect 7887 4024 7922 4058
rect 7956 4024 7991 4058
rect 8025 4024 8060 4058
rect 8094 4024 8129 4058
rect 8163 4024 8198 4058
rect 8232 4024 8267 4058
rect 8301 4024 8336 4058
rect 8370 4024 8405 4058
rect 8439 4024 8474 4058
rect 8508 4024 8543 4058
rect 8577 4024 8612 4058
rect 8646 4024 8681 4058
rect 8715 4024 8750 4058
rect 8784 4024 8819 4058
rect 8853 4024 8888 4058
rect 8922 4024 8957 4058
rect 8991 4024 9026 4058
rect 9060 4024 9095 4058
rect 9129 4024 9164 4058
rect 9198 4024 9233 4058
rect 9267 4024 9302 4058
rect 9336 4024 9371 4058
rect 9405 4024 9440 4058
rect 9474 4024 9509 4058
rect 9543 4024 9578 4058
rect 9612 4024 9647 4058
rect 9681 4024 9716 4058
rect 9750 4024 9785 4058
rect 9819 4024 9854 4058
rect 9888 4024 9922 4058
rect 9956 4024 9990 4058
rect 10024 4024 10058 4058
rect 10092 4024 10126 4058
rect 10160 4024 10194 4058
rect 10228 4024 10262 4058
rect 10296 4024 10330 4058
rect 10364 4024 10398 4058
rect 10432 4024 10466 4058
rect 10500 4024 10534 4058
rect 10568 4024 10602 4058
rect 10636 4024 10670 4058
rect 10704 4024 10738 4058
rect 10772 4024 10806 4058
rect 10840 4024 10874 4058
rect 10908 4024 10942 4058
rect 10976 4024 11010 4058
rect 11044 4024 11078 4058
rect 11112 4024 11146 4058
rect 11180 4024 11214 4058
rect 11248 4024 11282 4058
rect 11316 4024 11350 4058
rect 11384 4024 11418 4058
rect 11452 4024 11486 4058
rect 11520 4024 11554 4058
rect 11588 4024 11622 4058
rect 11656 4024 11690 4058
rect 11724 4024 11758 4058
rect 11792 4024 11826 4058
rect 11860 4024 11894 4058
rect 11928 4024 11962 4058
rect 11996 4024 12030 4058
rect 12064 4024 12098 4058
rect 12132 4024 12166 4058
rect 12200 4024 12234 4058
rect 12268 4024 12302 4058
rect 12336 4024 12370 4058
rect 12404 4024 12438 4058
rect 12472 4024 12506 4058
rect 12540 4024 12574 4058
rect 12608 4024 12642 4058
rect 12676 4024 12710 4058
rect 12744 4024 12778 4058
rect 12812 4024 12846 4058
rect 12880 4024 12914 4058
rect 12948 4024 12982 4058
rect 13016 4024 13050 4058
rect 13084 4024 13118 4058
rect 13152 4024 13186 4058
rect 13220 4024 13254 4058
rect 13288 4024 13322 4058
rect 13356 4024 13390 4058
rect 13424 4024 13458 4058
rect 13492 4024 13526 4058
rect 13560 4024 13594 4058
rect 13628 4024 13662 4058
rect 13696 4024 13730 4058
rect 13764 4024 13798 4058
rect 13832 4024 13866 4058
rect 13900 4024 13934 4058
rect 13968 4024 14002 4058
rect 14036 4024 14070 4058
rect 14104 4024 14138 4058
rect 14172 4024 14206 4058
rect 14240 4024 14274 4058
rect 14308 4024 14342 4058
rect 14376 4024 14410 4058
rect 14444 4024 14478 4058
rect 14512 4024 14546 4058
rect 14580 4024 14614 4058
rect 14648 4024 14682 4058
rect 14716 4024 14750 4058
rect 14784 4024 14818 4058
rect 14852 4024 14886 4058
rect 14920 4024 14954 4058
rect 14988 4024 15022 4058
rect 15056 4024 15090 4058
rect 15124 4024 15158 4058
rect 15192 4024 15226 4058
rect 15260 4024 15294 4058
rect 15328 4024 15362 4058
rect 15396 4024 15430 4058
rect 15464 4024 15498 4058
rect 15532 4024 15566 4058
rect 15600 4024 15634 4058
rect 15668 4024 15702 4058
rect 15736 4024 15770 4058
rect 15804 4024 15838 4058
rect 15872 4024 15906 4058
rect 15940 4024 15974 4058
rect 16008 4024 16042 4058
rect 16076 4024 16110 4058
rect 16144 4024 16178 4058
rect 16212 4024 16246 4058
rect 16280 4024 16314 4058
rect 16348 4024 16382 4058
rect 16416 4024 16450 4058
rect 16484 4024 16518 4058
rect 16552 4024 16586 4058
rect 16620 4024 16654 4058
rect 16688 4024 16722 4058
rect 16756 4024 16790 4058
rect 16824 4024 16858 4058
rect 16892 4024 16926 4058
rect 16960 4024 16994 4058
rect 17028 4024 17062 4058
rect 17096 4024 17130 4058
rect 17164 4024 17198 4058
rect 17232 4024 17266 4058
rect 17300 4024 17334 4058
rect 17368 4024 17402 4058
rect 17436 4024 17470 4058
rect 17504 4024 17538 4058
rect 17572 4024 17606 4058
rect 17640 4024 17674 4058
rect 17708 4024 17742 4058
rect 17776 4024 17810 4058
rect 17844 4024 17878 4058
rect 17912 4024 17946 4058
rect 17980 4024 18014 4058
rect 18048 4024 18082 4058
rect 18116 4024 18150 4058
rect 18184 4024 18218 4058
rect 18252 4024 18286 4058
rect 18320 4024 18354 4058
rect 18388 4024 18422 4058
rect 18456 4024 18490 4058
rect 18524 4024 18558 4058
rect 18592 4024 18626 4058
rect 18660 4024 18694 4058
rect 18728 4024 18762 4058
rect 18796 4024 18830 4058
rect 18864 4024 18898 4058
rect 18932 4024 18966 4058
rect 19000 4024 19034 4058
rect 19068 4024 19102 4058
rect 19136 4024 19170 4058
rect 19204 4024 19238 4058
rect 19272 4024 19306 4058
rect 19340 4024 19374 4058
rect 19408 4024 19442 4058
rect 19476 4024 19510 4058
rect 19544 4024 19578 4058
rect 19612 4024 19646 4058
rect 19680 4024 19714 4058
rect 19748 4024 19782 4058
rect 19816 4024 19850 4058
rect 19884 4024 19918 4058
rect 19952 4024 19986 4058
rect 20020 4024 20054 4058
rect 20088 4024 20122 4058
rect 20156 4024 20190 4058
rect 20224 4024 20258 4058
rect 20292 4024 20326 4058
rect 20360 4024 20394 4058
rect 20428 4024 20462 4058
rect 20496 4024 20530 4058
rect 20564 4024 20598 4058
rect 20632 4024 20666 4058
rect 20700 4024 20734 4058
rect 20768 4024 20802 4058
rect 20836 4024 20870 4058
rect 20904 4024 20938 4058
rect 20972 4024 21006 4058
rect 21040 4024 21074 4058
rect 21108 4024 21142 4058
rect 21176 4024 21210 4058
rect 21244 4024 21278 4058
rect 21312 4024 21346 4058
rect 21380 4024 21414 4058
rect 21448 4024 21482 4058
rect 21516 4024 21550 4058
rect 21584 4024 21618 4058
rect 21652 4024 21686 4058
rect 21720 4024 21754 4058
rect 21788 4024 21822 4058
rect 21856 4024 21890 4058
rect 21924 4024 21958 4058
rect 21992 4024 22026 4058
rect 22060 4024 22094 4058
rect 22128 4024 22162 4058
rect 22196 4024 22230 4058
rect 22264 4024 22298 4058
rect 22332 4024 22366 4058
rect 22400 4024 22434 4058
rect 22468 4024 22502 4058
rect 22536 4024 22570 4058
rect 22604 4024 22638 4058
rect 22672 4024 22706 4058
rect 22740 4024 22774 4058
rect 22808 4024 22842 4058
rect 22876 4024 22910 4058
rect 22944 4024 22978 4058
rect 23012 4024 23046 4058
rect 23080 4024 23114 4058
rect 23148 4024 23182 4058
rect 23216 4024 23250 4058
rect 23284 4024 23318 4058
rect 23352 4024 23386 4058
rect 23420 4024 23454 4058
rect 23488 4024 23522 4058
rect 23556 4024 23590 4058
rect 23624 4024 23658 4058
rect 23692 4024 23726 4058
rect 23760 4024 23794 4058
rect 23828 4024 23862 4058
rect 23896 4024 23930 4058
rect 23964 4024 23998 4058
rect 24032 4024 24066 4058
rect 24100 4024 24134 4058
rect 24168 4024 24202 4058
rect 24236 4024 24270 4058
rect 24304 4024 24338 4058
rect 24372 4024 24406 4058
rect 24440 4024 24474 4058
rect 24508 4024 24542 4058
rect 24576 4024 24610 4058
rect 24644 4024 24678 4058
rect 24712 4024 24746 4058
rect 24780 4024 24814 4058
rect 24848 4024 24882 4058
rect 24916 4024 24950 4058
rect 24984 4024 25018 4058
rect 25052 4024 25086 4058
rect 25120 4024 25154 4058
rect 25188 4024 25222 4058
rect 25256 4024 25290 4058
rect 25324 4024 25358 4058
rect 25392 4024 25426 4058
rect 25460 4024 25494 4058
rect 25528 4024 25562 4058
rect 25596 4024 25630 4058
rect 25664 4024 25698 4058
rect 25732 4024 25766 4058
rect 25800 4024 25834 4058
rect 25868 4024 25902 4058
rect 25936 4024 25970 4058
rect 26004 4024 26038 4058
rect 26072 4024 26106 4058
rect 26140 4024 26174 4058
rect 26208 4024 26242 4058
rect 26276 4024 26310 4058
rect 26344 4024 26378 4058
rect 26412 4024 26446 4058
rect 26480 4024 26514 4058
rect 26548 4024 26582 4058
rect 26616 4024 26650 4058
rect 26684 4024 26718 4058
rect 26752 4024 26786 4058
rect 26820 4024 26854 4058
rect 26888 4024 26922 4058
rect 26956 4024 26990 4058
rect 27024 4024 27058 4058
rect 27092 4024 27126 4058
rect 27160 4024 27194 4058
rect 27228 4024 27262 4058
rect 27296 4024 27330 4058
rect 27364 4024 27398 4058
rect 27432 4024 27466 4058
rect 27500 4024 27534 4058
rect 27568 4024 27602 4058
rect 27636 4024 27670 4058
rect 27704 4024 27738 4058
rect 27772 4024 27806 4058
rect 27840 4024 27874 4058
rect 27908 4024 27942 4058
rect 27976 4024 28000 4058
rect 6415 3984 28000 4024
rect 6415 3950 6473 3984
rect 6507 3950 6542 3984
rect 6576 3950 6611 3984
rect 6645 3950 6680 3984
rect 6714 3950 6749 3984
rect 6783 3950 6818 3984
rect 6852 3950 6887 3984
rect 6921 3950 6956 3984
rect 6990 3950 7025 3984
rect 7059 3950 7094 3984
rect 7128 3950 7163 3984
rect 7197 3950 7232 3984
rect 7266 3950 7301 3984
rect 7335 3950 7370 3984
rect 7404 3950 7439 3984
rect 7473 3950 7508 3984
rect 7542 3950 7577 3984
rect 7611 3950 7646 3984
rect 7680 3950 7715 3984
rect 7749 3950 7784 3984
rect 7818 3950 7853 3984
rect 7887 3950 7922 3984
rect 7956 3950 7991 3984
rect 8025 3950 8060 3984
rect 8094 3950 8129 3984
rect 8163 3950 8198 3984
rect 8232 3950 8267 3984
rect 8301 3950 8336 3984
rect 8370 3950 8405 3984
rect 8439 3950 8474 3984
rect 8508 3950 8543 3984
rect 8577 3950 8612 3984
rect 8646 3950 8681 3984
rect 8715 3950 8750 3984
rect 8784 3950 8819 3984
rect 8853 3950 8888 3984
rect 8922 3950 8957 3984
rect 8991 3950 9026 3984
rect 9060 3950 9095 3984
rect 9129 3950 9164 3984
rect 9198 3950 9233 3984
rect 9267 3950 9302 3984
rect 9336 3950 9371 3984
rect 9405 3950 9440 3984
rect 9474 3950 9509 3984
rect 9543 3950 9578 3984
rect 9612 3950 9647 3984
rect 9681 3950 9716 3984
rect 9750 3950 9785 3984
rect 9819 3950 9854 3984
rect 9888 3950 9922 3984
rect 9956 3950 9990 3984
rect 10024 3950 10058 3984
rect 10092 3950 10126 3984
rect 10160 3950 10194 3984
rect 10228 3950 10262 3984
rect 10296 3950 10330 3984
rect 10364 3950 10398 3984
rect 10432 3950 10466 3984
rect 10500 3950 10534 3984
rect 10568 3950 10602 3984
rect 10636 3950 10670 3984
rect 10704 3950 10738 3984
rect 10772 3950 10806 3984
rect 10840 3950 10874 3984
rect 10908 3950 10942 3984
rect 10976 3950 11010 3984
rect 11044 3950 11078 3984
rect 11112 3950 11146 3984
rect 11180 3950 11214 3984
rect 11248 3950 11282 3984
rect 11316 3950 11350 3984
rect 11384 3950 11418 3984
rect 11452 3950 11486 3984
rect 11520 3950 11554 3984
rect 11588 3950 11622 3984
rect 11656 3950 11690 3984
rect 11724 3950 11758 3984
rect 11792 3950 11826 3984
rect 11860 3950 11894 3984
rect 11928 3950 11962 3984
rect 11996 3950 12030 3984
rect 12064 3950 12098 3984
rect 12132 3950 12166 3984
rect 12200 3950 12234 3984
rect 12268 3950 12302 3984
rect 12336 3950 12370 3984
rect 12404 3950 12438 3984
rect 12472 3950 12506 3984
rect 12540 3950 12574 3984
rect 12608 3950 12642 3984
rect 12676 3950 12710 3984
rect 12744 3950 12778 3984
rect 12812 3950 12846 3984
rect 12880 3950 12914 3984
rect 12948 3950 12982 3984
rect 13016 3950 13050 3984
rect 13084 3950 13118 3984
rect 13152 3950 13186 3984
rect 13220 3950 13254 3984
rect 13288 3950 13322 3984
rect 13356 3950 13390 3984
rect 13424 3950 13458 3984
rect 13492 3950 13526 3984
rect 13560 3950 13594 3984
rect 13628 3950 13662 3984
rect 13696 3950 13730 3984
rect 13764 3950 13798 3984
rect 13832 3950 13866 3984
rect 13900 3950 13934 3984
rect 13968 3950 14002 3984
rect 14036 3950 14070 3984
rect 14104 3950 14138 3984
rect 14172 3950 14206 3984
rect 14240 3950 14274 3984
rect 14308 3950 14342 3984
rect 14376 3950 14410 3984
rect 14444 3950 14478 3984
rect 14512 3950 14546 3984
rect 14580 3950 14614 3984
rect 14648 3950 14682 3984
rect 14716 3950 14750 3984
rect 14784 3950 14818 3984
rect 14852 3950 14886 3984
rect 14920 3950 14954 3984
rect 14988 3950 15022 3984
rect 15056 3950 15090 3984
rect 15124 3950 15158 3984
rect 15192 3950 15226 3984
rect 15260 3950 15294 3984
rect 15328 3950 15362 3984
rect 15396 3950 15430 3984
rect 15464 3950 15498 3984
rect 15532 3950 15566 3984
rect 15600 3950 15634 3984
rect 15668 3950 15702 3984
rect 15736 3950 15770 3984
rect 15804 3950 15838 3984
rect 15872 3950 15906 3984
rect 15940 3950 15974 3984
rect 16008 3950 16042 3984
rect 16076 3950 16110 3984
rect 16144 3950 16178 3984
rect 16212 3950 16246 3984
rect 16280 3950 16314 3984
rect 16348 3950 16382 3984
rect 16416 3950 16450 3984
rect 16484 3950 16518 3984
rect 16552 3950 16586 3984
rect 16620 3950 16654 3984
rect 16688 3950 16722 3984
rect 16756 3950 16790 3984
rect 16824 3950 16858 3984
rect 16892 3950 16926 3984
rect 16960 3950 16994 3984
rect 17028 3950 17062 3984
rect 17096 3950 17130 3984
rect 17164 3950 17198 3984
rect 17232 3950 17266 3984
rect 17300 3950 17334 3984
rect 17368 3950 17402 3984
rect 17436 3950 17470 3984
rect 17504 3950 17538 3984
rect 17572 3950 17606 3984
rect 17640 3950 17674 3984
rect 17708 3950 17742 3984
rect 17776 3950 17810 3984
rect 17844 3950 17878 3984
rect 17912 3950 17946 3984
rect 17980 3950 18014 3984
rect 18048 3950 18082 3984
rect 18116 3950 18150 3984
rect 18184 3950 18218 3984
rect 18252 3950 18286 3984
rect 18320 3950 18354 3984
rect 18388 3950 18422 3984
rect 18456 3950 18490 3984
rect 18524 3950 18558 3984
rect 18592 3950 18626 3984
rect 18660 3950 18694 3984
rect 18728 3950 18762 3984
rect 18796 3950 18830 3984
rect 18864 3950 18898 3984
rect 18932 3950 18966 3984
rect 19000 3950 19034 3984
rect 19068 3950 19102 3984
rect 19136 3950 19170 3984
rect 19204 3950 19238 3984
rect 19272 3950 19306 3984
rect 19340 3950 19374 3984
rect 19408 3950 19442 3984
rect 19476 3950 19510 3984
rect 19544 3950 19578 3984
rect 19612 3950 19646 3984
rect 19680 3950 19714 3984
rect 19748 3950 19782 3984
rect 19816 3950 19850 3984
rect 19884 3950 19918 3984
rect 19952 3950 19986 3984
rect 20020 3950 20054 3984
rect 20088 3950 20122 3984
rect 20156 3950 20190 3984
rect 20224 3950 20258 3984
rect 20292 3950 20326 3984
rect 20360 3950 20394 3984
rect 20428 3950 20462 3984
rect 20496 3950 20530 3984
rect 20564 3950 20598 3984
rect 20632 3950 20666 3984
rect 20700 3950 20734 3984
rect 20768 3950 20802 3984
rect 20836 3950 20870 3984
rect 20904 3950 20938 3984
rect 20972 3950 21006 3984
rect 21040 3950 21074 3984
rect 21108 3950 21142 3984
rect 21176 3950 21210 3984
rect 21244 3950 21278 3984
rect 21312 3950 21346 3984
rect 21380 3950 21414 3984
rect 21448 3950 21482 3984
rect 21516 3950 21550 3984
rect 21584 3950 21618 3984
rect 21652 3950 21686 3984
rect 21720 3950 21754 3984
rect 21788 3950 21822 3984
rect 21856 3950 21890 3984
rect 21924 3950 21958 3984
rect 21992 3950 22026 3984
rect 22060 3950 22094 3984
rect 22128 3950 22162 3984
rect 22196 3950 22230 3984
rect 22264 3950 22298 3984
rect 22332 3950 22366 3984
rect 22400 3950 22434 3984
rect 22468 3950 22502 3984
rect 22536 3950 22570 3984
rect 22604 3950 22638 3984
rect 22672 3950 22706 3984
rect 22740 3950 22774 3984
rect 22808 3950 22842 3984
rect 22876 3950 22910 3984
rect 22944 3950 22978 3984
rect 23012 3950 23046 3984
rect 23080 3950 23114 3984
rect 23148 3950 23182 3984
rect 23216 3950 23250 3984
rect 23284 3950 23318 3984
rect 23352 3950 23386 3984
rect 23420 3950 23454 3984
rect 23488 3950 23522 3984
rect 23556 3950 23590 3984
rect 23624 3950 23658 3984
rect 23692 3950 23726 3984
rect 23760 3950 23794 3984
rect 23828 3950 23862 3984
rect 23896 3950 23930 3984
rect 23964 3950 23998 3984
rect 24032 3950 24066 3984
rect 24100 3950 24134 3984
rect 24168 3950 24202 3984
rect 24236 3950 24270 3984
rect 24304 3950 24338 3984
rect 24372 3950 24406 3984
rect 24440 3950 24474 3984
rect 24508 3950 24542 3984
rect 24576 3950 24610 3984
rect 24644 3950 24678 3984
rect 24712 3950 24746 3984
rect 24780 3950 24814 3984
rect 24848 3950 24882 3984
rect 24916 3950 24950 3984
rect 24984 3950 25018 3984
rect 25052 3950 25086 3984
rect 25120 3950 25154 3984
rect 25188 3950 25222 3984
rect 25256 3950 25290 3984
rect 25324 3950 25358 3984
rect 25392 3950 25426 3984
rect 25460 3950 25494 3984
rect 25528 3950 25562 3984
rect 25596 3950 25630 3984
rect 25664 3950 25698 3984
rect 25732 3950 25766 3984
rect 25800 3950 25834 3984
rect 25868 3950 25902 3984
rect 25936 3950 25970 3984
rect 26004 3950 26038 3984
rect 26072 3950 26106 3984
rect 26140 3950 26174 3984
rect 26208 3950 26242 3984
rect 26276 3950 26310 3984
rect 26344 3950 26378 3984
rect 26412 3950 26446 3984
rect 26480 3950 26514 3984
rect 26548 3950 26582 3984
rect 26616 3950 26650 3984
rect 26684 3950 26718 3984
rect 26752 3950 26786 3984
rect 26820 3950 26854 3984
rect 26888 3950 26922 3984
rect 26956 3950 26990 3984
rect 27024 3950 27058 3984
rect 27092 3950 27126 3984
rect 27160 3950 27194 3984
rect 27228 3950 27262 3984
rect 27296 3950 27330 3984
rect 27364 3950 27398 3984
rect 27432 3950 27466 3984
rect 27500 3950 27534 3984
rect 27568 3950 27602 3984
rect 27636 3950 27670 3984
rect 27704 3950 27738 3984
rect 27772 3950 27806 3984
rect 27840 3950 27874 3984
rect 27908 3950 27942 3984
rect 27976 3950 28000 3984
rect 6415 3910 28000 3950
rect 6415 3876 6473 3910
rect 6507 3876 6542 3910
rect 6576 3876 6611 3910
rect 6645 3876 6680 3910
rect 6714 3876 6749 3910
rect 6783 3876 6818 3910
rect 6852 3876 6887 3910
rect 6921 3876 6956 3910
rect 6990 3876 7025 3910
rect 7059 3876 7094 3910
rect 7128 3876 7163 3910
rect 7197 3876 7232 3910
rect 7266 3876 7301 3910
rect 7335 3876 7370 3910
rect 7404 3876 7439 3910
rect 7473 3876 7508 3910
rect 7542 3876 7577 3910
rect 7611 3876 7646 3910
rect 7680 3876 7715 3910
rect 7749 3876 7784 3910
rect 7818 3876 7853 3910
rect 7887 3876 7922 3910
rect 7956 3876 7991 3910
rect 8025 3876 8060 3910
rect 8094 3876 8129 3910
rect 8163 3876 8198 3910
rect 8232 3876 8267 3910
rect 8301 3876 8336 3910
rect 8370 3876 8405 3910
rect 8439 3876 8474 3910
rect 8508 3876 8543 3910
rect 8577 3876 8612 3910
rect 8646 3876 8681 3910
rect 8715 3876 8750 3910
rect 8784 3876 8819 3910
rect 8853 3876 8888 3910
rect 8922 3876 8957 3910
rect 8991 3876 9026 3910
rect 9060 3876 9095 3910
rect 9129 3876 9164 3910
rect 9198 3876 9233 3910
rect 9267 3876 9302 3910
rect 9336 3876 9371 3910
rect 9405 3876 9440 3910
rect 9474 3876 9509 3910
rect 9543 3876 9578 3910
rect 9612 3876 9647 3910
rect 9681 3876 9716 3910
rect 9750 3876 9785 3910
rect 9819 3876 9854 3910
rect 9888 3876 9922 3910
rect 9956 3876 9990 3910
rect 10024 3876 10058 3910
rect 10092 3876 10126 3910
rect 10160 3876 10194 3910
rect 10228 3876 10262 3910
rect 10296 3876 10330 3910
rect 10364 3876 10398 3910
rect 10432 3876 10466 3910
rect 10500 3876 10534 3910
rect 10568 3876 10602 3910
rect 10636 3876 10670 3910
rect 10704 3876 10738 3910
rect 10772 3876 10806 3910
rect 10840 3876 10874 3910
rect 10908 3876 10942 3910
rect 10976 3876 11010 3910
rect 11044 3876 11078 3910
rect 11112 3876 11146 3910
rect 11180 3876 11214 3910
rect 11248 3876 11282 3910
rect 11316 3876 11350 3910
rect 11384 3876 11418 3910
rect 11452 3876 11486 3910
rect 11520 3876 11554 3910
rect 11588 3876 11622 3910
rect 11656 3876 11690 3910
rect 11724 3876 11758 3910
rect 11792 3876 11826 3910
rect 11860 3876 11894 3910
rect 11928 3876 11962 3910
rect 11996 3876 12030 3910
rect 12064 3876 12098 3910
rect 12132 3876 12166 3910
rect 12200 3876 12234 3910
rect 12268 3876 12302 3910
rect 12336 3876 12370 3910
rect 12404 3876 12438 3910
rect 12472 3876 12506 3910
rect 12540 3876 12574 3910
rect 12608 3876 12642 3910
rect 12676 3876 12710 3910
rect 12744 3876 12778 3910
rect 12812 3876 12846 3910
rect 12880 3876 12914 3910
rect 12948 3876 12982 3910
rect 13016 3876 13050 3910
rect 13084 3876 13118 3910
rect 13152 3876 13186 3910
rect 13220 3876 13254 3910
rect 13288 3876 13322 3910
rect 13356 3876 13390 3910
rect 13424 3876 13458 3910
rect 13492 3876 13526 3910
rect 13560 3876 13594 3910
rect 13628 3876 13662 3910
rect 13696 3876 13730 3910
rect 13764 3876 13798 3910
rect 13832 3876 13866 3910
rect 13900 3876 13934 3910
rect 13968 3876 14002 3910
rect 14036 3876 14070 3910
rect 14104 3876 14138 3910
rect 14172 3876 14206 3910
rect 14240 3876 14274 3910
rect 14308 3876 14342 3910
rect 14376 3876 14410 3910
rect 14444 3876 14478 3910
rect 14512 3876 14546 3910
rect 14580 3876 14614 3910
rect 14648 3876 14682 3910
rect 14716 3876 14750 3910
rect 14784 3876 14818 3910
rect 14852 3876 14886 3910
rect 14920 3876 14954 3910
rect 14988 3876 15022 3910
rect 15056 3876 15090 3910
rect 15124 3876 15158 3910
rect 15192 3876 15226 3910
rect 15260 3876 15294 3910
rect 15328 3876 15362 3910
rect 15396 3876 15430 3910
rect 15464 3876 15498 3910
rect 15532 3876 15566 3910
rect 15600 3876 15634 3910
rect 15668 3876 15702 3910
rect 15736 3876 15770 3910
rect 15804 3876 15838 3910
rect 15872 3876 15906 3910
rect 15940 3876 15974 3910
rect 16008 3876 16042 3910
rect 16076 3876 16110 3910
rect 16144 3876 16178 3910
rect 16212 3876 16246 3910
rect 16280 3876 16314 3910
rect 16348 3876 16382 3910
rect 16416 3876 16450 3910
rect 16484 3876 16518 3910
rect 16552 3876 16586 3910
rect 16620 3876 16654 3910
rect 16688 3876 16722 3910
rect 16756 3876 16790 3910
rect 16824 3876 16858 3910
rect 16892 3876 16926 3910
rect 16960 3876 16994 3910
rect 17028 3876 17062 3910
rect 17096 3876 17130 3910
rect 17164 3876 17198 3910
rect 17232 3876 17266 3910
rect 17300 3876 17334 3910
rect 17368 3876 17402 3910
rect 17436 3876 17470 3910
rect 17504 3876 17538 3910
rect 17572 3876 17606 3910
rect 17640 3876 17674 3910
rect 17708 3876 17742 3910
rect 17776 3876 17810 3910
rect 17844 3876 17878 3910
rect 17912 3876 17946 3910
rect 17980 3876 18014 3910
rect 18048 3876 18082 3910
rect 18116 3876 18150 3910
rect 18184 3876 18218 3910
rect 18252 3876 18286 3910
rect 18320 3876 18354 3910
rect 18388 3876 18422 3910
rect 18456 3876 18490 3910
rect 18524 3876 18558 3910
rect 18592 3876 18626 3910
rect 18660 3876 18694 3910
rect 18728 3876 18762 3910
rect 18796 3876 18830 3910
rect 18864 3876 18898 3910
rect 18932 3876 18966 3910
rect 19000 3876 19034 3910
rect 19068 3876 19102 3910
rect 19136 3876 19170 3910
rect 19204 3876 19238 3910
rect 19272 3876 19306 3910
rect 19340 3876 19374 3910
rect 19408 3876 19442 3910
rect 19476 3876 19510 3910
rect 19544 3876 19578 3910
rect 19612 3876 19646 3910
rect 19680 3876 19714 3910
rect 19748 3876 19782 3910
rect 19816 3876 19850 3910
rect 19884 3876 19918 3910
rect 19952 3876 19986 3910
rect 20020 3876 20054 3910
rect 20088 3876 20122 3910
rect 20156 3876 20190 3910
rect 20224 3876 20258 3910
rect 20292 3876 20326 3910
rect 20360 3876 20394 3910
rect 20428 3876 20462 3910
rect 20496 3876 20530 3910
rect 20564 3876 20598 3910
rect 20632 3876 20666 3910
rect 20700 3876 20734 3910
rect 20768 3876 20802 3910
rect 20836 3876 20870 3910
rect 20904 3876 20938 3910
rect 20972 3876 21006 3910
rect 21040 3876 21074 3910
rect 21108 3876 21142 3910
rect 21176 3876 21210 3910
rect 21244 3876 21278 3910
rect 21312 3876 21346 3910
rect 21380 3876 21414 3910
rect 21448 3876 21482 3910
rect 21516 3876 21550 3910
rect 21584 3876 21618 3910
rect 21652 3876 21686 3910
rect 21720 3876 21754 3910
rect 21788 3876 21822 3910
rect 21856 3876 21890 3910
rect 21924 3876 21958 3910
rect 21992 3876 22026 3910
rect 22060 3876 22094 3910
rect 22128 3876 22162 3910
rect 22196 3876 22230 3910
rect 22264 3876 22298 3910
rect 22332 3876 22366 3910
rect 22400 3876 22434 3910
rect 22468 3876 22502 3910
rect 22536 3876 22570 3910
rect 22604 3876 22638 3910
rect 22672 3876 22706 3910
rect 22740 3876 22774 3910
rect 22808 3876 22842 3910
rect 22876 3876 22910 3910
rect 22944 3876 22978 3910
rect 23012 3876 23046 3910
rect 23080 3876 23114 3910
rect 23148 3876 23182 3910
rect 23216 3876 23250 3910
rect 23284 3876 23318 3910
rect 23352 3876 23386 3910
rect 23420 3876 23454 3910
rect 23488 3876 23522 3910
rect 23556 3876 23590 3910
rect 23624 3876 23658 3910
rect 23692 3876 23726 3910
rect 23760 3876 23794 3910
rect 23828 3876 23862 3910
rect 23896 3876 23930 3910
rect 23964 3876 23998 3910
rect 24032 3876 24066 3910
rect 24100 3876 24134 3910
rect 24168 3876 24202 3910
rect 24236 3876 24270 3910
rect 24304 3876 24338 3910
rect 24372 3876 24406 3910
rect 24440 3876 24474 3910
rect 24508 3876 24542 3910
rect 24576 3876 24610 3910
rect 24644 3876 24678 3910
rect 24712 3876 24746 3910
rect 24780 3876 24814 3910
rect 24848 3876 24882 3910
rect 24916 3876 24950 3910
rect 24984 3876 25018 3910
rect 25052 3876 25086 3910
rect 25120 3876 25154 3910
rect 25188 3876 25222 3910
rect 25256 3876 25290 3910
rect 25324 3876 25358 3910
rect 25392 3876 25426 3910
rect 25460 3876 25494 3910
rect 25528 3876 25562 3910
rect 25596 3876 25630 3910
rect 25664 3876 25698 3910
rect 25732 3876 25766 3910
rect 25800 3876 25834 3910
rect 25868 3876 25902 3910
rect 25936 3876 25970 3910
rect 26004 3876 26038 3910
rect 26072 3876 26106 3910
rect 26140 3876 26174 3910
rect 26208 3876 26242 3910
rect 26276 3876 26310 3910
rect 26344 3876 26378 3910
rect 26412 3876 26446 3910
rect 26480 3876 26514 3910
rect 26548 3876 26582 3910
rect 26616 3876 26650 3910
rect 26684 3876 26718 3910
rect 26752 3876 26786 3910
rect 26820 3876 26854 3910
rect 26888 3876 26922 3910
rect 26956 3876 26990 3910
rect 27024 3876 27058 3910
rect 27092 3876 27126 3910
rect 27160 3876 27194 3910
rect 27228 3876 27262 3910
rect 27296 3876 27330 3910
rect 27364 3876 27398 3910
rect 27432 3876 27466 3910
rect 27500 3876 27534 3910
rect 27568 3876 27602 3910
rect 27636 3876 27670 3910
rect 27704 3876 27738 3910
rect 27772 3876 27806 3910
rect 27840 3876 27874 3910
rect 27908 3876 27942 3910
rect 27976 3876 28000 3910
rect 6415 3836 28000 3876
rect 6415 3802 6473 3836
rect 6507 3802 6542 3836
rect 6576 3802 6611 3836
rect 6645 3802 6680 3836
rect 6714 3802 6749 3836
rect 6783 3802 6818 3836
rect 6852 3802 6887 3836
rect 6921 3802 6956 3836
rect 6990 3802 7025 3836
rect 7059 3802 7094 3836
rect 7128 3802 7163 3836
rect 7197 3802 7232 3836
rect 7266 3802 7301 3836
rect 7335 3802 7370 3836
rect 7404 3802 7439 3836
rect 7473 3802 7508 3836
rect 7542 3802 7577 3836
rect 7611 3802 7646 3836
rect 7680 3802 7715 3836
rect 7749 3802 7784 3836
rect 7818 3802 7853 3836
rect 7887 3802 7922 3836
rect 7956 3802 7991 3836
rect 8025 3802 8060 3836
rect 8094 3802 8129 3836
rect 8163 3802 8198 3836
rect 8232 3802 8267 3836
rect 8301 3802 8336 3836
rect 8370 3802 8405 3836
rect 8439 3802 8474 3836
rect 8508 3802 8543 3836
rect 8577 3802 8612 3836
rect 8646 3802 8681 3836
rect 8715 3802 8750 3836
rect 8784 3802 8819 3836
rect 8853 3802 8888 3836
rect 8922 3802 8957 3836
rect 8991 3802 9026 3836
rect 9060 3802 9095 3836
rect 9129 3802 9164 3836
rect 9198 3802 9233 3836
rect 9267 3802 9302 3836
rect 9336 3802 9371 3836
rect 9405 3802 9440 3836
rect 9474 3802 9509 3836
rect 9543 3802 9578 3836
rect 9612 3802 9647 3836
rect 9681 3802 9716 3836
rect 9750 3802 9785 3836
rect 9819 3802 9854 3836
rect 9888 3802 9922 3836
rect 9956 3802 9990 3836
rect 10024 3802 10058 3836
rect 10092 3802 10126 3836
rect 10160 3802 10194 3836
rect 10228 3802 10262 3836
rect 10296 3802 10330 3836
rect 10364 3802 10398 3836
rect 10432 3802 10466 3836
rect 10500 3802 10534 3836
rect 10568 3802 10602 3836
rect 10636 3802 10670 3836
rect 10704 3802 10738 3836
rect 10772 3802 10806 3836
rect 10840 3802 10874 3836
rect 10908 3802 10942 3836
rect 10976 3802 11010 3836
rect 11044 3802 11078 3836
rect 11112 3802 11146 3836
rect 11180 3802 11214 3836
rect 11248 3802 11282 3836
rect 11316 3802 11350 3836
rect 11384 3802 11418 3836
rect 11452 3802 11486 3836
rect 11520 3802 11554 3836
rect 11588 3802 11622 3836
rect 11656 3802 11690 3836
rect 11724 3802 11758 3836
rect 11792 3802 11826 3836
rect 11860 3802 11894 3836
rect 11928 3802 11962 3836
rect 11996 3802 12030 3836
rect 12064 3802 12098 3836
rect 12132 3802 12166 3836
rect 12200 3802 12234 3836
rect 12268 3802 12302 3836
rect 12336 3802 12370 3836
rect 12404 3802 12438 3836
rect 12472 3802 12506 3836
rect 12540 3802 12574 3836
rect 12608 3802 12642 3836
rect 12676 3802 12710 3836
rect 12744 3802 12778 3836
rect 12812 3802 12846 3836
rect 12880 3802 12914 3836
rect 12948 3802 12982 3836
rect 13016 3802 13050 3836
rect 13084 3802 13118 3836
rect 13152 3802 13186 3836
rect 13220 3802 13254 3836
rect 13288 3802 13322 3836
rect 13356 3802 13390 3836
rect 13424 3802 13458 3836
rect 13492 3802 13526 3836
rect 13560 3802 13594 3836
rect 13628 3802 13662 3836
rect 13696 3802 13730 3836
rect 13764 3802 13798 3836
rect 13832 3802 13866 3836
rect 13900 3802 13934 3836
rect 13968 3802 14002 3836
rect 14036 3802 14070 3836
rect 14104 3802 14138 3836
rect 14172 3802 14206 3836
rect 14240 3802 14274 3836
rect 14308 3802 14342 3836
rect 14376 3802 14410 3836
rect 14444 3802 14478 3836
rect 14512 3802 14546 3836
rect 14580 3802 14614 3836
rect 14648 3802 14682 3836
rect 14716 3802 14750 3836
rect 14784 3802 14818 3836
rect 14852 3802 14886 3836
rect 14920 3802 14954 3836
rect 14988 3802 15022 3836
rect 15056 3802 15090 3836
rect 15124 3802 15158 3836
rect 15192 3802 15226 3836
rect 15260 3802 15294 3836
rect 15328 3802 15362 3836
rect 15396 3802 15430 3836
rect 15464 3802 15498 3836
rect 15532 3802 15566 3836
rect 15600 3802 15634 3836
rect 15668 3802 15702 3836
rect 15736 3802 15770 3836
rect 15804 3802 15838 3836
rect 15872 3802 15906 3836
rect 15940 3802 15974 3836
rect 16008 3802 16042 3836
rect 16076 3802 16110 3836
rect 16144 3802 16178 3836
rect 16212 3802 16246 3836
rect 16280 3802 16314 3836
rect 16348 3802 16382 3836
rect 16416 3802 16450 3836
rect 16484 3802 16518 3836
rect 16552 3802 16586 3836
rect 16620 3802 16654 3836
rect 16688 3802 16722 3836
rect 16756 3802 16790 3836
rect 16824 3802 16858 3836
rect 16892 3802 16926 3836
rect 16960 3802 16994 3836
rect 17028 3802 17062 3836
rect 17096 3802 17130 3836
rect 17164 3802 17198 3836
rect 17232 3802 17266 3836
rect 17300 3802 17334 3836
rect 17368 3802 17402 3836
rect 17436 3802 17470 3836
rect 17504 3802 17538 3836
rect 17572 3802 17606 3836
rect 17640 3802 17674 3836
rect 17708 3802 17742 3836
rect 17776 3802 17810 3836
rect 17844 3802 17878 3836
rect 17912 3802 17946 3836
rect 17980 3802 18014 3836
rect 18048 3802 18082 3836
rect 18116 3802 18150 3836
rect 18184 3802 18218 3836
rect 18252 3802 18286 3836
rect 18320 3802 18354 3836
rect 18388 3802 18422 3836
rect 18456 3802 18490 3836
rect 18524 3802 18558 3836
rect 18592 3802 18626 3836
rect 18660 3802 18694 3836
rect 18728 3802 18762 3836
rect 18796 3802 18830 3836
rect 18864 3802 18898 3836
rect 18932 3802 18966 3836
rect 19000 3802 19034 3836
rect 19068 3802 19102 3836
rect 19136 3802 19170 3836
rect 19204 3802 19238 3836
rect 19272 3802 19306 3836
rect 19340 3802 19374 3836
rect 19408 3802 19442 3836
rect 19476 3802 19510 3836
rect 19544 3802 19578 3836
rect 19612 3802 19646 3836
rect 19680 3802 19714 3836
rect 19748 3802 19782 3836
rect 19816 3802 19850 3836
rect 19884 3802 19918 3836
rect 19952 3802 19986 3836
rect 20020 3802 20054 3836
rect 20088 3802 20122 3836
rect 20156 3802 20190 3836
rect 20224 3802 20258 3836
rect 20292 3802 20326 3836
rect 20360 3802 20394 3836
rect 20428 3802 20462 3836
rect 20496 3802 20530 3836
rect 20564 3802 20598 3836
rect 20632 3802 20666 3836
rect 20700 3802 20734 3836
rect 20768 3802 20802 3836
rect 20836 3802 20870 3836
rect 20904 3802 20938 3836
rect 20972 3802 21006 3836
rect 21040 3802 21074 3836
rect 21108 3802 21142 3836
rect 21176 3802 21210 3836
rect 21244 3802 21278 3836
rect 21312 3802 21346 3836
rect 21380 3802 21414 3836
rect 21448 3802 21482 3836
rect 21516 3802 21550 3836
rect 21584 3802 21618 3836
rect 21652 3802 21686 3836
rect 21720 3802 21754 3836
rect 21788 3802 21822 3836
rect 21856 3802 21890 3836
rect 21924 3802 21958 3836
rect 21992 3802 22026 3836
rect 22060 3802 22094 3836
rect 22128 3802 22162 3836
rect 22196 3802 22230 3836
rect 22264 3802 22298 3836
rect 22332 3802 22366 3836
rect 22400 3802 22434 3836
rect 22468 3802 22502 3836
rect 22536 3802 22570 3836
rect 22604 3802 22638 3836
rect 22672 3802 22706 3836
rect 22740 3802 22774 3836
rect 22808 3802 22842 3836
rect 22876 3802 22910 3836
rect 22944 3802 22978 3836
rect 23012 3802 23046 3836
rect 23080 3802 23114 3836
rect 23148 3802 23182 3836
rect 23216 3802 23250 3836
rect 23284 3802 23318 3836
rect 23352 3802 23386 3836
rect 23420 3802 23454 3836
rect 23488 3802 23522 3836
rect 23556 3802 23590 3836
rect 23624 3802 23658 3836
rect 23692 3802 23726 3836
rect 23760 3802 23794 3836
rect 23828 3802 23862 3836
rect 23896 3802 23930 3836
rect 23964 3802 23998 3836
rect 24032 3802 24066 3836
rect 24100 3802 24134 3836
rect 24168 3802 24202 3836
rect 24236 3802 24270 3836
rect 24304 3802 24338 3836
rect 24372 3802 24406 3836
rect 24440 3802 24474 3836
rect 24508 3802 24542 3836
rect 24576 3802 24610 3836
rect 24644 3802 24678 3836
rect 24712 3802 24746 3836
rect 24780 3802 24814 3836
rect 24848 3802 24882 3836
rect 24916 3802 24950 3836
rect 24984 3802 25018 3836
rect 25052 3802 25086 3836
rect 25120 3802 25154 3836
rect 25188 3802 25222 3836
rect 25256 3802 25290 3836
rect 25324 3802 25358 3836
rect 25392 3802 25426 3836
rect 25460 3802 25494 3836
rect 25528 3802 25562 3836
rect 25596 3802 25630 3836
rect 25664 3802 25698 3836
rect 25732 3802 25766 3836
rect 25800 3802 25834 3836
rect 25868 3802 25902 3836
rect 25936 3802 25970 3836
rect 26004 3802 26038 3836
rect 26072 3802 26106 3836
rect 26140 3802 26174 3836
rect 26208 3802 26242 3836
rect 26276 3802 26310 3836
rect 26344 3802 26378 3836
rect 26412 3802 26446 3836
rect 26480 3802 26514 3836
rect 26548 3802 26582 3836
rect 26616 3802 26650 3836
rect 26684 3802 26718 3836
rect 26752 3802 26786 3836
rect 26820 3802 26854 3836
rect 26888 3802 26922 3836
rect 26956 3802 26990 3836
rect 27024 3802 27058 3836
rect 27092 3802 27126 3836
rect 27160 3802 27194 3836
rect 27228 3802 27262 3836
rect 27296 3802 27330 3836
rect 27364 3802 27398 3836
rect 27432 3802 27466 3836
rect 27500 3802 27534 3836
rect 27568 3802 27602 3836
rect 27636 3802 27670 3836
rect 27704 3802 27738 3836
rect 27772 3802 27806 3836
rect 27840 3802 27874 3836
rect 27908 3802 27942 3836
rect 27976 3802 28000 3836
rect 6415 3762 28000 3802
rect 6415 3754 6473 3762
rect 3292 3728 3316 3754
rect 2320 3692 3316 3728
rect 2320 3688 2532 3692
rect 2566 3688 2624 3692
rect 2658 3688 2716 3692
rect 2750 3688 3316 3692
rect 2320 3654 2344 3688
rect 2378 3654 2415 3688
rect 2449 3654 2486 3688
rect 2520 3658 2532 3688
rect 2591 3658 2624 3688
rect 2520 3654 2557 3658
rect 2591 3654 2628 3658
rect 2662 3654 2698 3688
rect 2750 3658 2768 3688
rect 2732 3654 2768 3658
rect 2802 3654 2838 3688
rect 2872 3654 2908 3688
rect 2942 3654 2978 3688
rect 3012 3654 3048 3688
rect 3082 3654 3118 3688
rect 3152 3654 3188 3688
rect 3222 3654 3258 3688
rect 3292 3654 3316 3688
rect 2320 3614 3316 3654
rect 2320 3580 2344 3614
rect 2378 3580 2415 3614
rect 2449 3580 2486 3614
rect 2520 3605 2557 3614
rect 2591 3605 2628 3614
rect 2520 3580 2532 3605
rect 2591 3580 2624 3605
rect 2662 3580 2698 3614
rect 2732 3605 2768 3614
rect 2750 3580 2768 3605
rect 2802 3580 2838 3614
rect 2872 3580 2908 3614
rect 2942 3580 2978 3614
rect 3012 3580 3048 3614
rect 3082 3580 3118 3614
rect 3152 3580 3188 3614
rect 3222 3580 3258 3614
rect 3292 3580 3316 3614
rect 2320 3571 2532 3580
rect 2566 3571 2624 3580
rect 2658 3571 2716 3580
rect 2750 3571 3316 3580
rect 2320 3540 3316 3571
rect 2320 3506 2344 3540
rect 2378 3506 2415 3540
rect 2449 3506 2486 3540
rect 2520 3518 2557 3540
rect 2591 3518 2628 3540
rect 2520 3506 2532 3518
rect 2591 3506 2624 3518
rect 2662 3506 2698 3540
rect 2732 3518 2768 3540
rect 2750 3506 2768 3518
rect 2802 3506 2838 3540
rect 2872 3506 2908 3540
rect 2942 3506 2978 3540
rect 3012 3506 3048 3540
rect 3082 3506 3118 3540
rect 3152 3506 3188 3540
rect 3222 3506 3258 3540
rect 3292 3506 3316 3540
rect 2320 3484 2532 3506
rect 2566 3484 2624 3506
rect 2658 3484 2716 3506
rect 2750 3484 3316 3506
rect 2320 3466 3316 3484
rect 2320 3432 2344 3466
rect 2378 3432 2415 3466
rect 2449 3432 2486 3466
rect 2520 3432 2557 3466
rect 2591 3432 2628 3466
rect 2662 3432 2698 3466
rect 2732 3432 2768 3466
rect 2802 3432 2838 3466
rect 2872 3432 2908 3466
rect 2942 3432 2978 3466
rect 3012 3432 3048 3466
rect 3082 3432 3118 3466
rect 3152 3432 3188 3466
rect 3222 3432 3258 3466
rect 3292 3432 3316 3466
rect 2320 3430 3316 3432
rect 6449 3728 6473 3754
rect 6507 3728 6542 3762
rect 6576 3728 6611 3762
rect 6645 3728 6680 3762
rect 6714 3728 6749 3762
rect 6783 3728 6818 3762
rect 6852 3728 6887 3762
rect 6921 3728 6956 3762
rect 6990 3728 7025 3762
rect 7059 3728 7094 3762
rect 7128 3728 7163 3762
rect 7197 3728 7232 3762
rect 7266 3728 7301 3762
rect 7335 3728 7370 3762
rect 7404 3728 7439 3762
rect 7473 3728 7508 3762
rect 7542 3728 7577 3762
rect 7611 3728 7646 3762
rect 7680 3728 7715 3762
rect 7749 3728 7784 3762
rect 7818 3728 7853 3762
rect 7887 3728 7922 3762
rect 7956 3728 7991 3762
rect 8025 3728 8060 3762
rect 8094 3728 8129 3762
rect 8163 3728 8198 3762
rect 8232 3728 8267 3762
rect 8301 3728 8336 3762
rect 8370 3728 8405 3762
rect 8439 3728 8474 3762
rect 8508 3728 8543 3762
rect 8577 3728 8612 3762
rect 8646 3728 8681 3762
rect 8715 3728 8750 3762
rect 8784 3728 8819 3762
rect 8853 3728 8888 3762
rect 8922 3728 8957 3762
rect 8991 3728 9026 3762
rect 9060 3728 9095 3762
rect 9129 3728 9164 3762
rect 9198 3728 9233 3762
rect 9267 3728 9302 3762
rect 9336 3728 9371 3762
rect 9405 3728 9440 3762
rect 9474 3728 9509 3762
rect 9543 3728 9578 3762
rect 9612 3728 9647 3762
rect 9681 3728 9716 3762
rect 9750 3728 9785 3762
rect 9819 3728 9854 3762
rect 9888 3728 9922 3762
rect 9956 3728 9990 3762
rect 10024 3728 10058 3762
rect 10092 3728 10126 3762
rect 10160 3728 10194 3762
rect 10228 3728 10262 3762
rect 10296 3728 10330 3762
rect 10364 3728 10398 3762
rect 10432 3728 10466 3762
rect 10500 3728 10534 3762
rect 10568 3728 10602 3762
rect 10636 3728 10670 3762
rect 10704 3728 10738 3762
rect 10772 3728 10806 3762
rect 10840 3728 10874 3762
rect 10908 3728 10942 3762
rect 10976 3728 11010 3762
rect 11044 3728 11078 3762
rect 11112 3728 11146 3762
rect 11180 3728 11214 3762
rect 11248 3728 11282 3762
rect 11316 3728 11350 3762
rect 11384 3728 11418 3762
rect 11452 3728 11486 3762
rect 11520 3728 11554 3762
rect 11588 3728 11622 3762
rect 11656 3728 11690 3762
rect 11724 3728 11758 3762
rect 11792 3728 11826 3762
rect 11860 3728 11894 3762
rect 11928 3728 11962 3762
rect 11996 3728 12030 3762
rect 12064 3728 12098 3762
rect 12132 3728 12166 3762
rect 12200 3728 12234 3762
rect 12268 3728 12302 3762
rect 12336 3728 12370 3762
rect 12404 3728 12438 3762
rect 12472 3728 12506 3762
rect 12540 3728 12574 3762
rect 12608 3728 12642 3762
rect 12676 3728 12710 3762
rect 12744 3728 12778 3762
rect 12812 3728 12846 3762
rect 12880 3728 12914 3762
rect 12948 3728 12982 3762
rect 13016 3728 13050 3762
rect 13084 3728 13118 3762
rect 13152 3728 13186 3762
rect 13220 3728 13254 3762
rect 13288 3728 13322 3762
rect 13356 3728 13390 3762
rect 13424 3728 13458 3762
rect 13492 3728 13526 3762
rect 13560 3728 13594 3762
rect 13628 3728 13662 3762
rect 13696 3728 13730 3762
rect 13764 3728 13798 3762
rect 13832 3728 13866 3762
rect 13900 3728 13934 3762
rect 13968 3728 14002 3762
rect 14036 3728 14070 3762
rect 14104 3728 14138 3762
rect 14172 3728 14206 3762
rect 14240 3728 14274 3762
rect 14308 3728 14342 3762
rect 14376 3728 14410 3762
rect 14444 3728 14478 3762
rect 14512 3728 14546 3762
rect 14580 3728 14614 3762
rect 14648 3728 14682 3762
rect 14716 3728 14750 3762
rect 14784 3728 14818 3762
rect 14852 3728 14886 3762
rect 14920 3728 14954 3762
rect 14988 3728 15022 3762
rect 15056 3728 15090 3762
rect 15124 3728 15158 3762
rect 15192 3728 15226 3762
rect 15260 3728 15294 3762
rect 15328 3728 15362 3762
rect 15396 3728 15430 3762
rect 15464 3728 15498 3762
rect 15532 3728 15566 3762
rect 15600 3728 15634 3762
rect 15668 3728 15702 3762
rect 15736 3728 15770 3762
rect 15804 3728 15838 3762
rect 15872 3728 15906 3762
rect 15940 3728 15974 3762
rect 16008 3728 16042 3762
rect 16076 3728 16110 3762
rect 16144 3728 16178 3762
rect 16212 3728 16246 3762
rect 16280 3728 16314 3762
rect 16348 3728 16382 3762
rect 16416 3728 16450 3762
rect 16484 3728 16518 3762
rect 16552 3728 16586 3762
rect 16620 3728 16654 3762
rect 16688 3728 16722 3762
rect 16756 3728 16790 3762
rect 16824 3728 16858 3762
rect 16892 3728 16926 3762
rect 16960 3728 16994 3762
rect 17028 3728 17062 3762
rect 17096 3728 17130 3762
rect 17164 3728 17198 3762
rect 17232 3728 17266 3762
rect 17300 3728 17334 3762
rect 17368 3728 17402 3762
rect 17436 3728 17470 3762
rect 17504 3728 17538 3762
rect 17572 3728 17606 3762
rect 17640 3728 17674 3762
rect 17708 3728 17742 3762
rect 17776 3728 17810 3762
rect 17844 3728 17878 3762
rect 17912 3728 17946 3762
rect 17980 3728 18014 3762
rect 18048 3728 18082 3762
rect 18116 3728 18150 3762
rect 18184 3728 18218 3762
rect 18252 3728 18286 3762
rect 18320 3728 18354 3762
rect 18388 3728 18422 3762
rect 18456 3728 18490 3762
rect 18524 3728 18558 3762
rect 18592 3728 18626 3762
rect 18660 3728 18694 3762
rect 18728 3728 18762 3762
rect 18796 3728 18830 3762
rect 18864 3728 18898 3762
rect 18932 3728 18966 3762
rect 19000 3728 19034 3762
rect 19068 3728 19102 3762
rect 19136 3728 19170 3762
rect 19204 3728 19238 3762
rect 19272 3728 19306 3762
rect 19340 3728 19374 3762
rect 19408 3728 19442 3762
rect 19476 3728 19510 3762
rect 19544 3728 19578 3762
rect 19612 3728 19646 3762
rect 19680 3728 19714 3762
rect 19748 3728 19782 3762
rect 19816 3728 19850 3762
rect 19884 3728 19918 3762
rect 19952 3728 19986 3762
rect 20020 3728 20054 3762
rect 20088 3728 20122 3762
rect 20156 3728 20190 3762
rect 20224 3728 20258 3762
rect 20292 3728 20326 3762
rect 20360 3728 20394 3762
rect 20428 3728 20462 3762
rect 20496 3728 20530 3762
rect 20564 3728 20598 3762
rect 20632 3728 20666 3762
rect 20700 3728 20734 3762
rect 20768 3728 20802 3762
rect 20836 3728 20870 3762
rect 20904 3728 20938 3762
rect 20972 3728 21006 3762
rect 21040 3728 21074 3762
rect 21108 3728 21142 3762
rect 21176 3728 21210 3762
rect 21244 3728 21278 3762
rect 21312 3728 21346 3762
rect 21380 3728 21414 3762
rect 21448 3728 21482 3762
rect 21516 3728 21550 3762
rect 21584 3728 21618 3762
rect 21652 3728 21686 3762
rect 21720 3728 21754 3762
rect 21788 3728 21822 3762
rect 21856 3728 21890 3762
rect 21924 3728 21958 3762
rect 21992 3728 22026 3762
rect 22060 3728 22094 3762
rect 22128 3728 22162 3762
rect 22196 3728 22230 3762
rect 22264 3728 22298 3762
rect 22332 3728 22366 3762
rect 22400 3728 22434 3762
rect 22468 3728 22502 3762
rect 22536 3728 22570 3762
rect 22604 3728 22638 3762
rect 22672 3728 22706 3762
rect 22740 3728 22774 3762
rect 22808 3728 22842 3762
rect 22876 3728 22910 3762
rect 22944 3728 22978 3762
rect 23012 3728 23046 3762
rect 23080 3728 23114 3762
rect 23148 3728 23182 3762
rect 23216 3728 23250 3762
rect 23284 3728 23318 3762
rect 23352 3728 23386 3762
rect 23420 3728 23454 3762
rect 23488 3728 23522 3762
rect 23556 3728 23590 3762
rect 23624 3728 23658 3762
rect 23692 3728 23726 3762
rect 23760 3728 23794 3762
rect 23828 3728 23862 3762
rect 23896 3728 23930 3762
rect 23964 3728 23998 3762
rect 24032 3728 24066 3762
rect 24100 3728 24134 3762
rect 24168 3728 24202 3762
rect 24236 3728 24270 3762
rect 24304 3728 24338 3762
rect 24372 3728 24406 3762
rect 24440 3728 24474 3762
rect 24508 3728 24542 3762
rect 24576 3728 24610 3762
rect 24644 3728 24678 3762
rect 24712 3728 24746 3762
rect 24780 3728 24814 3762
rect 24848 3728 24882 3762
rect 24916 3728 24950 3762
rect 24984 3728 25018 3762
rect 25052 3728 25086 3762
rect 25120 3728 25154 3762
rect 25188 3728 25222 3762
rect 25256 3728 25290 3762
rect 25324 3728 25358 3762
rect 25392 3728 25426 3762
rect 25460 3728 25494 3762
rect 25528 3728 25562 3762
rect 25596 3728 25630 3762
rect 25664 3728 25698 3762
rect 25732 3728 25766 3762
rect 25800 3728 25834 3762
rect 25868 3728 25902 3762
rect 25936 3728 25970 3762
rect 26004 3728 26038 3762
rect 26072 3728 26106 3762
rect 26140 3728 26174 3762
rect 26208 3728 26242 3762
rect 26276 3728 26310 3762
rect 26344 3728 26378 3762
rect 26412 3728 26446 3762
rect 26480 3728 26514 3762
rect 26548 3728 26582 3762
rect 26616 3728 26650 3762
rect 26684 3728 26718 3762
rect 26752 3728 26786 3762
rect 26820 3728 26854 3762
rect 26888 3728 26922 3762
rect 26956 3728 26990 3762
rect 27024 3728 27058 3762
rect 27092 3728 27126 3762
rect 27160 3728 27194 3762
rect 27228 3728 27262 3762
rect 27296 3728 27330 3762
rect 27364 3728 27398 3762
rect 27432 3728 27466 3762
rect 27500 3728 27534 3762
rect 27568 3728 27602 3762
rect 27636 3728 27670 3762
rect 27704 3728 27738 3762
rect 27772 3728 27806 3762
rect 27840 3728 27874 3762
rect 27908 3728 27942 3762
rect 27976 3728 28000 3762
rect 6449 3688 28000 3728
rect 6449 3654 6473 3688
rect 6507 3654 6542 3688
rect 6576 3654 6611 3688
rect 6645 3654 6680 3688
rect 6714 3654 6749 3688
rect 6783 3654 6818 3688
rect 6852 3654 6887 3688
rect 6921 3654 6956 3688
rect 6990 3654 7025 3688
rect 7059 3654 7094 3688
rect 7128 3654 7163 3688
rect 7197 3654 7232 3688
rect 7266 3654 7301 3688
rect 7335 3654 7370 3688
rect 7404 3654 7439 3688
rect 7473 3654 7508 3688
rect 7542 3654 7577 3688
rect 7611 3654 7646 3688
rect 7680 3654 7715 3688
rect 7749 3654 7784 3688
rect 7818 3654 7853 3688
rect 7887 3654 7922 3688
rect 7956 3654 7991 3688
rect 8025 3654 8060 3688
rect 8094 3654 8129 3688
rect 8163 3654 8198 3688
rect 8232 3654 8267 3688
rect 8301 3654 8336 3688
rect 8370 3654 8405 3688
rect 8439 3654 8474 3688
rect 8508 3654 8543 3688
rect 8577 3654 8612 3688
rect 8646 3654 8681 3688
rect 8715 3654 8750 3688
rect 8784 3654 8819 3688
rect 8853 3654 8888 3688
rect 8922 3654 8957 3688
rect 8991 3654 9026 3688
rect 9060 3654 9095 3688
rect 9129 3654 9164 3688
rect 9198 3654 9233 3688
rect 9267 3654 9302 3688
rect 9336 3654 9371 3688
rect 9405 3654 9440 3688
rect 9474 3654 9509 3688
rect 9543 3654 9578 3688
rect 9612 3654 9647 3688
rect 9681 3654 9716 3688
rect 9750 3654 9785 3688
rect 9819 3654 9854 3688
rect 9888 3654 9922 3688
rect 9956 3654 9990 3688
rect 10024 3654 10058 3688
rect 10092 3654 10126 3688
rect 10160 3654 10194 3688
rect 10228 3654 10262 3688
rect 10296 3654 10330 3688
rect 10364 3654 10398 3688
rect 10432 3654 10466 3688
rect 10500 3654 10534 3688
rect 10568 3654 10602 3688
rect 10636 3654 10670 3688
rect 10704 3654 10738 3688
rect 10772 3654 10806 3688
rect 10840 3654 10874 3688
rect 10908 3654 10942 3688
rect 10976 3654 11010 3688
rect 11044 3654 11078 3688
rect 11112 3654 11146 3688
rect 11180 3654 11214 3688
rect 11248 3654 11282 3688
rect 11316 3654 11350 3688
rect 11384 3654 11418 3688
rect 11452 3654 11486 3688
rect 11520 3654 11554 3688
rect 11588 3654 11622 3688
rect 11656 3654 11690 3688
rect 11724 3654 11758 3688
rect 11792 3654 11826 3688
rect 11860 3654 11894 3688
rect 11928 3654 11962 3688
rect 11996 3654 12030 3688
rect 12064 3654 12098 3688
rect 12132 3654 12166 3688
rect 12200 3654 12234 3688
rect 12268 3654 12302 3688
rect 12336 3654 12370 3688
rect 12404 3654 12438 3688
rect 12472 3654 12506 3688
rect 12540 3654 12574 3688
rect 12608 3654 12642 3688
rect 12676 3654 12710 3688
rect 12744 3654 12778 3688
rect 12812 3654 12846 3688
rect 12880 3654 12914 3688
rect 12948 3654 12982 3688
rect 13016 3654 13050 3688
rect 13084 3654 13118 3688
rect 13152 3654 13186 3688
rect 13220 3654 13254 3688
rect 13288 3654 13322 3688
rect 13356 3654 13390 3688
rect 13424 3654 13458 3688
rect 13492 3654 13526 3688
rect 13560 3654 13594 3688
rect 13628 3654 13662 3688
rect 13696 3654 13730 3688
rect 13764 3654 13798 3688
rect 13832 3654 13866 3688
rect 13900 3654 13934 3688
rect 13968 3654 14002 3688
rect 14036 3654 14070 3688
rect 14104 3654 14138 3688
rect 14172 3654 14206 3688
rect 14240 3654 14274 3688
rect 14308 3654 14342 3688
rect 14376 3654 14410 3688
rect 14444 3654 14478 3688
rect 14512 3654 14546 3688
rect 14580 3654 14614 3688
rect 14648 3654 14682 3688
rect 14716 3654 14750 3688
rect 14784 3654 14818 3688
rect 14852 3654 14886 3688
rect 14920 3654 14954 3688
rect 14988 3654 15022 3688
rect 15056 3654 15090 3688
rect 15124 3654 15158 3688
rect 15192 3654 15226 3688
rect 15260 3654 15294 3688
rect 15328 3654 15362 3688
rect 15396 3654 15430 3688
rect 15464 3654 15498 3688
rect 15532 3654 15566 3688
rect 15600 3654 15634 3688
rect 15668 3654 15702 3688
rect 15736 3654 15770 3688
rect 15804 3654 15838 3688
rect 15872 3654 15906 3688
rect 15940 3654 15974 3688
rect 16008 3654 16042 3688
rect 16076 3654 16110 3688
rect 16144 3654 16178 3688
rect 16212 3654 16246 3688
rect 16280 3654 16314 3688
rect 16348 3654 16382 3688
rect 16416 3654 16450 3688
rect 16484 3654 16518 3688
rect 16552 3654 16586 3688
rect 16620 3654 16654 3688
rect 16688 3654 16722 3688
rect 16756 3654 16790 3688
rect 16824 3654 16858 3688
rect 16892 3654 16926 3688
rect 16960 3654 16994 3688
rect 17028 3654 17062 3688
rect 17096 3654 17130 3688
rect 17164 3654 17198 3688
rect 17232 3654 17266 3688
rect 17300 3654 17334 3688
rect 17368 3654 17402 3688
rect 17436 3654 17470 3688
rect 17504 3654 17538 3688
rect 17572 3654 17606 3688
rect 17640 3654 17674 3688
rect 17708 3654 17742 3688
rect 17776 3654 17810 3688
rect 17844 3654 17878 3688
rect 17912 3654 17946 3688
rect 17980 3654 18014 3688
rect 18048 3654 18082 3688
rect 18116 3654 18150 3688
rect 18184 3654 18218 3688
rect 18252 3654 18286 3688
rect 18320 3654 18354 3688
rect 18388 3654 18422 3688
rect 18456 3654 18490 3688
rect 18524 3654 18558 3688
rect 18592 3654 18626 3688
rect 18660 3654 18694 3688
rect 18728 3654 18762 3688
rect 18796 3654 18830 3688
rect 18864 3654 18898 3688
rect 18932 3654 18966 3688
rect 19000 3654 19034 3688
rect 19068 3654 19102 3688
rect 19136 3654 19170 3688
rect 19204 3654 19238 3688
rect 19272 3654 19306 3688
rect 19340 3654 19374 3688
rect 19408 3654 19442 3688
rect 19476 3654 19510 3688
rect 19544 3654 19578 3688
rect 19612 3654 19646 3688
rect 19680 3654 19714 3688
rect 19748 3654 19782 3688
rect 19816 3654 19850 3688
rect 19884 3654 19918 3688
rect 19952 3654 19986 3688
rect 20020 3654 20054 3688
rect 20088 3654 20122 3688
rect 20156 3654 20190 3688
rect 20224 3654 20258 3688
rect 20292 3654 20326 3688
rect 20360 3654 20394 3688
rect 20428 3654 20462 3688
rect 20496 3654 20530 3688
rect 20564 3654 20598 3688
rect 20632 3654 20666 3688
rect 20700 3654 20734 3688
rect 20768 3654 20802 3688
rect 20836 3654 20870 3688
rect 20904 3654 20938 3688
rect 20972 3654 21006 3688
rect 21040 3654 21074 3688
rect 21108 3654 21142 3688
rect 21176 3654 21210 3688
rect 21244 3654 21278 3688
rect 21312 3654 21346 3688
rect 21380 3654 21414 3688
rect 21448 3654 21482 3688
rect 21516 3654 21550 3688
rect 21584 3654 21618 3688
rect 21652 3654 21686 3688
rect 21720 3654 21754 3688
rect 21788 3654 21822 3688
rect 21856 3654 21890 3688
rect 21924 3654 21958 3688
rect 21992 3654 22026 3688
rect 22060 3654 22094 3688
rect 22128 3654 22162 3688
rect 22196 3654 22230 3688
rect 22264 3654 22298 3688
rect 22332 3654 22366 3688
rect 22400 3654 22434 3688
rect 22468 3654 22502 3688
rect 22536 3654 22570 3688
rect 22604 3654 22638 3688
rect 22672 3654 22706 3688
rect 22740 3654 22774 3688
rect 22808 3654 22842 3688
rect 22876 3654 22910 3688
rect 22944 3654 22978 3688
rect 23012 3654 23046 3688
rect 23080 3654 23114 3688
rect 23148 3654 23182 3688
rect 23216 3654 23250 3688
rect 23284 3654 23318 3688
rect 23352 3654 23386 3688
rect 23420 3654 23454 3688
rect 23488 3654 23522 3688
rect 23556 3654 23590 3688
rect 23624 3654 23658 3688
rect 23692 3654 23726 3688
rect 23760 3654 23794 3688
rect 23828 3654 23862 3688
rect 23896 3654 23930 3688
rect 23964 3654 23998 3688
rect 24032 3654 24066 3688
rect 24100 3654 24134 3688
rect 24168 3654 24202 3688
rect 24236 3654 24270 3688
rect 24304 3654 24338 3688
rect 24372 3654 24406 3688
rect 24440 3654 24474 3688
rect 24508 3654 24542 3688
rect 24576 3654 24610 3688
rect 24644 3654 24678 3688
rect 24712 3654 24746 3688
rect 24780 3654 24814 3688
rect 24848 3654 24882 3688
rect 24916 3654 24950 3688
rect 24984 3654 25018 3688
rect 25052 3654 25086 3688
rect 25120 3654 25154 3688
rect 25188 3654 25222 3688
rect 25256 3654 25290 3688
rect 25324 3654 25358 3688
rect 25392 3654 25426 3688
rect 25460 3654 25494 3688
rect 25528 3654 25562 3688
rect 25596 3654 25630 3688
rect 25664 3654 25698 3688
rect 25732 3654 25766 3688
rect 25800 3654 25834 3688
rect 25868 3654 25902 3688
rect 25936 3654 25970 3688
rect 26004 3654 26038 3688
rect 26072 3654 26106 3688
rect 26140 3654 26174 3688
rect 26208 3654 26242 3688
rect 26276 3654 26310 3688
rect 26344 3654 26378 3688
rect 26412 3654 26446 3688
rect 26480 3654 26514 3688
rect 26548 3654 26582 3688
rect 26616 3654 26650 3688
rect 26684 3654 26718 3688
rect 26752 3654 26786 3688
rect 26820 3654 26854 3688
rect 26888 3654 26922 3688
rect 26956 3654 26990 3688
rect 27024 3654 27058 3688
rect 27092 3654 27126 3688
rect 27160 3654 27194 3688
rect 27228 3654 27262 3688
rect 27296 3654 27330 3688
rect 27364 3654 27398 3688
rect 27432 3654 27466 3688
rect 27500 3654 27534 3688
rect 27568 3654 27602 3688
rect 27636 3654 27670 3688
rect 27704 3654 27738 3688
rect 27772 3654 27806 3688
rect 27840 3654 27874 3688
rect 27908 3654 27942 3688
rect 27976 3654 28000 3688
rect 6449 3614 28000 3654
rect 6449 3580 6473 3614
rect 6507 3580 6542 3614
rect 6576 3580 6611 3614
rect 6645 3580 6680 3614
rect 6714 3580 6749 3614
rect 6783 3580 6818 3614
rect 6852 3580 6887 3614
rect 6921 3580 6956 3614
rect 6990 3580 7025 3614
rect 7059 3580 7094 3614
rect 7128 3580 7163 3614
rect 7197 3580 7232 3614
rect 7266 3580 7301 3614
rect 7335 3580 7370 3614
rect 7404 3580 7439 3614
rect 7473 3580 7508 3614
rect 7542 3580 7577 3614
rect 7611 3580 7646 3614
rect 7680 3580 7715 3614
rect 7749 3580 7784 3614
rect 7818 3580 7853 3614
rect 7887 3580 7922 3614
rect 7956 3580 7991 3614
rect 8025 3580 8060 3614
rect 8094 3580 8129 3614
rect 8163 3580 8198 3614
rect 8232 3580 8267 3614
rect 8301 3580 8336 3614
rect 8370 3580 8405 3614
rect 8439 3580 8474 3614
rect 8508 3580 8543 3614
rect 8577 3580 8612 3614
rect 8646 3580 8681 3614
rect 8715 3580 8750 3614
rect 8784 3580 8819 3614
rect 8853 3580 8888 3614
rect 8922 3580 8957 3614
rect 8991 3580 9026 3614
rect 9060 3580 9095 3614
rect 9129 3580 9164 3614
rect 9198 3580 9233 3614
rect 9267 3580 9302 3614
rect 9336 3580 9371 3614
rect 9405 3580 9440 3614
rect 9474 3580 9509 3614
rect 9543 3580 9578 3614
rect 9612 3580 9647 3614
rect 9681 3580 9716 3614
rect 9750 3580 9785 3614
rect 9819 3580 9854 3614
rect 9888 3580 9922 3614
rect 9956 3580 9990 3614
rect 10024 3580 10058 3614
rect 10092 3580 10126 3614
rect 10160 3580 10194 3614
rect 10228 3580 10262 3614
rect 10296 3580 10330 3614
rect 10364 3580 10398 3614
rect 10432 3580 10466 3614
rect 10500 3580 10534 3614
rect 10568 3580 10602 3614
rect 10636 3580 10670 3614
rect 10704 3580 10738 3614
rect 10772 3580 10806 3614
rect 10840 3580 10874 3614
rect 10908 3580 10942 3614
rect 10976 3580 11010 3614
rect 11044 3580 11078 3614
rect 11112 3580 11146 3614
rect 11180 3580 11214 3614
rect 11248 3580 11282 3614
rect 11316 3580 11350 3614
rect 11384 3580 11418 3614
rect 11452 3580 11486 3614
rect 11520 3580 11554 3614
rect 11588 3580 11622 3614
rect 11656 3580 11690 3614
rect 11724 3580 11758 3614
rect 11792 3580 11826 3614
rect 11860 3580 11894 3614
rect 11928 3580 11962 3614
rect 11996 3580 12030 3614
rect 12064 3580 12098 3614
rect 12132 3580 12166 3614
rect 12200 3580 12234 3614
rect 12268 3580 12302 3614
rect 12336 3580 12370 3614
rect 12404 3580 12438 3614
rect 12472 3580 12506 3614
rect 12540 3580 12574 3614
rect 12608 3580 12642 3614
rect 12676 3580 12710 3614
rect 12744 3580 12778 3614
rect 12812 3580 12846 3614
rect 12880 3580 12914 3614
rect 12948 3580 12982 3614
rect 13016 3580 13050 3614
rect 13084 3580 13118 3614
rect 13152 3580 13186 3614
rect 13220 3580 13254 3614
rect 13288 3580 13322 3614
rect 13356 3580 13390 3614
rect 13424 3580 13458 3614
rect 13492 3580 13526 3614
rect 13560 3580 13594 3614
rect 13628 3580 13662 3614
rect 13696 3580 13730 3614
rect 13764 3580 13798 3614
rect 13832 3580 13866 3614
rect 13900 3580 13934 3614
rect 13968 3580 14002 3614
rect 14036 3580 14070 3614
rect 14104 3580 14138 3614
rect 14172 3580 14206 3614
rect 14240 3580 14274 3614
rect 14308 3580 14342 3614
rect 14376 3580 14410 3614
rect 14444 3580 14478 3614
rect 14512 3580 14546 3614
rect 14580 3580 14614 3614
rect 14648 3580 14682 3614
rect 14716 3580 14750 3614
rect 14784 3580 14818 3614
rect 14852 3580 14886 3614
rect 14920 3580 14954 3614
rect 14988 3580 15022 3614
rect 15056 3580 15090 3614
rect 15124 3580 15158 3614
rect 15192 3580 15226 3614
rect 15260 3580 15294 3614
rect 15328 3580 15362 3614
rect 15396 3580 15430 3614
rect 15464 3580 15498 3614
rect 15532 3580 15566 3614
rect 15600 3580 15634 3614
rect 15668 3580 15702 3614
rect 15736 3580 15770 3614
rect 15804 3580 15838 3614
rect 15872 3580 15906 3614
rect 15940 3580 15974 3614
rect 16008 3580 16042 3614
rect 16076 3580 16110 3614
rect 16144 3580 16178 3614
rect 16212 3580 16246 3614
rect 16280 3580 16314 3614
rect 16348 3580 16382 3614
rect 16416 3580 16450 3614
rect 16484 3580 16518 3614
rect 16552 3580 16586 3614
rect 16620 3580 16654 3614
rect 16688 3580 16722 3614
rect 16756 3580 16790 3614
rect 16824 3580 16858 3614
rect 16892 3580 16926 3614
rect 16960 3580 16994 3614
rect 17028 3580 17062 3614
rect 17096 3580 17130 3614
rect 17164 3580 17198 3614
rect 17232 3580 17266 3614
rect 17300 3580 17334 3614
rect 17368 3580 17402 3614
rect 17436 3580 17470 3614
rect 17504 3580 17538 3614
rect 17572 3580 17606 3614
rect 17640 3580 17674 3614
rect 17708 3580 17742 3614
rect 17776 3580 17810 3614
rect 17844 3580 17878 3614
rect 17912 3580 17946 3614
rect 17980 3580 18014 3614
rect 18048 3580 18082 3614
rect 18116 3580 18150 3614
rect 18184 3580 18218 3614
rect 18252 3580 18286 3614
rect 18320 3580 18354 3614
rect 18388 3580 18422 3614
rect 18456 3580 18490 3614
rect 18524 3580 18558 3614
rect 18592 3580 18626 3614
rect 18660 3580 18694 3614
rect 18728 3580 18762 3614
rect 18796 3580 18830 3614
rect 18864 3580 18898 3614
rect 18932 3580 18966 3614
rect 19000 3580 19034 3614
rect 19068 3580 19102 3614
rect 19136 3580 19170 3614
rect 19204 3580 19238 3614
rect 19272 3580 19306 3614
rect 19340 3580 19374 3614
rect 19408 3580 19442 3614
rect 19476 3580 19510 3614
rect 19544 3580 19578 3614
rect 19612 3580 19646 3614
rect 19680 3580 19714 3614
rect 19748 3580 19782 3614
rect 19816 3580 19850 3614
rect 19884 3580 19918 3614
rect 19952 3580 19986 3614
rect 20020 3580 20054 3614
rect 20088 3580 20122 3614
rect 20156 3580 20190 3614
rect 20224 3580 20258 3614
rect 20292 3580 20326 3614
rect 20360 3580 20394 3614
rect 20428 3580 20462 3614
rect 20496 3580 20530 3614
rect 20564 3580 20598 3614
rect 20632 3580 20666 3614
rect 20700 3580 20734 3614
rect 20768 3580 20802 3614
rect 20836 3580 20870 3614
rect 20904 3580 20938 3614
rect 20972 3580 21006 3614
rect 21040 3580 21074 3614
rect 21108 3580 21142 3614
rect 21176 3580 21210 3614
rect 21244 3580 21278 3614
rect 21312 3580 21346 3614
rect 21380 3580 21414 3614
rect 21448 3580 21482 3614
rect 21516 3580 21550 3614
rect 21584 3580 21618 3614
rect 21652 3580 21686 3614
rect 21720 3580 21754 3614
rect 21788 3580 21822 3614
rect 21856 3580 21890 3614
rect 21924 3580 21958 3614
rect 21992 3580 22026 3614
rect 22060 3580 22094 3614
rect 22128 3580 22162 3614
rect 22196 3580 22230 3614
rect 22264 3580 22298 3614
rect 22332 3580 22366 3614
rect 22400 3580 22434 3614
rect 22468 3580 22502 3614
rect 22536 3580 22570 3614
rect 22604 3580 22638 3614
rect 22672 3580 22706 3614
rect 22740 3580 22774 3614
rect 22808 3580 22842 3614
rect 22876 3580 22910 3614
rect 22944 3580 22978 3614
rect 23012 3580 23046 3614
rect 23080 3580 23114 3614
rect 23148 3580 23182 3614
rect 23216 3580 23250 3614
rect 23284 3580 23318 3614
rect 23352 3580 23386 3614
rect 23420 3580 23454 3614
rect 23488 3580 23522 3614
rect 23556 3580 23590 3614
rect 23624 3580 23658 3614
rect 23692 3580 23726 3614
rect 23760 3580 23794 3614
rect 23828 3580 23862 3614
rect 23896 3580 23930 3614
rect 23964 3580 23998 3614
rect 24032 3580 24066 3614
rect 24100 3580 24134 3614
rect 24168 3580 24202 3614
rect 24236 3580 24270 3614
rect 24304 3580 24338 3614
rect 24372 3580 24406 3614
rect 24440 3580 24474 3614
rect 24508 3580 24542 3614
rect 24576 3580 24610 3614
rect 24644 3580 24678 3614
rect 24712 3580 24746 3614
rect 24780 3580 24814 3614
rect 24848 3580 24882 3614
rect 24916 3580 24950 3614
rect 24984 3580 25018 3614
rect 25052 3580 25086 3614
rect 25120 3580 25154 3614
rect 25188 3580 25222 3614
rect 25256 3580 25290 3614
rect 25324 3580 25358 3614
rect 25392 3580 25426 3614
rect 25460 3580 25494 3614
rect 25528 3580 25562 3614
rect 25596 3580 25630 3614
rect 25664 3580 25698 3614
rect 25732 3580 25766 3614
rect 25800 3580 25834 3614
rect 25868 3580 25902 3614
rect 25936 3580 25970 3614
rect 26004 3580 26038 3614
rect 26072 3580 26106 3614
rect 26140 3580 26174 3614
rect 26208 3580 26242 3614
rect 26276 3580 26310 3614
rect 26344 3580 26378 3614
rect 26412 3580 26446 3614
rect 26480 3580 26514 3614
rect 26548 3580 26582 3614
rect 26616 3580 26650 3614
rect 26684 3580 26718 3614
rect 26752 3580 26786 3614
rect 26820 3580 26854 3614
rect 26888 3580 26922 3614
rect 26956 3580 26990 3614
rect 27024 3580 27058 3614
rect 27092 3580 27126 3614
rect 27160 3580 27194 3614
rect 27228 3580 27262 3614
rect 27296 3580 27330 3614
rect 27364 3580 27398 3614
rect 27432 3580 27466 3614
rect 27500 3580 27534 3614
rect 27568 3580 27602 3614
rect 27636 3580 27670 3614
rect 27704 3580 27738 3614
rect 27772 3580 27806 3614
rect 27840 3580 27874 3614
rect 27908 3580 27942 3614
rect 27976 3580 28000 3614
rect 6449 3561 28000 3580
rect 6449 3540 12119 3561
rect 12153 3540 12193 3561
rect 12227 3540 12267 3561
rect 12301 3540 12341 3561
rect 12375 3540 12415 3561
rect 12449 3540 12489 3561
rect 12523 3540 12563 3561
rect 12597 3540 12637 3561
rect 12671 3540 12711 3561
rect 12745 3540 12785 3561
rect 12819 3540 12859 3561
rect 12893 3540 12933 3561
rect 12967 3540 13006 3561
rect 13040 3540 13079 3561
rect 13113 3540 13152 3561
rect 6449 3506 6473 3540
rect 6507 3506 6542 3540
rect 6576 3506 6611 3540
rect 6645 3506 6680 3540
rect 6714 3506 6749 3540
rect 6783 3506 6818 3540
rect 6852 3506 6887 3540
rect 6921 3506 6956 3540
rect 6990 3506 7025 3540
rect 7059 3506 7094 3540
rect 7128 3506 7163 3540
rect 7197 3506 7232 3540
rect 7266 3506 7301 3540
rect 7335 3506 7370 3540
rect 7404 3506 7439 3540
rect 7473 3506 7508 3540
rect 7542 3506 7577 3540
rect 7611 3506 7646 3540
rect 7680 3506 7715 3540
rect 7749 3506 7784 3540
rect 7818 3506 7853 3540
rect 7887 3506 7922 3540
rect 7956 3506 7991 3540
rect 8025 3506 8060 3540
rect 8094 3506 8129 3540
rect 8163 3506 8198 3540
rect 8232 3506 8267 3540
rect 8301 3506 8336 3540
rect 8370 3506 8405 3540
rect 8439 3506 8474 3540
rect 8508 3506 8543 3540
rect 8577 3506 8612 3540
rect 8646 3506 8681 3540
rect 8715 3506 8750 3540
rect 8784 3506 8819 3540
rect 8853 3506 8888 3540
rect 8922 3506 8957 3540
rect 8991 3506 9026 3540
rect 9060 3506 9095 3540
rect 9129 3506 9164 3540
rect 9198 3506 9233 3540
rect 9267 3506 9302 3540
rect 9336 3506 9371 3540
rect 9405 3506 9440 3540
rect 9474 3506 9509 3540
rect 9543 3506 9578 3540
rect 9612 3506 9647 3540
rect 9681 3506 9716 3540
rect 9750 3506 9785 3540
rect 9819 3506 9854 3540
rect 9888 3506 9922 3540
rect 9956 3506 9990 3540
rect 10024 3506 10058 3540
rect 10092 3506 10126 3540
rect 10160 3506 10194 3540
rect 10228 3506 10262 3540
rect 10296 3506 10330 3540
rect 10364 3506 10398 3540
rect 10432 3506 10466 3540
rect 10500 3506 10534 3540
rect 10568 3506 10602 3540
rect 10636 3506 10670 3540
rect 10704 3506 10738 3540
rect 10772 3506 10806 3540
rect 10840 3506 10874 3540
rect 10908 3506 10942 3540
rect 10976 3506 11010 3540
rect 11044 3506 11078 3540
rect 11112 3506 11146 3540
rect 11180 3506 11214 3540
rect 11248 3506 11282 3540
rect 11316 3506 11350 3540
rect 11384 3506 11418 3540
rect 11452 3506 11486 3540
rect 11520 3506 11554 3540
rect 11588 3506 11622 3540
rect 11656 3506 11690 3540
rect 11724 3506 11758 3540
rect 11792 3506 11826 3540
rect 11860 3506 11894 3540
rect 11928 3506 11962 3540
rect 11996 3506 12030 3540
rect 12064 3506 12098 3540
rect 12153 3527 12166 3540
rect 12227 3527 12234 3540
rect 12301 3527 12302 3540
rect 12132 3506 12166 3527
rect 12200 3506 12234 3527
rect 12268 3506 12302 3527
rect 12336 3527 12341 3540
rect 12404 3527 12415 3540
rect 12472 3527 12489 3540
rect 12540 3527 12563 3540
rect 12608 3527 12637 3540
rect 12336 3506 12370 3527
rect 12404 3506 12438 3527
rect 12472 3506 12506 3527
rect 12540 3506 12574 3527
rect 12608 3506 12642 3527
rect 12676 3506 12710 3540
rect 12745 3527 12778 3540
rect 12819 3527 12846 3540
rect 12893 3527 12914 3540
rect 12967 3527 12982 3540
rect 13040 3527 13050 3540
rect 13113 3527 13118 3540
rect 12744 3506 12778 3527
rect 12812 3506 12846 3527
rect 12880 3506 12914 3527
rect 12948 3506 12982 3527
rect 13016 3506 13050 3527
rect 13084 3506 13118 3527
rect 13186 3540 13225 3561
rect 13259 3540 13298 3561
rect 13332 3540 13371 3561
rect 13405 3540 13444 3561
rect 13478 3540 13517 3561
rect 13551 3540 13590 3561
rect 13624 3540 13663 3561
rect 13697 3540 13736 3561
rect 13770 3540 13809 3561
rect 13843 3540 13882 3561
rect 13916 3540 13955 3561
rect 13989 3540 14028 3561
rect 14062 3540 14101 3561
rect 14135 3540 14174 3561
rect 14208 3540 14247 3561
rect 14281 3540 14320 3561
rect 14354 3540 14393 3561
rect 14427 3540 14466 3561
rect 14500 3540 14539 3561
rect 14573 3540 14612 3561
rect 14646 3540 14685 3561
rect 14719 3540 14758 3561
rect 14792 3540 28000 3561
rect 13152 3506 13186 3527
rect 13220 3527 13225 3540
rect 13288 3527 13298 3540
rect 13356 3527 13371 3540
rect 13424 3527 13444 3540
rect 13492 3527 13517 3540
rect 13560 3527 13590 3540
rect 13220 3506 13254 3527
rect 13288 3506 13322 3527
rect 13356 3506 13390 3527
rect 13424 3506 13458 3527
rect 13492 3506 13526 3527
rect 13560 3506 13594 3527
rect 13628 3506 13662 3540
rect 13697 3527 13730 3540
rect 13770 3527 13798 3540
rect 13843 3527 13866 3540
rect 13916 3527 13934 3540
rect 13989 3527 14002 3540
rect 14062 3527 14070 3540
rect 14135 3527 14138 3540
rect 13696 3506 13730 3527
rect 13764 3506 13798 3527
rect 13832 3506 13866 3527
rect 13900 3506 13934 3527
rect 13968 3506 14002 3527
rect 14036 3506 14070 3527
rect 14104 3506 14138 3527
rect 14172 3527 14174 3540
rect 14240 3527 14247 3540
rect 14308 3527 14320 3540
rect 14376 3527 14393 3540
rect 14444 3527 14466 3540
rect 14512 3527 14539 3540
rect 14580 3527 14612 3540
rect 14172 3506 14206 3527
rect 14240 3506 14274 3527
rect 14308 3506 14342 3527
rect 14376 3506 14410 3527
rect 14444 3506 14478 3527
rect 14512 3506 14546 3527
rect 14580 3506 14614 3527
rect 14648 3506 14682 3540
rect 14719 3527 14750 3540
rect 14792 3527 14818 3540
rect 14716 3506 14750 3527
rect 14784 3506 14818 3527
rect 14852 3506 14886 3540
rect 14920 3506 14954 3540
rect 14988 3506 15022 3540
rect 15056 3506 15090 3540
rect 15124 3506 15158 3540
rect 15192 3506 15226 3540
rect 15260 3506 15294 3540
rect 15328 3506 15362 3540
rect 15396 3506 15430 3540
rect 15464 3506 15498 3540
rect 15532 3506 15566 3540
rect 15600 3506 15634 3540
rect 15668 3506 15702 3540
rect 15736 3506 15770 3540
rect 15804 3506 15838 3540
rect 15872 3506 15906 3540
rect 15940 3506 15974 3540
rect 16008 3506 16042 3540
rect 16076 3506 16110 3540
rect 16144 3506 16178 3540
rect 16212 3506 16246 3540
rect 16280 3506 16314 3540
rect 16348 3506 16382 3540
rect 16416 3506 16450 3540
rect 16484 3506 16518 3540
rect 16552 3506 16586 3540
rect 16620 3506 16654 3540
rect 16688 3506 16722 3540
rect 16756 3506 16790 3540
rect 16824 3506 16858 3540
rect 16892 3506 16926 3540
rect 16960 3506 16994 3540
rect 17028 3506 17062 3540
rect 17124 3506 17130 3540
rect 17164 3506 17166 3540
rect 17232 3506 17242 3540
rect 17300 3506 17318 3540
rect 17368 3506 17394 3540
rect 17436 3506 17470 3540
rect 17504 3506 17538 3540
rect 17579 3506 17606 3540
rect 17654 3506 17674 3540
rect 17729 3506 17742 3540
rect 17804 3506 17810 3540
rect 17844 3506 17845 3540
rect 17912 3506 17920 3540
rect 17980 3506 17995 3540
rect 18048 3506 18070 3540
rect 18116 3506 18145 3540
rect 18184 3506 18218 3540
rect 18254 3506 18286 3540
rect 18329 3506 18354 3540
rect 18404 3506 18422 3540
rect 18479 3506 18490 3540
rect 18554 3506 18558 3540
rect 18592 3506 18595 3540
rect 18660 3506 18670 3540
rect 18728 3506 18762 3540
rect 18796 3506 18830 3540
rect 18864 3506 18898 3540
rect 18932 3506 18966 3540
rect 19000 3506 19034 3540
rect 19068 3506 19102 3540
rect 19136 3506 19170 3540
rect 19204 3506 19238 3540
rect 19272 3506 19306 3540
rect 19340 3506 19374 3540
rect 19408 3506 19442 3540
rect 19476 3506 19510 3540
rect 19544 3506 19578 3540
rect 19612 3506 19646 3540
rect 19680 3506 19714 3540
rect 19748 3506 19782 3540
rect 19816 3506 19850 3540
rect 19884 3506 19918 3540
rect 19952 3506 19986 3540
rect 20020 3506 20054 3540
rect 20088 3506 20122 3540
rect 20156 3506 20190 3540
rect 20224 3506 20258 3540
rect 20292 3506 20326 3540
rect 20360 3506 20394 3540
rect 20428 3506 20462 3540
rect 20496 3506 20530 3540
rect 20564 3506 20598 3540
rect 20632 3506 20666 3540
rect 20700 3506 20734 3540
rect 20768 3506 20802 3540
rect 20836 3506 20870 3540
rect 20904 3506 20938 3540
rect 20972 3506 21006 3540
rect 21040 3506 21074 3540
rect 21108 3506 21142 3540
rect 21176 3506 21210 3540
rect 21244 3506 21278 3540
rect 21312 3506 21346 3540
rect 21380 3506 21414 3540
rect 21448 3506 21482 3540
rect 21516 3506 21550 3540
rect 21584 3506 21618 3540
rect 21652 3506 21686 3540
rect 21720 3506 21754 3540
rect 21788 3506 21822 3540
rect 21856 3506 21890 3540
rect 21924 3506 21958 3540
rect 21992 3506 22026 3540
rect 22060 3506 22094 3540
rect 22128 3506 22162 3540
rect 22196 3506 22230 3540
rect 22264 3506 22298 3540
rect 22332 3506 22366 3540
rect 22400 3506 22434 3540
rect 22468 3506 22502 3540
rect 22536 3506 22570 3540
rect 22604 3506 22638 3540
rect 22672 3506 22706 3540
rect 22740 3506 22774 3540
rect 22808 3506 22842 3540
rect 22876 3506 22910 3540
rect 22944 3506 22978 3540
rect 23012 3506 23046 3540
rect 23080 3506 23114 3540
rect 23148 3506 23182 3540
rect 23216 3506 23250 3540
rect 23284 3506 23318 3540
rect 23352 3506 23386 3540
rect 23420 3506 23454 3540
rect 23488 3506 23522 3540
rect 23556 3506 23590 3540
rect 23624 3506 23658 3540
rect 23692 3506 23726 3540
rect 23760 3506 23794 3540
rect 23828 3506 23862 3540
rect 23896 3506 23930 3540
rect 23964 3506 23998 3540
rect 24032 3506 24066 3540
rect 24100 3506 24134 3540
rect 24168 3506 24202 3540
rect 24236 3506 24270 3540
rect 24304 3506 24338 3540
rect 24372 3506 24406 3540
rect 24440 3506 24474 3540
rect 24508 3506 24542 3540
rect 24576 3506 24610 3540
rect 24644 3506 24678 3540
rect 24712 3506 24746 3540
rect 24780 3506 24814 3540
rect 24848 3506 24882 3540
rect 24916 3506 24950 3540
rect 24984 3506 25018 3540
rect 25052 3506 25086 3540
rect 25120 3506 25154 3540
rect 25188 3506 25222 3540
rect 25256 3506 25290 3540
rect 25324 3506 25358 3540
rect 25392 3506 25426 3540
rect 25460 3506 25494 3540
rect 25528 3506 25562 3540
rect 25596 3506 25630 3540
rect 25664 3506 25698 3540
rect 25732 3506 25766 3540
rect 25800 3506 25834 3540
rect 25868 3506 25902 3540
rect 25936 3506 25970 3540
rect 26004 3506 26038 3540
rect 26072 3506 26106 3540
rect 26140 3506 26174 3540
rect 26208 3506 26242 3540
rect 26276 3506 26310 3540
rect 26344 3506 26378 3540
rect 26412 3506 26446 3540
rect 26480 3506 26514 3540
rect 26548 3506 26582 3540
rect 26616 3506 26650 3540
rect 26684 3506 26718 3540
rect 26752 3506 26786 3540
rect 26820 3506 26854 3540
rect 26888 3506 26922 3540
rect 26956 3506 26990 3540
rect 27024 3506 27058 3540
rect 27092 3506 27126 3540
rect 27160 3506 27194 3540
rect 27228 3506 27262 3540
rect 27296 3506 27330 3540
rect 27364 3506 27398 3540
rect 27432 3506 27466 3540
rect 27500 3506 27534 3540
rect 27568 3506 27602 3540
rect 27636 3506 27670 3540
rect 27704 3506 27738 3540
rect 27772 3506 27806 3540
rect 27840 3506 27874 3540
rect 27908 3506 27942 3540
rect 27976 3506 28000 3540
rect 6449 3483 28000 3506
rect 6449 3466 12119 3483
rect 12153 3466 12193 3483
rect 12227 3466 12267 3483
rect 12301 3466 12341 3483
rect 12375 3466 12415 3483
rect 12449 3466 12489 3483
rect 12523 3466 12563 3483
rect 12597 3466 12637 3483
rect 12671 3466 12711 3483
rect 12745 3466 12785 3483
rect 12819 3466 12859 3483
rect 12893 3466 12933 3483
rect 12967 3466 13006 3483
rect 13040 3466 13079 3483
rect 13113 3466 13152 3483
rect 6449 3432 6473 3466
rect 6507 3432 6542 3466
rect 6576 3432 6611 3466
rect 6645 3432 6680 3466
rect 6714 3432 6749 3466
rect 6783 3432 6818 3466
rect 6852 3432 6887 3466
rect 6921 3432 6956 3466
rect 6990 3432 7025 3466
rect 7059 3432 7094 3466
rect 7128 3432 7163 3466
rect 7197 3432 7232 3466
rect 7266 3432 7301 3466
rect 7335 3432 7370 3466
rect 7404 3432 7439 3466
rect 7473 3432 7508 3466
rect 7542 3432 7577 3466
rect 7611 3432 7646 3466
rect 7680 3432 7715 3466
rect 7749 3432 7784 3466
rect 7818 3432 7853 3466
rect 7887 3432 7922 3466
rect 7956 3432 7991 3466
rect 8025 3432 8060 3466
rect 8094 3432 8129 3466
rect 8163 3432 8198 3466
rect 8232 3432 8267 3466
rect 8301 3432 8336 3466
rect 8370 3432 8405 3466
rect 8439 3432 8474 3466
rect 8508 3432 8543 3466
rect 8577 3432 8612 3466
rect 8646 3432 8681 3466
rect 8715 3432 8750 3466
rect 8784 3432 8819 3466
rect 8853 3432 8888 3466
rect 8922 3432 8957 3466
rect 8991 3432 9026 3466
rect 9060 3432 9095 3466
rect 9129 3432 9164 3466
rect 9198 3432 9233 3466
rect 9267 3432 9302 3466
rect 9336 3432 9371 3466
rect 9405 3432 9440 3466
rect 9474 3432 9509 3466
rect 9543 3432 9578 3466
rect 9612 3432 9647 3466
rect 9681 3432 9716 3466
rect 9750 3432 9785 3466
rect 9819 3432 9854 3466
rect 9888 3432 9922 3466
rect 9956 3432 9990 3466
rect 10024 3432 10058 3466
rect 10092 3432 10126 3466
rect 10160 3432 10194 3466
rect 10228 3432 10262 3466
rect 10296 3432 10330 3466
rect 10364 3432 10398 3466
rect 10432 3432 10466 3466
rect 10500 3432 10534 3466
rect 10568 3432 10602 3466
rect 10636 3432 10670 3466
rect 10704 3432 10738 3466
rect 10772 3432 10806 3466
rect 10840 3432 10874 3466
rect 10908 3432 10942 3466
rect 10976 3432 11010 3466
rect 11044 3432 11078 3466
rect 11112 3432 11146 3466
rect 11180 3432 11214 3466
rect 11248 3432 11282 3466
rect 11316 3432 11350 3466
rect 11384 3432 11418 3466
rect 11452 3432 11486 3466
rect 11520 3432 11554 3466
rect 11588 3432 11622 3466
rect 11656 3432 11690 3466
rect 11724 3432 11758 3466
rect 11792 3432 11826 3466
rect 11860 3432 11894 3466
rect 11928 3432 11962 3466
rect 11996 3432 12030 3466
rect 12064 3432 12098 3466
rect 12153 3449 12166 3466
rect 12227 3449 12234 3466
rect 12301 3449 12302 3466
rect 12132 3432 12166 3449
rect 12200 3432 12234 3449
rect 12268 3432 12302 3449
rect 12336 3449 12341 3466
rect 12404 3449 12415 3466
rect 12472 3449 12489 3466
rect 12540 3449 12563 3466
rect 12608 3449 12637 3466
rect 12336 3432 12370 3449
rect 12404 3432 12438 3449
rect 12472 3432 12506 3449
rect 12540 3432 12574 3449
rect 12608 3432 12642 3449
rect 12676 3432 12710 3466
rect 12745 3449 12778 3466
rect 12819 3449 12846 3466
rect 12893 3449 12914 3466
rect 12967 3449 12982 3466
rect 13040 3449 13050 3466
rect 13113 3449 13118 3466
rect 12744 3432 12778 3449
rect 12812 3432 12846 3449
rect 12880 3432 12914 3449
rect 12948 3432 12982 3449
rect 13016 3432 13050 3449
rect 13084 3432 13118 3449
rect 13186 3466 13225 3483
rect 13259 3466 13298 3483
rect 13332 3466 13371 3483
rect 13405 3466 13444 3483
rect 13478 3466 13517 3483
rect 13551 3466 13590 3483
rect 13624 3466 13663 3483
rect 13697 3466 13736 3483
rect 13770 3466 13809 3483
rect 13843 3466 13882 3483
rect 13916 3466 13955 3483
rect 13989 3466 14028 3483
rect 14062 3466 14101 3483
rect 14135 3466 14174 3483
rect 14208 3466 14247 3483
rect 14281 3466 14320 3483
rect 14354 3466 14393 3483
rect 14427 3466 14466 3483
rect 14500 3466 14539 3483
rect 14573 3466 14612 3483
rect 14646 3466 14685 3483
rect 14719 3466 14758 3483
rect 14792 3466 28000 3483
rect 13152 3432 13186 3449
rect 13220 3449 13225 3466
rect 13288 3449 13298 3466
rect 13356 3449 13371 3466
rect 13424 3449 13444 3466
rect 13492 3449 13517 3466
rect 13560 3449 13590 3466
rect 13220 3432 13254 3449
rect 13288 3432 13322 3449
rect 13356 3432 13390 3449
rect 13424 3432 13458 3449
rect 13492 3432 13526 3449
rect 13560 3432 13594 3449
rect 13628 3432 13662 3466
rect 13697 3449 13730 3466
rect 13770 3449 13798 3466
rect 13843 3449 13866 3466
rect 13916 3449 13934 3466
rect 13989 3449 14002 3466
rect 14062 3449 14070 3466
rect 14135 3449 14138 3466
rect 13696 3432 13730 3449
rect 13764 3432 13798 3449
rect 13832 3432 13866 3449
rect 13900 3432 13934 3449
rect 13968 3432 14002 3449
rect 14036 3432 14070 3449
rect 14104 3432 14138 3449
rect 14172 3449 14174 3466
rect 14240 3449 14247 3466
rect 14308 3449 14320 3466
rect 14376 3449 14393 3466
rect 14444 3449 14466 3466
rect 14512 3449 14539 3466
rect 14580 3449 14612 3466
rect 14172 3432 14206 3449
rect 14240 3432 14274 3449
rect 14308 3432 14342 3449
rect 14376 3432 14410 3449
rect 14444 3432 14478 3449
rect 14512 3432 14546 3449
rect 14580 3432 14614 3449
rect 14648 3432 14682 3466
rect 14719 3449 14750 3466
rect 14792 3449 14818 3466
rect 14716 3432 14750 3449
rect 14784 3432 14818 3449
rect 14852 3432 14886 3466
rect 14920 3432 14954 3466
rect 14988 3432 15022 3466
rect 15056 3432 15090 3466
rect 15124 3432 15158 3466
rect 15192 3432 15226 3466
rect 15260 3432 15294 3466
rect 15328 3432 15362 3466
rect 15396 3432 15430 3466
rect 15464 3432 15498 3466
rect 15532 3432 15566 3466
rect 15600 3432 15634 3466
rect 15668 3432 15702 3466
rect 15736 3432 15770 3466
rect 15804 3432 15838 3466
rect 15872 3432 15906 3466
rect 15940 3432 15974 3466
rect 16008 3432 16042 3466
rect 16076 3432 16110 3466
rect 16144 3432 16178 3466
rect 16212 3432 16246 3466
rect 16280 3432 16314 3466
rect 16348 3432 16382 3466
rect 16416 3432 16450 3466
rect 16484 3432 16518 3466
rect 16552 3432 16586 3466
rect 16620 3432 16654 3466
rect 16688 3432 16722 3466
rect 16756 3432 16790 3466
rect 16824 3432 16858 3466
rect 16892 3432 16926 3466
rect 16960 3432 16994 3466
rect 17028 3432 17062 3466
rect 17096 3432 17130 3466
rect 17164 3432 17198 3466
rect 17232 3432 17266 3466
rect 17300 3432 17334 3466
rect 17368 3432 17402 3466
rect 17436 3432 17470 3466
rect 17504 3432 17538 3466
rect 17572 3432 17606 3466
rect 17640 3432 17674 3466
rect 17708 3432 17742 3466
rect 17776 3432 17810 3466
rect 17844 3432 17878 3466
rect 17912 3432 17946 3466
rect 17980 3432 18014 3466
rect 18048 3432 18082 3466
rect 18116 3432 18150 3466
rect 18184 3432 18218 3466
rect 18252 3432 18286 3466
rect 18320 3432 18354 3466
rect 18388 3432 18422 3466
rect 18456 3432 18490 3466
rect 18524 3432 18558 3466
rect 18592 3432 18626 3466
rect 18660 3432 18694 3466
rect 18728 3432 18762 3466
rect 18796 3432 18830 3466
rect 18864 3432 18898 3466
rect 18932 3432 18966 3466
rect 19000 3432 19034 3466
rect 19068 3432 19102 3466
rect 19136 3432 19170 3466
rect 19204 3432 19238 3466
rect 19272 3432 19306 3466
rect 19340 3432 19374 3466
rect 19408 3432 19442 3466
rect 19476 3432 19510 3466
rect 19544 3432 19578 3466
rect 19612 3432 19646 3466
rect 19680 3432 19714 3466
rect 19748 3432 19782 3466
rect 19816 3432 19850 3466
rect 19884 3432 19918 3466
rect 19952 3432 19986 3466
rect 20020 3432 20054 3466
rect 20088 3432 20122 3466
rect 20156 3432 20190 3466
rect 20224 3432 20258 3466
rect 20292 3432 20326 3466
rect 20360 3432 20394 3466
rect 20428 3432 20462 3466
rect 20496 3432 20530 3466
rect 20564 3432 20598 3466
rect 20632 3432 20666 3466
rect 20700 3432 20734 3466
rect 20768 3432 20802 3466
rect 20836 3432 20870 3466
rect 20904 3432 20938 3466
rect 20972 3432 21006 3466
rect 21040 3432 21074 3466
rect 21108 3432 21142 3466
rect 21176 3432 21210 3466
rect 21244 3432 21278 3466
rect 21312 3432 21346 3466
rect 21380 3432 21414 3466
rect 21448 3432 21482 3466
rect 21516 3432 21550 3466
rect 21584 3432 21618 3466
rect 21652 3432 21686 3466
rect 21720 3432 21754 3466
rect 21788 3432 21822 3466
rect 21856 3432 21890 3466
rect 21924 3432 21958 3466
rect 21992 3432 22026 3466
rect 22060 3432 22094 3466
rect 22128 3432 22162 3466
rect 22196 3432 22230 3466
rect 22264 3432 22298 3466
rect 22332 3432 22366 3466
rect 22400 3432 22434 3466
rect 22468 3432 22502 3466
rect 22536 3432 22570 3466
rect 22604 3432 22638 3466
rect 22672 3432 22706 3466
rect 22740 3432 22774 3466
rect 22808 3432 22842 3466
rect 22876 3432 22910 3466
rect 22944 3432 22978 3466
rect 23012 3432 23046 3466
rect 23080 3432 23114 3466
rect 23148 3432 23182 3466
rect 23216 3432 23250 3466
rect 23284 3432 23318 3466
rect 23352 3432 23386 3466
rect 23420 3432 23454 3466
rect 23488 3432 23522 3466
rect 23556 3432 23590 3466
rect 23624 3432 23658 3466
rect 23692 3432 23726 3466
rect 23760 3432 23794 3466
rect 23828 3432 23862 3466
rect 23896 3432 23930 3466
rect 23964 3432 23998 3466
rect 24032 3432 24066 3466
rect 24100 3432 24134 3466
rect 24168 3432 24202 3466
rect 24236 3432 24270 3466
rect 24304 3432 24338 3466
rect 24372 3432 24406 3466
rect 24440 3432 24474 3466
rect 24508 3432 24542 3466
rect 24576 3432 24610 3466
rect 24644 3432 24678 3466
rect 24712 3432 24746 3466
rect 24780 3432 24814 3466
rect 24848 3432 24882 3466
rect 24916 3432 24950 3466
rect 24984 3432 25018 3466
rect 25052 3432 25086 3466
rect 25120 3432 25154 3466
rect 25188 3432 25222 3466
rect 25256 3432 25290 3466
rect 25324 3432 25358 3466
rect 25392 3432 25426 3466
rect 25460 3432 25494 3466
rect 25528 3432 25562 3466
rect 25596 3432 25630 3466
rect 25664 3432 25698 3466
rect 25732 3432 25766 3466
rect 25800 3432 25834 3466
rect 25868 3432 25902 3466
rect 25936 3432 25970 3466
rect 26004 3432 26038 3466
rect 26072 3432 26106 3466
rect 26140 3432 26174 3466
rect 26208 3432 26242 3466
rect 26276 3432 26310 3466
rect 26344 3432 26378 3466
rect 26412 3432 26446 3466
rect 26480 3432 26514 3466
rect 26548 3432 26582 3466
rect 26616 3432 26650 3466
rect 26684 3432 26718 3466
rect 26752 3432 26786 3466
rect 26820 3432 26854 3466
rect 26888 3432 26922 3466
rect 26956 3432 26990 3466
rect 27024 3432 27058 3466
rect 27092 3432 27126 3466
rect 27160 3432 27194 3466
rect 27228 3432 27262 3466
rect 27296 3432 27330 3466
rect 27364 3432 27398 3466
rect 27432 3432 27466 3466
rect 27500 3432 27534 3466
rect 27568 3432 27602 3466
rect 27636 3432 27670 3466
rect 27704 3432 27738 3466
rect 27772 3432 27806 3466
rect 27840 3432 27874 3466
rect 27908 3432 27942 3466
rect 27976 3432 28000 3466
rect 6449 3430 28000 3432
rect 3601 2043 3635 2081
<< viali >>
rect 27219 37566 27253 37600
rect 27292 37585 27321 37614
rect 27321 37585 27326 37614
rect 27365 37585 27389 37614
rect 27389 37585 27399 37614
rect 27439 37585 27457 37614
rect 27457 37585 27473 37614
rect 27513 37585 27525 37614
rect 27525 37585 27547 37614
rect 27292 37580 27326 37585
rect 27365 37580 27399 37585
rect 27439 37580 27473 37585
rect 27513 37580 27547 37585
rect 27363 37435 27397 37469
rect 27435 37435 27469 37469
rect 27219 37321 27253 37333
rect 27219 37299 27253 37321
rect 27585 37517 27619 37542
rect 27585 37508 27619 37517
rect 27585 37449 27619 37470
rect 27585 37436 27619 37449
rect 27585 37381 27619 37398
rect 27585 37364 27619 37381
rect 27585 37291 27619 37325
rect 27291 37219 27325 37253
rect 27365 37219 27381 37253
rect 27381 37219 27399 37253
rect 27439 37219 27449 37253
rect 27449 37219 27473 37253
rect 27512 37219 27517 37253
rect 27517 37219 27546 37253
rect 2256 34506 2290 34540
rect 2333 34506 2367 34540
rect 2410 34506 2444 34540
rect 2487 34506 2521 34540
rect 2564 34506 2598 34540
rect 2641 34506 2675 34540
rect 2718 34506 2752 34540
rect 2795 34506 2829 34540
rect 2872 34506 2906 34540
rect 2949 34506 2983 34540
rect 3026 34506 3060 34540
rect 3103 34506 3137 34540
rect 2256 34434 2290 34468
rect 2333 34434 2367 34468
rect 2410 34434 2444 34468
rect 2487 34434 2521 34468
rect 2564 34434 2598 34468
rect 2641 34434 2675 34468
rect 2718 34434 2752 34468
rect 2795 34434 2829 34468
rect 2872 34434 2906 34468
rect 2949 34434 2983 34468
rect 3026 34434 3060 34468
rect 3103 34434 3137 34468
rect 2256 34362 2290 34396
rect 2333 34362 2367 34396
rect 2410 34362 2444 34396
rect 2487 34362 2521 34396
rect 2564 34362 2598 34396
rect 2641 34362 2675 34396
rect 2718 34362 2752 34396
rect 2795 34362 2829 34396
rect 2872 34362 2906 34396
rect 2949 34362 2983 34396
rect 3026 34362 3060 34396
rect 3103 34362 3137 34396
rect 2279 32543 2601 32649
rect 2783 32543 3105 32649
rect 23806 23283 23840 23284
rect 23879 23283 23913 23284
rect 23952 23283 23986 23284
rect 24025 23283 24059 23284
rect 24098 23283 24132 23284
rect 24171 23283 24205 23284
rect 24244 23283 24278 23284
rect 24317 23283 24351 23284
rect 24390 23283 24424 23284
rect 24462 23283 24496 23284
rect 24534 23283 24568 23284
rect 24606 23283 24640 23284
rect 23806 23250 23816 23283
rect 23816 23250 23840 23283
rect 23879 23250 23885 23283
rect 23885 23250 23913 23283
rect 23952 23250 23954 23283
rect 23954 23250 23986 23283
rect 24025 23250 24057 23283
rect 24057 23250 24059 23283
rect 24098 23250 24126 23283
rect 24126 23250 24132 23283
rect 24171 23250 24195 23283
rect 24195 23250 24205 23283
rect 24244 23250 24264 23283
rect 24264 23250 24278 23283
rect 24317 23250 24333 23283
rect 24333 23250 24351 23283
rect 24390 23250 24402 23283
rect 24402 23250 24424 23283
rect 24462 23250 24471 23283
rect 24471 23250 24496 23283
rect 24534 23250 24540 23283
rect 24540 23250 24568 23283
rect 24606 23250 24609 23283
rect 24609 23250 24640 23283
rect 24678 23250 24712 23284
rect 24750 23283 24784 23284
rect 24822 23283 24856 23284
rect 24894 23283 24928 23284
rect 24966 23283 25000 23284
rect 25038 23283 25072 23284
rect 25110 23283 25144 23284
rect 25182 23283 25216 23284
rect 25254 23283 25288 23284
rect 25326 23283 25360 23284
rect 25398 23283 25432 23284
rect 25470 23283 25504 23284
rect 25542 23283 25576 23284
rect 25614 23283 25648 23284
rect 25686 23283 25720 23284
rect 25758 23283 25792 23284
rect 25830 23283 25864 23284
rect 25902 23283 25936 23284
rect 25974 23283 26008 23284
rect 26046 23283 26080 23284
rect 26118 23283 26152 23284
rect 26190 23283 26224 23284
rect 26262 23283 26296 23284
rect 24750 23250 24782 23283
rect 24782 23250 24784 23283
rect 24822 23250 24851 23283
rect 24851 23250 24856 23283
rect 24894 23250 24920 23283
rect 24920 23250 24928 23283
rect 24966 23250 24989 23283
rect 24989 23250 25000 23283
rect 25038 23250 25058 23283
rect 25058 23250 25072 23283
rect 25110 23250 25127 23283
rect 25127 23250 25144 23283
rect 25182 23250 25196 23283
rect 25196 23250 25216 23283
rect 25254 23250 25265 23283
rect 25265 23250 25288 23283
rect 25326 23250 25334 23283
rect 25334 23250 25360 23283
rect 25398 23250 25403 23283
rect 25403 23250 25432 23283
rect 25470 23250 25472 23283
rect 25472 23250 25504 23283
rect 25542 23250 25575 23283
rect 25575 23250 25576 23283
rect 25614 23250 25644 23283
rect 25644 23250 25648 23283
rect 25686 23250 25713 23283
rect 25713 23250 25720 23283
rect 25758 23250 25782 23283
rect 25782 23250 25792 23283
rect 25830 23250 25851 23283
rect 25851 23250 25864 23283
rect 25902 23250 25920 23283
rect 25920 23250 25936 23283
rect 25974 23250 25989 23283
rect 25989 23250 26008 23283
rect 26046 23250 26058 23283
rect 26058 23250 26080 23283
rect 26118 23250 26127 23283
rect 26127 23250 26152 23283
rect 26190 23250 26196 23283
rect 26196 23250 26224 23283
rect 26262 23250 26265 23283
rect 26265 23250 26296 23283
rect 26334 23250 26368 23284
rect 26406 23283 26440 23284
rect 26478 23283 26512 23284
rect 26550 23283 26584 23284
rect 26622 23283 26656 23284
rect 26694 23283 26728 23284
rect 26766 23283 26800 23284
rect 26838 23283 26872 23284
rect 26910 23283 26944 23284
rect 26982 23283 27016 23284
rect 27054 23283 27088 23284
rect 27126 23283 27160 23284
rect 27198 23283 27232 23284
rect 27270 23283 27304 23284
rect 27342 23283 27376 23284
rect 27414 23283 27448 23284
rect 27486 23283 27520 23284
rect 26406 23250 26436 23283
rect 26436 23250 26440 23283
rect 26478 23250 26504 23283
rect 26504 23250 26512 23283
rect 26550 23250 26572 23283
rect 26572 23250 26584 23283
rect 26622 23250 26640 23283
rect 26640 23250 26656 23283
rect 26694 23250 26708 23283
rect 26708 23250 26728 23283
rect 26766 23250 26776 23283
rect 26776 23250 26800 23283
rect 26838 23250 26844 23283
rect 26844 23250 26872 23283
rect 26910 23250 26912 23283
rect 26912 23250 26944 23283
rect 26982 23250 27014 23283
rect 27014 23250 27016 23283
rect 27054 23250 27082 23283
rect 27082 23250 27088 23283
rect 27126 23250 27150 23283
rect 27150 23250 27160 23283
rect 27198 23250 27218 23283
rect 27218 23250 27232 23283
rect 27270 23250 27286 23283
rect 27286 23250 27304 23283
rect 27342 23250 27354 23283
rect 27354 23250 27376 23283
rect 27414 23250 27422 23283
rect 27422 23250 27448 23283
rect 27486 23250 27490 23283
rect 27490 23250 27520 23283
rect 27558 23250 27592 23284
rect 27630 23283 27664 23284
rect 27702 23283 27736 23284
rect 27774 23283 27808 23284
rect 27846 23283 27880 23284
rect 27918 23283 27952 23284
rect 27630 23250 27660 23283
rect 27660 23250 27664 23283
rect 27702 23250 27728 23283
rect 27728 23250 27736 23283
rect 27774 23250 27796 23283
rect 27796 23250 27808 23283
rect 27846 23250 27864 23283
rect 27864 23250 27880 23283
rect 27918 23250 27932 23283
rect 27932 23250 27952 23283
rect 23806 23179 23816 23198
rect 23816 23179 23840 23198
rect 23879 23179 23885 23198
rect 23885 23179 23913 23198
rect 23952 23179 23954 23198
rect 23954 23179 23986 23198
rect 24025 23179 24057 23198
rect 24057 23179 24059 23198
rect 24098 23179 24126 23198
rect 24126 23179 24132 23198
rect 24171 23179 24195 23198
rect 24195 23179 24205 23198
rect 24244 23179 24264 23198
rect 24264 23179 24278 23198
rect 24317 23179 24333 23198
rect 24333 23179 24351 23198
rect 24390 23179 24402 23198
rect 24402 23179 24424 23198
rect 24462 23179 24471 23198
rect 24471 23179 24496 23198
rect 24534 23179 24540 23198
rect 24540 23179 24568 23198
rect 24606 23179 24609 23198
rect 24609 23179 24640 23198
rect 23806 23164 23840 23179
rect 23879 23164 23913 23179
rect 23952 23164 23986 23179
rect 24025 23164 24059 23179
rect 24098 23164 24132 23179
rect 24171 23164 24205 23179
rect 24244 23164 24278 23179
rect 24317 23164 24351 23179
rect 24390 23164 24424 23179
rect 24462 23164 24496 23179
rect 24534 23164 24568 23179
rect 24606 23164 24640 23179
rect 24678 23164 24712 23198
rect 24750 23179 24782 23198
rect 24782 23179 24784 23198
rect 24822 23179 24851 23198
rect 24851 23179 24856 23198
rect 24894 23179 24920 23198
rect 24920 23179 24928 23198
rect 24966 23179 24989 23198
rect 24989 23179 25000 23198
rect 25038 23179 25058 23198
rect 25058 23179 25072 23198
rect 25110 23179 25127 23198
rect 25127 23179 25144 23198
rect 25182 23179 25196 23198
rect 25196 23179 25216 23198
rect 25254 23179 25265 23198
rect 25265 23179 25288 23198
rect 25326 23179 25334 23198
rect 25334 23179 25360 23198
rect 25398 23179 25403 23198
rect 25403 23179 25432 23198
rect 25470 23179 25472 23198
rect 25472 23179 25504 23198
rect 25542 23179 25575 23198
rect 25575 23179 25576 23198
rect 25614 23179 25644 23198
rect 25644 23179 25648 23198
rect 25686 23179 25713 23198
rect 25713 23179 25720 23198
rect 25758 23179 25782 23198
rect 25782 23179 25792 23198
rect 25830 23179 25851 23198
rect 25851 23179 25864 23198
rect 25902 23179 25920 23198
rect 25920 23179 25936 23198
rect 25974 23179 25989 23198
rect 25989 23179 26008 23198
rect 26046 23179 26058 23198
rect 26058 23179 26080 23198
rect 26118 23179 26127 23198
rect 26127 23179 26152 23198
rect 26190 23179 26196 23198
rect 26196 23179 26224 23198
rect 26262 23179 26265 23198
rect 26265 23179 26296 23198
rect 24750 23164 24784 23179
rect 24822 23164 24856 23179
rect 24894 23164 24928 23179
rect 24966 23164 25000 23179
rect 25038 23164 25072 23179
rect 25110 23164 25144 23179
rect 25182 23164 25216 23179
rect 25254 23164 25288 23179
rect 25326 23164 25360 23179
rect 25398 23164 25432 23179
rect 25470 23164 25504 23179
rect 25542 23164 25576 23179
rect 25614 23164 25648 23179
rect 25686 23164 25720 23179
rect 25758 23164 25792 23179
rect 25830 23164 25864 23179
rect 25902 23164 25936 23179
rect 25974 23164 26008 23179
rect 26046 23164 26080 23179
rect 26118 23164 26152 23179
rect 26190 23164 26224 23179
rect 26262 23164 26296 23179
rect 26334 23164 26368 23198
rect 26406 23179 26436 23198
rect 26436 23179 26440 23198
rect 26478 23179 26504 23198
rect 26504 23179 26512 23198
rect 26550 23179 26572 23198
rect 26572 23179 26584 23198
rect 26622 23179 26640 23198
rect 26640 23179 26656 23198
rect 26694 23179 26708 23198
rect 26708 23179 26728 23198
rect 26766 23179 26776 23198
rect 26776 23179 26800 23198
rect 26838 23179 26844 23198
rect 26844 23179 26872 23198
rect 26910 23179 26912 23198
rect 26912 23179 26944 23198
rect 26982 23179 27014 23198
rect 27014 23179 27016 23198
rect 27054 23179 27082 23198
rect 27082 23179 27088 23198
rect 27126 23179 27150 23198
rect 27150 23179 27160 23198
rect 27198 23179 27218 23198
rect 27218 23179 27232 23198
rect 27270 23179 27286 23198
rect 27286 23179 27304 23198
rect 27342 23179 27354 23198
rect 27354 23179 27376 23198
rect 27414 23179 27422 23198
rect 27422 23179 27448 23198
rect 27486 23179 27490 23198
rect 27490 23179 27520 23198
rect 26406 23164 26440 23179
rect 26478 23164 26512 23179
rect 26550 23164 26584 23179
rect 26622 23164 26656 23179
rect 26694 23164 26728 23179
rect 26766 23164 26800 23179
rect 26838 23164 26872 23179
rect 26910 23164 26944 23179
rect 26982 23164 27016 23179
rect 27054 23164 27088 23179
rect 27126 23164 27160 23179
rect 27198 23164 27232 23179
rect 27270 23164 27304 23179
rect 27342 23164 27376 23179
rect 27414 23164 27448 23179
rect 27486 23164 27520 23179
rect 27558 23164 27592 23198
rect 27630 23179 27660 23198
rect 27660 23179 27664 23198
rect 27702 23179 27728 23198
rect 27728 23179 27736 23198
rect 27774 23179 27796 23198
rect 27796 23179 27808 23198
rect 27846 23179 27864 23198
rect 27864 23179 27880 23198
rect 27918 23179 27932 23198
rect 27932 23179 27952 23198
rect 27630 23164 27664 23179
rect 27702 23164 27736 23179
rect 27774 23164 27808 23179
rect 27846 23164 27880 23179
rect 27918 23164 27952 23179
rect 23806 23109 23816 23112
rect 23816 23109 23840 23112
rect 23879 23109 23885 23112
rect 23885 23109 23913 23112
rect 23952 23109 23954 23112
rect 23954 23109 23986 23112
rect 24025 23109 24057 23112
rect 24057 23109 24059 23112
rect 24098 23109 24126 23112
rect 24126 23109 24132 23112
rect 24171 23109 24195 23112
rect 24195 23109 24205 23112
rect 24244 23109 24264 23112
rect 24264 23109 24278 23112
rect 24317 23109 24333 23112
rect 24333 23109 24351 23112
rect 24390 23109 24402 23112
rect 24402 23109 24424 23112
rect 24462 23109 24471 23112
rect 24471 23109 24496 23112
rect 24534 23109 24540 23112
rect 24540 23109 24568 23112
rect 24606 23109 24609 23112
rect 24609 23109 24640 23112
rect 23806 23078 23840 23109
rect 23879 23078 23913 23109
rect 23952 23078 23986 23109
rect 24025 23078 24059 23109
rect 24098 23078 24132 23109
rect 24171 23078 24205 23109
rect 24244 23078 24278 23109
rect 24317 23078 24351 23109
rect 24390 23078 24424 23109
rect 24462 23078 24496 23109
rect 24534 23078 24568 23109
rect 24606 23078 24640 23109
rect 24678 23078 24712 23112
rect 24750 23109 24782 23112
rect 24782 23109 24784 23112
rect 24822 23109 24851 23112
rect 24851 23109 24856 23112
rect 24894 23109 24920 23112
rect 24920 23109 24928 23112
rect 24966 23109 24989 23112
rect 24989 23109 25000 23112
rect 25038 23109 25058 23112
rect 25058 23109 25072 23112
rect 25110 23109 25127 23112
rect 25127 23109 25144 23112
rect 25182 23109 25196 23112
rect 25196 23109 25216 23112
rect 25254 23109 25265 23112
rect 25265 23109 25288 23112
rect 25326 23109 25334 23112
rect 25334 23109 25360 23112
rect 25398 23109 25403 23112
rect 25403 23109 25432 23112
rect 25470 23109 25472 23112
rect 25472 23109 25504 23112
rect 25542 23109 25575 23112
rect 25575 23109 25576 23112
rect 25614 23109 25644 23112
rect 25644 23109 25648 23112
rect 25686 23109 25713 23112
rect 25713 23109 25720 23112
rect 25758 23109 25782 23112
rect 25782 23109 25792 23112
rect 25830 23109 25851 23112
rect 25851 23109 25864 23112
rect 25902 23109 25920 23112
rect 25920 23109 25936 23112
rect 25974 23109 25989 23112
rect 25989 23109 26008 23112
rect 26046 23109 26058 23112
rect 26058 23109 26080 23112
rect 26118 23109 26127 23112
rect 26127 23109 26152 23112
rect 26190 23109 26196 23112
rect 26196 23109 26224 23112
rect 26262 23109 26265 23112
rect 26265 23109 26296 23112
rect 24750 23078 24784 23109
rect 24822 23078 24856 23109
rect 24894 23078 24928 23109
rect 24966 23078 25000 23109
rect 25038 23078 25072 23109
rect 25110 23078 25144 23109
rect 25182 23078 25216 23109
rect 25254 23078 25288 23109
rect 25326 23078 25360 23109
rect 25398 23078 25432 23109
rect 25470 23078 25504 23109
rect 25542 23078 25576 23109
rect 25614 23078 25648 23109
rect 25686 23078 25720 23109
rect 25758 23078 25792 23109
rect 25830 23078 25864 23109
rect 25902 23078 25936 23109
rect 25974 23078 26008 23109
rect 26046 23078 26080 23109
rect 26118 23078 26152 23109
rect 26190 23078 26224 23109
rect 26262 23078 26296 23109
rect 26334 23078 26368 23112
rect 26406 23109 26436 23112
rect 26436 23109 26440 23112
rect 26478 23109 26504 23112
rect 26504 23109 26512 23112
rect 26550 23109 26572 23112
rect 26572 23109 26584 23112
rect 26622 23109 26640 23112
rect 26640 23109 26656 23112
rect 26694 23109 26708 23112
rect 26708 23109 26728 23112
rect 26766 23109 26776 23112
rect 26776 23109 26800 23112
rect 26838 23109 26844 23112
rect 26844 23109 26872 23112
rect 26910 23109 26912 23112
rect 26912 23109 26944 23112
rect 26982 23109 27014 23112
rect 27014 23109 27016 23112
rect 27054 23109 27082 23112
rect 27082 23109 27088 23112
rect 27126 23109 27150 23112
rect 27150 23109 27160 23112
rect 27198 23109 27218 23112
rect 27218 23109 27232 23112
rect 27270 23109 27286 23112
rect 27286 23109 27304 23112
rect 27342 23109 27354 23112
rect 27354 23109 27376 23112
rect 27414 23109 27422 23112
rect 27422 23109 27448 23112
rect 27486 23109 27490 23112
rect 27490 23109 27520 23112
rect 26406 23078 26440 23109
rect 26478 23078 26512 23109
rect 26550 23078 26584 23109
rect 26622 23078 26656 23109
rect 26694 23078 26728 23109
rect 26766 23078 26800 23109
rect 26838 23078 26872 23109
rect 26910 23078 26944 23109
rect 26982 23078 27016 23109
rect 27054 23078 27088 23109
rect 27126 23078 27160 23109
rect 27198 23078 27232 23109
rect 27270 23078 27304 23109
rect 27342 23078 27376 23109
rect 27414 23078 27448 23109
rect 27486 23078 27520 23109
rect 27558 23078 27592 23112
rect 27630 23109 27660 23112
rect 27660 23109 27664 23112
rect 27702 23109 27728 23112
rect 27728 23109 27736 23112
rect 27774 23109 27796 23112
rect 27796 23109 27808 23112
rect 27846 23109 27864 23112
rect 27864 23109 27880 23112
rect 27918 23109 27932 23112
rect 27932 23109 27952 23112
rect 27630 23078 27664 23109
rect 27702 23078 27736 23109
rect 27774 23078 27808 23109
rect 27846 23078 27880 23109
rect 27918 23078 27952 23109
rect 23806 23003 23840 23026
rect 23879 23003 23913 23026
rect 23952 23003 23986 23026
rect 24025 23003 24059 23026
rect 24098 23003 24132 23026
rect 24171 23003 24205 23026
rect 24244 23003 24278 23026
rect 24317 23003 24351 23026
rect 24390 23003 24424 23026
rect 24462 23003 24496 23026
rect 24534 23003 24568 23026
rect 24606 23003 24640 23026
rect 23806 22992 23816 23003
rect 23816 22992 23840 23003
rect 23879 22992 23885 23003
rect 23885 22992 23913 23003
rect 23952 22992 23954 23003
rect 23954 22992 23986 23003
rect 24025 22992 24057 23003
rect 24057 22992 24059 23003
rect 24098 22992 24126 23003
rect 24126 22992 24132 23003
rect 24171 22992 24195 23003
rect 24195 22992 24205 23003
rect 24244 22992 24264 23003
rect 24264 22992 24278 23003
rect 24317 22992 24333 23003
rect 24333 22992 24351 23003
rect 24390 22992 24402 23003
rect 24402 22992 24424 23003
rect 24462 22992 24471 23003
rect 24471 22992 24496 23003
rect 24534 22992 24540 23003
rect 24540 22992 24568 23003
rect 24606 22992 24609 23003
rect 24609 22992 24640 23003
rect 24678 22992 24712 23026
rect 24750 23003 24784 23026
rect 24822 23003 24856 23026
rect 24894 23003 24928 23026
rect 24966 23003 25000 23026
rect 25038 23003 25072 23026
rect 25110 23003 25144 23026
rect 25182 23003 25216 23026
rect 25254 23003 25288 23026
rect 25326 23003 25360 23026
rect 25398 23003 25432 23026
rect 25470 23003 25504 23026
rect 25542 23003 25576 23026
rect 25614 23003 25648 23026
rect 25686 23003 25720 23026
rect 25758 23003 25792 23026
rect 25830 23003 25864 23026
rect 25902 23003 25936 23026
rect 25974 23003 26008 23026
rect 26046 23003 26080 23026
rect 26118 23003 26152 23026
rect 26190 23003 26224 23026
rect 26262 23003 26296 23026
rect 24750 22992 24782 23003
rect 24782 22992 24784 23003
rect 24822 22992 24851 23003
rect 24851 22992 24856 23003
rect 24894 22992 24920 23003
rect 24920 22992 24928 23003
rect 24966 22992 24989 23003
rect 24989 22992 25000 23003
rect 25038 22992 25058 23003
rect 25058 22992 25072 23003
rect 25110 22992 25127 23003
rect 25127 22992 25144 23003
rect 25182 22992 25196 23003
rect 25196 22992 25216 23003
rect 25254 22992 25265 23003
rect 25265 22992 25288 23003
rect 25326 22992 25334 23003
rect 25334 22992 25360 23003
rect 25398 22992 25403 23003
rect 25403 22992 25432 23003
rect 25470 22992 25472 23003
rect 25472 22992 25504 23003
rect 25542 22992 25575 23003
rect 25575 22992 25576 23003
rect 25614 22992 25644 23003
rect 25644 22992 25648 23003
rect 25686 22992 25713 23003
rect 25713 22992 25720 23003
rect 25758 22992 25782 23003
rect 25782 22992 25792 23003
rect 25830 22992 25851 23003
rect 25851 22992 25864 23003
rect 25902 22992 25920 23003
rect 25920 22992 25936 23003
rect 25974 22992 25989 23003
rect 25989 22992 26008 23003
rect 26046 22992 26058 23003
rect 26058 22992 26080 23003
rect 26118 22992 26127 23003
rect 26127 22992 26152 23003
rect 26190 22992 26196 23003
rect 26196 22992 26224 23003
rect 26262 22992 26265 23003
rect 26265 22992 26296 23003
rect 26334 22992 26368 23026
rect 26406 23003 26440 23026
rect 26478 23003 26512 23026
rect 26550 23003 26584 23026
rect 26622 23003 26656 23026
rect 26694 23003 26728 23026
rect 26766 23003 26800 23026
rect 26838 23003 26872 23026
rect 26910 23003 26944 23026
rect 26982 23003 27016 23026
rect 27054 23003 27088 23026
rect 27126 23003 27160 23026
rect 27198 23003 27232 23026
rect 27270 23003 27304 23026
rect 27342 23003 27376 23026
rect 27414 23003 27448 23026
rect 27486 23003 27520 23026
rect 26406 22992 26436 23003
rect 26436 22992 26440 23003
rect 26478 22992 26504 23003
rect 26504 22992 26512 23003
rect 26550 22992 26572 23003
rect 26572 22992 26584 23003
rect 26622 22992 26640 23003
rect 26640 22992 26656 23003
rect 26694 22992 26708 23003
rect 26708 22992 26728 23003
rect 26766 22992 26776 23003
rect 26776 22992 26800 23003
rect 26838 22992 26844 23003
rect 26844 22992 26872 23003
rect 26910 22992 26912 23003
rect 26912 22992 26944 23003
rect 26982 22992 27014 23003
rect 27014 22992 27016 23003
rect 27054 22992 27082 23003
rect 27082 22992 27088 23003
rect 27126 22992 27150 23003
rect 27150 22992 27160 23003
rect 27198 22992 27218 23003
rect 27218 22992 27232 23003
rect 27270 22992 27286 23003
rect 27286 22992 27304 23003
rect 27342 22992 27354 23003
rect 27354 22992 27376 23003
rect 27414 22992 27422 23003
rect 27422 22992 27448 23003
rect 27486 22992 27490 23003
rect 27490 22992 27520 23003
rect 27558 22992 27592 23026
rect 27630 23003 27664 23026
rect 27702 23003 27736 23026
rect 27774 23003 27808 23026
rect 27846 23003 27880 23026
rect 27918 23003 27952 23026
rect 27630 22992 27660 23003
rect 27660 22992 27664 23003
rect 27702 22992 27728 23003
rect 27728 22992 27736 23003
rect 27774 22992 27796 23003
rect 27796 22992 27808 23003
rect 27846 22992 27864 23003
rect 27864 22992 27880 23003
rect 27918 22992 27932 23003
rect 27932 22992 27952 23003
rect 26434 22856 26468 22890
rect 26509 22856 26543 22890
rect 26584 22856 26618 22890
rect 26659 22856 26693 22890
rect 26734 22856 26768 22890
rect 26808 22856 26842 22890
rect 26882 22856 26916 22890
rect 26956 22856 26990 22890
rect 27030 22856 27064 22890
rect 27104 22856 27138 22890
rect 27178 22856 27212 22890
rect 27252 22856 27286 22890
rect 27326 22856 27360 22890
rect 27400 22856 27434 22890
rect 27474 22856 27508 22890
rect 27548 22856 27582 22890
rect 27622 22856 27656 22890
rect 27696 22856 27730 22890
rect 27770 22856 27804 22890
rect 27844 22856 27878 22890
rect 27918 22856 27952 22890
rect 26434 22784 26468 22818
rect 26509 22784 26543 22818
rect 26584 22784 26618 22818
rect 26659 22784 26693 22818
rect 26734 22784 26768 22818
rect 26808 22784 26842 22818
rect 26882 22784 26916 22818
rect 26956 22784 26990 22818
rect 27030 22784 27064 22818
rect 27104 22784 27138 22818
rect 27178 22784 27212 22818
rect 27252 22784 27286 22818
rect 27326 22784 27360 22818
rect 27400 22784 27434 22818
rect 27474 22784 27508 22818
rect 27548 22784 27582 22818
rect 27622 22784 27656 22818
rect 27696 22784 27730 22818
rect 27770 22784 27804 22818
rect 27844 22784 27878 22818
rect 27918 22784 27952 22818
rect 26434 22712 26468 22746
rect 26509 22712 26543 22746
rect 26584 22712 26618 22746
rect 26659 22712 26693 22746
rect 26734 22712 26768 22746
rect 26808 22712 26842 22746
rect 26882 22712 26916 22746
rect 26956 22712 26990 22746
rect 27030 22712 27064 22746
rect 27104 22712 27138 22746
rect 27178 22712 27212 22746
rect 27252 22712 27286 22746
rect 27326 22712 27360 22746
rect 27400 22712 27434 22746
rect 27474 22712 27508 22746
rect 27548 22712 27582 22746
rect 27622 22712 27656 22746
rect 27696 22712 27730 22746
rect 27770 22712 27804 22746
rect 27844 22712 27878 22746
rect 27918 22712 27952 22746
rect 26434 22640 26468 22674
rect 26509 22640 26543 22674
rect 26584 22640 26618 22674
rect 26659 22640 26693 22674
rect 26734 22640 26768 22674
rect 26808 22640 26842 22674
rect 26882 22640 26916 22674
rect 26956 22640 26990 22674
rect 27030 22640 27064 22674
rect 27104 22640 27138 22674
rect 27178 22640 27212 22674
rect 27252 22640 27286 22674
rect 27326 22640 27360 22674
rect 27400 22640 27434 22674
rect 27474 22640 27508 22674
rect 27548 22640 27582 22674
rect 27622 22640 27656 22674
rect 27696 22640 27730 22674
rect 27770 22640 27804 22674
rect 27844 22640 27878 22674
rect 27918 22640 27952 22674
rect 26434 22600 26451 22602
rect 26451 22600 26468 22602
rect 26509 22600 26522 22602
rect 26522 22600 26543 22602
rect 26584 22600 26593 22602
rect 26593 22600 26618 22602
rect 26659 22600 26664 22602
rect 26664 22600 26693 22602
rect 26734 22600 26735 22602
rect 26735 22600 26768 22602
rect 26808 22600 26840 22602
rect 26840 22600 26842 22602
rect 26882 22600 26911 22602
rect 26911 22600 26916 22602
rect 26956 22600 26982 22602
rect 26982 22600 26990 22602
rect 27030 22600 27053 22602
rect 27053 22600 27064 22602
rect 27104 22600 27124 22602
rect 27124 22600 27138 22602
rect 27178 22600 27195 22602
rect 27195 22600 27212 22602
rect 27252 22600 27266 22602
rect 27266 22600 27286 22602
rect 27326 22600 27336 22602
rect 27336 22600 27360 22602
rect 27400 22600 27406 22602
rect 27406 22600 27434 22602
rect 27474 22600 27476 22602
rect 27476 22600 27508 22602
rect 26434 22568 26468 22600
rect 26509 22568 26543 22600
rect 26584 22568 26618 22600
rect 26659 22568 26693 22600
rect 26734 22568 26768 22600
rect 26808 22568 26842 22600
rect 26882 22568 26916 22600
rect 26956 22568 26990 22600
rect 27030 22568 27064 22600
rect 27104 22568 27138 22600
rect 27178 22568 27212 22600
rect 27252 22568 27286 22600
rect 27326 22568 27360 22600
rect 27400 22568 27434 22600
rect 27474 22568 27508 22600
rect 27548 22568 27582 22602
rect 27622 22600 27652 22602
rect 27652 22600 27656 22602
rect 27696 22600 27722 22602
rect 27722 22600 27730 22602
rect 27770 22600 27792 22602
rect 27792 22600 27804 22602
rect 27844 22600 27862 22602
rect 27862 22600 27878 22602
rect 27918 22600 27932 22602
rect 27932 22600 27952 22602
rect 27622 22568 27656 22600
rect 27696 22568 27730 22600
rect 27770 22568 27804 22600
rect 27844 22568 27878 22600
rect 27918 22568 27952 22600
rect 26434 22526 26451 22530
rect 26451 22526 26468 22530
rect 26509 22526 26522 22530
rect 26522 22526 26543 22530
rect 26584 22526 26593 22530
rect 26593 22526 26618 22530
rect 26659 22526 26664 22530
rect 26664 22526 26693 22530
rect 26734 22526 26735 22530
rect 26735 22526 26768 22530
rect 26808 22526 26840 22530
rect 26840 22526 26842 22530
rect 26882 22526 26911 22530
rect 26911 22526 26916 22530
rect 26956 22526 26982 22530
rect 26982 22526 26990 22530
rect 27030 22526 27053 22530
rect 27053 22526 27064 22530
rect 27104 22526 27124 22530
rect 27124 22526 27138 22530
rect 27178 22526 27195 22530
rect 27195 22526 27212 22530
rect 27252 22526 27266 22530
rect 27266 22526 27286 22530
rect 27326 22526 27336 22530
rect 27336 22526 27360 22530
rect 27400 22526 27406 22530
rect 27406 22526 27434 22530
rect 27474 22526 27476 22530
rect 27476 22526 27508 22530
rect 26434 22496 26468 22526
rect 26509 22496 26543 22526
rect 26584 22496 26618 22526
rect 26659 22496 26693 22526
rect 26734 22496 26768 22526
rect 26808 22496 26842 22526
rect 26882 22496 26916 22526
rect 26956 22496 26990 22526
rect 27030 22496 27064 22526
rect 27104 22496 27138 22526
rect 27178 22496 27212 22526
rect 27252 22496 27286 22526
rect 27326 22496 27360 22526
rect 27400 22496 27434 22526
rect 27474 22496 27508 22526
rect 27548 22496 27582 22530
rect 27622 22526 27652 22530
rect 27652 22526 27656 22530
rect 27696 22526 27722 22530
rect 27722 22526 27730 22530
rect 27770 22526 27792 22530
rect 27792 22526 27804 22530
rect 27844 22526 27862 22530
rect 27862 22526 27878 22530
rect 27918 22526 27932 22530
rect 27932 22526 27952 22530
rect 27622 22496 27656 22526
rect 27696 22496 27730 22526
rect 27770 22496 27804 22526
rect 27844 22496 27878 22526
rect 27918 22496 27952 22526
rect 26434 22452 26451 22458
rect 26451 22452 26468 22458
rect 26509 22452 26522 22458
rect 26522 22452 26543 22458
rect 26584 22452 26593 22458
rect 26593 22452 26618 22458
rect 26659 22452 26664 22458
rect 26664 22452 26693 22458
rect 26734 22452 26735 22458
rect 26735 22452 26768 22458
rect 26808 22452 26840 22458
rect 26840 22452 26842 22458
rect 26882 22452 26911 22458
rect 26911 22452 26916 22458
rect 26956 22452 26982 22458
rect 26982 22452 26990 22458
rect 27030 22452 27053 22458
rect 27053 22452 27064 22458
rect 27104 22452 27124 22458
rect 27124 22452 27138 22458
rect 27178 22452 27195 22458
rect 27195 22452 27212 22458
rect 27252 22452 27266 22458
rect 27266 22452 27286 22458
rect 27326 22452 27336 22458
rect 27336 22452 27360 22458
rect 27400 22452 27406 22458
rect 27406 22452 27434 22458
rect 27474 22452 27476 22458
rect 27476 22452 27508 22458
rect 26434 22424 26468 22452
rect 26509 22424 26543 22452
rect 26584 22424 26618 22452
rect 26659 22424 26693 22452
rect 26734 22424 26768 22452
rect 26808 22424 26842 22452
rect 26882 22424 26916 22452
rect 26956 22424 26990 22452
rect 27030 22424 27064 22452
rect 27104 22424 27138 22452
rect 27178 22424 27212 22452
rect 27252 22424 27286 22452
rect 27326 22424 27360 22452
rect 27400 22424 27434 22452
rect 27474 22424 27508 22452
rect 27548 22424 27582 22458
rect 27622 22452 27652 22458
rect 27652 22452 27656 22458
rect 27696 22452 27722 22458
rect 27722 22452 27730 22458
rect 27770 22452 27792 22458
rect 27792 22452 27804 22458
rect 27844 22452 27862 22458
rect 27862 22452 27878 22458
rect 27918 22452 27932 22458
rect 27932 22452 27952 22458
rect 27622 22424 27656 22452
rect 27696 22424 27730 22452
rect 27770 22424 27804 22452
rect 27844 22424 27878 22452
rect 27918 22424 27952 22452
rect 26434 22378 26451 22386
rect 26451 22378 26468 22386
rect 26509 22378 26522 22386
rect 26522 22378 26543 22386
rect 26584 22378 26593 22386
rect 26593 22378 26618 22386
rect 26659 22378 26664 22386
rect 26664 22378 26693 22386
rect 26734 22378 26735 22386
rect 26735 22378 26768 22386
rect 26808 22378 26840 22386
rect 26840 22378 26842 22386
rect 26882 22378 26911 22386
rect 26911 22378 26916 22386
rect 26956 22378 26982 22386
rect 26982 22378 26990 22386
rect 27030 22378 27053 22386
rect 27053 22378 27064 22386
rect 27104 22378 27124 22386
rect 27124 22378 27138 22386
rect 27178 22378 27195 22386
rect 27195 22378 27212 22386
rect 27252 22378 27266 22386
rect 27266 22378 27286 22386
rect 27326 22378 27336 22386
rect 27336 22378 27360 22386
rect 27400 22378 27406 22386
rect 27406 22378 27434 22386
rect 27474 22378 27476 22386
rect 27476 22378 27508 22386
rect 26434 22352 26468 22378
rect 26509 22352 26543 22378
rect 26584 22352 26618 22378
rect 26659 22352 26693 22378
rect 26734 22352 26768 22378
rect 26808 22352 26842 22378
rect 26882 22352 26916 22378
rect 26956 22352 26990 22378
rect 27030 22352 27064 22378
rect 27104 22352 27138 22378
rect 27178 22352 27212 22378
rect 27252 22352 27286 22378
rect 27326 22352 27360 22378
rect 27400 22352 27434 22378
rect 27474 22352 27508 22378
rect 27548 22352 27582 22386
rect 27622 22378 27652 22386
rect 27652 22378 27656 22386
rect 27696 22378 27722 22386
rect 27722 22378 27730 22386
rect 27770 22378 27792 22386
rect 27792 22378 27804 22386
rect 27844 22378 27862 22386
rect 27862 22378 27878 22386
rect 27918 22378 27932 22386
rect 27932 22378 27952 22386
rect 27622 22352 27656 22378
rect 27696 22352 27730 22378
rect 27770 22352 27804 22378
rect 27844 22352 27878 22378
rect 27918 22352 27952 22378
rect 26434 22304 26451 22314
rect 26451 22304 26468 22314
rect 26509 22304 26522 22314
rect 26522 22304 26543 22314
rect 26584 22304 26593 22314
rect 26593 22304 26618 22314
rect 26659 22304 26664 22314
rect 26664 22304 26693 22314
rect 26734 22304 26735 22314
rect 26735 22304 26768 22314
rect 26808 22304 26840 22314
rect 26840 22304 26842 22314
rect 26882 22304 26911 22314
rect 26911 22304 26916 22314
rect 26956 22304 26982 22314
rect 26982 22304 26990 22314
rect 27030 22304 27053 22314
rect 27053 22304 27064 22314
rect 27104 22304 27124 22314
rect 27124 22304 27138 22314
rect 27178 22304 27195 22314
rect 27195 22304 27212 22314
rect 27252 22304 27266 22314
rect 27266 22304 27286 22314
rect 27326 22304 27336 22314
rect 27336 22304 27360 22314
rect 27400 22304 27406 22314
rect 27406 22304 27434 22314
rect 27474 22304 27476 22314
rect 27476 22304 27508 22314
rect 26434 22280 26468 22304
rect 26509 22280 26543 22304
rect 26584 22280 26618 22304
rect 26659 22280 26693 22304
rect 26734 22280 26768 22304
rect 26808 22280 26842 22304
rect 26882 22280 26916 22304
rect 26956 22280 26990 22304
rect 27030 22280 27064 22304
rect 27104 22280 27138 22304
rect 27178 22280 27212 22304
rect 27252 22280 27286 22304
rect 27326 22280 27360 22304
rect 27400 22280 27434 22304
rect 27474 22280 27508 22304
rect 27548 22280 27582 22314
rect 27622 22304 27652 22314
rect 27652 22304 27656 22314
rect 27696 22304 27722 22314
rect 27722 22304 27730 22314
rect 27770 22304 27792 22314
rect 27792 22304 27804 22314
rect 27844 22304 27862 22314
rect 27862 22304 27878 22314
rect 27918 22304 27932 22314
rect 27932 22304 27952 22314
rect 27622 22280 27656 22304
rect 27696 22280 27730 22304
rect 27770 22280 27804 22304
rect 27844 22280 27878 22304
rect 27918 22280 27952 22304
rect 26434 22230 26451 22242
rect 26451 22230 26468 22242
rect 26509 22230 26522 22242
rect 26522 22230 26543 22242
rect 26584 22230 26593 22242
rect 26593 22230 26618 22242
rect 26659 22230 26664 22242
rect 26664 22230 26693 22242
rect 26734 22230 26735 22242
rect 26735 22230 26768 22242
rect 26808 22230 26840 22242
rect 26840 22230 26842 22242
rect 26882 22230 26911 22242
rect 26911 22230 26916 22242
rect 26956 22230 26982 22242
rect 26982 22230 26990 22242
rect 27030 22230 27053 22242
rect 27053 22230 27064 22242
rect 27104 22230 27124 22242
rect 27124 22230 27138 22242
rect 27178 22230 27195 22242
rect 27195 22230 27212 22242
rect 27252 22230 27266 22242
rect 27266 22230 27286 22242
rect 27326 22230 27336 22242
rect 27336 22230 27360 22242
rect 27400 22230 27406 22242
rect 27406 22230 27434 22242
rect 27474 22230 27476 22242
rect 27476 22230 27508 22242
rect 26434 22208 26468 22230
rect 26509 22208 26543 22230
rect 26584 22208 26618 22230
rect 26659 22208 26693 22230
rect 26734 22208 26768 22230
rect 26808 22208 26842 22230
rect 26882 22208 26916 22230
rect 26956 22208 26990 22230
rect 27030 22208 27064 22230
rect 27104 22208 27138 22230
rect 27178 22208 27212 22230
rect 27252 22208 27286 22230
rect 27326 22208 27360 22230
rect 27400 22208 27434 22230
rect 27474 22208 27508 22230
rect 27548 22208 27582 22242
rect 27622 22230 27652 22242
rect 27652 22230 27656 22242
rect 27696 22230 27722 22242
rect 27722 22230 27730 22242
rect 27770 22230 27792 22242
rect 27792 22230 27804 22242
rect 27844 22230 27862 22242
rect 27862 22230 27878 22242
rect 27918 22230 27932 22242
rect 27932 22230 27952 22242
rect 27622 22208 27656 22230
rect 27696 22208 27730 22230
rect 27770 22208 27804 22230
rect 27844 22208 27878 22230
rect 27918 22208 27952 22230
rect 26434 22156 26451 22170
rect 26451 22156 26468 22170
rect 26509 22156 26522 22170
rect 26522 22156 26543 22170
rect 26584 22156 26593 22170
rect 26593 22156 26618 22170
rect 26659 22156 26664 22170
rect 26664 22156 26693 22170
rect 26734 22156 26735 22170
rect 26735 22156 26768 22170
rect 26808 22156 26840 22170
rect 26840 22156 26842 22170
rect 26882 22156 26911 22170
rect 26911 22156 26916 22170
rect 26956 22156 26982 22170
rect 26982 22156 26990 22170
rect 27030 22156 27053 22170
rect 27053 22156 27064 22170
rect 27104 22156 27124 22170
rect 27124 22156 27138 22170
rect 27178 22156 27195 22170
rect 27195 22156 27212 22170
rect 27252 22156 27266 22170
rect 27266 22156 27286 22170
rect 27326 22156 27336 22170
rect 27336 22156 27360 22170
rect 27400 22156 27406 22170
rect 27406 22156 27434 22170
rect 27474 22156 27476 22170
rect 27476 22156 27508 22170
rect 26434 22136 26468 22156
rect 26509 22136 26543 22156
rect 26584 22136 26618 22156
rect 26659 22136 26693 22156
rect 26734 22136 26768 22156
rect 26808 22136 26842 22156
rect 26882 22136 26916 22156
rect 26956 22136 26990 22156
rect 27030 22136 27064 22156
rect 27104 22136 27138 22156
rect 27178 22136 27212 22156
rect 27252 22136 27286 22156
rect 27326 22136 27360 22156
rect 27400 22136 27434 22156
rect 27474 22136 27508 22156
rect 27548 22136 27582 22170
rect 27622 22156 27652 22170
rect 27652 22156 27656 22170
rect 27696 22156 27722 22170
rect 27722 22156 27730 22170
rect 27770 22156 27792 22170
rect 27792 22156 27804 22170
rect 27844 22156 27862 22170
rect 27862 22156 27878 22170
rect 27918 22156 27932 22170
rect 27932 22156 27952 22170
rect 27622 22136 27656 22156
rect 27696 22136 27730 22156
rect 27770 22136 27804 22156
rect 27844 22136 27878 22156
rect 27918 22136 27952 22156
rect 2832 3802 2838 3831
rect 2838 3802 2866 3831
rect 2915 3802 2942 3831
rect 2942 3802 2949 3831
rect 2998 3802 3012 3831
rect 3012 3802 3032 3831
rect 3081 3802 3082 3831
rect 3082 3802 3115 3831
rect 3164 3802 3188 3831
rect 3188 3802 3198 3831
rect 2832 3797 2866 3802
rect 2915 3797 2949 3802
rect 2998 3797 3032 3802
rect 3081 3797 3115 3802
rect 3164 3797 3198 3802
rect 2532 3762 2566 3779
rect 2624 3762 2658 3779
rect 2716 3762 2750 3779
rect 2532 3745 2557 3762
rect 2557 3745 2566 3762
rect 2624 3745 2628 3762
rect 2628 3745 2658 3762
rect 2716 3745 2732 3762
rect 2732 3745 2750 3762
rect 2532 3688 2566 3692
rect 2624 3688 2658 3692
rect 2716 3688 2750 3692
rect 2532 3658 2557 3688
rect 2557 3658 2566 3688
rect 2624 3658 2628 3688
rect 2628 3658 2658 3688
rect 2716 3658 2732 3688
rect 2732 3658 2750 3688
rect 2532 3580 2557 3605
rect 2557 3580 2566 3605
rect 2624 3580 2628 3605
rect 2628 3580 2658 3605
rect 2716 3580 2732 3605
rect 2732 3580 2750 3605
rect 2532 3571 2566 3580
rect 2624 3571 2658 3580
rect 2716 3571 2750 3580
rect 2532 3506 2557 3518
rect 2557 3506 2566 3518
rect 2624 3506 2628 3518
rect 2628 3506 2658 3518
rect 2716 3506 2732 3518
rect 2732 3506 2750 3518
rect 2532 3484 2566 3506
rect 2624 3484 2658 3506
rect 2716 3484 2750 3506
rect 12119 3540 12153 3561
rect 12193 3540 12227 3561
rect 12267 3540 12301 3561
rect 12341 3540 12375 3561
rect 12415 3540 12449 3561
rect 12489 3540 12523 3561
rect 12563 3540 12597 3561
rect 12637 3540 12671 3561
rect 12711 3540 12745 3561
rect 12785 3540 12819 3561
rect 12859 3540 12893 3561
rect 12933 3540 12967 3561
rect 13006 3540 13040 3561
rect 13079 3540 13113 3561
rect 12119 3527 12132 3540
rect 12132 3527 12153 3540
rect 12193 3527 12200 3540
rect 12200 3527 12227 3540
rect 12267 3527 12268 3540
rect 12268 3527 12301 3540
rect 12341 3527 12370 3540
rect 12370 3527 12375 3540
rect 12415 3527 12438 3540
rect 12438 3527 12449 3540
rect 12489 3527 12506 3540
rect 12506 3527 12523 3540
rect 12563 3527 12574 3540
rect 12574 3527 12597 3540
rect 12637 3527 12642 3540
rect 12642 3527 12671 3540
rect 12711 3527 12744 3540
rect 12744 3527 12745 3540
rect 12785 3527 12812 3540
rect 12812 3527 12819 3540
rect 12859 3527 12880 3540
rect 12880 3527 12893 3540
rect 12933 3527 12948 3540
rect 12948 3527 12967 3540
rect 13006 3527 13016 3540
rect 13016 3527 13040 3540
rect 13079 3527 13084 3540
rect 13084 3527 13113 3540
rect 13152 3527 13186 3561
rect 13225 3540 13259 3561
rect 13298 3540 13332 3561
rect 13371 3540 13405 3561
rect 13444 3540 13478 3561
rect 13517 3540 13551 3561
rect 13590 3540 13624 3561
rect 13663 3540 13697 3561
rect 13736 3540 13770 3561
rect 13809 3540 13843 3561
rect 13882 3540 13916 3561
rect 13955 3540 13989 3561
rect 14028 3540 14062 3561
rect 14101 3540 14135 3561
rect 14174 3540 14208 3561
rect 14247 3540 14281 3561
rect 14320 3540 14354 3561
rect 14393 3540 14427 3561
rect 14466 3540 14500 3561
rect 14539 3540 14573 3561
rect 14612 3540 14646 3561
rect 14685 3540 14719 3561
rect 14758 3540 14792 3561
rect 13225 3527 13254 3540
rect 13254 3527 13259 3540
rect 13298 3527 13322 3540
rect 13322 3527 13332 3540
rect 13371 3527 13390 3540
rect 13390 3527 13405 3540
rect 13444 3527 13458 3540
rect 13458 3527 13478 3540
rect 13517 3527 13526 3540
rect 13526 3527 13551 3540
rect 13590 3527 13594 3540
rect 13594 3527 13624 3540
rect 13663 3527 13696 3540
rect 13696 3527 13697 3540
rect 13736 3527 13764 3540
rect 13764 3527 13770 3540
rect 13809 3527 13832 3540
rect 13832 3527 13843 3540
rect 13882 3527 13900 3540
rect 13900 3527 13916 3540
rect 13955 3527 13968 3540
rect 13968 3527 13989 3540
rect 14028 3527 14036 3540
rect 14036 3527 14062 3540
rect 14101 3527 14104 3540
rect 14104 3527 14135 3540
rect 14174 3527 14206 3540
rect 14206 3527 14208 3540
rect 14247 3527 14274 3540
rect 14274 3527 14281 3540
rect 14320 3527 14342 3540
rect 14342 3527 14354 3540
rect 14393 3527 14410 3540
rect 14410 3527 14427 3540
rect 14466 3527 14478 3540
rect 14478 3527 14500 3540
rect 14539 3527 14546 3540
rect 14546 3527 14573 3540
rect 14612 3527 14614 3540
rect 14614 3527 14646 3540
rect 14685 3527 14716 3540
rect 14716 3527 14719 3540
rect 14758 3527 14784 3540
rect 14784 3527 14792 3540
rect 17090 3506 17096 3540
rect 17096 3506 17124 3540
rect 17166 3506 17198 3540
rect 17198 3506 17200 3540
rect 17242 3506 17266 3540
rect 17266 3506 17276 3540
rect 17318 3506 17334 3540
rect 17334 3506 17352 3540
rect 17394 3506 17402 3540
rect 17402 3506 17428 3540
rect 17470 3506 17504 3540
rect 17545 3506 17572 3540
rect 17572 3506 17579 3540
rect 17620 3506 17640 3540
rect 17640 3506 17654 3540
rect 17695 3506 17708 3540
rect 17708 3506 17729 3540
rect 17770 3506 17776 3540
rect 17776 3506 17804 3540
rect 17845 3506 17878 3540
rect 17878 3506 17879 3540
rect 17920 3506 17946 3540
rect 17946 3506 17954 3540
rect 17995 3506 18014 3540
rect 18014 3506 18029 3540
rect 18070 3506 18082 3540
rect 18082 3506 18104 3540
rect 18145 3506 18150 3540
rect 18150 3506 18179 3540
rect 18220 3506 18252 3540
rect 18252 3506 18254 3540
rect 18295 3506 18320 3540
rect 18320 3506 18329 3540
rect 18370 3506 18388 3540
rect 18388 3506 18404 3540
rect 18445 3506 18456 3540
rect 18456 3506 18479 3540
rect 18520 3506 18524 3540
rect 18524 3506 18554 3540
rect 18595 3506 18626 3540
rect 18626 3506 18629 3540
rect 18670 3506 18694 3540
rect 18694 3506 18704 3540
rect 12119 3466 12153 3483
rect 12193 3466 12227 3483
rect 12267 3466 12301 3483
rect 12341 3466 12375 3483
rect 12415 3466 12449 3483
rect 12489 3466 12523 3483
rect 12563 3466 12597 3483
rect 12637 3466 12671 3483
rect 12711 3466 12745 3483
rect 12785 3466 12819 3483
rect 12859 3466 12893 3483
rect 12933 3466 12967 3483
rect 13006 3466 13040 3483
rect 13079 3466 13113 3483
rect 12119 3449 12132 3466
rect 12132 3449 12153 3466
rect 12193 3449 12200 3466
rect 12200 3449 12227 3466
rect 12267 3449 12268 3466
rect 12268 3449 12301 3466
rect 12341 3449 12370 3466
rect 12370 3449 12375 3466
rect 12415 3449 12438 3466
rect 12438 3449 12449 3466
rect 12489 3449 12506 3466
rect 12506 3449 12523 3466
rect 12563 3449 12574 3466
rect 12574 3449 12597 3466
rect 12637 3449 12642 3466
rect 12642 3449 12671 3466
rect 12711 3449 12744 3466
rect 12744 3449 12745 3466
rect 12785 3449 12812 3466
rect 12812 3449 12819 3466
rect 12859 3449 12880 3466
rect 12880 3449 12893 3466
rect 12933 3449 12948 3466
rect 12948 3449 12967 3466
rect 13006 3449 13016 3466
rect 13016 3449 13040 3466
rect 13079 3449 13084 3466
rect 13084 3449 13113 3466
rect 13152 3449 13186 3483
rect 13225 3466 13259 3483
rect 13298 3466 13332 3483
rect 13371 3466 13405 3483
rect 13444 3466 13478 3483
rect 13517 3466 13551 3483
rect 13590 3466 13624 3483
rect 13663 3466 13697 3483
rect 13736 3466 13770 3483
rect 13809 3466 13843 3483
rect 13882 3466 13916 3483
rect 13955 3466 13989 3483
rect 14028 3466 14062 3483
rect 14101 3466 14135 3483
rect 14174 3466 14208 3483
rect 14247 3466 14281 3483
rect 14320 3466 14354 3483
rect 14393 3466 14427 3483
rect 14466 3466 14500 3483
rect 14539 3466 14573 3483
rect 14612 3466 14646 3483
rect 14685 3466 14719 3483
rect 14758 3466 14792 3483
rect 13225 3449 13254 3466
rect 13254 3449 13259 3466
rect 13298 3449 13322 3466
rect 13322 3449 13332 3466
rect 13371 3449 13390 3466
rect 13390 3449 13405 3466
rect 13444 3449 13458 3466
rect 13458 3449 13478 3466
rect 13517 3449 13526 3466
rect 13526 3449 13551 3466
rect 13590 3449 13594 3466
rect 13594 3449 13624 3466
rect 13663 3449 13696 3466
rect 13696 3449 13697 3466
rect 13736 3449 13764 3466
rect 13764 3449 13770 3466
rect 13809 3449 13832 3466
rect 13832 3449 13843 3466
rect 13882 3449 13900 3466
rect 13900 3449 13916 3466
rect 13955 3449 13968 3466
rect 13968 3449 13989 3466
rect 14028 3449 14036 3466
rect 14036 3449 14062 3466
rect 14101 3449 14104 3466
rect 14104 3449 14135 3466
rect 14174 3449 14206 3466
rect 14206 3449 14208 3466
rect 14247 3449 14274 3466
rect 14274 3449 14281 3466
rect 14320 3449 14342 3466
rect 14342 3449 14354 3466
rect 14393 3449 14410 3466
rect 14410 3449 14427 3466
rect 14466 3449 14478 3466
rect 14478 3449 14500 3466
rect 14539 3449 14546 3466
rect 14546 3449 14573 3466
rect 14612 3449 14614 3466
rect 14614 3449 14646 3466
rect 14685 3449 14716 3466
rect 14716 3449 14719 3466
rect 14758 3449 14784 3466
rect 14784 3449 14792 3466
rect 3601 2081 3635 2115
rect 3601 2009 3635 2043
<< metal1 >>
tri 19968 38962 20058 39052 sw
rect 11998 38680 12004 38732
rect 12056 38680 12073 38732
rect 12125 38680 12142 38732
rect 12194 38680 12211 38732
rect 12263 38680 12280 38732
rect 12332 38680 12348 38732
rect 12400 38680 12406 38732
rect 11998 38660 12406 38680
rect 11998 38608 12004 38660
rect 12056 38608 12073 38660
rect 12125 38608 12142 38660
rect 12194 38608 12211 38660
rect 12263 38608 12280 38660
rect 12332 38608 12348 38660
rect 12400 38608 12406 38660
rect 11998 38588 12406 38608
rect 11998 38536 12004 38588
rect 12056 38536 12073 38588
rect 12125 38536 12142 38588
rect 12194 38536 12211 38588
rect 12263 38536 12280 38588
rect 12332 38536 12348 38588
rect 12400 38536 12406 38588
rect 19968 38596 20169 38607
rect 19968 38536 19997 38596
tri 19997 38536 20057 38596 nw
tri 19968 38507 19997 38536 nw
rect 25737 37825 25743 37877
rect 25795 37825 25807 37877
rect 25859 37867 26534 37877
tri 26534 37867 26544 37877 sw
rect 25859 37825 26544 37867
tri 26544 37825 26586 37867 sw
tri 26512 37793 26544 37825 ne
rect 26544 37793 26586 37825
tri 26586 37793 26618 37825 sw
tri 26544 37741 26596 37793 ne
rect 26596 37741 27625 37793
tri 27116 37644 27213 37741 ne
rect 26764 37572 26770 37624
rect 26822 37572 26834 37624
rect 26886 37614 26972 37624
tri 26972 37614 26982 37624 sw
rect 27213 37614 27625 37741
rect 26886 37607 26982 37614
tri 26982 37607 26989 37614 sw
rect 26886 37600 26989 37607
tri 26989 37600 26996 37607 sw
rect 27213 37600 27292 37614
rect 26886 37572 26996 37600
tri 26958 37566 26964 37572 ne
rect 26964 37566 26996 37572
tri 26996 37566 27030 37600 sw
rect 27213 37566 27219 37600
rect 27253 37580 27292 37600
rect 27326 37580 27365 37614
rect 27399 37580 27439 37614
rect 27473 37580 27513 37614
rect 27547 37580 27625 37614
rect 27253 37574 27625 37580
rect 27253 37566 27259 37574
tri 26964 37542 26988 37566 ne
rect 26988 37542 27030 37566
tri 27030 37542 27054 37566 sw
tri 26988 37541 26989 37542 ne
rect 26989 37541 27054 37542
tri 27054 37541 27055 37542 sw
tri 26989 37508 27022 37541 ne
rect 27022 37514 27055 37541
tri 27055 37514 27082 37541 sw
rect 27213 37514 27259 37566
rect 27579 37542 27625 37574
rect 27022 37508 27082 37514
tri 27082 37508 27088 37514 sw
rect 27579 37508 27585 37542
rect 27619 37508 27625 37542
tri 27022 37475 27055 37508 ne
rect 27055 37475 27088 37508
tri 27088 37475 27121 37508 sw
tri 27055 37470 27060 37475 ne
rect 27060 37470 27481 37475
tri 27060 37469 27061 37470 ne
rect 27061 37469 27481 37470
tri 27061 37435 27095 37469 ne
rect 27095 37435 27363 37469
rect 27397 37435 27435 37469
rect 27469 37435 27481 37469
tri 27095 37429 27101 37435 ne
rect 27101 37429 27481 37435
rect 27579 37470 27625 37508
rect 27579 37436 27585 37470
rect 27619 37436 27625 37470
rect 27579 37398 27625 37436
rect 27213 37333 27259 37379
rect 27213 37299 27219 37333
rect 27253 37299 27259 37333
rect 27213 37259 27259 37299
rect 27579 37364 27585 37398
rect 27619 37364 27625 37398
rect 27579 37325 27625 37364
rect 27579 37291 27585 37325
rect 27619 37291 27625 37325
rect 27579 37259 27625 37291
rect 27213 37253 27625 37259
rect 27213 37219 27291 37253
rect 27325 37219 27365 37253
rect 27399 37219 27439 37253
rect 27473 37219 27512 37253
rect 27546 37219 27625 37253
rect 27213 37213 27625 37219
rect 2244 34540 3189 34546
rect 2244 34506 2256 34540
rect 2290 34506 2333 34540
rect 2367 34506 2410 34540
rect 2444 34506 2487 34540
rect 2521 34506 2564 34540
rect 2598 34506 2641 34540
rect 2675 34506 2718 34540
rect 2752 34506 2795 34540
rect 2829 34506 2872 34540
rect 2906 34506 2949 34540
rect 2983 34506 3026 34540
rect 3060 34506 3103 34540
rect 3137 34506 3189 34540
rect 2244 34477 3189 34506
tri 3189 34477 3258 34546 sw
rect 2244 34468 3258 34477
rect 2244 34434 2256 34468
rect 2290 34434 2333 34468
rect 2367 34434 2410 34468
rect 2444 34434 2487 34468
rect 2521 34434 2564 34468
rect 2598 34434 2641 34468
rect 2675 34434 2718 34468
rect 2752 34434 2795 34468
rect 2829 34434 2872 34468
rect 2906 34434 2949 34468
rect 2983 34434 3026 34468
rect 3060 34434 3103 34468
rect 3137 34434 3258 34468
rect 2244 34396 3258 34434
rect 2244 34362 2256 34396
rect 2290 34362 2333 34396
rect 2367 34362 2410 34396
rect 2444 34362 2487 34396
rect 2521 34362 2564 34396
rect 2598 34362 2641 34396
rect 2675 34362 2718 34396
rect 2752 34362 2795 34396
rect 2829 34362 2872 34396
rect 2906 34362 2949 34396
rect 2983 34362 3026 34396
rect 3060 34362 3103 34396
rect 3137 34362 3258 34396
rect 2244 34356 3258 34362
tri 2914 34148 3122 34356 ne
rect 3122 33178 3258 34356
tri 3258 33178 3329 33249 sw
rect 3122 33126 3128 33178
rect 3180 33126 3199 33178
rect 3251 33126 3271 33178
rect 3323 33126 3329 33178
rect 3122 33110 3329 33126
rect 3122 33058 3128 33110
rect 3180 33058 3199 33110
rect 3251 33058 3271 33110
rect 3323 33058 3329 33110
rect 2215 32649 2613 32658
rect 2215 32543 2279 32649
rect 2601 32543 2613 32649
rect 2215 32537 2613 32543
rect 2771 32654 3117 32655
rect 2771 32649 2885 32654
rect 2937 32649 2972 32654
rect 3024 32649 3059 32654
rect 2771 32543 2783 32649
rect 3111 32602 3117 32654
rect 3105 32590 3117 32602
rect 2771 32538 2885 32543
rect 2937 32538 2972 32543
rect 3024 32538 3059 32543
rect 3111 32538 3117 32590
rect 2771 32537 3117 32538
tri 2036 32079 2215 32258 se
rect 2215 32162 2382 32537
tri 2382 32459 2460 32537 nw
rect 2215 32079 2299 32162
tri 2299 32079 2382 32162 nw
rect 2036 31950 2204 32079
tri 2204 31984 2299 32079 nw
rect 2088 31898 2140 31950
rect 2192 31898 2204 31950
rect 2036 31882 2204 31898
rect 2088 31830 2140 31882
rect 2192 31830 2204 31882
rect 2036 31814 2204 31830
rect 2088 31762 2140 31814
rect 2192 31762 2204 31814
rect 2036 31756 2204 31762
rect 1666 31115 1888 31121
rect 1666 31063 1667 31115
rect 1719 31063 1751 31115
rect 1803 31063 1835 31115
rect 1887 31063 1888 31115
rect 1666 31036 1888 31063
rect 1666 30984 1667 31036
rect 1719 30984 1751 31036
rect 1803 30984 1835 31036
rect 1887 30984 1888 31036
rect 1666 30957 1888 30984
rect 1666 30905 1667 30957
rect 1719 30905 1751 30957
rect 1803 30905 1835 30957
rect 1887 30905 1888 30957
rect 1666 30878 1888 30905
rect 1666 30826 1667 30878
rect 1719 30826 1751 30878
rect 1803 30826 1835 30878
rect 1887 30826 1888 30878
rect 1666 30820 1888 30826
rect 23794 23284 28000 23290
rect 23794 23250 23806 23284
rect 23840 23250 23879 23284
rect 23913 23250 23952 23284
rect 23986 23250 24025 23284
rect 24059 23250 24098 23284
rect 24132 23250 24171 23284
rect 24205 23250 24244 23284
rect 24278 23250 24317 23284
rect 24351 23250 24390 23284
rect 24424 23250 24462 23284
rect 24496 23250 24534 23284
rect 24568 23250 24606 23284
rect 24640 23250 24678 23284
rect 24712 23250 24750 23284
rect 24784 23250 24822 23284
rect 24856 23250 24894 23284
rect 24928 23250 24966 23284
rect 25000 23250 25038 23284
rect 25072 23250 25110 23284
rect 25144 23250 25182 23284
rect 25216 23250 25254 23284
rect 25288 23250 25326 23284
rect 25360 23250 25398 23284
rect 25432 23250 25470 23284
rect 25504 23250 25542 23284
rect 25576 23250 25614 23284
rect 25648 23250 25686 23284
rect 25720 23250 25758 23284
rect 25792 23250 25830 23284
rect 25864 23250 25902 23284
rect 25936 23250 25974 23284
rect 26008 23250 26046 23284
rect 26080 23250 26118 23284
rect 26152 23250 26190 23284
rect 26224 23250 26262 23284
rect 26296 23250 26334 23284
rect 26368 23250 26406 23284
rect 26440 23250 26478 23284
rect 26512 23250 26550 23284
rect 26584 23250 26622 23284
rect 26656 23250 26694 23284
rect 26728 23250 26766 23284
rect 26800 23250 26838 23284
rect 26872 23250 26910 23284
rect 26944 23250 26982 23284
rect 27016 23276 27054 23284
rect 27088 23276 27126 23284
rect 27160 23276 27198 23284
rect 27232 23276 27270 23284
rect 27304 23276 27342 23284
rect 27376 23276 27414 23284
rect 27448 23276 27486 23284
rect 27520 23276 27558 23284
rect 27592 23276 27630 23284
rect 27016 23250 27050 23276
rect 23794 23224 27050 23250
rect 27102 23224 27121 23276
rect 27173 23224 27192 23276
rect 27244 23224 27262 23276
rect 27314 23224 27332 23276
rect 27384 23224 27402 23276
rect 27454 23224 27472 23276
rect 27524 23224 27542 23276
rect 27594 23224 27612 23276
rect 27664 23250 27702 23284
rect 27736 23250 27774 23284
rect 27808 23250 27846 23284
rect 27880 23250 27918 23284
rect 27952 23250 28000 23284
rect 27664 23224 28000 23250
rect 23794 23210 28000 23224
rect 23794 23198 27050 23210
rect 23794 23164 23806 23198
rect 23840 23164 23879 23198
rect 23913 23164 23952 23198
rect 23986 23164 24025 23198
rect 24059 23164 24098 23198
rect 24132 23164 24171 23198
rect 24205 23164 24244 23198
rect 24278 23164 24317 23198
rect 24351 23164 24390 23198
rect 24424 23164 24462 23198
rect 24496 23164 24534 23198
rect 24568 23164 24606 23198
rect 24640 23164 24678 23198
rect 24712 23164 24750 23198
rect 24784 23164 24822 23198
rect 24856 23164 24894 23198
rect 24928 23164 24966 23198
rect 25000 23164 25038 23198
rect 25072 23164 25110 23198
rect 25144 23164 25182 23198
rect 25216 23164 25254 23198
rect 25288 23164 25326 23198
rect 25360 23164 25398 23198
rect 25432 23164 25470 23198
rect 25504 23164 25542 23198
rect 25576 23164 25614 23198
rect 25648 23164 25686 23198
rect 25720 23164 25758 23198
rect 25792 23164 25830 23198
rect 25864 23164 25902 23198
rect 25936 23164 25974 23198
rect 26008 23164 26046 23198
rect 26080 23164 26118 23198
rect 26152 23164 26190 23198
rect 26224 23164 26262 23198
rect 26296 23164 26334 23198
rect 26368 23164 26406 23198
rect 26440 23164 26478 23198
rect 26512 23164 26550 23198
rect 26584 23164 26622 23198
rect 26656 23164 26694 23198
rect 26728 23164 26766 23198
rect 26800 23164 26838 23198
rect 26872 23164 26910 23198
rect 26944 23164 26982 23198
rect 27016 23164 27050 23198
rect 23794 23158 27050 23164
rect 27102 23158 27121 23210
rect 27173 23158 27192 23210
rect 27244 23158 27262 23210
rect 27314 23158 27332 23210
rect 27384 23158 27402 23210
rect 27454 23158 27472 23210
rect 27524 23158 27542 23210
rect 27594 23158 27612 23210
rect 27664 23198 28000 23210
rect 27664 23164 27702 23198
rect 27736 23164 27774 23198
rect 27808 23164 27846 23198
rect 27880 23164 27918 23198
rect 27952 23164 28000 23198
rect 27664 23158 28000 23164
rect 23794 23144 28000 23158
rect 23794 23112 27050 23144
rect 23794 23078 23806 23112
rect 23840 23078 23879 23112
rect 23913 23078 23952 23112
rect 23986 23078 24025 23112
rect 24059 23078 24098 23112
rect 24132 23078 24171 23112
rect 24205 23078 24244 23112
rect 24278 23078 24317 23112
rect 24351 23078 24390 23112
rect 24424 23078 24462 23112
rect 24496 23078 24534 23112
rect 24568 23078 24606 23112
rect 24640 23078 24678 23112
rect 24712 23078 24750 23112
rect 24784 23078 24822 23112
rect 24856 23078 24894 23112
rect 24928 23078 24966 23112
rect 25000 23078 25038 23112
rect 25072 23078 25110 23112
rect 25144 23078 25182 23112
rect 25216 23078 25254 23112
rect 25288 23078 25326 23112
rect 25360 23078 25398 23112
rect 25432 23078 25470 23112
rect 25504 23078 25542 23112
rect 25576 23078 25614 23112
rect 25648 23078 25686 23112
rect 25720 23078 25758 23112
rect 25792 23078 25830 23112
rect 25864 23078 25902 23112
rect 25936 23078 25974 23112
rect 26008 23078 26046 23112
rect 26080 23078 26118 23112
rect 26152 23078 26190 23112
rect 26224 23078 26262 23112
rect 26296 23078 26334 23112
rect 26368 23078 26406 23112
rect 26440 23078 26478 23112
rect 26512 23078 26550 23112
rect 26584 23078 26622 23112
rect 26656 23078 26694 23112
rect 26728 23078 26766 23112
rect 26800 23078 26838 23112
rect 26872 23078 26910 23112
rect 26944 23078 26982 23112
rect 27016 23092 27050 23112
rect 27102 23092 27121 23144
rect 27173 23092 27192 23144
rect 27244 23092 27262 23144
rect 27314 23092 27332 23144
rect 27384 23092 27402 23144
rect 27454 23092 27472 23144
rect 27524 23092 27542 23144
rect 27594 23092 27612 23144
rect 27664 23112 28000 23144
rect 27016 23078 27054 23092
rect 27088 23078 27126 23092
rect 27160 23078 27198 23092
rect 27232 23078 27270 23092
rect 27304 23078 27342 23092
rect 27376 23078 27414 23092
rect 27448 23078 27486 23092
rect 27520 23078 27558 23092
rect 27592 23078 27630 23092
rect 27664 23078 27702 23112
rect 27736 23078 27774 23112
rect 27808 23078 27846 23112
rect 27880 23078 27918 23112
rect 27952 23078 28000 23112
rect 23794 23026 27050 23078
rect 27102 23026 27121 23078
rect 27173 23026 27192 23078
rect 27244 23026 27262 23078
rect 27314 23026 27332 23078
rect 27384 23026 27402 23078
rect 27454 23026 27472 23078
rect 27524 23026 27542 23078
rect 27594 23026 27612 23078
rect 27664 23026 28000 23078
rect 23794 22992 23806 23026
rect 23840 22992 23879 23026
rect 23913 22992 23952 23026
rect 23986 22992 24025 23026
rect 24059 22992 24098 23026
rect 24132 22992 24171 23026
rect 24205 22992 24244 23026
rect 24278 22992 24317 23026
rect 24351 22992 24390 23026
rect 24424 22992 24462 23026
rect 24496 22992 24534 23026
rect 24568 22992 24606 23026
rect 24640 22992 24678 23026
rect 24712 22992 24750 23026
rect 24784 22992 24822 23026
rect 24856 22992 24894 23026
rect 24928 22992 24966 23026
rect 25000 22992 25038 23026
rect 25072 22992 25110 23026
rect 25144 22992 25182 23026
rect 25216 22992 25254 23026
rect 25288 22992 25326 23026
rect 25360 22992 25398 23026
rect 25432 22992 25470 23026
rect 25504 22992 25542 23026
rect 25576 22992 25614 23026
rect 25648 22992 25686 23026
rect 25720 22992 25758 23026
rect 25792 22992 25830 23026
rect 25864 22992 25902 23026
rect 25936 22992 25974 23026
rect 26008 22992 26046 23026
rect 26080 22992 26118 23026
rect 26152 22992 26190 23026
rect 26224 22992 26262 23026
rect 26296 22992 26334 23026
rect 26368 22992 26406 23026
rect 26440 22992 26478 23026
rect 26512 22992 26550 23026
rect 26584 22992 26622 23026
rect 26656 22992 26694 23026
rect 26728 22992 26766 23026
rect 26800 22992 26838 23026
rect 26872 22992 26910 23026
rect 26944 22992 26982 23026
rect 27016 23012 27054 23026
rect 27088 23012 27126 23026
rect 27160 23012 27198 23026
rect 27232 23012 27270 23026
rect 27304 23012 27342 23026
rect 27376 23012 27414 23026
rect 27448 23012 27486 23026
rect 27520 23012 27558 23026
rect 27592 23012 27630 23026
rect 27016 22992 27050 23012
rect 23794 22986 27050 22992
tri 26332 22896 26422 22986 ne
rect 26422 22960 27050 22986
rect 27102 22960 27121 23012
rect 27173 22960 27192 23012
rect 27244 22960 27262 23012
rect 27314 22960 27332 23012
rect 27384 22960 27402 23012
rect 27454 22960 27472 23012
rect 27524 22960 27542 23012
rect 27594 22960 27612 23012
rect 27664 22992 27702 23026
rect 27736 22992 27774 23026
rect 27808 22992 27846 23026
rect 27880 22992 27918 23026
rect 27952 22992 28000 23026
rect 27664 22960 28000 22992
rect 26422 22946 28000 22960
rect 26422 22894 27050 22946
rect 27102 22894 27121 22946
rect 27173 22894 27192 22946
rect 27244 22894 27262 22946
rect 27314 22894 27332 22946
rect 27384 22894 27402 22946
rect 27454 22894 27472 22946
rect 27524 22894 27542 22946
rect 27594 22894 27612 22946
rect 27664 22894 28000 22946
rect 26422 22890 28000 22894
rect 26422 22856 26434 22890
rect 26468 22856 26509 22890
rect 26543 22856 26584 22890
rect 26618 22856 26659 22890
rect 26693 22856 26734 22890
rect 26768 22856 26808 22890
rect 26842 22856 26882 22890
rect 26916 22856 26956 22890
rect 26990 22856 27030 22890
rect 27064 22856 27104 22890
rect 27138 22856 27178 22890
rect 27212 22856 27252 22890
rect 27286 22856 27326 22890
rect 27360 22861 27400 22890
rect 27434 22861 27474 22890
rect 27508 22861 27548 22890
rect 27582 22861 27622 22890
rect 27656 22861 27696 22890
rect 27471 22856 27474 22861
rect 26422 22818 27355 22856
rect 27407 22818 27419 22856
rect 27471 22818 27483 22856
rect 26422 22784 26434 22818
rect 26468 22784 26509 22818
rect 26543 22784 26584 22818
rect 26618 22784 26659 22818
rect 26693 22784 26734 22818
rect 26768 22784 26808 22818
rect 26842 22784 26882 22818
rect 26916 22784 26956 22818
rect 26990 22784 27030 22818
rect 27064 22784 27104 22818
rect 27138 22784 27178 22818
rect 27212 22784 27252 22818
rect 27286 22784 27326 22818
rect 27471 22809 27474 22818
rect 27535 22809 27547 22861
rect 27599 22809 27611 22861
rect 27663 22856 27696 22861
rect 27730 22856 27770 22890
rect 27804 22856 27844 22890
rect 27878 22856 27918 22890
rect 27952 22856 28000 22890
rect 27663 22818 28000 22856
rect 27663 22809 27696 22818
rect 27360 22794 27400 22809
rect 27434 22794 27474 22809
rect 27508 22794 27548 22809
rect 27582 22794 27622 22809
rect 27656 22794 27696 22809
rect 27471 22784 27474 22794
rect 26422 22746 27355 22784
rect 27407 22746 27419 22784
rect 27471 22746 27483 22784
rect 26422 22712 26434 22746
rect 26468 22712 26509 22746
rect 26543 22712 26584 22746
rect 26618 22712 26659 22746
rect 26693 22712 26734 22746
rect 26768 22712 26808 22746
rect 26842 22712 26882 22746
rect 26916 22712 26956 22746
rect 26990 22712 27030 22746
rect 27064 22712 27104 22746
rect 27138 22712 27178 22746
rect 27212 22712 27252 22746
rect 27286 22712 27326 22746
rect 27471 22742 27474 22746
rect 27535 22742 27547 22794
rect 27599 22742 27611 22794
rect 27663 22784 27696 22794
rect 27730 22784 27770 22818
rect 27804 22784 27844 22818
rect 27878 22784 27918 22818
rect 27952 22784 28000 22818
rect 27663 22746 28000 22784
rect 27663 22742 27696 22746
rect 27360 22727 27400 22742
rect 27434 22727 27474 22742
rect 27508 22727 27548 22742
rect 27582 22727 27622 22742
rect 27656 22727 27696 22742
rect 27471 22712 27474 22727
rect 26422 22675 27355 22712
rect 27407 22675 27419 22712
rect 27471 22675 27483 22712
rect 27535 22675 27547 22727
rect 27599 22675 27611 22727
rect 27663 22712 27696 22727
rect 27730 22712 27770 22746
rect 27804 22712 27844 22746
rect 27878 22712 27918 22746
rect 27952 22712 28000 22746
rect 27663 22675 28000 22712
rect 26422 22674 28000 22675
rect 26422 22640 26434 22674
rect 26468 22640 26509 22674
rect 26543 22640 26584 22674
rect 26618 22640 26659 22674
rect 26693 22640 26734 22674
rect 26768 22640 26808 22674
rect 26842 22640 26882 22674
rect 26916 22640 26956 22674
rect 26990 22640 27030 22674
rect 27064 22640 27104 22674
rect 27138 22640 27178 22674
rect 27212 22640 27252 22674
rect 27286 22640 27326 22674
rect 27360 22660 27400 22674
rect 27434 22660 27474 22674
rect 27508 22660 27548 22674
rect 27582 22660 27622 22674
rect 27656 22660 27696 22674
rect 27471 22640 27474 22660
rect 26422 22608 27355 22640
rect 27407 22608 27419 22640
rect 27471 22608 27483 22640
rect 27535 22608 27547 22660
rect 27599 22608 27611 22660
rect 27663 22640 27696 22660
rect 27730 22640 27770 22674
rect 27804 22640 27844 22674
rect 27878 22640 27918 22674
rect 27952 22640 28000 22674
rect 27663 22608 28000 22640
rect 26422 22602 28000 22608
rect 26422 22568 26434 22602
rect 26468 22568 26509 22602
rect 26543 22568 26584 22602
rect 26618 22568 26659 22602
rect 26693 22568 26734 22602
rect 26768 22568 26808 22602
rect 26842 22568 26882 22602
rect 26916 22568 26956 22602
rect 26990 22568 27030 22602
rect 27064 22568 27104 22602
rect 27138 22568 27178 22602
rect 27212 22568 27252 22602
rect 27286 22568 27326 22602
rect 27360 22593 27400 22602
rect 27434 22593 27474 22602
rect 27508 22593 27548 22602
rect 27582 22593 27622 22602
rect 27656 22593 27696 22602
rect 27471 22568 27474 22593
rect 26422 22541 27355 22568
rect 27407 22541 27419 22568
rect 27471 22541 27483 22568
rect 27535 22541 27547 22593
rect 27599 22541 27611 22593
rect 27663 22568 27696 22593
rect 27730 22568 27770 22602
rect 27804 22568 27844 22602
rect 27878 22568 27918 22602
rect 27952 22568 28000 22602
rect 27663 22541 28000 22568
rect 26422 22530 28000 22541
rect 26422 22496 26434 22530
rect 26468 22496 26509 22530
rect 26543 22496 26584 22530
rect 26618 22496 26659 22530
rect 26693 22496 26734 22530
rect 26768 22496 26808 22530
rect 26842 22496 26882 22530
rect 26916 22496 26956 22530
rect 26990 22496 27030 22530
rect 27064 22496 27104 22530
rect 27138 22496 27178 22530
rect 27212 22496 27252 22530
rect 27286 22496 27326 22530
rect 27360 22526 27400 22530
rect 27434 22526 27474 22530
rect 27508 22526 27548 22530
rect 27582 22526 27622 22530
rect 27656 22526 27696 22530
rect 27471 22496 27474 22526
rect 26422 22474 27355 22496
rect 27407 22474 27419 22496
rect 27471 22474 27483 22496
rect 27535 22474 27547 22526
rect 27599 22474 27611 22526
rect 27663 22496 27696 22526
rect 27730 22496 27770 22530
rect 27804 22496 27844 22530
rect 27878 22496 27918 22530
rect 27952 22496 28000 22530
rect 27663 22474 28000 22496
rect 26422 22459 28000 22474
rect 26422 22458 27355 22459
rect 27407 22458 27419 22459
rect 27471 22458 27483 22459
rect 26422 22424 26434 22458
rect 26468 22424 26509 22458
rect 26543 22424 26584 22458
rect 26618 22424 26659 22458
rect 26693 22424 26734 22458
rect 26768 22424 26808 22458
rect 26842 22424 26882 22458
rect 26916 22424 26956 22458
rect 26990 22424 27030 22458
rect 27064 22424 27104 22458
rect 27138 22424 27178 22458
rect 27212 22424 27252 22458
rect 27286 22424 27326 22458
rect 27471 22424 27474 22458
rect 26422 22407 27355 22424
rect 27407 22407 27419 22424
rect 27471 22407 27483 22424
rect 27535 22407 27547 22459
rect 27599 22407 27611 22459
rect 27663 22458 28000 22459
rect 27663 22424 27696 22458
rect 27730 22424 27770 22458
rect 27804 22424 27844 22458
rect 27878 22424 27918 22458
rect 27952 22424 28000 22458
rect 27663 22407 28000 22424
rect 26422 22392 28000 22407
rect 26422 22386 27355 22392
rect 27407 22386 27419 22392
rect 27471 22386 27483 22392
rect 26422 22352 26434 22386
rect 26468 22352 26509 22386
rect 26543 22352 26584 22386
rect 26618 22352 26659 22386
rect 26693 22352 26734 22386
rect 26768 22352 26808 22386
rect 26842 22352 26882 22386
rect 26916 22352 26956 22386
rect 26990 22352 27030 22386
rect 27064 22352 27104 22386
rect 27138 22352 27178 22386
rect 27212 22352 27252 22386
rect 27286 22352 27326 22386
rect 27471 22352 27474 22386
rect 26422 22340 27355 22352
rect 27407 22340 27419 22352
rect 27471 22340 27483 22352
rect 27535 22340 27547 22392
rect 27599 22340 27611 22392
rect 27663 22386 28000 22392
rect 27663 22352 27696 22386
rect 27730 22352 27770 22386
rect 27804 22352 27844 22386
rect 27878 22352 27918 22386
rect 27952 22352 28000 22386
rect 27663 22340 28000 22352
rect 26422 22324 28000 22340
rect 26422 22314 27355 22324
rect 27407 22314 27419 22324
rect 27471 22314 27483 22324
rect 26422 22280 26434 22314
rect 26468 22280 26509 22314
rect 26543 22280 26584 22314
rect 26618 22280 26659 22314
rect 26693 22280 26734 22314
rect 26768 22280 26808 22314
rect 26842 22280 26882 22314
rect 26916 22280 26956 22314
rect 26990 22280 27030 22314
rect 27064 22280 27104 22314
rect 27138 22280 27178 22314
rect 27212 22280 27252 22314
rect 27286 22280 27326 22314
rect 27471 22280 27474 22314
rect 26422 22272 27355 22280
rect 27407 22272 27419 22280
rect 27471 22272 27483 22280
rect 27535 22272 27547 22324
rect 27599 22272 27611 22324
rect 27663 22314 28000 22324
rect 27663 22280 27696 22314
rect 27730 22280 27770 22314
rect 27804 22280 27844 22314
rect 27878 22280 27918 22314
rect 27952 22280 28000 22314
rect 27663 22272 28000 22280
rect 26422 22256 28000 22272
rect 26422 22242 27355 22256
rect 27407 22242 27419 22256
rect 27471 22242 27483 22256
rect 26422 22208 26434 22242
rect 26468 22208 26509 22242
rect 26543 22208 26584 22242
rect 26618 22208 26659 22242
rect 26693 22208 26734 22242
rect 26768 22208 26808 22242
rect 26842 22208 26882 22242
rect 26916 22208 26956 22242
rect 26990 22208 27030 22242
rect 27064 22208 27104 22242
rect 27138 22208 27178 22242
rect 27212 22208 27252 22242
rect 27286 22208 27326 22242
rect 27471 22208 27474 22242
rect 26422 22204 27355 22208
rect 27407 22204 27419 22208
rect 27471 22204 27483 22208
rect 27535 22204 27547 22256
rect 27599 22204 27611 22256
rect 27663 22242 28000 22256
rect 27663 22208 27696 22242
rect 27730 22208 27770 22242
rect 27804 22208 27844 22242
rect 27878 22208 27918 22242
rect 27952 22208 28000 22242
rect 27663 22204 28000 22208
rect 26422 22188 28000 22204
rect 26422 22170 27355 22188
rect 27407 22170 27419 22188
rect 27471 22170 27483 22188
rect 26422 22136 26434 22170
rect 26468 22136 26509 22170
rect 26543 22136 26584 22170
rect 26618 22136 26659 22170
rect 26693 22136 26734 22170
rect 26768 22136 26808 22170
rect 26842 22136 26882 22170
rect 26916 22136 26956 22170
rect 26990 22136 27030 22170
rect 27064 22136 27104 22170
rect 27138 22136 27178 22170
rect 27212 22136 27252 22170
rect 27286 22136 27326 22170
rect 27471 22136 27474 22170
rect 27535 22136 27547 22188
rect 27599 22136 27611 22188
rect 27663 22170 28000 22188
rect 27663 22136 27696 22170
rect 27730 22136 27770 22170
rect 27804 22136 27844 22170
rect 27878 22136 27918 22170
rect 27952 22136 28000 22170
rect 26422 22130 28000 22136
rect 1836 21364 1960 21370
rect 1888 21312 1908 21364
rect 1836 21300 1960 21312
rect 1888 21248 1908 21300
rect 1836 21236 1960 21248
rect 1888 21184 1908 21236
rect 27341 21323 27364 21375
rect 27416 21323 27428 21375
rect 27480 21323 27503 21375
rect 27341 21269 27503 21323
rect 27341 21217 27364 21269
rect 27416 21217 27428 21269
rect 27480 21217 27503 21269
rect 27515 21367 27673 21373
rect 27567 21315 27621 21367
rect 27515 21288 27673 21315
rect 27567 21236 27621 21288
rect 1836 21172 1960 21184
rect 1888 21120 1908 21172
rect 27515 21209 27673 21236
rect 27567 21157 27621 21209
rect 27515 21151 27673 21157
rect 1836 21108 1960 21120
rect 1888 21056 1908 21108
rect 1836 21044 1960 21056
rect 1888 20992 1908 21044
rect 1836 20980 1960 20992
rect 1888 20928 1908 20980
rect 1836 20916 1960 20928
rect 1888 20864 1908 20916
rect 1836 20852 1960 20864
rect 1888 20800 1908 20852
rect 1836 20788 1960 20800
rect 1888 20736 1908 20788
rect 1836 20724 1960 20736
rect 1888 20672 1908 20724
rect 1836 20660 1960 20672
rect 1888 20608 1908 20660
rect 1836 20596 1960 20608
rect 1888 20544 1908 20596
rect 1836 20532 1960 20544
rect 1888 20480 1908 20532
rect 1836 20468 1960 20480
rect 1888 20416 1908 20468
rect 1836 20404 1960 20416
rect 1888 20352 1908 20404
rect 1836 20340 1960 20352
rect 1888 20288 1908 20340
rect 1836 20276 1960 20288
rect 1888 20224 1908 20276
rect 1836 20212 1960 20224
rect 1888 20160 1908 20212
rect 1836 20148 1960 20160
rect 1888 20096 1908 20148
rect 1836 20084 1960 20096
rect 1888 20032 1908 20084
rect 1836 20020 1960 20032
rect 1888 19968 1908 20020
rect 1836 19956 1960 19968
rect 1888 19904 1908 19956
rect 1836 19892 1960 19904
rect 1888 19840 1908 19892
rect 1836 19828 1960 19840
rect 1888 19776 1908 19828
rect 1836 19764 1960 19776
rect 1888 19712 1908 19764
rect 1836 19700 1960 19712
rect 1888 19648 1908 19700
rect 1836 19636 1960 19648
rect 1888 19584 1908 19636
rect 1836 19572 1960 19584
rect 1888 19520 1908 19572
rect 1836 19507 1960 19520
rect 1888 19455 1908 19507
rect 1836 19442 1960 19455
rect 1888 19390 1908 19442
rect 1836 19377 1960 19390
rect 1888 19325 1908 19377
rect 1836 19312 1960 19325
rect 1888 19260 1908 19312
rect 1836 19247 1960 19260
rect 1888 19195 1908 19247
rect 1836 19182 1960 19195
rect 1888 19130 1908 19182
rect 1836 19117 1960 19130
rect 1888 19065 1908 19117
rect 1836 19052 1960 19065
rect 1888 19000 1908 19052
rect 1836 18987 1960 19000
rect 1888 18935 1908 18987
rect 1836 18922 1960 18935
rect 1888 18870 1908 18922
rect 1836 18857 1960 18870
rect 1888 18805 1908 18857
rect 1836 18792 1960 18805
rect 1888 18740 1908 18792
rect 1836 18727 1960 18740
rect 1888 18675 1908 18727
rect 1836 18662 1960 18675
rect 1888 18610 1908 18662
rect 1836 18597 1960 18610
rect 1888 18545 1908 18597
rect 1836 18532 1960 18545
rect 1888 18480 1908 18532
rect 1836 18474 1960 18480
rect 1796 18192 1984 18198
rect 1848 18140 1864 18192
rect 1916 18140 1932 18192
rect 1796 18120 1984 18140
rect 1848 18068 1864 18120
rect 1916 18068 1932 18120
rect 1796 18047 1984 18068
rect 1848 17995 1864 18047
rect 1916 17995 1932 18047
rect 1796 17974 1984 17995
rect 1848 17922 1864 17974
rect 1916 17922 1932 17974
rect 1796 17901 1984 17922
rect 1848 17849 1864 17901
rect 1916 17849 1932 17901
rect 1796 17828 1984 17849
rect 1848 17776 1864 17828
rect 1916 17776 1932 17828
rect 1796 17755 1984 17776
rect 1848 17703 1864 17755
rect 1916 17703 1932 17755
rect 1796 17697 1984 17703
rect 1796 17518 1984 17524
rect 1848 17466 1864 17518
rect 1916 17466 1932 17518
rect 1796 17453 1984 17466
rect 1848 17401 1864 17453
rect 1916 17401 1932 17453
rect 1796 17387 1984 17401
rect 1848 17335 1864 17387
rect 1916 17335 1932 17387
rect 1796 17321 1984 17335
rect 1848 17269 1864 17321
rect 1916 17269 1932 17321
rect 1796 17255 1984 17269
rect 1848 17203 1864 17255
rect 1916 17203 1932 17255
rect 1796 17189 1984 17203
rect 1848 17137 1864 17189
rect 1916 17137 1932 17189
rect 1796 17123 1984 17137
rect 1848 17071 1864 17123
rect 1916 17071 1932 17123
rect 1796 17065 1984 17071
rect 1796 16313 1984 16319
rect 1848 16261 1864 16313
rect 1916 16261 1932 16313
rect 1796 16249 1984 16261
rect 1848 16197 1864 16249
rect 1916 16197 1932 16249
rect 1796 16185 1984 16197
rect 1848 16133 1864 16185
rect 1916 16133 1932 16185
rect 1796 16121 1984 16133
rect 1848 16069 1864 16121
rect 1916 16069 1932 16121
rect 1796 16057 1984 16069
rect 1848 16005 1864 16057
rect 1916 16005 1932 16057
rect 1796 15993 1984 16005
rect 1848 15941 1864 15993
rect 1916 15941 1932 15993
rect 1796 15929 1984 15941
rect 1848 15877 1864 15929
rect 1916 15877 1932 15929
rect 1796 15864 1984 15877
rect 1848 15812 1864 15864
rect 1916 15812 1932 15864
rect 1796 15799 1984 15812
rect 1848 15747 1864 15799
rect 1916 15747 1932 15799
rect 1796 15734 1984 15747
rect 1848 15682 1864 15734
rect 1916 15682 1932 15734
rect 1796 15669 1984 15682
rect 1848 15617 1864 15669
rect 1916 15617 1932 15669
rect 1796 15604 1984 15617
rect 1848 15552 1864 15604
rect 1916 15552 1932 15604
rect 1796 15539 1984 15552
rect 1848 15487 1864 15539
rect 1916 15487 1932 15539
rect 1796 15481 1984 15487
rect 1796 14640 1984 14646
rect 1848 14588 1864 14640
rect 1916 14588 1932 14640
rect 1796 14568 1984 14588
rect 1848 14516 1864 14568
rect 1916 14516 1932 14568
rect 1796 14496 1984 14516
tri 26220 14496 26275 14551 se
rect 26275 14499 26814 14551
rect 26866 14499 26878 14551
rect 26930 14499 26936 14551
rect 26275 14496 26293 14499
tri 26293 14496 26296 14499 nw
rect 1848 14444 1864 14496
rect 1916 14444 1932 14496
rect 3382 14444 3388 14496
rect 3440 14444 3452 14496
rect 3504 14466 26263 14496
tri 26263 14466 26293 14496 nw
rect 3504 14456 3522 14466
tri 3522 14456 3532 14466 nw
rect 3504 14444 3510 14456
tri 3510 14444 3522 14456 nw
tri 26339 14444 26351 14456 se
rect 26351 14444 26357 14456
rect 1796 14424 1984 14444
tri 26333 14438 26339 14444 se
rect 26339 14438 26357 14444
rect 1848 14372 1864 14424
rect 1916 14372 1932 14424
tri 3567 14422 3583 14438 se
rect 3583 14422 26357 14438
rect 1796 14351 1984 14372
rect 3214 14370 3220 14422
rect 3272 14370 3284 14422
rect 3336 14404 3342 14422
tri 3342 14404 3360 14422 sw
tri 3549 14404 3567 14422 se
rect 3567 14404 26357 14422
rect 26409 14404 26421 14456
rect 26473 14404 26479 14456
rect 3336 14370 3617 14404
tri 3617 14370 3651 14404 nw
rect 1848 14299 1864 14351
rect 1916 14299 1932 14351
rect 1796 14278 1984 14299
rect 1848 14226 1864 14278
rect 1916 14226 1932 14278
rect 1796 14205 1984 14226
rect 1848 14153 1864 14205
rect 1916 14153 1932 14205
rect 1796 14132 1984 14153
rect 1848 14080 1864 14132
rect 1916 14080 1932 14132
rect 1796 14074 1984 14080
rect 27562 13627 27690 13628
rect 27105 13623 27302 13624
rect 27105 13571 27111 13623
rect 27163 13571 27178 13623
rect 27230 13571 27244 13623
rect 27296 13571 27302 13623
rect 27105 13553 27302 13571
rect 27105 13501 27111 13553
rect 27163 13501 27178 13553
rect 27230 13501 27244 13553
rect 27296 13501 27302 13553
rect 27105 13483 27302 13501
rect 27105 13431 27111 13483
rect 27163 13431 27178 13483
rect 27230 13431 27244 13483
rect 27296 13431 27302 13483
rect 27562 13575 27568 13627
rect 27620 13575 27632 13627
rect 27684 13575 27690 13627
rect 27562 13557 27690 13575
rect 27562 13505 27568 13557
rect 27620 13505 27632 13557
rect 27684 13505 27690 13557
rect 27562 13487 27690 13505
rect 27562 13435 27568 13487
rect 27620 13435 27632 13487
rect 27684 13435 27690 13487
rect 27562 13434 27690 13435
rect 27105 13430 27302 13431
rect 27968 12936 28032 12937
rect 27105 12934 27302 12935
rect 27105 12882 27111 12934
rect 27163 12882 27178 12934
rect 27230 12882 27244 12934
rect 27296 12882 27302 12934
tri 1398 12862 1406 12870 se
rect 1406 12862 1811 12870
rect 826 12856 1811 12862
rect 878 12804 890 12856
rect 942 12804 954 12856
rect 1006 12804 1811 12856
rect 826 12781 1811 12804
rect 878 12729 890 12781
rect 942 12729 954 12781
rect 1006 12729 1811 12781
rect 27105 12864 27302 12882
rect 27105 12812 27111 12864
rect 27163 12812 27178 12864
rect 27230 12812 27244 12864
rect 27296 12812 27302 12864
rect 27105 12794 27302 12812
rect 27105 12742 27111 12794
rect 27163 12742 27178 12794
rect 27230 12742 27244 12794
rect 27296 12742 27302 12794
rect 27105 12741 27302 12742
rect 27365 12934 27562 12935
rect 27365 12882 27371 12934
rect 27423 12882 27438 12934
rect 27490 12882 27504 12934
rect 27556 12882 27562 12934
rect 27365 12864 27562 12882
rect 27365 12812 27371 12864
rect 27423 12812 27438 12864
rect 27490 12812 27504 12864
rect 27556 12812 27562 12864
rect 27365 12794 27562 12812
rect 27365 12742 27371 12794
rect 27423 12742 27438 12794
rect 27490 12742 27504 12794
rect 27556 12742 27562 12794
rect 27968 12884 27974 12936
rect 28026 12884 28032 12936
rect 27968 12866 28032 12884
rect 27968 12814 27974 12866
rect 28026 12814 28032 12866
rect 27968 12796 28032 12814
rect 27968 12744 27974 12796
rect 28026 12744 28032 12796
rect 27968 12743 28032 12744
rect 27365 12741 27562 12742
rect 826 12705 1811 12729
rect 878 12653 890 12705
rect 942 12653 954 12705
rect 1006 12653 1811 12705
rect 826 12629 1811 12653
rect 878 12577 890 12629
rect 942 12577 954 12629
rect 1006 12577 1811 12629
rect 826 12571 1811 12577
tri 1357 12522 1406 12571 ne
rect 1406 12380 1811 12571
rect 25801 11368 25807 11420
rect 25859 11368 25871 11420
rect 25923 11368 25929 11420
rect 27471 11095 27617 11101
rect 27523 11043 27565 11095
rect 27471 11000 27617 11043
rect 13662 10935 13668 10987
rect 13720 10935 13732 10987
rect 13784 10981 13790 10987
rect 13784 10935 13965 10981
rect 27523 10948 27565 11000
rect 27471 10942 27617 10948
rect 102 10920 154 10926
rect 707 10920 759 10926
rect 154 10868 707 10907
rect 102 10856 759 10868
rect 154 10848 707 10856
rect 102 10798 154 10804
rect 707 10798 759 10804
rect 226 10785 278 10791
rect 226 10730 278 10733
rect 1153 10757 1205 10763
rect 226 10721 1153 10730
rect 278 10705 1153 10721
rect 10493 10738 10540 10920
rect 278 10693 1205 10705
rect 278 10671 1153 10693
rect 226 10663 278 10669
rect 1153 10635 1205 10641
rect 10336 10692 10540 10738
rect 24614 10742 24794 10748
rect 10336 10647 10388 10692
rect 10336 10583 10388 10595
rect 24666 10690 24678 10742
rect 24730 10690 24742 10742
rect 24614 10676 24794 10690
rect 24666 10624 24678 10676
rect 24730 10624 24742 10676
rect 27905 10645 28070 10791
rect 24614 10610 24794 10624
rect 24666 10558 24678 10610
rect 24730 10558 24742 10610
rect 24614 10551 24794 10558
rect 27284 10595 27433 10644
tri 27433 10595 27470 10632 sw
rect 27284 10589 27617 10595
rect 10336 10525 10388 10531
tri 24558 10525 24584 10551 ne
rect 24584 10543 24828 10551
rect 24584 10525 24614 10543
tri 24584 10495 24614 10525 ne
rect 24666 10491 24678 10543
rect 24730 10491 24742 10543
rect 24794 10535 24828 10543
tri 24828 10535 24844 10551 sw
rect 24614 10476 24794 10491
tri 24794 10485 24844 10535 nw
rect 27284 10537 27471 10589
rect 27523 10537 27565 10589
rect 27284 10494 27617 10537
rect 24666 10424 24678 10476
rect 24730 10424 24742 10476
rect 27284 10470 27471 10494
tri 27284 10436 27318 10470 ne
rect 27318 10442 27471 10470
rect 27523 10442 27565 10494
rect 27318 10436 27617 10442
rect 24614 10409 24794 10424
rect 24666 10357 24678 10409
rect 24730 10357 24742 10409
rect 24614 10351 24794 10357
rect 14195 10281 14201 10288
rect 13667 10241 14201 10281
rect 13667 10115 13707 10241
rect 14195 10236 14201 10241
rect 14253 10236 14265 10288
rect 14317 10236 14323 10288
rect 24635 9238 24641 9290
rect 24693 9238 24705 9290
rect 24757 9238 24763 9290
tri 23361 8128 23429 8196 ne
rect 23429 8128 23601 8196
tri 23601 8128 23669 8196 nw
tri 25677 8128 25745 8196 ne
rect 25745 8128 25896 8196
rect 22385 8099 22391 8128
rect 22263 8076 22391 8099
rect 22443 8076 22463 8128
rect 22515 8076 22535 8128
rect 22587 8076 22606 8128
rect 22658 8076 22677 8128
rect 22729 8076 22748 8128
rect 22800 8076 22819 8128
rect 22871 8076 22890 8128
rect 22942 8099 22948 8128
tri 23429 8121 23436 8128 ne
rect 23436 8121 23594 8128
tri 23594 8121 23601 8128 nw
tri 25745 8121 25752 8128 ne
rect 25752 8121 25896 8128
rect 22951 8099 23003 8121
tri 23003 8099 23025 8121 nw
tri 23436 8107 23450 8121 ne
rect 23450 8107 23580 8121
tri 23580 8107 23594 8121 nw
tri 25752 8107 25766 8121 ne
rect 25766 8107 25896 8121
tri 25896 8107 25985 8196 nw
rect 22942 8076 22952 8099
rect 22263 8054 22952 8076
rect 22263 8002 22391 8054
rect 22443 8002 22463 8054
rect 22515 8002 22535 8054
rect 22587 8002 22606 8054
rect 22658 8002 22677 8054
rect 22729 8002 22748 8054
rect 22800 8002 22819 8054
rect 22871 8002 22890 8054
rect 22942 8002 22952 8054
tri 22952 8048 23003 8099 nw
rect 14040 7870 14154 7988
rect 22263 7980 22952 8002
rect 22263 7928 22391 7980
rect 22443 7928 22463 7980
rect 22515 7928 22535 7980
rect 22587 7928 22606 7980
rect 22658 7928 22677 7980
rect 22729 7928 22748 7980
rect 22800 7928 22819 7980
rect 22871 7928 22890 7980
rect 22942 7928 22952 7980
tri 14064 7830 14104 7870 ne
rect 3815 7087 3821 7139
rect 3873 7087 3885 7139
rect 3937 7087 3943 7139
tri 12994 7038 13014 7058 se
rect 13014 7038 13142 7058
rect 12965 7006 13142 7038
tri 12986 6978 13014 7006 ne
rect 13014 6978 13142 7006
tri 13076 6953 13101 6978 ne
rect 2924 6402 2930 6454
rect 2982 6402 2995 6454
rect 2924 6390 2995 6402
rect 2924 6338 2930 6390
rect 2982 6338 2995 6390
rect 3239 6338 3245 6454
rect 258 6319 720 6323
tri 720 6319 724 6323 sw
rect 258 6285 724 6319
tri 724 6285 758 6319 sw
tri 13067 6285 13101 6319 se
rect 13101 6285 13142 6978
rect 14104 6390 14154 7870
rect 14026 6338 14032 6390
rect 14084 6338 14096 6390
rect 14148 6338 14154 6390
tri 13142 6285 13176 6319 sw
rect 258 6233 758 6285
tri 758 6233 810 6285 sw
rect 13059 6233 13065 6285
rect 13117 6233 13129 6285
rect 13181 6233 13187 6285
tri 23584 6276 23585 6277 se
rect 23585 6276 23591 6277
rect 258 6224 810 6233
tri 810 6224 819 6233 sw
rect 15635 6224 15641 6276
rect 15693 6224 15705 6276
rect 15757 6273 15763 6276
tri 15763 6273 15766 6276 sw
tri 23581 6273 23584 6276 se
rect 23584 6273 23591 6276
rect 15757 6227 23591 6273
rect 15757 6225 15764 6227
tri 15764 6225 15766 6227 nw
tri 23581 6225 23583 6227 ne
rect 23583 6225 23591 6227
rect 23643 6225 23655 6277
rect 23707 6225 23713 6277
rect 15757 6224 15763 6225
tri 15763 6224 15764 6225 nw
rect 258 6196 819 6224
tri 819 6196 847 6224 sw
rect 258 6175 847 6196
tri 847 6175 868 6196 sw
rect 5940 6195 6540 6196
rect 258 5956 720 6175
rect 5940 6143 5946 6195
rect 5998 6143 6013 6195
rect 6065 6143 6080 6195
rect 6132 6143 6147 6195
rect 6199 6143 6214 6195
rect 6266 6143 6281 6195
rect 6333 6143 6348 6195
rect 6400 6143 6415 6195
rect 6467 6143 6482 6195
rect 6534 6143 6540 6195
rect 5940 6121 6540 6143
rect 5940 6069 5946 6121
rect 5998 6069 6013 6121
rect 6065 6069 6080 6121
rect 6132 6069 6147 6121
rect 6199 6069 6214 6121
rect 6266 6069 6281 6121
rect 6333 6069 6348 6121
rect 6400 6069 6415 6121
rect 6467 6069 6482 6121
rect 6534 6069 6540 6121
rect 5940 6047 6540 6069
rect 5940 5995 5946 6047
rect 5998 5995 6013 6047
rect 6065 5995 6080 6047
rect 6132 5995 6147 6047
rect 6199 5995 6214 6047
rect 6266 5995 6281 6047
rect 6333 5995 6348 6047
rect 6400 5995 6415 6047
rect 6467 5995 6482 6047
rect 6534 5995 6540 6047
rect 12225 6195 12825 6196
rect 12225 6143 12231 6195
rect 12283 6143 12298 6195
rect 12350 6143 12365 6195
rect 12417 6143 12432 6195
rect 12484 6143 12499 6195
rect 12551 6143 12566 6195
rect 12618 6143 12633 6195
rect 12685 6143 12700 6195
rect 12752 6143 12767 6195
rect 12819 6143 12825 6195
rect 12225 6121 12825 6143
rect 12225 6069 12231 6121
rect 12283 6069 12298 6121
rect 12350 6069 12365 6121
rect 12417 6069 12432 6121
rect 12484 6069 12499 6121
rect 12551 6069 12566 6121
rect 12618 6069 12633 6121
rect 12685 6069 12700 6121
rect 12752 6069 12767 6121
rect 12819 6069 12825 6121
rect 12225 6047 12825 6069
rect 12225 5995 12231 6047
rect 12283 5995 12298 6047
rect 12350 5995 12365 6047
rect 12417 5995 12432 6047
rect 12484 5995 12499 6047
rect 12551 5995 12566 6047
rect 12618 5995 12633 6047
rect 12685 5995 12700 6047
rect 12752 5995 12767 6047
rect 12819 5995 12825 6047
rect 16057 6195 16657 6196
rect 16057 6143 16076 6195
rect 16128 6143 16142 6195
rect 16194 6143 16208 6195
rect 16260 6143 16274 6195
rect 16326 6143 16339 6195
rect 16391 6143 16404 6195
rect 16456 6143 16469 6195
rect 16521 6143 16534 6195
rect 16586 6143 16599 6195
rect 16651 6143 16657 6195
rect 16057 6121 16657 6143
rect 16057 6069 16076 6121
rect 16128 6069 16142 6121
rect 16194 6069 16208 6121
rect 16260 6069 16274 6121
rect 16326 6069 16339 6121
rect 16391 6069 16404 6121
rect 16456 6069 16469 6121
rect 16521 6069 16534 6121
rect 16586 6069 16599 6121
rect 16651 6069 16657 6121
rect 16057 6047 16657 6069
rect 16057 5995 16076 6047
rect 16128 5995 16142 6047
rect 16194 5995 16208 6047
rect 16260 5995 16274 6047
rect 16326 5995 16339 6047
rect 16391 5995 16404 6047
rect 16456 5995 16469 6047
rect 16521 5995 16534 6047
rect 16586 5995 16599 6047
rect 16651 5995 16657 6047
rect 20292 6195 20892 6196
rect 20292 6143 20298 6195
rect 20350 6143 20365 6195
rect 20417 6143 20432 6195
rect 20484 6143 20499 6195
rect 20551 6143 20566 6195
rect 20618 6143 20633 6195
rect 20685 6143 20700 6195
rect 20752 6143 20767 6195
rect 20819 6143 20834 6195
rect 20886 6143 20892 6195
rect 20292 6121 20892 6143
rect 20292 6069 20298 6121
rect 20350 6069 20365 6121
rect 20417 6069 20432 6121
rect 20484 6069 20499 6121
rect 20551 6069 20566 6121
rect 20618 6069 20633 6121
rect 20685 6069 20700 6121
rect 20752 6069 20767 6121
rect 20819 6069 20834 6121
rect 20886 6069 20892 6121
rect 20292 6047 20892 6069
rect 20292 5995 20298 6047
rect 20350 5995 20365 6047
rect 20417 5995 20432 6047
rect 20484 5995 20499 6047
rect 20551 5995 20566 6047
rect 20618 5995 20633 6047
rect 20685 5995 20700 6047
rect 20752 5995 20767 6047
rect 20819 5995 20834 6047
rect 20886 5995 20892 6047
rect 4040 5658 4314 5664
rect 4092 5606 4314 5658
rect 4040 5594 4314 5606
rect 4092 5542 4314 5594
rect 4040 5534 4314 5542
rect 7436 5496 8036 5498
rect 7436 5444 7442 5496
rect 7494 5444 7509 5496
rect 7561 5444 7576 5496
rect 7628 5444 7643 5496
rect 7695 5444 7710 5496
rect 7762 5444 7777 5496
rect 7829 5444 7844 5496
rect 7896 5444 7911 5496
rect 7963 5444 7978 5496
rect 8030 5444 8036 5496
rect 7436 5424 8036 5444
rect 7436 5372 7442 5424
rect 7494 5372 7509 5424
rect 7561 5372 7576 5424
rect 7628 5372 7643 5424
rect 7695 5372 7710 5424
rect 7762 5372 7777 5424
rect 7829 5372 7844 5424
rect 7896 5372 7911 5424
rect 7963 5372 7978 5424
rect 8030 5372 8036 5424
rect 7436 5352 8036 5372
rect 7436 5300 7442 5352
rect 7494 5300 7509 5352
rect 7561 5300 7576 5352
rect 7628 5300 7643 5352
rect 7695 5300 7710 5352
rect 7762 5300 7777 5352
rect 7829 5300 7844 5352
rect 7896 5300 7911 5352
rect 7963 5300 7978 5352
rect 8030 5300 8036 5352
rect 7436 5299 8036 5300
rect 11505 5496 12105 5498
rect 11505 5444 11511 5496
rect 11563 5444 11578 5496
rect 11630 5444 11645 5496
rect 11697 5444 11712 5496
rect 11764 5444 11779 5496
rect 11831 5444 11846 5496
rect 11898 5444 11913 5496
rect 11965 5444 11980 5496
rect 12032 5444 12047 5496
rect 12099 5444 12105 5496
rect 11505 5424 12105 5444
rect 11505 5372 11511 5424
rect 11563 5372 11578 5424
rect 11630 5372 11645 5424
rect 11697 5372 11712 5424
rect 11764 5372 11779 5424
rect 11831 5372 11846 5424
rect 11898 5372 11913 5424
rect 11965 5372 11980 5424
rect 12032 5372 12047 5424
rect 12099 5372 12105 5424
rect 11505 5352 12105 5372
rect 11505 5300 11511 5352
rect 11563 5300 11578 5352
rect 11630 5300 11645 5352
rect 11697 5300 11712 5352
rect 11764 5300 11779 5352
rect 11831 5300 11846 5352
rect 11898 5300 11913 5352
rect 11965 5300 11980 5352
rect 12032 5300 12047 5352
rect 12099 5300 12105 5352
rect 11505 5299 12105 5300
rect 14527 5496 15127 5498
rect 14527 5444 14533 5496
rect 14585 5444 14603 5496
rect 14655 5444 14672 5496
rect 14724 5444 14741 5496
rect 14793 5444 14810 5496
rect 14862 5444 14879 5496
rect 14931 5444 14948 5496
rect 15000 5444 15127 5496
rect 14527 5424 15127 5444
rect 14527 5372 14533 5424
rect 14585 5372 14603 5424
rect 14655 5372 14672 5424
rect 14724 5372 14741 5424
rect 14793 5372 14810 5424
rect 14862 5372 14879 5424
rect 14931 5372 14948 5424
rect 15000 5372 15127 5424
rect 14527 5352 15127 5372
rect 14527 5300 14533 5352
rect 14585 5300 14603 5352
rect 14655 5300 14672 5352
rect 14724 5300 14741 5352
rect 14793 5300 14810 5352
rect 14862 5300 14879 5352
rect 14931 5300 14948 5352
rect 15000 5300 15127 5352
rect 14527 5299 15127 5300
rect 16890 4433 16896 4485
rect 16948 4433 16975 4485
rect 17027 4433 17053 4485
rect 17105 4433 17131 4485
rect 17183 4433 17189 4485
rect 16890 4361 17189 4433
rect 16890 4309 16896 4361
rect 16948 4309 16975 4361
rect 17027 4309 17053 4361
rect 17105 4309 17131 4361
rect 17183 4309 17189 4361
rect 2820 4145 2826 4197
rect 2878 4145 2892 4197
rect 2944 4145 2957 4197
rect 3009 4145 3022 4197
rect 3074 4145 3087 4197
rect 3139 4145 3152 4197
rect 3204 4145 3210 4197
rect 2525 3779 2757 3791
rect 2820 3788 2826 3840
rect 2878 3788 2892 3840
rect 2944 3831 2957 3840
rect 3009 3831 3022 3840
rect 3074 3831 3087 3840
rect 2949 3797 2957 3831
rect 3074 3797 3081 3831
rect 2944 3788 2957 3797
rect 3009 3788 3022 3797
rect 3074 3788 3087 3797
rect 3139 3788 3152 3840
rect 3204 3788 3210 3840
rect 4040 3788 4046 3840
rect 4098 3788 4110 3840
rect 4162 3788 26139 3840
rect 26191 3788 26203 3840
rect 26255 3788 27827 3840
rect 2525 3745 2532 3779
rect 2566 3756 2624 3779
rect 2658 3756 2716 3779
rect 2750 3756 2757 3779
rect 2566 3745 2595 3756
rect 2658 3745 2705 3756
rect 2525 3704 2595 3745
rect 2647 3704 2705 3745
tri 3053 3708 3105 3760 se
rect 3105 3708 22552 3760
rect 22604 3708 22616 3760
rect 22668 3708 22674 3760
rect 22847 3708 23149 3760
rect 23201 3708 23213 3760
rect 23265 3708 26605 3760
rect 26657 3708 26669 3760
rect 26721 3708 27827 3760
rect 2525 3692 2757 3704
rect 2525 3658 2532 3692
rect 2566 3679 2624 3692
rect 2658 3679 2716 3692
rect 2750 3679 2757 3692
tri 3031 3686 3053 3708 se
rect 3053 3686 3105 3708
tri 3105 3686 3127 3708 nw
tri 3025 3680 3031 3686 se
rect 3031 3680 3099 3686
tri 3099 3680 3105 3686 nw
rect 2566 3658 2595 3679
rect 2658 3658 2705 3679
rect 2525 3627 2595 3658
rect 2647 3627 2705 3658
tri 2973 3628 3025 3680 se
rect 3025 3628 3047 3680
tri 3047 3628 3099 3680 nw
tri 3133 3628 3182 3677 se
rect 3182 3628 7609 3677
tri 7609 3628 7658 3677 sw
rect 7701 3628 7707 3680
rect 7759 3628 7771 3680
rect 7823 3628 20914 3680
rect 20966 3628 20978 3680
rect 21030 3628 21036 3680
rect 22847 3628 24059 3680
rect 24111 3628 24123 3680
rect 24175 3628 26731 3680
rect 26783 3628 26795 3680
rect 26847 3628 27827 3680
rect 2525 3605 2757 3627
tri 2957 3612 2973 3628 se
rect 2973 3612 3031 3628
tri 3031 3612 3047 3628 nw
tri 3117 3612 3133 3628 se
rect 3133 3625 7658 3628
rect 3133 3612 3182 3625
rect 2525 3571 2532 3605
rect 2566 3602 2624 3605
rect 2658 3602 2716 3605
rect 2750 3602 2757 3605
rect 2566 3571 2595 3602
rect 2658 3571 2705 3602
tri 2945 3600 2957 3612 se
rect 2957 3600 3019 3612
tri 3019 3600 3031 3612 nw
tri 3108 3603 3117 3612 se
rect 3117 3603 3182 3612
tri 3182 3603 3204 3625 nw
tri 7581 3603 7603 3625 ne
rect 7603 3612 7658 3625
tri 7658 3612 7674 3628 sw
rect 7603 3603 7674 3612
tri 3105 3600 3108 3603 se
rect 3108 3600 3179 3603
tri 3179 3600 3182 3603 nw
tri 7603 3600 7606 3603 ne
rect 7606 3600 7674 3603
tri 7674 3600 7686 3612 sw
rect 2525 3550 2595 3571
rect 2647 3550 2705 3571
tri 2906 3561 2945 3600 se
rect 2945 3561 2980 3600
tri 2980 3561 3019 3600 nw
tri 3066 3561 3105 3600 se
rect 3105 3597 3176 3600
tri 3176 3597 3179 3600 nw
tri 7606 3597 7609 3600 ne
rect 7609 3597 10415 3600
rect 3105 3563 3142 3597
tri 3142 3563 3176 3597 nw
tri 3182 3563 3216 3597 se
rect 3216 3585 7544 3597
tri 7544 3585 7556 3597 sw
tri 7609 3585 7621 3597 ne
rect 7621 3585 10415 3597
rect 3216 3563 7556 3585
rect 3105 3561 3140 3563
tri 3140 3561 3142 3563 nw
tri 3180 3561 3182 3563 se
rect 3182 3561 7556 3563
tri 7556 3561 7580 3585 sw
tri 7621 3561 7645 3585 ne
rect 7645 3561 10415 3585
rect 2525 3518 2757 3550
tri 2893 3548 2906 3561 se
rect 2906 3548 2967 3561
tri 2967 3548 2980 3561 nw
tri 3053 3548 3066 3561 se
rect 3066 3548 3127 3561
tri 3127 3548 3140 3561 nw
tri 3167 3548 3180 3561 se
rect 3180 3555 7580 3561
rect 3180 3548 3220 3555
tri 2883 3538 2893 3548 se
rect 2893 3538 2957 3548
tri 2957 3538 2967 3548 nw
tri 3043 3538 3053 3548 se
rect 3053 3538 3111 3548
tri 2877 3532 2883 3538 se
rect 2883 3532 2951 3538
tri 2951 3532 2957 3538 nw
tri 3037 3532 3043 3538 se
rect 3043 3532 3111 3538
tri 3111 3532 3127 3548 nw
tri 3151 3532 3167 3548 se
rect 3167 3532 3220 3548
tri 2872 3527 2877 3532 se
rect 2877 3527 2946 3532
tri 2946 3527 2951 3532 nw
tri 3034 3529 3037 3532 se
rect 3037 3529 3108 3532
tri 3108 3529 3111 3532 nw
tri 3148 3529 3151 3532 se
rect 3151 3529 3220 3532
tri 3032 3527 3034 3529 se
rect 3034 3527 3106 3529
tri 3106 3527 3108 3529 nw
tri 3146 3527 3148 3529 se
rect 3148 3527 3220 3529
tri 3220 3527 3248 3555 nw
tri 7506 3527 7534 3555 ne
rect 7534 3548 7580 3555
tri 7580 3548 7593 3561 sw
tri 7645 3548 7658 3561 ne
rect 7658 3548 10415 3561
rect 10467 3548 10479 3600
rect 10531 3548 10537 3600
rect 12107 3561 14804 3567
rect 7534 3532 7593 3548
tri 7593 3532 7609 3548 sw
rect 7534 3529 7609 3532
tri 7609 3529 7612 3532 sw
rect 7534 3527 7612 3529
tri 7612 3527 7614 3529 sw
rect 12107 3527 12119 3561
rect 12153 3527 12193 3561
rect 12227 3527 12267 3561
rect 12301 3527 12341 3561
rect 12375 3527 12415 3561
rect 12449 3527 12489 3561
rect 12523 3527 12563 3561
rect 12597 3527 12637 3561
rect 12671 3527 12711 3561
rect 12745 3527 12785 3561
rect 12819 3527 12859 3561
rect 12893 3527 12933 3561
rect 12967 3527 13006 3561
rect 13040 3527 13079 3561
rect 13113 3527 13152 3561
rect 13186 3527 13225 3561
rect 13259 3527 13298 3561
rect 13332 3527 13371 3561
rect 13405 3527 13444 3561
rect 13478 3527 13517 3561
rect 13551 3527 13590 3561
rect 13624 3527 13663 3561
rect 13697 3527 13736 3561
rect 13770 3527 13809 3561
rect 13843 3527 13882 3561
rect 13916 3527 13955 3561
rect 13989 3527 14028 3561
rect 14062 3527 14101 3561
rect 14135 3527 14174 3561
rect 14208 3527 14247 3561
rect 14281 3527 14320 3561
rect 14354 3527 14393 3561
rect 14427 3527 14466 3561
rect 14500 3527 14539 3561
rect 14573 3527 14612 3561
rect 14646 3527 14685 3561
rect 14719 3527 14758 3561
rect 14792 3527 14804 3561
tri 2865 3520 2872 3527 se
rect 2872 3520 2939 3527
tri 2939 3520 2946 3527 nw
tri 3025 3520 3032 3527 se
rect 3032 3523 3102 3527
tri 3102 3523 3106 3527 nw
tri 3142 3523 3146 3527 se
rect 3146 3523 3216 3527
tri 3216 3523 3220 3527 nw
tri 7534 3523 7538 3527 ne
rect 7538 3523 7614 3527
rect 3032 3520 3099 3523
tri 3099 3520 3102 3523 nw
tri 3139 3520 3142 3523 se
rect 3142 3520 3213 3523
tri 3213 3520 3216 3523 nw
tri 7538 3520 7541 3523 ne
rect 7541 3520 7614 3523
tri 7614 3520 7621 3527 sw
rect 2525 3484 2532 3518
rect 2566 3484 2624 3518
rect 2658 3484 2716 3518
rect 2750 3484 2757 3518
tri 2851 3506 2865 3520 se
rect 2865 3506 2925 3520
tri 2925 3506 2939 3520 nw
tri 3011 3506 3025 3520 se
rect 3025 3506 3085 3520
tri 3085 3506 3099 3520 nw
tri 3125 3506 3139 3520 se
rect 3139 3506 3199 3520
tri 3199 3506 3213 3520 nw
tri 7541 3517 7544 3520 ne
rect 7544 3517 11198 3520
tri 7544 3506 7555 3517 ne
rect 7555 3506 11198 3517
tri 2848 3503 2851 3506 se
rect 2851 3503 2922 3506
tri 2922 3503 2925 3506 nw
tri 3008 3503 3011 3506 se
rect 3011 3503 3082 3506
tri 3082 3503 3085 3506 nw
tri 3122 3503 3125 3506 se
rect 3125 3503 3196 3506
tri 3196 3503 3199 3506 nw
tri 7555 3503 7558 3506 ne
rect 7558 3503 11198 3506
rect 2525 3472 2757 3484
tri 2828 3483 2848 3503 se
rect 2848 3483 2902 3503
tri 2902 3483 2922 3503 nw
tri 2988 3483 3008 3503 se
rect 3008 3489 3068 3503
tri 3068 3489 3082 3503 nw
tri 3108 3489 3122 3503 se
rect 3122 3489 3176 3503
rect 3008 3483 3062 3489
tri 3062 3483 3068 3489 nw
tri 3102 3483 3108 3489 se
rect 3108 3483 3176 3489
tri 3176 3483 3196 3503 nw
rect 3337 3497 3595 3503
tri 2817 3472 2828 3483 se
rect 2828 3472 2883 3483
tri 2809 3464 2817 3472 se
rect 2817 3464 2883 3472
tri 2883 3464 2902 3483 nw
tri 2969 3464 2988 3483 se
rect 2988 3464 3034 3483
tri 2794 3449 2809 3464 se
rect 2809 3449 2868 3464
tri 2868 3449 2883 3464 nw
tri 2960 3455 2969 3464 se
rect 2969 3455 3034 3464
tri 3034 3455 3062 3483 nw
tri 3074 3455 3102 3483 se
rect 3102 3455 3142 3483
tri 2954 3449 2960 3455 se
rect 2960 3449 3028 3455
tri 3028 3449 3034 3455 nw
tri 3068 3449 3074 3455 se
rect 3074 3449 3142 3455
tri 3142 3449 3176 3483 nw
tri 2755 3410 2794 3449 se
rect 2794 3410 2829 3449
tri 2829 3410 2868 3449 nw
tri 2915 3410 2954 3449 se
rect 2954 3415 2994 3449
tri 2994 3415 3028 3449 nw
tri 3034 3415 3068 3449 se
rect 2954 3410 2960 3415
rect 904 3358 910 3410
rect 962 3358 974 3410
rect 1026 3381 2800 3410
tri 2800 3381 2829 3410 nw
tri 2886 3381 2915 3410 se
rect 2915 3381 2960 3410
tri 2960 3381 2994 3415 nw
tri 3000 3381 3034 3415 se
rect 3034 3381 3068 3415
rect 1026 3358 2777 3381
tri 2777 3358 2800 3381 nw
tri 2863 3358 2886 3381 se
rect 2886 3375 2954 3381
tri 2954 3375 2960 3381 nw
tri 2994 3375 3000 3381 se
rect 3000 3375 3068 3381
tri 3068 3375 3142 3449 nw
rect 3337 3445 3351 3497
rect 3403 3445 3415 3497
rect 3467 3445 3479 3497
rect 3531 3445 3543 3497
tri 7558 3483 7578 3503 ne
rect 7578 3483 11198 3503
tri 7578 3468 7593 3483 ne
rect 7593 3468 11198 3483
rect 11250 3468 11262 3520
rect 11314 3468 11917 3520
rect 11969 3468 11981 3520
rect 12033 3468 12039 3520
rect 12107 3483 14804 3527
rect 3337 3432 3595 3445
rect 12107 3449 12119 3483
rect 12153 3449 12193 3483
rect 12227 3449 12267 3483
rect 12301 3449 12341 3483
rect 12375 3449 12415 3483
rect 12449 3449 12489 3483
rect 12523 3449 12563 3483
rect 12597 3449 12637 3483
rect 12671 3449 12711 3483
rect 12745 3449 12785 3483
rect 12819 3449 12859 3483
rect 12893 3449 12933 3483
rect 12967 3449 13006 3483
rect 13040 3449 13079 3483
rect 13113 3449 13152 3483
rect 13186 3449 13225 3483
rect 13259 3449 13298 3483
rect 13332 3449 13371 3483
rect 13405 3449 13444 3483
rect 13478 3449 13517 3483
rect 13551 3449 13590 3483
rect 13624 3449 13663 3483
rect 13697 3449 13736 3483
rect 13770 3449 13809 3483
rect 13843 3449 13882 3483
rect 13916 3449 13955 3483
rect 13989 3449 14028 3483
rect 14062 3449 14101 3483
rect 14135 3449 14174 3483
rect 14208 3449 14247 3483
rect 14281 3449 14320 3483
rect 14354 3449 14393 3483
rect 14427 3449 14466 3483
rect 14500 3449 14539 3483
rect 14573 3449 14612 3483
rect 14646 3449 14685 3483
rect 14719 3449 14758 3483
rect 14792 3449 14804 3483
rect 14927 3480 14933 3532
rect 14985 3480 14997 3532
rect 15049 3520 16884 3532
tri 16884 3520 16896 3532 sw
rect 15049 3506 16896 3520
tri 16896 3506 16910 3520 sw
rect 15049 3480 16910 3506
tri 16910 3480 16936 3506 sw
rect 17074 3498 17080 3550
rect 17132 3498 17147 3550
rect 17199 3540 17214 3550
rect 17266 3540 17281 3550
rect 17333 3540 17348 3550
rect 17400 3540 17415 3550
rect 17467 3540 17482 3550
rect 17534 3540 17549 3550
rect 17200 3506 17214 3540
rect 17276 3506 17281 3540
rect 17467 3506 17470 3540
rect 17534 3506 17545 3540
rect 17199 3498 17214 3506
rect 17266 3498 17281 3506
rect 17333 3498 17348 3506
rect 17400 3498 17415 3506
rect 17467 3498 17482 3506
rect 17534 3498 17549 3506
rect 17601 3498 17616 3550
rect 17668 3498 17682 3550
rect 17734 3498 17748 3550
rect 17800 3540 17814 3550
rect 17866 3540 17880 3550
rect 17932 3540 17946 3550
rect 17998 3540 18012 3550
rect 18064 3540 18078 3550
rect 17804 3506 17814 3540
rect 17879 3506 17880 3540
rect 18064 3506 18070 3540
rect 17800 3498 17814 3506
rect 17866 3498 17880 3506
rect 17932 3498 17946 3506
rect 17998 3498 18012 3506
rect 18064 3498 18078 3506
rect 18130 3498 18144 3550
rect 18196 3498 18210 3550
rect 18262 3498 18276 3550
rect 18328 3540 18342 3550
rect 18394 3540 18408 3550
rect 18460 3540 18474 3550
rect 18526 3540 18540 3550
rect 18592 3540 18606 3550
rect 18658 3540 18672 3550
rect 18329 3506 18342 3540
rect 18404 3506 18408 3540
rect 18592 3506 18595 3540
rect 18658 3506 18670 3540
rect 18328 3498 18342 3506
rect 18394 3498 18408 3506
rect 18460 3498 18474 3506
rect 18526 3498 18540 3506
rect 18592 3498 18606 3506
rect 18658 3498 18672 3506
rect 18724 3498 18730 3550
rect 20279 3548 20285 3600
rect 20337 3548 20349 3600
rect 20401 3548 22414 3600
rect 22466 3548 22478 3600
rect 22530 3548 22640 3600
rect 26289 3548 26898 3600
rect 26950 3548 26962 3600
rect 27014 3548 27295 3600
rect 27347 3548 27359 3600
rect 27411 3548 27827 3600
tri 16826 3452 16854 3480 ne
rect 16854 3468 16936 3480
tri 16936 3468 16948 3480 sw
rect 18997 3468 19003 3520
rect 19055 3468 19067 3520
rect 19119 3468 22310 3520
rect 22362 3468 22374 3520
rect 22426 3468 22432 3520
rect 22847 3468 22853 3520
rect 22905 3468 22917 3520
rect 22969 3468 26227 3520
rect 26279 3468 26291 3520
rect 26343 3468 27827 3520
rect 16854 3452 16948 3468
tri 16948 3452 16964 3468 sw
rect 3337 3380 3351 3432
rect 3403 3380 3415 3432
rect 3467 3380 3479 3432
rect 3531 3380 3543 3432
rect 2886 3358 2920 3375
tri 2833 3328 2863 3358 se
rect 2863 3341 2920 3358
tri 2920 3341 2954 3375 nw
tri 2960 3341 2994 3375 se
rect 2863 3328 2886 3341
rect 703 3322 755 3328
tri 669 3250 703 3284 se
tri 2812 3307 2833 3328 se
rect 2833 3307 2886 3328
tri 2886 3307 2920 3341 nw
tri 2926 3307 2960 3341 se
rect 2960 3307 2994 3341
tri 2789 3284 2812 3307 se
rect 2812 3301 2880 3307
tri 2880 3301 2886 3307 nw
tri 2920 3301 2926 3307 se
rect 2926 3301 2994 3307
tri 2994 3301 3068 3375 nw
rect 3337 3367 3595 3380
rect 3337 3315 3351 3367
rect 3403 3315 3415 3367
rect 3467 3315 3479 3367
rect 3531 3315 3543 3367
rect 3337 3302 3595 3315
rect 7670 3341 7676 3393
rect 7728 3341 7740 3393
rect 7792 3388 7798 3393
tri 7798 3388 7803 3393 sw
rect 8070 3388 8076 3440
rect 8128 3388 8140 3440
rect 8192 3388 10711 3440
rect 10763 3388 10775 3440
rect 10827 3388 10833 3440
tri 11376 3388 11418 3430 se
rect 11418 3388 11621 3430
rect 7792 3378 7803 3388
tri 7803 3378 7813 3388 sw
tri 11366 3378 11376 3388 se
rect 11376 3378 11621 3388
rect 11673 3378 11685 3430
rect 11737 3378 11743 3430
rect 7792 3360 7813 3378
tri 7813 3360 7831 3378 sw
tri 11348 3360 11366 3378 se
rect 11366 3360 11422 3378
tri 11422 3360 11440 3378 nw
rect 12107 3360 14804 3449
rect 14927 3400 15843 3452
rect 15895 3400 15907 3452
rect 15959 3440 16778 3452
tri 16778 3440 16790 3452 sw
tri 16854 3440 16866 3452 ne
rect 16866 3440 16964 3452
tri 16964 3440 16976 3452 sw
rect 15959 3422 16790 3440
tri 16790 3422 16808 3440 sw
tri 16866 3422 16884 3440 ne
rect 16884 3422 22204 3440
rect 15959 3400 16808 3422
tri 16723 3374 16749 3400 ne
rect 16749 3388 16808 3400
tri 16808 3388 16842 3422 sw
tri 16884 3388 16918 3422 ne
rect 16918 3388 22204 3422
rect 22256 3388 22268 3440
rect 22320 3388 22326 3440
rect 22676 3388 24355 3440
rect 24407 3388 24419 3440
rect 24471 3388 26353 3440
rect 26405 3388 26417 3440
rect 26469 3388 27730 3440
rect 27782 3388 27794 3440
rect 27846 3388 27852 3440
rect 16749 3374 16842 3388
tri 14804 3360 14818 3374 sw
tri 16749 3360 16763 3374 ne
rect 16763 3360 16842 3374
tri 16842 3360 16870 3388 sw
rect 7792 3345 11407 3360
tri 11407 3345 11422 3360 nw
rect 12107 3345 14818 3360
tri 14818 3345 14833 3360 sw
tri 16763 3345 16778 3360 ne
rect 16778 3345 22096 3360
rect 7792 3341 11374 3345
rect 7670 3312 11374 3341
tri 11374 3312 11407 3345 nw
tri 12075 3312 12107 3344 se
rect 12107 3312 14833 3345
tri 14833 3312 14866 3345 sw
tri 16778 3312 16811 3345 ne
rect 16811 3312 22096 3345
rect 7670 3308 11370 3312
tri 11370 3308 11374 3312 nw
tri 12071 3308 12075 3312 se
rect 12075 3308 14866 3312
tri 14866 3308 14870 3312 sw
tri 22085 3308 22089 3312 ne
rect 22089 3308 22096 3312
rect 22148 3308 22160 3360
rect 22212 3308 22218 3360
rect 26513 3308 26520 3360
rect 26572 3308 26584 3360
rect 26636 3308 27495 3360
rect 27547 3308 27559 3360
rect 27611 3308 27617 3360
rect 2812 3284 2846 3301
rect 703 3258 755 3270
rect 622 3206 703 3250
tri 755 3250 789 3284 sw
tri 2755 3250 2789 3284 se
rect 2789 3267 2846 3284
tri 2846 3267 2880 3301 nw
tri 2886 3267 2920 3301 se
rect 2789 3250 2829 3267
tri 2829 3250 2846 3267 nw
tri 2869 3250 2886 3267 se
rect 2886 3250 2920 3267
rect 755 3227 2806 3250
tri 2806 3227 2829 3250 nw
tri 2846 3227 2869 3250 se
rect 2869 3227 2920 3250
tri 2920 3227 2994 3301 nw
rect 3337 3250 3351 3302
rect 3403 3250 3415 3302
rect 3467 3250 3479 3302
rect 3531 3250 3543 3302
tri 12043 3280 12071 3308 se
rect 12071 3280 14870 3308
rect 14741 3279 14870 3280
tri 14870 3279 14899 3308 sw
rect 3337 3237 3595 3250
rect 755 3210 2789 3227
tri 2789 3210 2806 3227 nw
tri 2829 3210 2846 3227 se
rect 2846 3210 2863 3227
rect 755 3206 2777 3210
rect 622 3198 2777 3206
tri 2777 3198 2789 3210 nw
tri 2817 3198 2829 3210 se
rect 2829 3198 2863 3210
tri 2789 3170 2817 3198 se
rect 2817 3170 2863 3198
tri 2863 3170 2920 3227 nw
rect 3337 3185 3351 3237
rect 3403 3185 3415 3237
rect 3467 3185 3479 3237
rect 3531 3185 3543 3237
rect 3337 3172 3595 3185
rect 463 3140 2811 3170
rect 463 3118 1760 3140
rect 1812 3118 2811 3140
tri 2811 3118 2863 3170 nw
rect 3337 3120 3351 3172
rect 3403 3120 3415 3172
rect 3467 3120 3479 3172
rect 3531 3120 3543 3172
rect 3337 3106 3595 3120
rect 1760 3076 1812 3088
rect 1165 3056 1217 3062
tri 1217 3018 1218 3019 sw
rect 1760 3018 1812 3024
rect 2547 3084 2599 3090
rect 2547 3020 2599 3032
tri 2546 3018 2547 3019 se
rect 1217 3004 1218 3018
rect 1165 2992 1218 3004
rect 1217 2985 1218 2992
tri 1218 2985 1251 3018 sw
tri 2513 2985 2546 3018 se
rect 2546 2985 2547 3018
rect 1217 2968 2547 2985
rect 1217 2962 2599 2968
rect 1217 2940 2571 2962
rect 1165 2934 2571 2940
tri 2571 2934 2599 2962 nw
rect 3337 3054 3351 3106
rect 3403 3054 3415 3106
rect 3467 3054 3479 3106
rect 3531 3054 3543 3106
rect 3337 3040 3595 3054
rect 3337 2988 3351 3040
rect 3403 2988 3415 3040
rect 3467 2988 3479 3040
rect 3531 2988 3543 3040
rect 3337 2974 3595 2988
rect 1165 2933 2570 2934
tri 2570 2933 2571 2934 nw
rect 3337 2922 3351 2974
rect 3403 2922 3415 2974
rect 3467 2922 3479 2974
rect 3531 2922 3543 2974
rect 3337 2908 3595 2922
rect 1217 2891 2600 2892
rect 1165 2839 1171 2891
rect 1223 2839 1235 2891
rect 1287 2886 2600 2891
rect 1287 2840 2548 2886
rect 1287 2839 1293 2840
tri 2514 2839 2515 2840 ne
rect 2515 2839 2548 2840
tri 2515 2806 2548 2839 ne
rect 2548 2822 2600 2834
rect 3337 2856 3351 2908
rect 3403 2856 3415 2908
rect 3467 2856 3479 2908
rect 3531 2856 3543 2908
rect 3337 2842 3595 2856
rect 3337 2790 3351 2842
rect 3403 2790 3415 2842
rect 3467 2790 3479 2842
rect 3531 2790 3543 2842
rect 3337 2784 3595 2790
rect 2548 2764 2600 2770
rect 3592 2121 3644 2127
rect 3592 2057 3644 2069
rect 3592 1999 3644 2005
rect 23253 2059 23447 2065
rect 23253 2007 23254 2059
rect 23306 2007 23324 2059
rect 23376 2007 23394 2059
rect 23446 2007 23447 2059
rect 3595 1997 3641 1999
rect 23253 1989 23447 2007
rect 23253 1937 23254 1989
rect 23306 1937 23324 1989
rect 23376 1937 23394 1989
rect 23446 1937 23447 1989
rect 23253 1919 23447 1937
rect 23253 1867 23254 1919
rect 23306 1867 23324 1919
rect 23376 1867 23394 1919
rect 23446 1867 23447 1919
rect 23253 1849 23447 1867
rect 1934 1835 2050 1841
rect 1986 1783 1998 1835
rect 1934 1770 2050 1783
rect 1986 1718 1998 1770
rect 23253 1797 23254 1849
rect 23306 1797 23324 1849
rect 23376 1797 23394 1849
rect 23446 1797 23447 1849
rect 23253 1778 23447 1797
rect 23253 1726 23254 1778
rect 23306 1726 23324 1778
rect 23376 1726 23394 1778
rect 23446 1726 23447 1778
rect 23253 1720 23447 1726
rect 1761 1705 1813 1711
rect 1761 1641 1813 1653
rect 1761 1583 1813 1589
rect 1934 1705 2050 1718
rect 1986 1653 1998 1705
rect 1934 1640 2050 1653
rect 1986 1588 1998 1640
rect 1934 1575 2050 1588
rect 1986 1523 1998 1575
rect 1934 1510 2050 1523
rect 1986 1458 1998 1510
rect 1934 1445 2050 1458
rect 1986 1393 1998 1445
rect 1934 1380 2050 1393
rect 1986 1328 1998 1380
rect 1934 1315 2050 1328
rect 1986 1263 1998 1315
rect 1934 1250 2050 1263
rect 1986 1198 1998 1250
rect 1934 1185 2050 1198
rect 1986 1133 1998 1185
rect 1934 1120 2050 1133
rect 1986 1068 1998 1120
rect 23782 1182 23788 1234
rect 23840 1182 23852 1234
rect 23904 1182 23916 1234
rect 23968 1182 23974 1234
rect 23782 1140 23974 1182
rect 23782 1088 23788 1140
rect 23840 1088 23852 1140
rect 23904 1088 23916 1140
rect 23968 1088 23974 1140
rect 1934 1055 2050 1068
rect 1986 1003 1998 1055
rect 1934 990 2050 1003
rect 1986 938 1998 990
rect 1934 925 2050 938
rect 1986 873 1998 925
rect 1934 860 2050 873
rect 1986 808 1998 860
rect 1934 795 2050 808
rect 1986 743 1998 795
rect 1934 730 2050 743
rect 1986 678 1998 730
rect 1934 664 2050 678
rect 1986 612 1998 664
rect 1934 598 2050 612
rect 1986 546 1998 598
rect 1934 532 2050 546
rect 1986 480 1998 532
rect 1934 466 2050 480
rect 1986 414 1998 466
rect 1934 408 2050 414
rect 4004 211 4056 217
rect 18259 178 18265 230
rect 18317 178 18336 230
rect 18388 178 18407 230
rect 18459 178 18477 230
rect 18529 178 18535 230
rect 4004 147 4056 159
rect 4004 89 4056 95
<< via1 >>
rect 12004 38680 12056 38732
rect 12073 38680 12125 38732
rect 12142 38680 12194 38732
rect 12211 38680 12263 38732
rect 12280 38680 12332 38732
rect 12348 38680 12400 38732
rect 12004 38608 12056 38660
rect 12073 38608 12125 38660
rect 12142 38608 12194 38660
rect 12211 38608 12263 38660
rect 12280 38608 12332 38660
rect 12348 38608 12400 38660
rect 12004 38536 12056 38588
rect 12073 38536 12125 38588
rect 12142 38536 12194 38588
rect 12211 38536 12263 38588
rect 12280 38536 12332 38588
rect 12348 38536 12400 38588
rect 25743 37825 25795 37877
rect 25807 37825 25859 37877
rect 26770 37572 26822 37624
rect 26834 37572 26886 37624
rect 3128 33126 3180 33178
rect 3199 33126 3251 33178
rect 3271 33126 3323 33178
rect 3128 33058 3180 33110
rect 3199 33058 3251 33110
rect 3271 33058 3323 33110
rect 2885 32649 2937 32654
rect 2972 32649 3024 32654
rect 3059 32649 3111 32654
rect 2885 32602 2937 32649
rect 2972 32602 3024 32649
rect 3059 32602 3105 32649
rect 3105 32602 3111 32649
rect 2885 32543 2937 32590
rect 2972 32543 3024 32590
rect 3059 32543 3105 32590
rect 3105 32543 3111 32590
rect 2885 32538 2937 32543
rect 2972 32538 3024 32543
rect 3059 32538 3111 32543
rect 2036 31898 2088 31950
rect 2140 31898 2192 31950
rect 2036 31830 2088 31882
rect 2140 31830 2192 31882
rect 2036 31762 2088 31814
rect 2140 31762 2192 31814
rect 1667 31063 1719 31115
rect 1751 31063 1803 31115
rect 1835 31063 1887 31115
rect 1667 30984 1719 31036
rect 1751 30984 1803 31036
rect 1835 30984 1887 31036
rect 1667 30905 1719 30957
rect 1751 30905 1803 30957
rect 1835 30905 1887 30957
rect 1667 30826 1719 30878
rect 1751 30826 1803 30878
rect 1835 30826 1887 30878
rect 27050 23250 27054 23276
rect 27054 23250 27088 23276
rect 27088 23250 27102 23276
rect 27050 23224 27102 23250
rect 27121 23250 27126 23276
rect 27126 23250 27160 23276
rect 27160 23250 27173 23276
rect 27121 23224 27173 23250
rect 27192 23250 27198 23276
rect 27198 23250 27232 23276
rect 27232 23250 27244 23276
rect 27192 23224 27244 23250
rect 27262 23250 27270 23276
rect 27270 23250 27304 23276
rect 27304 23250 27314 23276
rect 27262 23224 27314 23250
rect 27332 23250 27342 23276
rect 27342 23250 27376 23276
rect 27376 23250 27384 23276
rect 27332 23224 27384 23250
rect 27402 23250 27414 23276
rect 27414 23250 27448 23276
rect 27448 23250 27454 23276
rect 27402 23224 27454 23250
rect 27472 23250 27486 23276
rect 27486 23250 27520 23276
rect 27520 23250 27524 23276
rect 27472 23224 27524 23250
rect 27542 23250 27558 23276
rect 27558 23250 27592 23276
rect 27592 23250 27594 23276
rect 27542 23224 27594 23250
rect 27612 23250 27630 23276
rect 27630 23250 27664 23276
rect 27612 23224 27664 23250
rect 27050 23198 27102 23210
rect 27050 23164 27054 23198
rect 27054 23164 27088 23198
rect 27088 23164 27102 23198
rect 27050 23158 27102 23164
rect 27121 23198 27173 23210
rect 27121 23164 27126 23198
rect 27126 23164 27160 23198
rect 27160 23164 27173 23198
rect 27121 23158 27173 23164
rect 27192 23198 27244 23210
rect 27192 23164 27198 23198
rect 27198 23164 27232 23198
rect 27232 23164 27244 23198
rect 27192 23158 27244 23164
rect 27262 23198 27314 23210
rect 27262 23164 27270 23198
rect 27270 23164 27304 23198
rect 27304 23164 27314 23198
rect 27262 23158 27314 23164
rect 27332 23198 27384 23210
rect 27332 23164 27342 23198
rect 27342 23164 27376 23198
rect 27376 23164 27384 23198
rect 27332 23158 27384 23164
rect 27402 23198 27454 23210
rect 27402 23164 27414 23198
rect 27414 23164 27448 23198
rect 27448 23164 27454 23198
rect 27402 23158 27454 23164
rect 27472 23198 27524 23210
rect 27472 23164 27486 23198
rect 27486 23164 27520 23198
rect 27520 23164 27524 23198
rect 27472 23158 27524 23164
rect 27542 23198 27594 23210
rect 27542 23164 27558 23198
rect 27558 23164 27592 23198
rect 27592 23164 27594 23198
rect 27542 23158 27594 23164
rect 27612 23198 27664 23210
rect 27612 23164 27630 23198
rect 27630 23164 27664 23198
rect 27612 23158 27664 23164
rect 27050 23112 27102 23144
rect 27050 23092 27054 23112
rect 27054 23092 27088 23112
rect 27088 23092 27102 23112
rect 27121 23112 27173 23144
rect 27121 23092 27126 23112
rect 27126 23092 27160 23112
rect 27160 23092 27173 23112
rect 27192 23112 27244 23144
rect 27192 23092 27198 23112
rect 27198 23092 27232 23112
rect 27232 23092 27244 23112
rect 27262 23112 27314 23144
rect 27262 23092 27270 23112
rect 27270 23092 27304 23112
rect 27304 23092 27314 23112
rect 27332 23112 27384 23144
rect 27332 23092 27342 23112
rect 27342 23092 27376 23112
rect 27376 23092 27384 23112
rect 27402 23112 27454 23144
rect 27402 23092 27414 23112
rect 27414 23092 27448 23112
rect 27448 23092 27454 23112
rect 27472 23112 27524 23144
rect 27472 23092 27486 23112
rect 27486 23092 27520 23112
rect 27520 23092 27524 23112
rect 27542 23112 27594 23144
rect 27542 23092 27558 23112
rect 27558 23092 27592 23112
rect 27592 23092 27594 23112
rect 27612 23112 27664 23144
rect 27612 23092 27630 23112
rect 27630 23092 27664 23112
rect 27050 23026 27102 23078
rect 27121 23026 27173 23078
rect 27192 23026 27244 23078
rect 27262 23026 27314 23078
rect 27332 23026 27384 23078
rect 27402 23026 27454 23078
rect 27472 23026 27524 23078
rect 27542 23026 27594 23078
rect 27612 23026 27664 23078
rect 27050 22992 27054 23012
rect 27054 22992 27088 23012
rect 27088 22992 27102 23012
rect 27050 22960 27102 22992
rect 27121 22992 27126 23012
rect 27126 22992 27160 23012
rect 27160 22992 27173 23012
rect 27121 22960 27173 22992
rect 27192 22992 27198 23012
rect 27198 22992 27232 23012
rect 27232 22992 27244 23012
rect 27192 22960 27244 22992
rect 27262 22992 27270 23012
rect 27270 22992 27304 23012
rect 27304 22992 27314 23012
rect 27262 22960 27314 22992
rect 27332 22992 27342 23012
rect 27342 22992 27376 23012
rect 27376 22992 27384 23012
rect 27332 22960 27384 22992
rect 27402 22992 27414 23012
rect 27414 22992 27448 23012
rect 27448 22992 27454 23012
rect 27402 22960 27454 22992
rect 27472 22992 27486 23012
rect 27486 22992 27520 23012
rect 27520 22992 27524 23012
rect 27472 22960 27524 22992
rect 27542 22992 27558 23012
rect 27558 22992 27592 23012
rect 27592 22992 27594 23012
rect 27542 22960 27594 22992
rect 27612 22992 27630 23012
rect 27630 22992 27664 23012
rect 27612 22960 27664 22992
rect 27050 22894 27102 22946
rect 27121 22894 27173 22946
rect 27192 22894 27244 22946
rect 27262 22894 27314 22946
rect 27332 22894 27384 22946
rect 27402 22894 27454 22946
rect 27472 22894 27524 22946
rect 27542 22894 27594 22946
rect 27612 22894 27664 22946
rect 27355 22856 27360 22861
rect 27360 22856 27400 22861
rect 27400 22856 27407 22861
rect 27419 22856 27434 22861
rect 27434 22856 27471 22861
rect 27483 22856 27508 22861
rect 27508 22856 27535 22861
rect 27355 22818 27407 22856
rect 27419 22818 27471 22856
rect 27483 22818 27535 22856
rect 27355 22809 27360 22818
rect 27360 22809 27400 22818
rect 27400 22809 27407 22818
rect 27419 22809 27434 22818
rect 27434 22809 27471 22818
rect 27483 22809 27508 22818
rect 27508 22809 27535 22818
rect 27547 22856 27548 22861
rect 27548 22856 27582 22861
rect 27582 22856 27599 22861
rect 27547 22818 27599 22856
rect 27547 22809 27548 22818
rect 27548 22809 27582 22818
rect 27582 22809 27599 22818
rect 27611 22856 27622 22861
rect 27622 22856 27656 22861
rect 27656 22856 27663 22861
rect 27611 22818 27663 22856
rect 27611 22809 27622 22818
rect 27622 22809 27656 22818
rect 27656 22809 27663 22818
rect 27355 22784 27360 22794
rect 27360 22784 27400 22794
rect 27400 22784 27407 22794
rect 27419 22784 27434 22794
rect 27434 22784 27471 22794
rect 27483 22784 27508 22794
rect 27508 22784 27535 22794
rect 27355 22746 27407 22784
rect 27419 22746 27471 22784
rect 27483 22746 27535 22784
rect 27355 22742 27360 22746
rect 27360 22742 27400 22746
rect 27400 22742 27407 22746
rect 27419 22742 27434 22746
rect 27434 22742 27471 22746
rect 27483 22742 27508 22746
rect 27508 22742 27535 22746
rect 27547 22784 27548 22794
rect 27548 22784 27582 22794
rect 27582 22784 27599 22794
rect 27547 22746 27599 22784
rect 27547 22742 27548 22746
rect 27548 22742 27582 22746
rect 27582 22742 27599 22746
rect 27611 22784 27622 22794
rect 27622 22784 27656 22794
rect 27656 22784 27663 22794
rect 27611 22746 27663 22784
rect 27611 22742 27622 22746
rect 27622 22742 27656 22746
rect 27656 22742 27663 22746
rect 27355 22712 27360 22727
rect 27360 22712 27400 22727
rect 27400 22712 27407 22727
rect 27419 22712 27434 22727
rect 27434 22712 27471 22727
rect 27483 22712 27508 22727
rect 27508 22712 27535 22727
rect 27355 22675 27407 22712
rect 27419 22675 27471 22712
rect 27483 22675 27535 22712
rect 27547 22712 27548 22727
rect 27548 22712 27582 22727
rect 27582 22712 27599 22727
rect 27547 22675 27599 22712
rect 27611 22712 27622 22727
rect 27622 22712 27656 22727
rect 27656 22712 27663 22727
rect 27611 22675 27663 22712
rect 27355 22640 27360 22660
rect 27360 22640 27400 22660
rect 27400 22640 27407 22660
rect 27419 22640 27434 22660
rect 27434 22640 27471 22660
rect 27483 22640 27508 22660
rect 27508 22640 27535 22660
rect 27355 22608 27407 22640
rect 27419 22608 27471 22640
rect 27483 22608 27535 22640
rect 27547 22640 27548 22660
rect 27548 22640 27582 22660
rect 27582 22640 27599 22660
rect 27547 22608 27599 22640
rect 27611 22640 27622 22660
rect 27622 22640 27656 22660
rect 27656 22640 27663 22660
rect 27611 22608 27663 22640
rect 27355 22568 27360 22593
rect 27360 22568 27400 22593
rect 27400 22568 27407 22593
rect 27419 22568 27434 22593
rect 27434 22568 27471 22593
rect 27483 22568 27508 22593
rect 27508 22568 27535 22593
rect 27355 22541 27407 22568
rect 27419 22541 27471 22568
rect 27483 22541 27535 22568
rect 27547 22568 27548 22593
rect 27548 22568 27582 22593
rect 27582 22568 27599 22593
rect 27547 22541 27599 22568
rect 27611 22568 27622 22593
rect 27622 22568 27656 22593
rect 27656 22568 27663 22593
rect 27611 22541 27663 22568
rect 27355 22496 27360 22526
rect 27360 22496 27400 22526
rect 27400 22496 27407 22526
rect 27419 22496 27434 22526
rect 27434 22496 27471 22526
rect 27483 22496 27508 22526
rect 27508 22496 27535 22526
rect 27355 22474 27407 22496
rect 27419 22474 27471 22496
rect 27483 22474 27535 22496
rect 27547 22496 27548 22526
rect 27548 22496 27582 22526
rect 27582 22496 27599 22526
rect 27547 22474 27599 22496
rect 27611 22496 27622 22526
rect 27622 22496 27656 22526
rect 27656 22496 27663 22526
rect 27611 22474 27663 22496
rect 27355 22458 27407 22459
rect 27419 22458 27471 22459
rect 27483 22458 27535 22459
rect 27355 22424 27360 22458
rect 27360 22424 27400 22458
rect 27400 22424 27407 22458
rect 27419 22424 27434 22458
rect 27434 22424 27471 22458
rect 27483 22424 27508 22458
rect 27508 22424 27535 22458
rect 27355 22407 27407 22424
rect 27419 22407 27471 22424
rect 27483 22407 27535 22424
rect 27547 22458 27599 22459
rect 27547 22424 27548 22458
rect 27548 22424 27582 22458
rect 27582 22424 27599 22458
rect 27547 22407 27599 22424
rect 27611 22458 27663 22459
rect 27611 22424 27622 22458
rect 27622 22424 27656 22458
rect 27656 22424 27663 22458
rect 27611 22407 27663 22424
rect 27355 22386 27407 22392
rect 27419 22386 27471 22392
rect 27483 22386 27535 22392
rect 27355 22352 27360 22386
rect 27360 22352 27400 22386
rect 27400 22352 27407 22386
rect 27419 22352 27434 22386
rect 27434 22352 27471 22386
rect 27483 22352 27508 22386
rect 27508 22352 27535 22386
rect 27355 22340 27407 22352
rect 27419 22340 27471 22352
rect 27483 22340 27535 22352
rect 27547 22386 27599 22392
rect 27547 22352 27548 22386
rect 27548 22352 27582 22386
rect 27582 22352 27599 22386
rect 27547 22340 27599 22352
rect 27611 22386 27663 22392
rect 27611 22352 27622 22386
rect 27622 22352 27656 22386
rect 27656 22352 27663 22386
rect 27611 22340 27663 22352
rect 27355 22314 27407 22324
rect 27419 22314 27471 22324
rect 27483 22314 27535 22324
rect 27355 22280 27360 22314
rect 27360 22280 27400 22314
rect 27400 22280 27407 22314
rect 27419 22280 27434 22314
rect 27434 22280 27471 22314
rect 27483 22280 27508 22314
rect 27508 22280 27535 22314
rect 27355 22272 27407 22280
rect 27419 22272 27471 22280
rect 27483 22272 27535 22280
rect 27547 22314 27599 22324
rect 27547 22280 27548 22314
rect 27548 22280 27582 22314
rect 27582 22280 27599 22314
rect 27547 22272 27599 22280
rect 27611 22314 27663 22324
rect 27611 22280 27622 22314
rect 27622 22280 27656 22314
rect 27656 22280 27663 22314
rect 27611 22272 27663 22280
rect 27355 22242 27407 22256
rect 27419 22242 27471 22256
rect 27483 22242 27535 22256
rect 27355 22208 27360 22242
rect 27360 22208 27400 22242
rect 27400 22208 27407 22242
rect 27419 22208 27434 22242
rect 27434 22208 27471 22242
rect 27483 22208 27508 22242
rect 27508 22208 27535 22242
rect 27355 22204 27407 22208
rect 27419 22204 27471 22208
rect 27483 22204 27535 22208
rect 27547 22242 27599 22256
rect 27547 22208 27548 22242
rect 27548 22208 27582 22242
rect 27582 22208 27599 22242
rect 27547 22204 27599 22208
rect 27611 22242 27663 22256
rect 27611 22208 27622 22242
rect 27622 22208 27656 22242
rect 27656 22208 27663 22242
rect 27611 22204 27663 22208
rect 27355 22170 27407 22188
rect 27419 22170 27471 22188
rect 27483 22170 27535 22188
rect 27355 22136 27360 22170
rect 27360 22136 27400 22170
rect 27400 22136 27407 22170
rect 27419 22136 27434 22170
rect 27434 22136 27471 22170
rect 27483 22136 27508 22170
rect 27508 22136 27535 22170
rect 27547 22170 27599 22188
rect 27547 22136 27548 22170
rect 27548 22136 27582 22170
rect 27582 22136 27599 22170
rect 27611 22170 27663 22188
rect 27611 22136 27622 22170
rect 27622 22136 27656 22170
rect 27656 22136 27663 22170
rect 1836 21312 1888 21364
rect 1908 21312 1960 21364
rect 1836 21248 1888 21300
rect 1908 21248 1960 21300
rect 1836 21184 1888 21236
rect 1908 21184 1960 21236
rect 27364 21323 27416 21375
rect 27428 21323 27480 21375
rect 27364 21217 27416 21269
rect 27428 21217 27480 21269
rect 27515 21315 27567 21367
rect 27621 21315 27673 21367
rect 27515 21236 27567 21288
rect 27621 21236 27673 21288
rect 1836 21120 1888 21172
rect 1908 21120 1960 21172
rect 27515 21157 27567 21209
rect 27621 21157 27673 21209
rect 1836 21056 1888 21108
rect 1908 21056 1960 21108
rect 1836 20992 1888 21044
rect 1908 20992 1960 21044
rect 1836 20928 1888 20980
rect 1908 20928 1960 20980
rect 1836 20864 1888 20916
rect 1908 20864 1960 20916
rect 1836 20800 1888 20852
rect 1908 20800 1960 20852
rect 1836 20736 1888 20788
rect 1908 20736 1960 20788
rect 1836 20672 1888 20724
rect 1908 20672 1960 20724
rect 1836 20608 1888 20660
rect 1908 20608 1960 20660
rect 1836 20544 1888 20596
rect 1908 20544 1960 20596
rect 1836 20480 1888 20532
rect 1908 20480 1960 20532
rect 1836 20416 1888 20468
rect 1908 20416 1960 20468
rect 1836 20352 1888 20404
rect 1908 20352 1960 20404
rect 1836 20288 1888 20340
rect 1908 20288 1960 20340
rect 1836 20224 1888 20276
rect 1908 20224 1960 20276
rect 1836 20160 1888 20212
rect 1908 20160 1960 20212
rect 1836 20096 1888 20148
rect 1908 20096 1960 20148
rect 1836 20032 1888 20084
rect 1908 20032 1960 20084
rect 1836 19968 1888 20020
rect 1908 19968 1960 20020
rect 1836 19904 1888 19956
rect 1908 19904 1960 19956
rect 1836 19840 1888 19892
rect 1908 19840 1960 19892
rect 1836 19776 1888 19828
rect 1908 19776 1960 19828
rect 1836 19712 1888 19764
rect 1908 19712 1960 19764
rect 1836 19648 1888 19700
rect 1908 19648 1960 19700
rect 1836 19584 1888 19636
rect 1908 19584 1960 19636
rect 1836 19520 1888 19572
rect 1908 19520 1960 19572
rect 1836 19455 1888 19507
rect 1908 19455 1960 19507
rect 1836 19390 1888 19442
rect 1908 19390 1960 19442
rect 1836 19325 1888 19377
rect 1908 19325 1960 19377
rect 1836 19260 1888 19312
rect 1908 19260 1960 19312
rect 1836 19195 1888 19247
rect 1908 19195 1960 19247
rect 1836 19130 1888 19182
rect 1908 19130 1960 19182
rect 1836 19065 1888 19117
rect 1908 19065 1960 19117
rect 1836 19000 1888 19052
rect 1908 19000 1960 19052
rect 1836 18935 1888 18987
rect 1908 18935 1960 18987
rect 1836 18870 1888 18922
rect 1908 18870 1960 18922
rect 1836 18805 1888 18857
rect 1908 18805 1960 18857
rect 1836 18740 1888 18792
rect 1908 18740 1960 18792
rect 1836 18675 1888 18727
rect 1908 18675 1960 18727
rect 1836 18610 1888 18662
rect 1908 18610 1960 18662
rect 1836 18545 1888 18597
rect 1908 18545 1960 18597
rect 1836 18480 1888 18532
rect 1908 18480 1960 18532
rect 1796 18140 1848 18192
rect 1864 18140 1916 18192
rect 1932 18140 1984 18192
rect 1796 18068 1848 18120
rect 1864 18068 1916 18120
rect 1932 18068 1984 18120
rect 1796 17995 1848 18047
rect 1864 17995 1916 18047
rect 1932 17995 1984 18047
rect 1796 17922 1848 17974
rect 1864 17922 1916 17974
rect 1932 17922 1984 17974
rect 1796 17849 1848 17901
rect 1864 17849 1916 17901
rect 1932 17849 1984 17901
rect 1796 17776 1848 17828
rect 1864 17776 1916 17828
rect 1932 17776 1984 17828
rect 1796 17703 1848 17755
rect 1864 17703 1916 17755
rect 1932 17703 1984 17755
rect 1796 17466 1848 17518
rect 1864 17466 1916 17518
rect 1932 17466 1984 17518
rect 1796 17401 1848 17453
rect 1864 17401 1916 17453
rect 1932 17401 1984 17453
rect 1796 17335 1848 17387
rect 1864 17335 1916 17387
rect 1932 17335 1984 17387
rect 1796 17269 1848 17321
rect 1864 17269 1916 17321
rect 1932 17269 1984 17321
rect 1796 17203 1848 17255
rect 1864 17203 1916 17255
rect 1932 17203 1984 17255
rect 1796 17137 1848 17189
rect 1864 17137 1916 17189
rect 1932 17137 1984 17189
rect 1796 17071 1848 17123
rect 1864 17071 1916 17123
rect 1932 17071 1984 17123
rect 1796 16261 1848 16313
rect 1864 16261 1916 16313
rect 1932 16261 1984 16313
rect 1796 16197 1848 16249
rect 1864 16197 1916 16249
rect 1932 16197 1984 16249
rect 1796 16133 1848 16185
rect 1864 16133 1916 16185
rect 1932 16133 1984 16185
rect 1796 16069 1848 16121
rect 1864 16069 1916 16121
rect 1932 16069 1984 16121
rect 1796 16005 1848 16057
rect 1864 16005 1916 16057
rect 1932 16005 1984 16057
rect 1796 15941 1848 15993
rect 1864 15941 1916 15993
rect 1932 15941 1984 15993
rect 1796 15877 1848 15929
rect 1864 15877 1916 15929
rect 1932 15877 1984 15929
rect 1796 15812 1848 15864
rect 1864 15812 1916 15864
rect 1932 15812 1984 15864
rect 1796 15747 1848 15799
rect 1864 15747 1916 15799
rect 1932 15747 1984 15799
rect 1796 15682 1848 15734
rect 1864 15682 1916 15734
rect 1932 15682 1984 15734
rect 1796 15617 1848 15669
rect 1864 15617 1916 15669
rect 1932 15617 1984 15669
rect 1796 15552 1848 15604
rect 1864 15552 1916 15604
rect 1932 15552 1984 15604
rect 1796 15487 1848 15539
rect 1864 15487 1916 15539
rect 1932 15487 1984 15539
rect 1796 14588 1848 14640
rect 1864 14588 1916 14640
rect 1932 14588 1984 14640
rect 1796 14516 1848 14568
rect 1864 14516 1916 14568
rect 1932 14516 1984 14568
rect 26814 14499 26866 14551
rect 26878 14499 26930 14551
rect 1796 14444 1848 14496
rect 1864 14444 1916 14496
rect 1932 14444 1984 14496
rect 3388 14444 3440 14496
rect 3452 14444 3504 14496
rect 1796 14372 1848 14424
rect 1864 14372 1916 14424
rect 1932 14372 1984 14424
rect 3220 14370 3272 14422
rect 3284 14370 3336 14422
rect 26357 14404 26409 14456
rect 26421 14404 26473 14456
rect 1796 14299 1848 14351
rect 1864 14299 1916 14351
rect 1932 14299 1984 14351
rect 1796 14226 1848 14278
rect 1864 14226 1916 14278
rect 1932 14226 1984 14278
rect 1796 14153 1848 14205
rect 1864 14153 1916 14205
rect 1932 14153 1984 14205
rect 1796 14080 1848 14132
rect 1864 14080 1916 14132
rect 1932 14080 1984 14132
rect 27111 13571 27163 13623
rect 27178 13571 27230 13623
rect 27244 13571 27296 13623
rect 27111 13501 27163 13553
rect 27178 13501 27230 13553
rect 27244 13501 27296 13553
rect 27111 13431 27163 13483
rect 27178 13431 27230 13483
rect 27244 13431 27296 13483
rect 27568 13575 27620 13627
rect 27632 13575 27684 13627
rect 27568 13505 27620 13557
rect 27632 13505 27684 13557
rect 27568 13435 27620 13487
rect 27632 13435 27684 13487
rect 27111 12882 27163 12934
rect 27178 12882 27230 12934
rect 27244 12882 27296 12934
rect 826 12804 878 12856
rect 890 12804 942 12856
rect 954 12804 1006 12856
rect 826 12729 878 12781
rect 890 12729 942 12781
rect 954 12729 1006 12781
rect 27111 12812 27163 12864
rect 27178 12812 27230 12864
rect 27244 12812 27296 12864
rect 27111 12742 27163 12794
rect 27178 12742 27230 12794
rect 27244 12742 27296 12794
rect 27371 12882 27423 12934
rect 27438 12882 27490 12934
rect 27504 12882 27556 12934
rect 27371 12812 27423 12864
rect 27438 12812 27490 12864
rect 27504 12812 27556 12864
rect 27371 12742 27423 12794
rect 27438 12742 27490 12794
rect 27504 12742 27556 12794
rect 27974 12884 28026 12936
rect 27974 12814 28026 12866
rect 27974 12744 28026 12796
rect 826 12653 878 12705
rect 890 12653 942 12705
rect 954 12653 1006 12705
rect 826 12577 878 12629
rect 890 12577 942 12629
rect 954 12577 1006 12629
rect 25807 11368 25859 11420
rect 25871 11368 25923 11420
rect 27471 11043 27523 11095
rect 27565 11043 27617 11095
rect 13668 10935 13720 10987
rect 13732 10935 13784 10987
rect 27471 10948 27523 11000
rect 27565 10948 27617 11000
rect 102 10868 154 10920
rect 707 10868 759 10920
rect 102 10804 154 10856
rect 707 10804 759 10856
rect 226 10733 278 10785
rect 226 10669 278 10721
rect 1153 10705 1205 10757
rect 1153 10641 1205 10693
rect 10336 10595 10388 10647
rect 10336 10531 10388 10583
rect 24614 10690 24666 10742
rect 24678 10690 24730 10742
rect 24742 10690 24794 10742
rect 24614 10624 24666 10676
rect 24678 10624 24730 10676
rect 24742 10624 24794 10676
rect 24614 10558 24666 10610
rect 24678 10558 24730 10610
rect 24742 10558 24794 10610
rect 24614 10491 24666 10543
rect 24678 10491 24730 10543
rect 24742 10491 24794 10543
rect 27471 10537 27523 10589
rect 27565 10537 27617 10589
rect 24614 10424 24666 10476
rect 24678 10424 24730 10476
rect 24742 10424 24794 10476
rect 27471 10442 27523 10494
rect 27565 10442 27617 10494
rect 24614 10357 24666 10409
rect 24678 10357 24730 10409
rect 24742 10357 24794 10409
rect 14201 10236 14253 10288
rect 14265 10236 14317 10288
rect 24641 9238 24693 9290
rect 24705 9238 24757 9290
rect 22391 8076 22443 8128
rect 22463 8076 22515 8128
rect 22535 8076 22587 8128
rect 22606 8076 22658 8128
rect 22677 8076 22729 8128
rect 22748 8076 22800 8128
rect 22819 8076 22871 8128
rect 22890 8076 22942 8128
rect 22391 8002 22443 8054
rect 22463 8002 22515 8054
rect 22535 8002 22587 8054
rect 22606 8002 22658 8054
rect 22677 8002 22729 8054
rect 22748 8002 22800 8054
rect 22819 8002 22871 8054
rect 22890 8002 22942 8054
rect 22391 7928 22443 7980
rect 22463 7928 22515 7980
rect 22535 7928 22587 7980
rect 22606 7928 22658 7980
rect 22677 7928 22729 7980
rect 22748 7928 22800 7980
rect 22819 7928 22871 7980
rect 22890 7928 22942 7980
rect 3821 7087 3873 7139
rect 3885 7087 3937 7139
rect 2930 6402 2982 6454
rect 2930 6338 2982 6390
rect 2995 6338 3239 6454
rect 14032 6338 14084 6390
rect 14096 6338 14148 6390
rect 13065 6233 13117 6285
rect 13129 6233 13181 6285
rect 15641 6224 15693 6276
rect 15705 6224 15757 6276
rect 23591 6225 23643 6277
rect 23655 6225 23707 6277
rect 5946 6143 5998 6195
rect 6013 6143 6065 6195
rect 6080 6143 6132 6195
rect 6147 6143 6199 6195
rect 6214 6143 6266 6195
rect 6281 6143 6333 6195
rect 6348 6143 6400 6195
rect 6415 6143 6467 6195
rect 6482 6143 6534 6195
rect 5946 6069 5998 6121
rect 6013 6069 6065 6121
rect 6080 6069 6132 6121
rect 6147 6069 6199 6121
rect 6214 6069 6266 6121
rect 6281 6069 6333 6121
rect 6348 6069 6400 6121
rect 6415 6069 6467 6121
rect 6482 6069 6534 6121
rect 5946 5995 5998 6047
rect 6013 5995 6065 6047
rect 6080 5995 6132 6047
rect 6147 5995 6199 6047
rect 6214 5995 6266 6047
rect 6281 5995 6333 6047
rect 6348 5995 6400 6047
rect 6415 5995 6467 6047
rect 6482 5995 6534 6047
rect 12231 6143 12283 6195
rect 12298 6143 12350 6195
rect 12365 6143 12417 6195
rect 12432 6143 12484 6195
rect 12499 6143 12551 6195
rect 12566 6143 12618 6195
rect 12633 6143 12685 6195
rect 12700 6143 12752 6195
rect 12767 6143 12819 6195
rect 12231 6069 12283 6121
rect 12298 6069 12350 6121
rect 12365 6069 12417 6121
rect 12432 6069 12484 6121
rect 12499 6069 12551 6121
rect 12566 6069 12618 6121
rect 12633 6069 12685 6121
rect 12700 6069 12752 6121
rect 12767 6069 12819 6121
rect 12231 5995 12283 6047
rect 12298 5995 12350 6047
rect 12365 5995 12417 6047
rect 12432 5995 12484 6047
rect 12499 5995 12551 6047
rect 12566 5995 12618 6047
rect 12633 5995 12685 6047
rect 12700 5995 12752 6047
rect 12767 5995 12819 6047
rect 16076 6143 16128 6195
rect 16142 6143 16194 6195
rect 16208 6143 16260 6195
rect 16274 6143 16326 6195
rect 16339 6143 16391 6195
rect 16404 6143 16456 6195
rect 16469 6143 16521 6195
rect 16534 6143 16586 6195
rect 16599 6143 16651 6195
rect 16076 6069 16128 6121
rect 16142 6069 16194 6121
rect 16208 6069 16260 6121
rect 16274 6069 16326 6121
rect 16339 6069 16391 6121
rect 16404 6069 16456 6121
rect 16469 6069 16521 6121
rect 16534 6069 16586 6121
rect 16599 6069 16651 6121
rect 16076 5995 16128 6047
rect 16142 5995 16194 6047
rect 16208 5995 16260 6047
rect 16274 5995 16326 6047
rect 16339 5995 16391 6047
rect 16404 5995 16456 6047
rect 16469 5995 16521 6047
rect 16534 5995 16586 6047
rect 16599 5995 16651 6047
rect 20298 6143 20350 6195
rect 20365 6143 20417 6195
rect 20432 6143 20484 6195
rect 20499 6143 20551 6195
rect 20566 6143 20618 6195
rect 20633 6143 20685 6195
rect 20700 6143 20752 6195
rect 20767 6143 20819 6195
rect 20834 6143 20886 6195
rect 20298 6069 20350 6121
rect 20365 6069 20417 6121
rect 20432 6069 20484 6121
rect 20499 6069 20551 6121
rect 20566 6069 20618 6121
rect 20633 6069 20685 6121
rect 20700 6069 20752 6121
rect 20767 6069 20819 6121
rect 20834 6069 20886 6121
rect 20298 5995 20350 6047
rect 20365 5995 20417 6047
rect 20432 5995 20484 6047
rect 20499 5995 20551 6047
rect 20566 5995 20618 6047
rect 20633 5995 20685 6047
rect 20700 5995 20752 6047
rect 20767 5995 20819 6047
rect 20834 5995 20886 6047
rect 4040 5606 4092 5658
rect 4040 5542 4092 5594
rect 7442 5444 7494 5496
rect 7509 5444 7561 5496
rect 7576 5444 7628 5496
rect 7643 5444 7695 5496
rect 7710 5444 7762 5496
rect 7777 5444 7829 5496
rect 7844 5444 7896 5496
rect 7911 5444 7963 5496
rect 7978 5444 8030 5496
rect 7442 5372 7494 5424
rect 7509 5372 7561 5424
rect 7576 5372 7628 5424
rect 7643 5372 7695 5424
rect 7710 5372 7762 5424
rect 7777 5372 7829 5424
rect 7844 5372 7896 5424
rect 7911 5372 7963 5424
rect 7978 5372 8030 5424
rect 7442 5300 7494 5352
rect 7509 5300 7561 5352
rect 7576 5300 7628 5352
rect 7643 5300 7695 5352
rect 7710 5300 7762 5352
rect 7777 5300 7829 5352
rect 7844 5300 7896 5352
rect 7911 5300 7963 5352
rect 7978 5300 8030 5352
rect 11511 5444 11563 5496
rect 11578 5444 11630 5496
rect 11645 5444 11697 5496
rect 11712 5444 11764 5496
rect 11779 5444 11831 5496
rect 11846 5444 11898 5496
rect 11913 5444 11965 5496
rect 11980 5444 12032 5496
rect 12047 5444 12099 5496
rect 11511 5372 11563 5424
rect 11578 5372 11630 5424
rect 11645 5372 11697 5424
rect 11712 5372 11764 5424
rect 11779 5372 11831 5424
rect 11846 5372 11898 5424
rect 11913 5372 11965 5424
rect 11980 5372 12032 5424
rect 12047 5372 12099 5424
rect 11511 5300 11563 5352
rect 11578 5300 11630 5352
rect 11645 5300 11697 5352
rect 11712 5300 11764 5352
rect 11779 5300 11831 5352
rect 11846 5300 11898 5352
rect 11913 5300 11965 5352
rect 11980 5300 12032 5352
rect 12047 5300 12099 5352
rect 14533 5444 14585 5496
rect 14603 5444 14655 5496
rect 14672 5444 14724 5496
rect 14741 5444 14793 5496
rect 14810 5444 14862 5496
rect 14879 5444 14931 5496
rect 14948 5444 15000 5496
rect 14533 5372 14585 5424
rect 14603 5372 14655 5424
rect 14672 5372 14724 5424
rect 14741 5372 14793 5424
rect 14810 5372 14862 5424
rect 14879 5372 14931 5424
rect 14948 5372 15000 5424
rect 14533 5300 14585 5352
rect 14603 5300 14655 5352
rect 14672 5300 14724 5352
rect 14741 5300 14793 5352
rect 14810 5300 14862 5352
rect 14879 5300 14931 5352
rect 14948 5300 15000 5352
rect 16896 4433 16948 4485
rect 16975 4433 17027 4485
rect 17053 4433 17105 4485
rect 17131 4433 17183 4485
rect 16896 4309 16948 4361
rect 16975 4309 17027 4361
rect 17053 4309 17105 4361
rect 17131 4309 17183 4361
rect 2826 4145 2878 4197
rect 2892 4145 2944 4197
rect 2957 4145 3009 4197
rect 3022 4145 3074 4197
rect 3087 4145 3139 4197
rect 3152 4145 3204 4197
rect 2826 3831 2878 3840
rect 2826 3797 2832 3831
rect 2832 3797 2866 3831
rect 2866 3797 2878 3831
rect 2826 3788 2878 3797
rect 2892 3831 2944 3840
rect 2957 3831 3009 3840
rect 3022 3831 3074 3840
rect 3087 3831 3139 3840
rect 2892 3797 2915 3831
rect 2915 3797 2944 3831
rect 2957 3797 2998 3831
rect 2998 3797 3009 3831
rect 3022 3797 3032 3831
rect 3032 3797 3074 3831
rect 3087 3797 3115 3831
rect 3115 3797 3139 3831
rect 2892 3788 2944 3797
rect 2957 3788 3009 3797
rect 3022 3788 3074 3797
rect 3087 3788 3139 3797
rect 3152 3831 3204 3840
rect 3152 3797 3164 3831
rect 3164 3797 3198 3831
rect 3198 3797 3204 3831
rect 3152 3788 3204 3797
rect 4046 3788 4098 3840
rect 4110 3788 4162 3840
rect 26139 3788 26191 3840
rect 26203 3788 26255 3840
rect 2595 3745 2624 3756
rect 2624 3745 2647 3756
rect 2705 3745 2716 3756
rect 2716 3745 2750 3756
rect 2750 3745 2757 3756
rect 2595 3704 2647 3745
rect 2705 3704 2757 3745
rect 22552 3708 22604 3760
rect 22616 3708 22668 3760
rect 23149 3708 23201 3760
rect 23213 3708 23265 3760
rect 26605 3708 26657 3760
rect 26669 3708 26721 3760
rect 2595 3658 2624 3679
rect 2624 3658 2647 3679
rect 2705 3658 2716 3679
rect 2716 3658 2750 3679
rect 2750 3658 2757 3679
rect 2595 3627 2647 3658
rect 2705 3627 2757 3658
rect 7707 3628 7759 3680
rect 7771 3628 7823 3680
rect 20914 3628 20966 3680
rect 20978 3628 21030 3680
rect 24059 3628 24111 3680
rect 24123 3628 24175 3680
rect 26731 3628 26783 3680
rect 26795 3628 26847 3680
rect 2595 3571 2624 3602
rect 2624 3571 2647 3602
rect 2705 3571 2716 3602
rect 2716 3571 2750 3602
rect 2750 3571 2757 3602
rect 2595 3550 2647 3571
rect 2705 3550 2757 3571
rect 10415 3548 10467 3600
rect 10479 3548 10531 3600
rect 910 3358 962 3410
rect 974 3358 1026 3410
rect 3351 3445 3403 3497
rect 3415 3445 3467 3497
rect 3479 3445 3531 3497
rect 3543 3445 3595 3497
rect 11198 3468 11250 3520
rect 11262 3468 11314 3520
rect 11917 3468 11969 3520
rect 11981 3468 12033 3520
rect 14933 3480 14985 3532
rect 14997 3480 15049 3532
rect 17080 3540 17132 3550
rect 17080 3506 17090 3540
rect 17090 3506 17124 3540
rect 17124 3506 17132 3540
rect 17080 3498 17132 3506
rect 17147 3540 17199 3550
rect 17214 3540 17266 3550
rect 17281 3540 17333 3550
rect 17348 3540 17400 3550
rect 17415 3540 17467 3550
rect 17482 3540 17534 3550
rect 17549 3540 17601 3550
rect 17147 3506 17166 3540
rect 17166 3506 17199 3540
rect 17214 3506 17242 3540
rect 17242 3506 17266 3540
rect 17281 3506 17318 3540
rect 17318 3506 17333 3540
rect 17348 3506 17352 3540
rect 17352 3506 17394 3540
rect 17394 3506 17400 3540
rect 17415 3506 17428 3540
rect 17428 3506 17467 3540
rect 17482 3506 17504 3540
rect 17504 3506 17534 3540
rect 17549 3506 17579 3540
rect 17579 3506 17601 3540
rect 17147 3498 17199 3506
rect 17214 3498 17266 3506
rect 17281 3498 17333 3506
rect 17348 3498 17400 3506
rect 17415 3498 17467 3506
rect 17482 3498 17534 3506
rect 17549 3498 17601 3506
rect 17616 3540 17668 3550
rect 17616 3506 17620 3540
rect 17620 3506 17654 3540
rect 17654 3506 17668 3540
rect 17616 3498 17668 3506
rect 17682 3540 17734 3550
rect 17682 3506 17695 3540
rect 17695 3506 17729 3540
rect 17729 3506 17734 3540
rect 17682 3498 17734 3506
rect 17748 3540 17800 3550
rect 17814 3540 17866 3550
rect 17880 3540 17932 3550
rect 17946 3540 17998 3550
rect 18012 3540 18064 3550
rect 18078 3540 18130 3550
rect 17748 3506 17770 3540
rect 17770 3506 17800 3540
rect 17814 3506 17845 3540
rect 17845 3506 17866 3540
rect 17880 3506 17920 3540
rect 17920 3506 17932 3540
rect 17946 3506 17954 3540
rect 17954 3506 17995 3540
rect 17995 3506 17998 3540
rect 18012 3506 18029 3540
rect 18029 3506 18064 3540
rect 18078 3506 18104 3540
rect 18104 3506 18130 3540
rect 17748 3498 17800 3506
rect 17814 3498 17866 3506
rect 17880 3498 17932 3506
rect 17946 3498 17998 3506
rect 18012 3498 18064 3506
rect 18078 3498 18130 3506
rect 18144 3540 18196 3550
rect 18144 3506 18145 3540
rect 18145 3506 18179 3540
rect 18179 3506 18196 3540
rect 18144 3498 18196 3506
rect 18210 3540 18262 3550
rect 18210 3506 18220 3540
rect 18220 3506 18254 3540
rect 18254 3506 18262 3540
rect 18210 3498 18262 3506
rect 18276 3540 18328 3550
rect 18342 3540 18394 3550
rect 18408 3540 18460 3550
rect 18474 3540 18526 3550
rect 18540 3540 18592 3550
rect 18606 3540 18658 3550
rect 18672 3540 18724 3550
rect 18276 3506 18295 3540
rect 18295 3506 18328 3540
rect 18342 3506 18370 3540
rect 18370 3506 18394 3540
rect 18408 3506 18445 3540
rect 18445 3506 18460 3540
rect 18474 3506 18479 3540
rect 18479 3506 18520 3540
rect 18520 3506 18526 3540
rect 18540 3506 18554 3540
rect 18554 3506 18592 3540
rect 18606 3506 18629 3540
rect 18629 3506 18658 3540
rect 18672 3506 18704 3540
rect 18704 3506 18724 3540
rect 18276 3498 18328 3506
rect 18342 3498 18394 3506
rect 18408 3498 18460 3506
rect 18474 3498 18526 3506
rect 18540 3498 18592 3506
rect 18606 3498 18658 3506
rect 18672 3498 18724 3506
rect 20285 3548 20337 3600
rect 20349 3548 20401 3600
rect 22414 3548 22466 3600
rect 22478 3548 22530 3600
rect 26898 3548 26950 3600
rect 26962 3548 27014 3600
rect 27295 3548 27347 3600
rect 27359 3548 27411 3600
rect 19003 3468 19055 3520
rect 19067 3468 19119 3520
rect 22310 3468 22362 3520
rect 22374 3468 22426 3520
rect 22853 3468 22905 3520
rect 22917 3468 22969 3520
rect 26227 3468 26279 3520
rect 26291 3468 26343 3520
rect 3351 3380 3403 3432
rect 3415 3380 3467 3432
rect 3479 3380 3531 3432
rect 3543 3380 3595 3432
rect 703 3270 755 3322
rect 3351 3315 3403 3367
rect 3415 3315 3467 3367
rect 3479 3315 3531 3367
rect 3543 3315 3595 3367
rect 7676 3341 7728 3393
rect 7740 3341 7792 3393
rect 8076 3388 8128 3440
rect 8140 3388 8192 3440
rect 10711 3388 10763 3440
rect 10775 3388 10827 3440
rect 11621 3378 11673 3430
rect 11685 3378 11737 3430
rect 15843 3400 15895 3452
rect 15907 3400 15959 3452
rect 22204 3388 22256 3440
rect 22268 3388 22320 3440
rect 24355 3388 24407 3440
rect 24419 3388 24471 3440
rect 26353 3388 26405 3440
rect 26417 3388 26469 3440
rect 27730 3388 27782 3440
rect 27794 3388 27846 3440
rect 22096 3308 22148 3360
rect 22160 3308 22212 3360
rect 26520 3308 26572 3360
rect 26584 3308 26636 3360
rect 27495 3308 27547 3360
rect 27559 3308 27611 3360
rect 703 3206 755 3258
rect 3351 3250 3403 3302
rect 3415 3250 3467 3302
rect 3479 3250 3531 3302
rect 3543 3250 3595 3302
rect 3351 3185 3403 3237
rect 3415 3185 3467 3237
rect 3479 3185 3531 3237
rect 3543 3185 3595 3237
rect 1760 3088 1812 3140
rect 3351 3120 3403 3172
rect 3415 3120 3467 3172
rect 3479 3120 3531 3172
rect 3543 3120 3595 3172
rect 1165 3004 1217 3056
rect 1760 3024 1812 3076
rect 2547 3032 2599 3084
rect 1165 2940 1217 2992
rect 2547 2968 2599 3020
rect 3351 3054 3403 3106
rect 3415 3054 3467 3106
rect 3479 3054 3531 3106
rect 3543 3054 3595 3106
rect 3351 2988 3403 3040
rect 3415 2988 3467 3040
rect 3479 2988 3531 3040
rect 3543 2988 3595 3040
rect 3351 2922 3403 2974
rect 3415 2922 3467 2974
rect 3479 2922 3531 2974
rect 3543 2922 3595 2974
rect 1171 2839 1223 2891
rect 1235 2839 1287 2891
rect 2548 2834 2600 2886
rect 2548 2770 2600 2822
rect 3351 2856 3403 2908
rect 3415 2856 3467 2908
rect 3479 2856 3531 2908
rect 3543 2856 3595 2908
rect 3351 2790 3403 2842
rect 3415 2790 3467 2842
rect 3479 2790 3531 2842
rect 3543 2790 3595 2842
rect 3592 2115 3644 2121
rect 3592 2081 3601 2115
rect 3601 2081 3635 2115
rect 3635 2081 3644 2115
rect 3592 2069 3644 2081
rect 3592 2043 3644 2057
rect 3592 2009 3601 2043
rect 3601 2009 3635 2043
rect 3635 2009 3644 2043
rect 3592 2005 3644 2009
rect 23254 2007 23306 2059
rect 23324 2007 23376 2059
rect 23394 2007 23446 2059
rect 23254 1937 23306 1989
rect 23324 1937 23376 1989
rect 23394 1937 23446 1989
rect 23254 1867 23306 1919
rect 23324 1867 23376 1919
rect 23394 1867 23446 1919
rect 1934 1783 1986 1835
rect 1998 1783 2050 1835
rect 1934 1718 1986 1770
rect 1998 1718 2050 1770
rect 23254 1797 23306 1849
rect 23324 1797 23376 1849
rect 23394 1797 23446 1849
rect 23254 1726 23306 1778
rect 23324 1726 23376 1778
rect 23394 1726 23446 1778
rect 1761 1653 1813 1705
rect 1761 1589 1813 1641
rect 1934 1653 1986 1705
rect 1998 1653 2050 1705
rect 1934 1588 1986 1640
rect 1998 1588 2050 1640
rect 1934 1523 1986 1575
rect 1998 1523 2050 1575
rect 1934 1458 1986 1510
rect 1998 1458 2050 1510
rect 1934 1393 1986 1445
rect 1998 1393 2050 1445
rect 1934 1328 1986 1380
rect 1998 1328 2050 1380
rect 1934 1263 1986 1315
rect 1998 1263 2050 1315
rect 1934 1198 1986 1250
rect 1998 1198 2050 1250
rect 1934 1133 1986 1185
rect 1998 1133 2050 1185
rect 1934 1068 1986 1120
rect 1998 1068 2050 1120
rect 23788 1182 23840 1234
rect 23852 1182 23904 1234
rect 23916 1182 23968 1234
rect 23788 1088 23840 1140
rect 23852 1088 23904 1140
rect 23916 1088 23968 1140
rect 1934 1003 1986 1055
rect 1998 1003 2050 1055
rect 1934 938 1986 990
rect 1998 938 2050 990
rect 1934 873 1986 925
rect 1998 873 2050 925
rect 1934 808 1986 860
rect 1998 808 2050 860
rect 1934 743 1986 795
rect 1998 743 2050 795
rect 1934 678 1986 730
rect 1998 678 2050 730
rect 1934 612 1986 664
rect 1998 612 2050 664
rect 1934 546 1986 598
rect 1998 546 2050 598
rect 1934 480 1986 532
rect 1998 480 2050 532
rect 1934 414 1986 466
rect 1998 414 2050 466
rect 4004 159 4056 211
rect 18265 178 18317 230
rect 18336 178 18388 230
rect 18407 178 18459 230
rect 18477 178 18529 230
rect 4004 95 4056 147
<< metal2 >>
tri 17261 39682 17267 39688 ne
rect 17267 39682 17398 39688
rect 16924 39058 17088 39114
rect 16924 39057 17031 39058
tri 17031 39057 17032 39058 nw
tri 16924 39029 16952 39057 ne
rect 16952 39029 17003 39057
tri 17003 39029 17031 39057 nw
rect 11998 38680 12004 38732
rect 12056 38729 12073 38732
rect 12125 38729 12142 38732
rect 12194 38729 12211 38732
rect 12263 38729 12280 38732
rect 12332 38729 12348 38732
rect 12064 38680 12073 38729
rect 12332 38680 12339 38729
rect 12400 38680 12406 38732
rect 11998 38673 12008 38680
rect 12064 38673 12091 38680
rect 12147 38673 12174 38680
rect 12230 38673 12257 38680
rect 12313 38673 12339 38680
rect 12395 38673 12406 38680
rect 11998 38660 12406 38673
rect 11998 38608 12004 38660
rect 12056 38608 12073 38660
rect 12125 38608 12142 38660
rect 12194 38608 12211 38660
rect 12263 38608 12280 38660
rect 12332 38608 12348 38660
rect 12400 38608 12406 38660
rect 11998 38595 12406 38608
rect 11998 38588 12008 38595
rect 12064 38588 12091 38595
rect 12147 38588 12174 38595
rect 12230 38588 12257 38595
rect 12313 38588 12339 38595
rect 12395 38588 12406 38595
rect 11998 38536 12004 38588
rect 12064 38539 12073 38588
rect 12332 38539 12339 38588
rect 12056 38536 12073 38539
rect 12125 38536 12142 38539
rect 12194 38536 12211 38539
rect 12263 38536 12280 38539
rect 12332 38536 12348 38539
rect 12400 38536 12406 38588
rect 25737 37825 25743 37877
rect 25795 37825 25807 37877
rect 25859 37825 25865 37877
tri 26692 37572 26744 37624 se
rect 26744 37572 26770 37624
rect 26822 37572 26834 37624
rect 26886 37572 26892 37624
tri 26650 37530 26692 37572 se
rect 26692 37530 26744 37572
tri 26744 37530 26786 37572 nw
tri 26556 37436 26650 37530 se
tri 26650 37436 26744 37530 nw
tri 26462 37342 26556 37436 se
tri 26556 37342 26650 37436 nw
tri 26368 37248 26462 37342 se
tri 26462 37248 26556 37342 nw
tri 26286 37166 26368 37248 se
rect 25870 37157 25926 37166
tri 26274 37154 26286 37166 se
rect 26286 37154 26368 37166
tri 26368 37154 26462 37248 nw
tri 26250 37130 26274 37154 se
rect 26274 37130 26344 37154
tri 26344 37130 26368 37154 nw
rect 25926 37101 26278 37130
rect 25870 37077 26278 37101
rect 25926 37064 26278 37077
tri 26278 37064 26344 37130 nw
rect 25870 37012 25926 37021
rect 23396 34369 24185 34378
rect 23396 34313 23398 34369
rect 23454 34313 23478 34369
rect 23534 34313 23558 34369
rect 23614 34313 23638 34369
rect 23694 34313 24185 34369
rect 23396 34287 24185 34313
rect 23396 34231 23398 34287
rect 23454 34231 23478 34287
rect 23534 34231 23558 34287
rect 23614 34231 23638 34287
rect 23694 34231 24185 34287
rect 23396 34205 24185 34231
rect 23396 34149 23398 34205
rect 23454 34149 23478 34205
rect 23534 34149 23558 34205
rect 23614 34149 23638 34205
rect 23694 34149 24185 34205
rect 23396 34123 24185 34149
rect 23396 34067 23398 34123
rect 23454 34067 23478 34123
rect 23534 34067 23558 34123
rect 23614 34067 23638 34123
rect 23694 34067 24185 34123
rect 23396 34040 24185 34067
rect 23396 33984 23398 34040
rect 23454 33984 23478 34040
rect 23534 33984 23558 34040
rect 23614 33984 23638 34040
rect 23694 33984 24185 34040
rect 23396 33957 24185 33984
rect 23396 33901 23398 33957
rect 23454 33901 23478 33957
rect 23534 33901 23558 33957
rect 23614 33901 23638 33957
rect 23694 33901 24185 33957
rect 23396 33891 24185 33901
rect 3122 33126 3128 33178
rect 3180 33126 3199 33178
rect 3251 33126 3271 33178
rect 3323 33126 3845 33178
rect 3122 33121 3845 33126
tri 3845 33121 3902 33178 sw
rect 3122 33110 3902 33121
rect 3122 33058 3128 33110
rect 3180 33058 3199 33110
rect 3251 33058 3271 33110
rect 3323 33106 3902 33110
rect 3323 33058 3732 33106
tri 3613 32939 3732 33058 ne
rect 3788 33050 3846 33106
rect 3732 33010 3902 33050
rect 3788 32954 3846 33010
rect 3732 32914 3902 32954
rect 3788 32858 3846 32914
rect 3732 32818 3902 32858
rect 3788 32762 3846 32818
rect 3732 32721 3902 32762
rect 3788 32665 3846 32721
rect 3732 32656 3902 32665
rect 23396 33023 24185 33032
rect 23396 32967 23398 33023
rect 23454 32967 23478 33023
rect 23534 32967 23558 33023
rect 23614 32967 23638 33023
rect 23694 32967 24185 33023
rect 23396 32941 24185 32967
rect 23396 32885 23398 32941
rect 23454 32885 23478 32941
rect 23534 32885 23558 32941
rect 23614 32885 23638 32941
rect 23694 32885 24185 32941
rect 23396 32859 24185 32885
rect 23396 32803 23398 32859
rect 23454 32803 23478 32859
rect 23534 32803 23558 32859
rect 23614 32803 23638 32859
rect 23694 32803 24185 32859
rect 23396 32776 24185 32803
rect 23396 32720 23398 32776
rect 23454 32720 23478 32776
rect 23534 32720 23558 32776
rect 23614 32720 23638 32776
rect 23694 32720 24185 32776
rect 23396 32693 24185 32720
rect 2879 32602 2885 32654
rect 2937 32602 2972 32654
rect 3024 32602 3059 32654
rect 3111 32602 3117 32654
rect 2879 32590 3117 32602
rect 2879 32538 2885 32590
rect 2937 32538 2972 32590
rect 3024 32538 3059 32590
rect 3111 32538 3117 32590
rect 23396 32637 23398 32693
rect 23454 32637 23478 32693
rect 23534 32637 23558 32693
rect 23614 32637 23638 32693
rect 23694 32637 24185 32693
rect 23396 32610 24185 32637
rect 23396 32554 23398 32610
rect 23454 32554 23478 32610
rect 23534 32554 23558 32610
rect 23614 32554 23638 32610
rect 23694 32554 24185 32610
rect 23396 32545 24185 32554
tri 2722 32189 2879 32346 se
rect 2879 32234 3117 32538
rect 2879 32189 3044 32234
rect 602 32180 692 32189
rect 602 32124 619 32180
rect 675 32124 692 32180
tri 2694 32161 2722 32189 se
rect 2722 32161 3044 32189
tri 3044 32161 3117 32234 nw
tri 1900 32139 1922 32161 se
rect 1922 32139 2994 32161
rect 602 32111 692 32124
tri 692 32111 720 32139 sw
tri 1872 32111 1900 32139 se
rect 1900 32111 2994 32139
tri 2994 32111 3044 32161 nw
rect 602 32100 2889 32111
rect 602 32044 619 32100
rect 675 32044 2889 32100
rect 602 32020 2889 32044
rect 602 31964 619 32020
rect 675 32006 2889 32020
tri 2889 32006 2994 32111 nw
rect 675 31964 1982 32006
rect 602 31955 1982 31964
tri 1982 31955 2033 32006 nw
tri 2032 31950 2036 31954 se
rect 2036 31950 2192 31956
tri 1994 31912 2032 31950 se
rect 2032 31912 2036 31950
rect 807 31903 2036 31912
rect 807 31847 829 31903
rect 885 31898 2036 31903
rect 2088 31898 2140 31950
rect 885 31882 2192 31898
rect 885 31847 2036 31882
rect 807 31830 2036 31847
rect 2088 31830 2140 31882
rect 807 31823 2192 31830
rect 807 31767 829 31823
rect 885 31814 2192 31823
rect 885 31767 2036 31814
rect 807 31762 2036 31767
rect 2088 31762 2140 31814
rect 807 31756 2192 31762
rect 807 31743 907 31756
rect 807 31687 829 31743
rect 885 31687 907 31743
tri 907 31707 956 31756 nw
rect 807 31678 907 31687
rect 1666 31115 1888 31121
rect 1666 31056 1667 31115
rect 1719 31112 1751 31115
rect 1803 31112 1835 31115
rect 1723 31056 1747 31112
rect 1803 31056 1827 31112
rect 1887 31063 1888 31115
rect 1883 31056 1888 31063
rect 1666 31036 1888 31056
rect 1666 30969 1667 31036
rect 1719 31025 1751 31036
rect 1803 31025 1835 31036
rect 1723 30969 1747 31025
rect 1803 30969 1827 31025
rect 1887 30984 1888 31036
rect 1883 30969 1888 30984
rect 1666 30957 1888 30969
rect 1666 30882 1667 30957
rect 1719 30938 1751 30957
rect 1803 30938 1835 30957
rect 1723 30882 1747 30938
rect 1803 30882 1827 30938
rect 1887 30905 1888 30957
rect 1883 30882 1888 30905
rect 1666 30878 1888 30882
rect 1666 30794 1667 30878
rect 1719 30850 1751 30878
rect 1803 30850 1835 30878
rect 1723 30794 1747 30850
rect 1803 30794 1827 30850
rect 1887 30826 1888 30878
rect 1883 30820 1888 30826
tri 23237 30845 23270 30878 sw
rect 1883 30794 1884 30820
rect 1666 30785 1884 30794
rect 23237 30793 23270 30845
rect 23237 30785 23262 30793
tri 23262 30785 23270 30793 nw
tri 23237 30760 23262 30785 nw
rect 18743 23746 19021 23755
rect 18743 23690 18744 23746
rect 18800 23690 18854 23746
rect 18910 23690 18964 23746
rect 19020 23690 19021 23746
rect 18743 23659 19021 23690
rect 18743 23603 18744 23659
rect 18800 23603 18854 23659
rect 18910 23603 18964 23659
rect 19020 23603 19021 23659
rect 18743 23572 19021 23603
rect 18743 23516 18744 23572
rect 18800 23516 18854 23572
rect 18910 23516 18964 23572
rect 19020 23516 19021 23572
rect 18743 23485 19021 23516
rect 18743 23429 18744 23485
rect 18800 23429 18854 23485
rect 18910 23429 18964 23485
rect 19020 23429 19021 23485
rect 18743 23398 19021 23429
rect 18743 23342 18744 23398
rect 18800 23342 18854 23398
rect 18910 23342 18964 23398
rect 19020 23342 19021 23398
rect 18743 23311 19021 23342
rect 18743 23255 18744 23311
rect 18800 23255 18854 23311
rect 18910 23255 18964 23311
rect 19020 23255 19021 23311
rect 18743 23223 19021 23255
rect 18743 23167 18744 23223
rect 18800 23167 18854 23223
rect 18910 23167 18964 23223
rect 19020 23167 19021 23223
rect 18743 23135 19021 23167
rect 18743 23079 18744 23135
rect 18800 23079 18854 23135
rect 18910 23079 18964 23135
rect 19020 23079 19021 23135
rect 18743 23047 19021 23079
rect 18743 22991 18744 23047
rect 18800 22991 18854 23047
rect 18910 22991 18964 23047
rect 19020 22991 19021 23047
rect 18743 22959 19021 22991
rect 18743 22903 18744 22959
rect 18800 22903 18854 22959
rect 18910 22903 18964 22959
rect 19020 22903 19021 22959
rect 18743 22871 19021 22903
rect 27044 23276 27673 23279
rect 27044 23224 27050 23276
rect 27102 23272 27121 23276
rect 27173 23272 27192 23276
rect 27244 23272 27262 23276
rect 27314 23272 27332 23276
rect 27384 23272 27402 23276
rect 27112 23224 27121 23272
rect 27384 23224 27392 23272
rect 27454 23224 27472 23276
rect 27524 23272 27542 23276
rect 27532 23224 27542 23272
rect 27594 23224 27612 23276
rect 27664 23224 27673 23276
rect 27044 23216 27056 23224
rect 27112 23216 27140 23224
rect 27196 23216 27224 23224
rect 27280 23216 27308 23224
rect 27364 23216 27392 23224
rect 27448 23216 27476 23224
rect 27532 23216 27673 23224
rect 27044 23210 27673 23216
rect 27044 23158 27050 23210
rect 27102 23192 27121 23210
rect 27173 23192 27192 23210
rect 27244 23192 27262 23210
rect 27314 23192 27332 23210
rect 27384 23192 27402 23210
rect 27112 23158 27121 23192
rect 27384 23158 27392 23192
rect 27454 23158 27472 23210
rect 27524 23192 27542 23210
rect 27532 23158 27542 23192
rect 27594 23158 27612 23210
rect 27664 23158 27673 23210
rect 27044 23144 27056 23158
rect 27112 23144 27140 23158
rect 27196 23144 27224 23158
rect 27280 23144 27308 23158
rect 27364 23144 27392 23158
rect 27448 23144 27476 23158
rect 27532 23144 27673 23158
rect 27044 23092 27050 23144
rect 27112 23136 27121 23144
rect 27384 23136 27392 23144
rect 27102 23112 27121 23136
rect 27173 23112 27192 23136
rect 27244 23112 27262 23136
rect 27314 23112 27332 23136
rect 27384 23112 27402 23136
rect 27112 23092 27121 23112
rect 27384 23092 27392 23112
rect 27454 23092 27472 23144
rect 27532 23136 27542 23144
rect 27524 23112 27542 23136
rect 27532 23092 27542 23112
rect 27594 23092 27612 23144
rect 27664 23092 27673 23144
rect 27044 23078 27056 23092
rect 27112 23078 27140 23092
rect 27196 23078 27224 23092
rect 27280 23078 27308 23092
rect 27364 23078 27392 23092
rect 27448 23078 27476 23092
rect 27532 23078 27673 23092
rect 27044 23026 27050 23078
rect 27112 23056 27121 23078
rect 27384 23056 27392 23078
rect 27102 23032 27121 23056
rect 27173 23032 27192 23056
rect 27244 23032 27262 23056
rect 27314 23032 27332 23056
rect 27384 23032 27402 23056
rect 27112 23026 27121 23032
rect 27384 23026 27392 23032
rect 27454 23026 27472 23078
rect 27532 23056 27542 23078
rect 27524 23032 27542 23056
rect 27532 23026 27542 23032
rect 27594 23026 27612 23078
rect 27664 23026 27673 23078
rect 27044 23012 27056 23026
rect 27112 23012 27140 23026
rect 27196 23012 27224 23026
rect 27280 23012 27308 23026
rect 27364 23012 27392 23026
rect 27448 23012 27476 23026
rect 27532 23012 27673 23026
rect 27044 22960 27050 23012
rect 27112 22976 27121 23012
rect 27384 22976 27392 23012
rect 27102 22960 27121 22976
rect 27173 22960 27192 22976
rect 27244 22960 27262 22976
rect 27314 22960 27332 22976
rect 27384 22960 27402 22976
rect 27454 22960 27472 23012
rect 27532 22976 27542 23012
rect 27524 22960 27542 22976
rect 27594 22960 27612 23012
rect 27664 22960 27673 23012
rect 27044 22952 27673 22960
rect 27044 22946 27056 22952
rect 27112 22946 27140 22952
rect 27196 22946 27224 22952
rect 27280 22946 27308 22952
rect 27364 22946 27392 22952
rect 27448 22946 27476 22952
rect 27532 22946 27673 22952
rect 27044 22894 27050 22946
rect 27112 22896 27121 22946
rect 27384 22896 27392 22946
rect 27102 22894 27121 22896
rect 27173 22894 27192 22896
rect 27244 22894 27262 22896
rect 27314 22894 27332 22896
rect 27384 22894 27402 22896
rect 27454 22894 27472 22946
rect 27532 22896 27542 22946
rect 27524 22894 27542 22896
rect 27594 22894 27612 22946
rect 27664 22894 27673 22946
rect 27044 22891 27673 22894
rect 18743 22815 18744 22871
rect 18800 22815 18854 22871
rect 18910 22815 18964 22871
rect 19020 22815 19021 22871
rect 18743 22806 19021 22815
rect 27341 22861 27673 22891
rect 27341 22858 27355 22861
rect 27341 22802 27345 22858
rect 27407 22809 27419 22861
rect 27471 22809 27483 22861
rect 27535 22858 27547 22861
rect 27539 22809 27547 22858
rect 27599 22809 27611 22861
rect 27663 22809 27673 22861
rect 27401 22802 27483 22809
rect 27539 22802 27673 22809
rect 27341 22794 27673 22802
rect 27341 22776 27355 22794
rect 27341 22720 27345 22776
rect 27407 22742 27419 22794
rect 27471 22742 27483 22794
rect 27535 22776 27547 22794
rect 27539 22742 27547 22776
rect 27599 22742 27611 22794
rect 27663 22742 27673 22794
rect 27401 22727 27483 22742
rect 27539 22727 27673 22742
rect 27341 22694 27355 22720
rect 27341 22638 27345 22694
rect 27407 22675 27419 22727
rect 27471 22675 27483 22727
rect 27539 22720 27547 22727
rect 27535 22694 27547 22720
rect 27539 22675 27547 22694
rect 27599 22675 27611 22727
rect 27663 22675 27673 22727
rect 27401 22660 27483 22675
rect 27539 22660 27673 22675
rect 27341 22612 27355 22638
rect 27341 22556 27345 22612
rect 27407 22608 27419 22660
rect 27471 22608 27483 22660
rect 27539 22638 27547 22660
rect 27535 22612 27547 22638
rect 27539 22608 27547 22612
rect 27599 22608 27611 22660
rect 27663 22608 27673 22660
rect 27401 22593 27483 22608
rect 27539 22593 27673 22608
rect 27341 22541 27355 22556
rect 27407 22541 27419 22593
rect 27471 22541 27483 22593
rect 27539 22556 27547 22593
rect 27535 22541 27547 22556
rect 27599 22541 27611 22593
rect 27663 22541 27673 22593
rect 27341 22530 27673 22541
rect 27341 22474 27345 22530
rect 27401 22526 27483 22530
rect 27539 22526 27673 22530
rect 27407 22474 27419 22526
rect 27471 22474 27483 22526
rect 27539 22474 27547 22526
rect 27599 22474 27611 22526
rect 27663 22474 27673 22526
rect 27341 22459 27673 22474
rect 27341 22448 27355 22459
rect 27341 22392 27345 22448
rect 27407 22407 27419 22459
rect 27471 22407 27483 22459
rect 27535 22448 27547 22459
rect 27539 22407 27547 22448
rect 27599 22407 27611 22459
rect 27663 22407 27673 22459
rect 27401 22392 27483 22407
rect 27539 22392 27673 22407
rect 27341 22366 27355 22392
rect 27341 22310 27345 22366
rect 27407 22340 27419 22392
rect 27471 22340 27483 22392
rect 27535 22366 27547 22392
rect 27539 22340 27547 22366
rect 27599 22340 27611 22392
rect 27663 22340 27673 22392
rect 27401 22324 27483 22340
rect 27539 22324 27673 22340
rect 27341 22284 27355 22310
rect 27341 22228 27345 22284
rect 27407 22272 27419 22324
rect 27471 22272 27483 22324
rect 27539 22310 27547 22324
rect 27535 22284 27547 22310
rect 27539 22272 27547 22284
rect 27599 22272 27611 22324
rect 27663 22272 27673 22324
rect 27401 22256 27483 22272
rect 27539 22256 27673 22272
rect 27341 22204 27355 22228
rect 27407 22204 27419 22256
rect 27471 22204 27483 22256
rect 27539 22228 27547 22256
rect 27535 22204 27547 22228
rect 27599 22204 27611 22256
rect 27663 22204 27673 22256
rect 27341 22202 27673 22204
rect 27341 22146 27345 22202
rect 27401 22188 27483 22202
rect 27539 22188 27673 22202
rect 27341 22136 27355 22146
rect 27407 22136 27419 22188
rect 27471 22136 27483 22188
rect 27539 22146 27547 22188
rect 27535 22136 27547 22146
rect 27599 22136 27611 22188
rect 27663 22136 27673 22188
rect 27341 22120 27673 22136
rect 27341 22064 27345 22120
rect 27401 22064 27483 22120
rect 27539 22064 27673 22120
rect 27341 22038 27673 22064
rect 27341 21982 27345 22038
rect 27401 21982 27483 22038
rect 27539 21982 27673 22038
rect 27341 21956 27673 21982
rect 27341 21900 27345 21956
rect 27401 21900 27483 21956
rect 27539 21900 27673 21956
rect 27341 21874 27673 21900
rect 27341 21818 27345 21874
rect 27401 21818 27483 21874
rect 27539 21818 27673 21874
rect 27341 21792 27673 21818
rect 27341 21736 27345 21792
rect 27401 21736 27483 21792
rect 27539 21736 27673 21792
rect 27341 21710 27673 21736
rect 27341 21654 27345 21710
rect 27401 21654 27483 21710
rect 27539 21654 27673 21710
rect 27341 21628 27673 21654
rect 27341 21572 27345 21628
rect 27401 21572 27483 21628
rect 27539 21572 27673 21628
rect 27341 21546 27673 21572
rect 27341 21490 27345 21546
rect 27401 21490 27483 21546
rect 27539 21490 27673 21546
rect 27341 21464 27673 21490
rect 27341 21408 27345 21464
rect 27401 21408 27483 21464
rect 27539 21408 27673 21464
rect 27341 21382 27673 21408
rect 1834 21364 1962 21371
rect 1834 21312 1836 21364
rect 1888 21362 1908 21364
rect 1960 21312 1962 21364
rect 1834 21306 1870 21312
rect 1926 21306 1962 21312
rect 1834 21300 1962 21306
rect 1834 21248 1836 21300
rect 1888 21282 1908 21300
rect 1960 21248 1962 21300
rect 1834 21236 1870 21248
rect 1926 21236 1962 21248
rect 1834 21184 1836 21236
rect 1888 21202 1908 21226
rect 1960 21184 1962 21236
rect 1834 21172 1870 21184
rect 1926 21172 1962 21184
rect 1834 21120 1836 21172
rect 1888 21122 1908 21146
rect 1960 21120 1962 21172
rect 27341 21326 27345 21382
rect 27401 21375 27483 21382
rect 27341 21323 27364 21326
rect 27416 21323 27428 21375
rect 27480 21326 27483 21375
rect 27539 21367 27673 21382
rect 27480 21323 27515 21326
rect 27341 21315 27515 21323
rect 27567 21315 27621 21367
rect 27341 21299 27673 21315
rect 27341 21243 27345 21299
rect 27401 21269 27483 21299
rect 27539 21288 27673 21299
rect 27341 21217 27364 21243
rect 27416 21217 27428 21269
rect 27480 21243 27483 21269
rect 27480 21236 27515 21243
rect 27567 21236 27621 21288
rect 27480 21217 27673 21236
rect 27341 21216 27673 21217
rect 27341 21160 27345 21216
rect 27401 21160 27483 21216
rect 27539 21209 27673 21216
rect 27341 21157 27515 21160
rect 27567 21157 27621 21209
rect 27341 21151 27673 21157
rect 1834 21108 1870 21120
rect 1926 21108 1962 21120
rect 1834 21056 1836 21108
rect 1888 21056 1908 21066
rect 1960 21056 1962 21108
rect 1834 21044 1962 21056
rect 1834 20992 1836 21044
rect 1888 21042 1908 21044
rect 1960 20992 1962 21044
rect 1834 20986 1870 20992
rect 1926 20986 1962 20992
rect 1834 20980 1962 20986
rect 1834 20928 1836 20980
rect 1888 20962 1908 20980
rect 1960 20928 1962 20980
rect 1834 20916 1870 20928
rect 1926 20916 1962 20928
rect 1834 20864 1836 20916
rect 1888 20882 1908 20906
rect 1960 20864 1962 20916
rect 1834 20852 1870 20864
rect 1926 20852 1962 20864
rect 1834 20800 1836 20852
rect 1888 20802 1908 20826
rect 1960 20800 1962 20852
rect 1834 20788 1870 20800
rect 1926 20788 1962 20800
rect 1834 20736 1836 20788
rect 1888 20736 1908 20746
rect 1960 20736 1962 20788
rect 1834 20724 1962 20736
rect 1834 20672 1836 20724
rect 1888 20722 1908 20724
rect 1960 20672 1962 20724
rect 1834 20666 1870 20672
rect 1926 20666 1962 20672
rect 1834 20660 1962 20666
rect 1834 20608 1836 20660
rect 1888 20642 1908 20660
rect 1960 20608 1962 20660
rect 2387 20793 2515 20802
rect 2387 20737 2423 20793
rect 2479 20737 2515 20793
rect 2387 20708 2515 20737
rect 2387 20652 2423 20708
rect 2479 20652 2515 20708
rect 2387 20643 2515 20652
rect 1834 20596 1870 20608
rect 1926 20596 1962 20608
rect 1834 20544 1836 20596
rect 1888 20562 1908 20586
rect 1960 20544 1962 20596
rect 1834 20532 1870 20544
rect 1926 20532 1962 20544
rect 1834 20480 1836 20532
rect 1888 20482 1908 20506
rect 1960 20480 1962 20532
rect 1834 20468 1870 20480
rect 1926 20468 1962 20480
rect 1834 20416 1836 20468
rect 1888 20416 1908 20426
rect 1960 20416 1962 20468
rect 1834 20404 1962 20416
rect 1834 20352 1836 20404
rect 1888 20401 1908 20404
rect 1960 20352 1962 20404
rect 1834 20345 1870 20352
rect 1926 20345 1962 20352
rect 1834 20340 1962 20345
rect 1834 20288 1836 20340
rect 1888 20320 1908 20340
rect 1960 20288 1962 20340
rect 1834 20276 1870 20288
rect 1926 20276 1962 20288
rect 1834 20224 1836 20276
rect 1888 20239 1908 20264
rect 1960 20224 1962 20276
rect 1834 20212 1870 20224
rect 1926 20212 1962 20224
rect 1834 20160 1836 20212
rect 1888 20160 1908 20183
rect 1960 20160 1962 20212
rect 1834 20158 1962 20160
rect 1834 20148 1870 20158
rect 1926 20148 1962 20158
rect 1834 20096 1836 20148
rect 1888 20096 1908 20102
rect 1960 20096 1962 20148
rect 1834 20084 1962 20096
rect 1834 20032 1836 20084
rect 1888 20077 1908 20084
rect 1960 20032 1962 20084
rect 1834 20021 1870 20032
rect 1926 20021 1962 20032
rect 1834 20020 1962 20021
rect 1834 19968 1836 20020
rect 1888 19996 1908 20020
rect 1960 19968 1962 20020
rect 1834 19956 1870 19968
rect 1926 19956 1962 19968
rect 1834 19904 1836 19956
rect 1888 19915 1908 19940
rect 1960 19904 1962 19956
rect 1834 19892 1870 19904
rect 1926 19892 1962 19904
rect 1834 19840 1836 19892
rect 1888 19840 1908 19859
rect 1960 19840 1962 19892
rect 1834 19834 1962 19840
rect 1834 19828 1870 19834
rect 1926 19828 1962 19834
rect 1834 19776 1836 19828
rect 1888 19776 1908 19778
rect 1960 19776 1962 19828
rect 1834 19764 1962 19776
rect 1834 19712 1836 19764
rect 1888 19753 1908 19764
rect 1960 19712 1962 19764
rect 1834 19700 1870 19712
rect 1926 19700 1962 19712
rect 1834 19648 1836 19700
rect 1888 19672 1908 19697
rect 1960 19648 1962 19700
rect 1834 19636 1870 19648
rect 1926 19636 1962 19648
rect 1834 19584 1836 19636
rect 1888 19591 1908 19616
rect 1960 19584 1962 19636
rect 1834 19572 1870 19584
rect 1926 19572 1962 19584
rect 1834 19520 1836 19572
rect 1888 19520 1908 19535
rect 1960 19520 1962 19572
rect 1834 19510 1962 19520
rect 1834 19507 1870 19510
rect 1926 19507 1962 19510
rect 1834 19455 1836 19507
rect 1960 19455 1962 19507
rect 1834 19454 1870 19455
rect 1926 19454 1962 19455
rect 1834 19442 1962 19454
rect 1834 19390 1836 19442
rect 1888 19429 1908 19442
rect 1960 19390 1962 19442
rect 1834 19377 1870 19390
rect 1926 19377 1962 19390
rect 1834 19325 1836 19377
rect 1888 19348 1908 19373
rect 1960 19325 1962 19377
rect 1834 19312 1870 19325
rect 1926 19312 1962 19325
rect 1834 19260 1836 19312
rect 1888 19267 1908 19292
rect 1960 19260 1962 19312
rect 1834 19247 1870 19260
rect 1926 19247 1962 19260
rect 1834 19195 1836 19247
rect 1888 19195 1908 19211
rect 1960 19195 1962 19247
rect 1834 19186 1962 19195
rect 1834 19182 1870 19186
rect 1926 19182 1962 19186
rect 1834 19130 1836 19182
rect 1960 19130 1962 19182
rect 1834 19117 1962 19130
rect 1834 19065 1836 19117
rect 1888 19105 1908 19117
rect 1960 19065 1962 19117
rect 1834 19052 1870 19065
rect 1926 19052 1962 19065
rect 1834 19000 1836 19052
rect 1888 19024 1908 19049
rect 1960 19000 1962 19052
rect 1834 18987 1870 19000
rect 1926 18987 1962 19000
rect 1834 18935 1836 18987
rect 1888 18943 1908 18968
rect 1960 18935 1962 18987
rect 1834 18922 1870 18935
rect 1926 18922 1962 18935
rect 1834 18870 1836 18922
rect 1888 18870 1908 18887
rect 1960 18870 1962 18922
rect 1834 18862 1962 18870
rect 1834 18857 1870 18862
rect 1926 18857 1962 18862
rect 1834 18805 1836 18857
rect 1888 18805 1908 18806
rect 1960 18805 1962 18857
rect 1834 18792 1962 18805
rect 1834 18740 1836 18792
rect 1888 18781 1908 18792
rect 1960 18740 1962 18792
rect 1834 18727 1870 18740
rect 1926 18727 1962 18740
rect 1834 18675 1836 18727
rect 1888 18700 1908 18725
rect 1960 18675 1962 18727
rect 1834 18662 1870 18675
rect 1926 18662 1962 18675
rect 1834 18610 1836 18662
rect 1888 18619 1908 18644
rect 1960 18610 1962 18662
rect 1834 18597 1870 18610
rect 1926 18597 1962 18610
rect 1834 18545 1836 18597
rect 1888 18545 1908 18563
rect 1960 18545 1962 18597
rect 1834 18538 1962 18545
rect 1834 18532 1870 18538
rect 1926 18532 1962 18538
rect 1834 18480 1836 18532
rect 1888 18480 1908 18482
rect 1960 18480 1962 18532
rect 1834 18473 1962 18480
rect 1771 18201 1987 18210
rect 1827 18192 1851 18201
rect 1907 18192 1931 18201
rect 1848 18145 1851 18192
rect 1916 18145 1931 18192
rect 1771 18140 1796 18145
rect 1848 18140 1864 18145
rect 1916 18140 1932 18145
rect 1984 18140 1987 18145
rect 1771 18120 1987 18140
rect 1771 18112 1796 18120
rect 1848 18112 1864 18120
rect 1916 18112 1932 18120
rect 1984 18112 1987 18120
rect 1848 18068 1851 18112
rect 1916 18068 1931 18112
rect 1827 18056 1851 18068
rect 1907 18056 1931 18068
rect 1771 18047 1987 18056
rect 1771 18023 1796 18047
rect 1848 18023 1864 18047
rect 1916 18023 1932 18047
rect 1984 18023 1987 18047
rect 1848 17995 1851 18023
rect 1916 17995 1931 18023
rect 1827 17974 1851 17995
rect 1907 17974 1931 17995
rect 1848 17967 1851 17974
rect 1916 17967 1931 17974
rect 1771 17934 1796 17967
rect 1848 17934 1864 17967
rect 1916 17934 1932 17967
rect 1984 17934 1987 17967
rect 1848 17922 1851 17934
rect 1916 17922 1931 17934
rect 1827 17901 1851 17922
rect 1907 17901 1931 17922
rect 1848 17878 1851 17901
rect 1916 17878 1931 17901
rect 1771 17849 1796 17878
rect 1848 17849 1864 17878
rect 1916 17849 1932 17878
rect 1984 17849 1987 17878
rect 1771 17845 1987 17849
rect 1827 17828 1851 17845
rect 1907 17828 1931 17845
rect 1848 17789 1851 17828
rect 1916 17789 1931 17828
rect 1771 17776 1796 17789
rect 1848 17776 1864 17789
rect 1916 17776 1932 17789
rect 1984 17776 1987 17789
rect 1771 17755 1987 17776
rect 1848 17703 1851 17755
rect 1916 17703 1931 17755
rect 1827 17699 1851 17703
rect 1907 17699 1931 17703
rect 1771 17690 1987 17699
rect 1771 17527 1987 17536
rect 1771 17387 1987 17391
rect 1771 17366 1796 17387
rect 1848 17366 1864 17387
rect 1916 17366 1932 17387
rect 1984 17366 1987 17387
rect 1848 17335 1851 17366
rect 1916 17335 1931 17366
rect 1827 17321 1851 17335
rect 1907 17321 1931 17335
rect 1848 17310 1851 17321
rect 1916 17310 1931 17321
rect 1771 17285 1796 17310
rect 1848 17285 1864 17310
rect 1916 17285 1932 17310
rect 1984 17285 1987 17310
rect 1848 17269 1851 17285
rect 1916 17269 1931 17285
rect 1827 17255 1851 17269
rect 1907 17255 1931 17269
rect 1848 17229 1851 17255
rect 1916 17229 1931 17255
rect 1771 17204 1796 17229
rect 1848 17204 1864 17229
rect 1916 17204 1932 17229
rect 1984 17204 1987 17229
rect 1848 17203 1851 17204
rect 1916 17203 1931 17204
rect 1827 17189 1851 17203
rect 1907 17189 1931 17203
rect 1848 17148 1851 17189
rect 1916 17148 1931 17189
rect 1771 17137 1796 17148
rect 1848 17137 1864 17148
rect 1916 17137 1932 17148
rect 1984 17137 1987 17148
rect 1771 17123 1987 17137
rect 1848 17071 1851 17123
rect 1916 17071 1931 17123
rect 1827 17067 1851 17071
rect 1907 17067 1931 17071
rect 1771 17058 1987 17067
rect 1771 16322 1987 16331
rect 1827 16313 1851 16322
rect 1907 16313 1931 16322
rect 1848 16266 1851 16313
rect 1916 16266 1931 16313
rect 1771 16261 1796 16266
rect 1848 16261 1864 16266
rect 1916 16261 1932 16266
rect 1984 16261 1987 16266
rect 1771 16249 1987 16261
rect 1771 16235 1796 16249
rect 1848 16235 1864 16249
rect 1916 16235 1932 16249
rect 1984 16235 1987 16249
rect 1848 16197 1851 16235
rect 1916 16197 1931 16235
rect 1827 16185 1851 16197
rect 1907 16185 1931 16197
rect 1848 16179 1851 16185
rect 1916 16179 1931 16185
rect 1771 16148 1796 16179
rect 1848 16148 1864 16179
rect 1916 16148 1932 16179
rect 1984 16148 1987 16179
rect 1848 16133 1851 16148
rect 1916 16133 1931 16148
rect 1827 16121 1851 16133
rect 1907 16121 1931 16133
rect 1848 16092 1851 16121
rect 1916 16092 1931 16121
rect 1771 16069 1796 16092
rect 1848 16069 1864 16092
rect 1916 16069 1932 16092
rect 1984 16069 1987 16092
rect 1771 16061 1987 16069
rect 1827 16057 1851 16061
rect 1907 16057 1931 16061
rect 1848 16005 1851 16057
rect 1916 16005 1931 16057
rect 1771 15993 1987 16005
rect 1771 15974 1796 15993
rect 1848 15974 1864 15993
rect 1916 15974 1932 15993
rect 1984 15974 1987 15993
rect 1848 15941 1851 15974
rect 1916 15941 1931 15974
rect 1827 15929 1851 15941
rect 1907 15929 1931 15941
rect 1848 15918 1851 15929
rect 1916 15918 1931 15929
rect 1771 15887 1796 15918
rect 1848 15887 1864 15918
rect 1916 15887 1932 15918
rect 1984 15887 1987 15918
rect 1848 15877 1851 15887
rect 1916 15877 1931 15887
rect 1827 15864 1851 15877
rect 1907 15864 1931 15877
rect 1848 15831 1851 15864
rect 1916 15831 1931 15864
rect 1771 15812 1796 15831
rect 1848 15812 1864 15831
rect 1916 15812 1932 15831
rect 1984 15812 1987 15831
rect 1771 15800 1987 15812
rect 1827 15799 1851 15800
rect 1907 15799 1931 15800
rect 1848 15747 1851 15799
rect 1916 15747 1931 15799
rect 1827 15744 1851 15747
rect 1907 15744 1931 15747
rect 1771 15734 1987 15744
rect 1771 15713 1796 15734
rect 1848 15713 1864 15734
rect 1916 15713 1932 15734
rect 1984 15713 1987 15734
rect 1848 15682 1851 15713
rect 1916 15682 1931 15713
rect 1827 15669 1851 15682
rect 1907 15669 1931 15682
rect 1848 15657 1851 15669
rect 1916 15657 1931 15669
rect 1771 15626 1796 15657
rect 1848 15626 1864 15657
rect 1916 15626 1932 15657
rect 1984 15626 1987 15657
rect 1848 15617 1851 15626
rect 1916 15617 1931 15626
rect 1827 15604 1851 15617
rect 1907 15604 1931 15617
rect 1848 15570 1851 15604
rect 1916 15570 1931 15604
rect 1771 15552 1796 15570
rect 1848 15552 1864 15570
rect 1916 15552 1932 15570
rect 1984 15552 1987 15570
rect 1771 15539 1987 15552
rect 1848 15487 1851 15539
rect 1916 15487 1931 15539
rect 1827 15483 1851 15487
rect 1907 15483 1931 15487
rect 1771 15474 1987 15483
rect 1771 14649 1987 14658
rect 1827 14640 1851 14649
rect 1907 14640 1931 14649
rect 1848 14593 1851 14640
rect 1916 14593 1931 14640
rect 1771 14588 1796 14593
rect 1848 14588 1864 14593
rect 1916 14588 1932 14593
rect 1984 14588 1987 14593
rect 1771 14568 1987 14588
rect 1771 14563 1796 14568
rect 1848 14563 1864 14568
rect 1916 14563 1932 14568
rect 1984 14563 1987 14568
rect 1848 14516 1851 14563
rect 1916 14516 1931 14563
rect 1827 14507 1851 14516
rect 1907 14507 1931 14516
rect 1771 14496 1987 14507
tri 26511 14505 26557 14551 se
rect 26557 14505 26814 14551
rect 26511 14499 26814 14505
rect 26866 14499 26878 14551
rect 26930 14499 26936 14551
rect 26511 14496 26635 14499
tri 26635 14496 26638 14499 nw
rect 1771 14477 1796 14496
rect 1848 14477 1864 14496
rect 1916 14477 1932 14496
rect 1984 14477 1987 14496
rect 1848 14444 1851 14477
rect 1916 14444 1931 14477
rect 1189 14434 1245 14443
rect 1189 14354 1245 14378
tri 1182 14205 1189 14212 se
rect 1189 14205 1245 14298
tri 1163 14186 1182 14205 se
rect 1182 14186 1245 14205
rect 98 14126 1245 14186
rect 1827 14424 1851 14444
rect 1907 14424 1931 14444
rect 1848 14421 1851 14424
rect 1916 14421 1931 14424
rect 3290 14422 3342 14456
rect 3382 14444 3388 14496
rect 3440 14444 3452 14496
rect 3504 14444 3510 14496
rect 26511 14456 26595 14496
tri 26595 14456 26635 14496 nw
rect 1771 14391 1796 14421
rect 1848 14391 1864 14421
rect 1916 14391 1932 14421
rect 1984 14391 1987 14421
rect 1848 14372 1851 14391
rect 1916 14372 1931 14391
rect 1827 14351 1851 14372
rect 1907 14351 1931 14372
rect 3214 14370 3220 14422
rect 3272 14370 3284 14422
rect 3336 14370 3342 14422
rect 26351 14404 26357 14456
rect 26409 14404 26421 14456
rect 26473 14404 26479 14456
rect 1848 14335 1851 14351
rect 1916 14335 1931 14351
rect 1771 14305 1796 14335
rect 1848 14305 1864 14335
rect 1916 14305 1932 14335
rect 1984 14305 1987 14335
rect 1848 14299 1851 14305
rect 1916 14299 1931 14305
rect 1827 14278 1851 14299
rect 1907 14278 1931 14299
rect 1848 14249 1851 14278
rect 1916 14249 1931 14278
rect 1771 14226 1796 14249
rect 1848 14226 1864 14249
rect 1916 14226 1932 14249
rect 1984 14226 1987 14249
rect 1771 14219 1987 14226
rect 1827 14205 1851 14219
rect 1907 14205 1931 14219
rect 1309 14173 1365 14182
tri 1307 14126 1309 14128 se
rect 98 14089 169 14126
tri 169 14089 206 14126 nw
tri 1270 14089 1307 14126 se
rect 1307 14117 1309 14126
rect 1307 14093 1365 14117
rect 1307 14089 1309 14093
rect 98 14080 160 14089
tri 160 14080 169 14089 nw
rect 98 10920 159 14080
tri 159 14079 160 14080 nw
rect 98 10868 102 10920
rect 154 10868 159 10920
rect 98 10856 159 10868
rect 98 10804 102 10856
rect 154 10804 159 10856
rect 98 10797 159 10804
rect 221 14037 1309 14089
rect 1848 14163 1851 14205
rect 1916 14163 1931 14205
rect 1771 14153 1796 14163
rect 1848 14153 1864 14163
rect 1916 14153 1932 14163
rect 1984 14153 1987 14163
rect 1771 14132 1987 14153
rect 1848 14080 1851 14132
rect 1916 14080 1931 14132
rect 1827 14076 1851 14080
rect 1907 14076 1931 14080
rect 2794 14224 2850 14233
rect 2794 14144 2850 14168
rect 2794 14079 2850 14088
rect 22097 14128 23448 14130
rect 1771 14067 1987 14076
rect 22097 14072 22106 14128
rect 22162 14072 22187 14128
rect 22243 14072 22268 14128
rect 22324 14072 22349 14128
rect 22405 14072 22430 14128
rect 22486 14072 22511 14128
rect 22567 14072 22592 14128
rect 22648 14072 22673 14128
rect 22729 14072 22753 14128
rect 22809 14072 22833 14128
rect 22889 14072 22913 14128
rect 22969 14121 23448 14128
rect 22969 14072 23254 14121
rect 221 14027 1365 14037
rect 22097 14065 23254 14072
rect 23310 14065 23392 14121
rect 221 10785 282 14027
tri 282 13986 323 14027 nw
rect 22097 14026 23448 14065
rect 22097 13970 22106 14026
rect 22162 13970 22187 14026
rect 22243 13970 22268 14026
rect 22324 13970 22349 14026
rect 22405 13970 22430 14026
rect 22486 13970 22511 14026
rect 22567 13970 22592 14026
rect 22648 13970 22673 14026
rect 22729 13970 22753 14026
rect 22809 13970 22833 14026
rect 22889 13970 22913 14026
rect 22969 14024 23448 14026
rect 22969 13970 23254 14024
rect 22097 13968 23254 13970
rect 23310 13968 23392 14024
rect 22097 13926 23448 13968
rect 22097 13924 23254 13926
rect 22097 13868 22106 13924
rect 22162 13868 22187 13924
rect 22243 13868 22268 13924
rect 22324 13868 22349 13924
rect 22405 13868 22430 13924
rect 22486 13868 22511 13924
rect 22567 13868 22592 13924
rect 22648 13868 22673 13924
rect 22729 13868 22753 13924
rect 22809 13868 22833 13924
rect 22889 13868 22913 13924
rect 22969 13870 23254 13924
rect 23310 13870 23392 13926
rect 22969 13868 23448 13870
rect 22097 13828 23448 13868
rect 22097 13822 23254 13828
rect 22097 13766 22106 13822
rect 22162 13766 22187 13822
rect 22243 13766 22268 13822
rect 22324 13766 22349 13822
rect 22405 13766 22430 13822
rect 22486 13766 22511 13822
rect 22567 13766 22592 13822
rect 22648 13766 22673 13822
rect 22729 13766 22753 13822
rect 22809 13766 22833 13822
rect 22889 13766 22913 13822
rect 22969 13772 23254 13822
rect 23310 13772 23392 13828
rect 22969 13766 23448 13772
rect 22097 13763 23448 13766
rect 818 12856 827 12865
rect 883 12856 949 12865
rect 1005 12856 1014 12865
rect 818 12804 826 12856
rect 883 12809 890 12856
rect 878 12804 890 12809
rect 942 12809 949 12856
rect 942 12804 954 12809
rect 1006 12804 1014 12856
rect 818 12785 1014 12804
rect 818 12781 827 12785
rect 883 12781 949 12785
rect 1005 12781 1014 12785
rect 818 12729 826 12781
rect 883 12729 890 12781
rect 942 12729 949 12781
rect 1006 12729 1014 12781
rect 818 12705 1014 12729
rect 818 12653 826 12705
rect 883 12653 890 12705
rect 942 12653 949 12705
rect 1006 12653 1014 12705
rect 818 12649 827 12653
rect 883 12649 949 12653
rect 1005 12649 1014 12653
rect 818 12629 1014 12649
rect 818 12577 826 12629
rect 878 12625 890 12629
rect 883 12577 890 12625
rect 942 12625 954 12629
rect 942 12577 949 12625
rect 1006 12577 1014 12629
rect 23777 12717 25385 12753
rect 23777 12661 23786 12717
rect 23842 12661 23868 12717
rect 23924 12661 23950 12717
rect 24006 12661 24031 12717
rect 24087 12661 24112 12717
rect 24168 12661 25385 12717
rect 23777 12625 25385 12661
rect 818 12569 827 12577
rect 883 12569 949 12577
rect 1005 12569 1014 12577
rect 15769 11531 15778 11587
rect 15834 11531 15858 11587
rect 15914 11531 15923 11587
rect 3491 11463 3500 11519
rect 3556 11463 3645 11519
rect 3701 11463 3710 11519
rect 3491 11439 3710 11463
rect 3491 11383 3500 11439
rect 3556 11383 3645 11439
rect 3701 11383 3710 11439
rect 20071 11496 20519 11536
rect 20071 11440 20132 11496
rect 20188 11440 20213 11496
rect 20269 11440 20294 11496
rect 20350 11440 20374 11496
rect 20430 11440 20454 11496
rect 20510 11440 20519 11496
tri 26374 11440 26383 11449 se
rect 26383 11440 26441 14404
rect 20071 11420 20519 11440
tri 26354 11420 26374 11440 se
rect 26374 11422 26441 11440
rect 26374 11420 26439 11422
tri 26439 11420 26441 11422 nw
rect 25801 11368 25807 11420
rect 25859 11368 25871 11420
rect 25923 11383 26402 11420
tri 26402 11383 26439 11420 nw
rect 25923 11368 26387 11383
tri 26387 11368 26402 11383 nw
rect 26511 11313 26569 14456
tri 26569 14430 26595 14456 nw
rect 27562 13627 28065 13628
rect 27105 13623 27302 13624
rect 27105 13571 27111 13623
rect 27163 13571 27178 13623
rect 27230 13571 27244 13623
rect 27296 13571 27302 13623
rect 27105 13553 27302 13571
rect 27105 13501 27111 13553
rect 27163 13501 27178 13553
rect 27230 13501 27244 13553
rect 27296 13501 27302 13553
rect 27105 13483 27302 13501
rect 27105 13431 27111 13483
rect 27163 13431 27178 13483
rect 27230 13431 27244 13483
rect 27296 13431 27302 13483
rect 27562 13575 27568 13627
rect 27620 13575 27632 13627
rect 27684 13575 28065 13627
rect 27562 13557 28065 13575
rect 27562 13505 27568 13557
rect 27620 13505 27632 13557
rect 27684 13505 28065 13557
rect 27562 13487 28065 13505
rect 27562 13435 27568 13487
rect 27620 13435 27632 13487
rect 27684 13435 28065 13487
rect 27562 13434 28065 13435
rect 27105 12934 27302 13431
tri 27866 13366 27934 13434 ne
rect 27934 12936 28065 13434
rect 27105 12882 27111 12934
rect 27163 12882 27178 12934
rect 27230 12882 27244 12934
rect 27296 12882 27302 12934
rect 27105 12864 27302 12882
rect 27105 12812 27111 12864
rect 27163 12812 27178 12864
rect 27230 12812 27244 12864
rect 27296 12812 27302 12864
rect 27105 12794 27302 12812
rect 27105 12742 27111 12794
rect 27163 12742 27178 12794
rect 27230 12742 27244 12794
rect 27296 12742 27302 12794
rect 27105 12741 27302 12742
rect 27365 12934 27562 12935
rect 27365 12882 27371 12934
rect 27423 12882 27438 12934
rect 27490 12882 27504 12934
rect 27556 12882 27562 12934
rect 27365 12864 27562 12882
rect 27365 12812 27371 12864
rect 27423 12812 27438 12864
rect 27490 12812 27504 12864
rect 27556 12812 27562 12864
rect 27365 12794 27562 12812
rect 27365 12742 27371 12794
rect 27423 12742 27438 12794
rect 27490 12742 27504 12794
rect 27556 12742 27562 12794
rect 27934 12884 27974 12936
rect 28026 12884 28065 12936
rect 27934 12866 28065 12884
rect 27934 12814 27974 12866
rect 28026 12814 28065 12866
rect 27934 12796 28065 12814
rect 27934 12744 27974 12796
rect 28026 12744 28065 12796
rect 27934 12743 28065 12744
rect 27365 12741 27562 12742
rect 14445 11282 14501 11291
rect 14445 11202 14501 11226
rect 14445 11137 14501 11146
rect 27471 11095 27832 11103
rect 27523 11043 27565 11095
rect 27617 11043 27832 11095
rect 27471 11000 27832 11043
tri 13425 10941 13471 10987 se
rect 13471 10941 13668 10987
rect 13425 10935 13668 10941
rect 13720 10935 13732 10987
rect 13784 10935 13790 10987
rect 27523 10948 27565 11000
rect 27617 10948 27832 11000
rect 13425 10930 13510 10935
tri 13510 10930 13515 10935 nw
rect 221 10733 226 10785
rect 278 10733 282 10785
rect 700 10926 756 10930
rect 13425 10926 13506 10930
tri 13506 10926 13510 10930 nw
rect 700 10921 759 10926
rect 756 10920 759 10921
rect 756 10865 759 10868
rect 700 10856 759 10865
rect 700 10841 707 10856
rect 756 10798 759 10804
rect 700 10776 756 10785
rect 221 10721 282 10733
rect 221 10669 226 10721
rect 278 10669 282 10721
rect 221 10662 282 10669
rect 1151 10765 1207 10774
rect 1151 10705 1153 10709
rect 1205 10705 1207 10709
rect 1151 10693 1207 10705
rect 1151 10685 1153 10693
rect 1205 10685 1207 10693
rect 1151 10620 1207 10629
rect 10336 10648 10392 10657
rect 10336 10583 10392 10592
rect 10388 10568 10392 10583
rect 10336 10503 10392 10512
rect 3309 10221 3318 10277
rect 3374 10221 3422 10277
rect 3478 10221 3526 10277
rect 3582 10221 3630 10277
rect 3686 10221 3695 10277
rect 3309 10197 3695 10221
rect 3309 10141 3318 10197
rect 3374 10141 3422 10197
rect 3478 10141 3526 10197
rect 3582 10141 3630 10197
rect 3686 10141 3695 10197
rect 9879 10121 10069 10130
rect 9935 10065 10013 10121
rect 9879 10025 10069 10065
rect 3309 9947 3318 10003
rect 3374 9947 3422 10003
rect 3478 9947 3526 10003
rect 3582 9947 3630 10003
rect 3686 9947 3695 10003
rect 3309 9923 3695 9947
rect 3309 9867 3318 9923
rect 3374 9867 3422 9923
rect 3478 9867 3526 9923
rect 3582 9867 3630 9923
rect 3686 9867 3695 9923
rect 9935 9969 10013 10025
tri 13400 10013 13425 10038 se
rect 13425 10013 13471 10926
tri 13471 10891 13506 10926 nw
rect 17875 10829 17884 10885
rect 17940 10829 18004 10885
rect 18060 10829 18123 10885
rect 18179 10829 18188 10885
rect 17875 10759 18188 10829
rect 17875 10703 17884 10759
rect 17940 10703 18004 10759
rect 18060 10703 18123 10759
rect 18179 10703 18188 10759
rect 24599 10843 24895 10852
rect 24655 10787 24679 10843
rect 24735 10787 24759 10843
rect 24815 10787 24839 10843
rect 24599 10758 24895 10787
rect 24655 10742 24679 10758
rect 24735 10742 24759 10758
rect 24599 10690 24614 10702
rect 24666 10690 24678 10742
rect 24735 10702 24742 10742
rect 24815 10702 24839 10758
rect 24730 10690 24742 10702
rect 24794 10690 24895 10702
rect 24599 10676 24895 10690
rect 24599 10673 24614 10676
rect 24666 10624 24678 10676
rect 24730 10673 24742 10676
rect 24794 10673 24895 10676
rect 24735 10624 24742 10673
rect 24655 10617 24679 10624
rect 24735 10617 24759 10624
rect 24815 10617 24839 10673
rect 24599 10610 24895 10617
rect 24599 10588 24614 10610
rect 24666 10558 24678 10610
rect 24730 10588 24742 10610
rect 24794 10588 24895 10610
rect 24735 10558 24742 10588
rect 24655 10543 24679 10558
rect 24735 10543 24759 10558
rect 24599 10502 24614 10532
rect 24666 10491 24678 10543
rect 24735 10532 24742 10543
rect 24815 10532 24839 10588
rect 24730 10502 24742 10532
rect 24794 10502 24895 10532
rect 24735 10491 24742 10502
rect 24655 10476 24679 10491
rect 24735 10476 24759 10491
rect 24599 10424 24614 10446
rect 24666 10424 24678 10476
rect 24735 10446 24742 10476
rect 24815 10446 24839 10502
rect 24730 10424 24742 10446
rect 24794 10424 24895 10446
rect 24599 10416 24895 10424
rect 24655 10409 24679 10416
rect 24735 10409 24759 10416
rect 24599 10357 24614 10360
rect 24666 10357 24678 10409
rect 24735 10360 24742 10409
rect 24815 10360 24839 10416
rect 24730 10357 24742 10360
rect 24794 10357 24895 10360
rect 24599 10351 24895 10357
rect 27471 10589 27832 10948
rect 27523 10537 27565 10589
rect 27617 10537 27832 10589
rect 27471 10494 27832 10537
rect 27523 10442 27565 10494
rect 27617 10442 27832 10494
tri 15566 10288 15570 10292 se
rect 15570 10288 15579 10292
rect 14195 10236 14201 10288
rect 14253 10236 14265 10288
rect 14317 10236 15579 10288
rect 15635 10236 15659 10292
rect 15715 10236 15724 10292
rect 9879 9929 10069 9969
rect 9935 9873 10013 9929
rect 9879 9833 10069 9873
rect 13223 10004 13471 10013
rect 13279 9964 13471 10004
rect 13223 9924 13279 9948
tri 13279 9943 13300 9964 nw
rect 13223 9859 13279 9868
rect 9935 9777 10013 9833
rect 9879 9768 10069 9777
rect 25285 9381 25341 9390
rect 25285 9301 25341 9325
rect 24635 9238 24641 9290
rect 24693 9238 24705 9290
rect 24757 9245 25285 9290
rect 24757 9238 25341 9245
rect 25285 9236 25341 9238
rect 27471 9052 27832 10442
rect 27243 9043 27832 9052
rect 27299 8987 27323 9043
rect 27379 8987 27403 9043
rect 27459 8987 27483 9043
rect 27539 8987 27832 9043
tri 573 8832 717 8976 ne
rect 717 8832 975 8976
tri 975 8832 1119 8976 nw
rect 27243 8954 27832 8987
rect 27299 8898 27323 8954
rect 27379 8898 27403 8954
rect 27459 8898 27483 8954
rect 27539 8898 27832 8954
rect 27243 8865 27832 8898
tri 717 8825 724 8832 ne
rect 724 6760 975 8832
rect 27299 8809 27323 8865
rect 27379 8809 27403 8865
rect 27459 8809 27483 8865
rect 27539 8809 27832 8865
rect 27243 8776 27832 8809
rect 27299 8720 27323 8776
rect 27379 8720 27403 8776
rect 27459 8720 27483 8776
rect 27539 8720 27832 8776
rect 27243 8686 27832 8720
rect 27299 8630 27323 8686
rect 27379 8630 27403 8686
rect 27459 8630 27483 8686
rect 27539 8630 27832 8686
rect 27243 8621 27832 8630
rect 2794 8138 2850 8147
tri 2850 8085 2862 8097 sw
rect 2850 8082 2862 8085
rect 2794 8076 2862 8082
tri 2862 8076 2871 8085 sw
rect 2794 8063 2871 8076
tri 2871 8063 2884 8076 sw
rect 2794 8058 5891 8063
rect 2850 8011 5891 8058
rect 2850 8002 2859 8011
tri 2859 8002 2868 8011 nw
tri 5805 8002 5814 8011 ne
rect 5814 8002 5891 8011
rect 2794 7993 2850 8002
tri 2850 7993 2859 8002 nw
tri 5814 7993 5823 8002 ne
rect 5823 7993 5891 8002
tri 5823 7980 5836 7993 ne
rect 5836 7980 5891 7993
tri 5836 7977 5839 7980 ne
rect 5839 7695 5891 7980
rect 9728 8033 12598 8085
rect 9728 8002 9783 8033
tri 9783 8002 9814 8033 nw
tri 12512 8002 12543 8033 ne
rect 12543 8002 12598 8033
tri 5891 7695 5925 7729 sw
tri 7385 7695 7419 7729 se
rect 7419 7726 8329 7778
rect 7419 7695 7471 7726
rect 5839 7643 7471 7695
tri 7471 7692 7505 7726 nw
tri 8243 7692 8277 7726 ne
rect 8277 7696 8329 7726
tri 8329 7696 8363 7730 sw
tri 8980 7696 9014 7730 se
rect 9014 7696 9589 7736
tri 9589 7696 9623 7730 sw
tri 9694 7696 9728 7730 se
rect 9728 7696 9780 8002
tri 9780 7999 9783 8002 nw
tri 12543 7999 12546 8002 ne
rect 12546 7942 12598 8002
rect 22385 8076 22391 8128
rect 22443 8123 22463 8128
rect 22515 8123 22535 8128
rect 22587 8123 22606 8128
rect 22658 8123 22677 8128
rect 22729 8123 22748 8128
rect 22800 8123 22819 8128
rect 22871 8123 22890 8128
rect 22450 8076 22463 8123
rect 22532 8076 22535 8123
rect 22800 8076 22802 8123
rect 22871 8076 22883 8123
rect 22942 8076 22948 8128
rect 22385 8067 22394 8076
rect 22450 8067 22476 8076
rect 22532 8067 22558 8076
rect 22614 8067 22640 8076
rect 22696 8067 22721 8076
rect 22777 8067 22802 8076
rect 22858 8067 22883 8076
rect 22939 8067 22948 8076
rect 22385 8054 22948 8067
rect 22385 8002 22391 8054
rect 22443 8002 22463 8054
rect 22515 8002 22535 8054
rect 22587 8002 22606 8054
rect 22658 8002 22677 8054
rect 22729 8002 22748 8054
rect 22800 8002 22819 8054
rect 22871 8002 22890 8054
rect 22942 8002 22948 8054
rect 22385 7999 22948 8002
rect 22385 7980 22394 7999
rect 22450 7980 22476 7999
rect 22532 7980 22558 7999
rect 22614 7980 22640 7999
rect 22696 7980 22721 7999
rect 22777 7980 22802 7999
rect 22858 7980 22883 7999
rect 22939 7980 22948 7999
tri 12598 7942 12626 7970 sw
rect 12546 7936 12626 7942
tri 12626 7936 12632 7942 sw
tri 13306 7936 13312 7942 se
rect 13312 7936 13368 7942
rect 12546 7933 13368 7936
rect 12546 7884 13312 7933
tri 13278 7850 13312 7884 ne
rect 22385 7928 22391 7980
rect 22450 7943 22463 7980
rect 22532 7943 22535 7980
rect 22800 7943 22802 7980
rect 22871 7943 22883 7980
rect 22443 7928 22463 7943
rect 22515 7928 22535 7943
rect 22587 7928 22606 7943
rect 22658 7928 22677 7943
rect 22729 7928 22748 7943
rect 22800 7928 22819 7943
rect 22871 7928 22890 7943
rect 22942 7928 22948 7980
rect 13312 7853 13368 7877
rect 13312 7788 13368 7797
rect 8277 7684 9780 7696
rect 8277 7644 9066 7684
tri 9066 7650 9100 7684 nw
tri 9503 7650 9537 7684 ne
rect 9537 7644 9780 7684
rect 14405 7552 14461 7561
tri 14368 7461 14405 7498 se
rect 14405 7472 14461 7496
rect 13273 7405 13282 7461
rect 13338 7405 13362 7461
rect 13418 7459 13427 7461
tri 13427 7459 13429 7461 sw
tri 14366 7459 14368 7461 se
rect 14368 7459 14405 7461
rect 13418 7416 14405 7459
rect 13418 7407 14461 7416
rect 13418 7405 13427 7407
tri 13427 7405 13429 7407 nw
rect 24139 7228 24196 7382
rect 3804 7083 3813 7139
rect 3873 7087 3885 7139
rect 3869 7083 3893 7087
rect 3949 7083 3958 7139
rect 24682 7026 24773 7157
tri 24682 7003 24705 7026 ne
rect 24705 7003 24773 7026
rect 1151 6987 1811 6996
rect 1207 6931 1755 6987
tri 15793 6949 15818 6974 se
rect 15818 6965 15874 6974
rect 1151 6907 1811 6931
rect 1207 6851 1755 6907
tri 13491 6891 13549 6949 se
rect 13549 6909 15818 6949
rect 13549 6908 15874 6909
tri 13549 6891 13566 6908 nw
tri 15784 6891 15801 6908 ne
rect 15801 6891 15874 6908
tri 13490 6890 13491 6891 se
rect 13491 6890 13508 6891
tri 975 6760 1063 6848 sw
rect 1151 6842 1811 6851
rect 2378 6834 2387 6890
rect 2443 6834 2467 6890
rect 2523 6834 3813 6890
rect 3869 6834 3893 6890
rect 3949 6834 3958 6890
tri 13450 6850 13490 6890 se
rect 13490 6850 13508 6890
tri 13508 6850 13549 6891 nw
tri 15801 6874 15818 6891 ne
rect 15818 6885 15874 6891
tri 13184 6834 13200 6850 se
rect 13200 6834 13478 6850
tri 13170 6820 13184 6834 se
rect 13184 6820 13478 6834
tri 13478 6820 13508 6850 nw
rect 15818 6820 15874 6829
rect 26164 6877 26220 6886
tri 13169 6819 13170 6820 se
rect 13170 6819 13477 6820
tri 13477 6819 13478 6820 nw
tri 10702 6760 10761 6819 se
rect 10761 6810 13468 6819
tri 13468 6810 13477 6819 nw
rect 10761 6778 13186 6810
tri 13186 6778 13218 6810 nw
rect 26164 6797 26220 6821
rect 724 6757 5555 6760
rect 724 6719 5216 6757
tri 724 6560 883 6719 ne
rect 883 6701 5216 6719
rect 5272 6701 5307 6757
rect 5363 6701 5397 6757
rect 5453 6701 5487 6757
rect 5543 6701 5555 6757
tri 10696 6754 10702 6760 se
rect 10702 6754 10761 6760
tri 10761 6754 10785 6778 nw
tri 10674 6732 10696 6754 se
rect 10696 6732 10739 6754
tri 10739 6732 10761 6754 nw
rect 26164 6732 26220 6741
rect 883 6619 5555 6701
tri 10631 6689 10674 6732 se
rect 10674 6689 10696 6732
tri 10696 6689 10739 6732 nw
tri 10566 6624 10631 6689 se
rect 10631 6668 10675 6689
tri 10675 6668 10696 6689 nw
rect 10631 6666 10673 6668
tri 10673 6666 10675 6668 nw
tri 10732 6666 10734 6668 se
rect 10734 6666 20452 6668
tri 10631 6624 10673 6666 nw
tri 10690 6624 10732 6666 se
rect 10732 6627 20452 6666
rect 10732 6624 10734 6627
rect 883 6563 5216 6619
rect 5272 6563 5307 6619
rect 5363 6563 5397 6619
rect 5453 6563 5487 6619
rect 5543 6563 5555 6619
rect 883 6560 5555 6563
tri 10502 6560 10566 6624 se
rect 10566 6607 10614 6624
tri 10614 6607 10631 6624 nw
tri 10673 6607 10690 6624 se
rect 10690 6607 10734 6624
tri 10734 6607 10754 6627 nw
rect 10566 6605 10612 6607
tri 10612 6605 10614 6607 nw
tri 10671 6605 10673 6607 se
tri 10501 6559 10502 6560 se
rect 10502 6559 10566 6560
tri 10566 6559 10612 6605 nw
tri 10625 6559 10671 6605 se
rect 10671 6559 10673 6605
tri 10465 6523 10501 6559 se
rect 10501 6546 10553 6559
tri 10553 6546 10566 6559 nw
tri 10612 6546 10625 6559 se
rect 10625 6546 10673 6559
tri 10673 6546 10734 6607 nw
rect 10501 6544 10551 6546
tri 10551 6544 10553 6546 nw
tri 10610 6544 10612 6546 se
rect 10501 6523 10530 6544
tri 10530 6523 10551 6544 nw
tri 10589 6523 10610 6544 se
rect 10610 6523 10612 6544
tri 1620 6520 1623 6523 se
rect 1623 6520 10527 6523
tri 10527 6520 10530 6523 nw
tri 10586 6520 10589 6523 se
rect 10589 6520 10612 6523
rect 1539 6464 1548 6520
rect 1604 6464 1628 6520
rect 1684 6485 10492 6520
tri 10492 6485 10527 6520 nw
tri 10551 6485 10586 6520 se
rect 10586 6485 10612 6520
tri 10612 6485 10673 6546 nw
rect 1684 6482 10489 6485
tri 10489 6482 10492 6485 nw
tri 10548 6482 10551 6485 se
rect 10551 6482 10577 6485
rect 1684 6464 1696 6482
tri 1696 6464 1714 6482 nw
tri 10530 6464 10548 6482 se
rect 10548 6464 10577 6482
tri 10520 6454 10530 6464 se
rect 10530 6454 10577 6464
rect 2924 6402 2930 6454
rect 2982 6403 2995 6454
rect 3239 6403 3245 6454
tri 10516 6450 10520 6454 se
rect 10520 6450 10577 6454
tri 10577 6450 10612 6485 nw
rect 2924 6390 2934 6402
rect 1398 6376 1454 6385
tri 1454 6369 1468 6383 sw
rect 2257 6376 2313 6385
rect 1454 6346 1468 6369
tri 1468 6346 1491 6369 sw
tri 2234 6346 2257 6369 se
rect 1454 6320 2257 6346
rect 2924 6338 2930 6390
rect 2990 6347 2995 6403
rect 3239 6347 3247 6403
rect 2982 6338 2995 6347
rect 3239 6338 3245 6347
rect 4138 6343 4147 6399
rect 4203 6343 4227 6399
rect 4283 6378 4292 6399
rect 4416 6394 4434 6450
rect 4490 6394 4514 6450
rect 4570 6409 10536 6450
tri 10536 6409 10577 6450 nw
rect 4570 6394 4579 6409
tri 4579 6394 4594 6409 nw
rect 14026 6378 14032 6390
rect 4283 6352 4314 6378
tri 4314 6352 4340 6378 sw
tri 4688 6352 4714 6378 se
rect 4714 6352 7400 6378
rect 4283 6350 7400 6352
tri 7400 6350 7428 6378 sw
tri 8178 6350 8206 6378 se
rect 8206 6350 14032 6378
rect 4283 6343 7428 6350
tri 7428 6343 7435 6350 sw
tri 8171 6343 8178 6350 se
rect 8178 6343 14032 6350
rect 4138 6338 7435 6343
tri 7435 6338 7440 6343 sw
tri 8166 6338 8171 6343 se
rect 8171 6338 14032 6343
rect 14084 6338 14096 6390
rect 14148 6338 14154 6390
rect 1398 6296 2313 6320
tri 4285 6312 4311 6338 ne
rect 4311 6312 4717 6338
tri 4717 6312 4743 6338 nw
tri 7387 6312 7413 6338 ne
rect 7413 6332 7440 6338
tri 7440 6332 7446 6338 sw
tri 8160 6332 8166 6338 se
rect 8166 6332 8213 6338
tri 8213 6332 8219 6338 nw
rect 7413 6325 7446 6332
tri 7446 6325 7453 6332 sw
tri 8153 6325 8160 6332 se
rect 8160 6325 8206 6332
tri 8206 6325 8213 6332 nw
rect 7413 6312 7453 6325
tri 7413 6297 7428 6312 ne
rect 7428 6311 7453 6312
tri 7453 6311 7467 6325 sw
tri 8139 6311 8153 6325 se
rect 8153 6311 8192 6325
tri 8192 6311 8206 6325 nw
rect 23986 6323 24042 6332
rect 7428 6297 7467 6311
tri 7467 6297 7481 6311 sw
tri 8125 6297 8139 6311 se
rect 8139 6297 8166 6311
rect 1454 6275 2257 6296
rect 1398 6231 1454 6240
tri 1454 6238 1491 6275 nw
tri 2229 6247 2257 6275 ne
tri 7428 6292 7433 6297 ne
rect 7433 6292 7481 6297
tri 3747 6285 3754 6292 se
rect 3754 6285 4265 6292
tri 4265 6285 4272 6292 sw
tri 4758 6285 4765 6292 se
rect 4765 6285 7363 6292
tri 7363 6285 7370 6292 sw
tri 7433 6285 7440 6292 ne
rect 7440 6285 7481 6292
tri 7481 6285 7493 6297 sw
tri 8113 6285 8125 6297 se
rect 8125 6285 8166 6297
tri 8166 6285 8192 6311 nw
tri 23967 6292 23986 6311 se
tri 8305 6285 8312 6292 se
rect 8312 6285 9520 6292
tri 9520 6285 9527 6292 sw
tri 23960 6285 23967 6292 se
rect 23967 6285 23986 6292
tri 3743 6281 3747 6285 se
rect 3747 6281 4272 6285
tri 4272 6281 4276 6285 sw
tri 4754 6281 4758 6285 se
rect 4758 6281 7370 6285
rect 2257 6231 2313 6240
tri 3700 6238 3743 6281 se
rect 3743 6244 7370 6281
tri 7370 6244 7411 6285 sw
tri 7440 6244 7481 6285 ne
rect 7481 6272 7493 6285
tri 7493 6272 7506 6285 sw
tri 8100 6272 8113 6285 se
rect 8113 6272 8153 6285
tri 8153 6272 8166 6285 nw
tri 8304 6284 8305 6285 se
rect 8305 6284 9527 6285
tri 9527 6284 9528 6285 sw
tri 10502 6284 10503 6285 se
rect 10503 6284 13065 6285
tri 8292 6272 8304 6284 se
rect 8304 6272 9528 6284
tri 9528 6272 9540 6284 sw
tri 10490 6272 10502 6284 se
rect 10502 6272 13065 6284
rect 7481 6244 7506 6272
tri 7506 6244 7534 6272 sw
tri 8072 6244 8100 6272 se
rect 8100 6244 8114 6272
rect 3743 6240 7411 6244
rect 3743 6238 3774 6240
tri 3774 6238 3776 6240 nw
tri 7341 6238 7343 6240 ne
rect 7343 6238 7411 6240
tri 7411 6238 7417 6244 sw
tri 7481 6238 7487 6244 ne
rect 7487 6238 7534 6244
tri 3695 6233 3700 6238 se
rect 3700 6233 3769 6238
tri 3769 6233 3774 6238 nw
tri 7343 6233 7348 6238 ne
rect 7348 6234 7417 6238
tri 7417 6234 7421 6238 sw
tri 7487 6234 7491 6238 ne
rect 7491 6234 7534 6238
rect 7348 6233 7421 6234
tri 7421 6233 7422 6234 sw
tri 7491 6233 7492 6234 ne
rect 7492 6233 7534 6234
tri 7534 6233 7545 6244 sw
tri 8061 6233 8072 6244 se
rect 8072 6233 8114 6244
tri 8114 6233 8153 6272 nw
tri 8253 6233 8292 6272 se
rect 8292 6240 9540 6272
rect 8292 6233 8327 6240
tri 8327 6233 8334 6240 nw
tri 9507 6233 9514 6240 ne
rect 9514 6233 9540 6240
tri 9540 6233 9579 6272 sw
tri 10451 6233 10490 6272 se
rect 10490 6233 13065 6272
rect 13117 6233 13129 6285
rect 13181 6233 13187 6285
tri 23954 6279 23960 6285 se
rect 23960 6279 23986 6285
tri 15636 6277 15638 6279 se
rect 15638 6277 15696 6279
tri 15696 6277 15698 6279 sw
tri 23952 6277 23954 6279 se
rect 23954 6277 23986 6279
tri 15635 6276 15636 6277 se
rect 15636 6276 15698 6277
tri 15698 6276 15699 6277 sw
rect 15635 6270 15641 6276
rect 15693 6270 15705 6276
tri 3693 6231 3695 6233 se
rect 3695 6231 3760 6233
tri 3686 6224 3693 6231 se
rect 3693 6224 3760 6231
tri 3760 6224 3769 6233 nw
tri 7348 6224 7357 6233 ne
rect 7357 6231 7422 6233
tri 7422 6231 7424 6233 sw
tri 7492 6231 7494 6233 ne
rect 7494 6231 7545 6233
tri 7545 6231 7547 6233 sw
tri 8059 6231 8061 6233 se
rect 8061 6231 8105 6233
rect 7357 6224 7424 6231
tri 7424 6224 7431 6231 sw
tri 7494 6224 7501 6231 ne
rect 7501 6224 7547 6231
tri 7547 6224 7554 6231 sw
tri 8052 6224 8059 6231 se
rect 8059 6224 8105 6231
tri 8105 6224 8114 6233 nw
tri 8244 6224 8253 6233 se
rect 8253 6224 8318 6233
tri 8318 6224 8327 6233 nw
tri 9514 6224 9523 6233 ne
rect 9523 6224 9579 6233
tri 9579 6224 9588 6233 sw
tri 10442 6224 10451 6233 se
rect 10451 6224 10516 6233
tri 10516 6224 10525 6233 nw
rect 15635 6224 15640 6270
rect 15696 6224 15705 6270
rect 15757 6224 15763 6276
rect 23585 6225 23591 6277
rect 23643 6225 23655 6277
rect 23707 6267 23986 6277
rect 23707 6243 24042 6267
rect 23707 6225 23986 6243
tri 23952 6224 23953 6225 ne
rect 23953 6224 23986 6225
tri 3680 6218 3686 6224 se
rect 3686 6218 3754 6224
tri 3754 6218 3760 6224 nw
tri 7357 6218 7363 6224 ne
rect 7363 6218 7431 6224
tri 3668 6206 3680 6218 se
rect 3680 6206 3742 6218
tri 3742 6206 3754 6218 nw
tri 7363 6206 7375 6218 ne
rect 7375 6206 7431 6218
rect 3668 6196 3732 6206
tri 3732 6196 3742 6206 nw
tri 7375 6196 7385 6206 ne
rect 7385 6196 7431 6206
tri 7431 6196 7459 6224 sw
tri 7501 6196 7529 6224 ne
rect 7529 6219 7554 6224
tri 7554 6219 7559 6224 sw
tri 8047 6219 8052 6224 se
rect 8052 6219 8100 6224
tri 8100 6219 8105 6224 nw
tri 8239 6219 8244 6224 se
rect 8244 6219 8313 6224
tri 8313 6219 8318 6224 nw
tri 9523 6219 9528 6224 ne
rect 9528 6219 9588 6224
tri 9588 6219 9593 6224 sw
tri 10437 6219 10442 6224 se
rect 10442 6219 10511 6224
tri 10511 6219 10516 6224 nw
tri 15635 6219 15640 6224 ne
rect 7529 6196 7559 6219
tri 7559 6196 7582 6219 sw
tri 8024 6196 8047 6219 se
rect 8047 6196 8077 6219
tri 8077 6196 8100 6219 nw
tri 8238 6218 8239 6219 se
rect 8239 6218 8312 6219
tri 8312 6218 8313 6219 nw
tri 9528 6218 9529 6219 ne
rect 9529 6218 10488 6219
tri 8216 6196 8238 6218 se
rect 8238 6196 8290 6218
tri 8290 6196 8312 6218 nw
tri 9529 6196 9551 6218 ne
rect 9551 6196 10488 6218
tri 10488 6196 10511 6219 nw
rect 15696 6214 15702 6224
rect 15640 6196 15702 6214
tri 15702 6196 15730 6224 nw
tri 23953 6196 23981 6224 ne
rect 23981 6196 23986 6224
rect 3668 6195 3731 6196
tri 3731 6195 3732 6196 nw
rect 5940 6195 6540 6196
tri 7385 6195 7386 6196 ne
rect 7386 6195 7459 6196
tri 7459 6195 7460 6196 sw
tri 7529 6195 7530 6196 ne
rect 7530 6195 7582 6196
tri 7582 6195 7583 6196 sw
tri 8023 6195 8024 6196 se
rect 8024 6195 8076 6196
tri 8076 6195 8077 6196 nw
tri 8215 6195 8216 6196 se
rect 8216 6195 8289 6196
tri 8289 6195 8290 6196 nw
tri 9551 6195 9552 6196 ne
rect 9552 6195 10487 6196
tri 10487 6195 10488 6196 nw
rect 12225 6195 12825 6196
rect 3668 5679 3720 6195
tri 3720 6184 3731 6195 nw
rect 4432 6166 4488 6175
rect 4432 6086 4488 6110
rect 4432 6021 4488 6030
rect 5940 6143 5946 6195
rect 6005 6143 6013 6195
rect 6199 6143 6213 6195
rect 6269 6143 6281 6195
rect 6467 6143 6475 6195
rect 6534 6143 6540 6195
tri 7386 6164 7417 6195 ne
rect 7417 6191 7460 6195
tri 7460 6191 7464 6195 sw
tri 7530 6191 7534 6195 ne
rect 7534 6191 7583 6195
tri 7583 6191 7587 6195 sw
tri 8019 6191 8023 6195 se
rect 8023 6191 8072 6195
tri 8072 6191 8076 6195 nw
tri 8211 6191 8215 6195 se
rect 8215 6191 8238 6195
rect 7417 6164 7464 6191
tri 7464 6164 7491 6191 sw
tri 7534 6164 7561 6191 ne
rect 7561 6164 8032 6191
tri 7417 6143 7438 6164 ne
rect 7438 6160 7491 6164
tri 7491 6160 7495 6164 sw
tri 7561 6160 7565 6164 ne
rect 7565 6160 8032 6164
rect 7438 6151 7495 6160
tri 7495 6151 7504 6160 sw
tri 7565 6151 7574 6160 ne
rect 7574 6151 8032 6160
tri 8032 6151 8072 6191 nw
tri 8171 6151 8211 6191 se
rect 8211 6151 8238 6191
rect 7438 6144 7504 6151
tri 7504 6144 7511 6151 sw
tri 8164 6144 8171 6151 se
rect 8171 6144 8238 6151
tri 8238 6144 8289 6195 nw
tri 9552 6167 9580 6195 ne
rect 9580 6167 10459 6195
tri 10459 6167 10487 6195 nw
rect 7438 6143 7511 6144
tri 7511 6143 7512 6144 sw
tri 8163 6143 8164 6144 se
rect 8164 6143 8237 6144
tri 8237 6143 8238 6144 nw
rect 12225 6143 12231 6195
rect 12290 6143 12298 6195
rect 12484 6143 12498 6195
rect 12554 6143 12566 6195
rect 12752 6143 12760 6195
rect 12819 6143 12825 6195
rect 5940 6139 5949 6143
rect 6005 6139 6037 6143
rect 6093 6139 6125 6143
rect 6181 6139 6213 6143
rect 6269 6139 6301 6143
rect 6357 6139 6388 6143
rect 6444 6139 6475 6143
rect 6531 6139 6540 6143
rect 5940 6121 6540 6139
tri 7438 6121 7460 6143 ne
rect 7460 6121 7512 6143
tri 7512 6121 7534 6143 sw
tri 8141 6121 8163 6143 se
rect 8163 6121 8215 6143
tri 8215 6121 8237 6143 nw
rect 12225 6139 12234 6143
rect 12290 6139 12322 6143
rect 12378 6139 12410 6143
rect 12466 6139 12498 6143
rect 12554 6139 12586 6143
rect 12642 6139 12673 6143
rect 12729 6139 12760 6143
rect 12816 6139 12825 6143
rect 12225 6121 12825 6139
rect 15640 6195 15701 6196
tri 15701 6195 15702 6196 nw
rect 16057 6195 16657 6196
rect 15640 6190 15696 6195
tri 15696 6190 15701 6195 nw
rect 15640 6125 15696 6134
rect 16057 6143 16076 6195
rect 16135 6143 16142 6195
rect 16326 6143 16337 6195
rect 16393 6143 16404 6195
rect 16586 6143 16592 6195
rect 16651 6143 16657 6195
rect 16057 6139 16079 6143
rect 16135 6139 16165 6143
rect 16221 6139 16251 6143
rect 16307 6139 16337 6143
rect 16393 6139 16422 6143
rect 16478 6139 16507 6143
rect 16563 6139 16592 6143
rect 16648 6139 16657 6143
rect 5940 6069 5946 6121
rect 5998 6069 6013 6121
rect 6065 6069 6080 6121
rect 6132 6069 6147 6121
rect 6199 6069 6214 6121
rect 6266 6069 6281 6121
rect 6333 6069 6348 6121
rect 6400 6069 6415 6121
rect 6467 6069 6482 6121
rect 6534 6069 6540 6121
tri 7460 6090 7491 6121 ne
rect 7491 6090 7534 6121
tri 7534 6090 7565 6121 sw
tri 8110 6090 8141 6121 se
rect 8141 6090 8184 6121
tri 8184 6090 8215 6121 nw
tri 7491 6069 7512 6090 ne
rect 7512 6069 8163 6090
tri 8163 6069 8184 6090 nw
rect 12225 6069 12231 6121
rect 12283 6069 12298 6121
rect 12350 6069 12365 6121
rect 12417 6069 12432 6121
rect 12484 6069 12499 6121
rect 12551 6069 12566 6121
rect 12618 6069 12633 6121
rect 12685 6069 12700 6121
rect 12752 6069 12767 6121
rect 12819 6069 12825 6121
rect 5940 6051 6540 6069
rect 5940 6047 5949 6051
rect 6005 6047 6037 6051
rect 6093 6047 6125 6051
rect 6181 6047 6213 6051
rect 6269 6047 6301 6051
rect 6357 6047 6388 6051
rect 6444 6047 6475 6051
rect 6531 6047 6540 6051
tri 7512 6047 7534 6069 ne
rect 7534 6047 8141 6069
tri 8141 6047 8163 6069 nw
rect 12225 6051 12825 6069
rect 12225 6047 12234 6051
rect 12290 6047 12322 6051
rect 12378 6047 12410 6051
rect 12466 6047 12498 6051
rect 12554 6047 12586 6051
rect 12642 6047 12673 6051
rect 12729 6047 12760 6051
rect 12816 6047 12825 6051
rect 5940 5995 5946 6047
rect 6005 5995 6013 6047
rect 6199 5995 6213 6047
rect 6269 5995 6281 6047
rect 6467 5995 6475 6047
rect 6534 5995 6540 6047
tri 7534 6038 7543 6047 ne
rect 7543 6038 8132 6047
tri 8132 6038 8141 6047 nw
rect 12225 5995 12231 6047
rect 12290 5995 12298 6047
rect 12484 5995 12498 6047
rect 12554 5995 12566 6047
rect 12752 5995 12760 6047
rect 12819 5995 12825 6047
rect 16057 6121 16657 6139
rect 16057 6069 16076 6121
rect 16128 6069 16142 6121
rect 16194 6069 16208 6121
rect 16260 6069 16274 6121
rect 16326 6069 16339 6121
rect 16391 6069 16404 6121
rect 16456 6069 16469 6121
rect 16521 6069 16534 6121
rect 16586 6069 16599 6121
rect 16651 6069 16657 6121
rect 16057 6051 16657 6069
rect 16057 6047 16079 6051
rect 16135 6047 16165 6051
rect 16221 6047 16251 6051
rect 16307 6047 16337 6051
rect 16393 6047 16422 6051
rect 16478 6047 16507 6051
rect 16563 6047 16592 6051
rect 16648 6047 16657 6051
rect 16057 5995 16076 6047
rect 16135 5995 16142 6047
rect 16326 5995 16337 6047
rect 16393 5995 16404 6047
rect 16586 5995 16592 6047
rect 16651 5995 16657 6047
rect 20292 6195 20892 6196
rect 20292 6143 20298 6195
rect 20357 6143 20365 6195
rect 20551 6143 20565 6195
rect 20621 6143 20633 6195
rect 20819 6143 20827 6195
rect 20886 6143 20892 6195
tri 23981 6191 23986 6196 ne
rect 23986 6178 24042 6187
rect 20292 6139 20301 6143
rect 20357 6139 20389 6143
rect 20445 6139 20477 6143
rect 20533 6139 20565 6143
rect 20621 6139 20653 6143
rect 20709 6139 20740 6143
rect 20796 6139 20827 6143
rect 20883 6139 20892 6143
rect 20292 6121 20892 6139
rect 20292 6069 20298 6121
rect 20350 6069 20365 6121
rect 20417 6069 20432 6121
rect 20484 6069 20499 6121
rect 20551 6069 20566 6121
rect 20618 6069 20633 6121
rect 20685 6069 20700 6121
rect 20752 6069 20767 6121
rect 20819 6069 20834 6121
rect 20886 6069 20892 6121
rect 20292 6051 20892 6069
rect 20292 6047 20301 6051
rect 20357 6047 20389 6051
rect 20445 6047 20477 6051
rect 20533 6047 20565 6051
rect 20621 6047 20653 6051
rect 20709 6047 20740 6051
rect 20796 6047 20827 6051
rect 20883 6047 20892 6051
rect 20292 5995 20298 6047
rect 20357 5995 20365 6047
rect 20551 5995 20565 6047
rect 20621 5995 20633 6047
rect 20819 5995 20827 6047
rect 20886 5995 20892 6047
tri 16062 5853 16204 5995 nw
rect 4040 5658 4092 5664
rect 4040 5594 4092 5606
tri 2806 4197 2820 4211 sw
rect 2806 4145 2826 4197
rect 2878 4145 2892 4197
rect 2944 4145 2957 4197
rect 3009 4145 3022 4197
rect 3074 4145 3087 4197
rect 3139 4145 3152 4197
rect 3204 4145 3210 4197
rect 964 3445 1016 4115
rect 1427 3926 1483 3935
rect 1427 3846 1483 3870
rect 1427 3781 1483 3790
rect 2595 3840 3210 4145
rect 2595 3788 2826 3840
rect 2878 3788 2892 3840
rect 2944 3788 2957 3840
rect 3009 3788 3022 3840
rect 3074 3788 3087 3840
rect 3139 3788 3152 3840
rect 3204 3788 3210 3840
rect 4040 3840 4092 5542
rect 7436 5497 8036 5498
rect 7436 5496 7445 5497
rect 7501 5496 7533 5497
rect 7589 5496 7621 5497
rect 7677 5496 7709 5497
rect 7765 5496 7797 5497
rect 7853 5496 7884 5497
rect 7940 5496 7971 5497
rect 8027 5496 8036 5497
rect 7436 5444 7442 5496
rect 7501 5444 7509 5496
rect 7695 5444 7709 5496
rect 7765 5444 7777 5496
rect 7963 5444 7971 5496
rect 8030 5444 8036 5496
rect 7436 5441 7445 5444
rect 7501 5441 7533 5444
rect 7589 5441 7621 5444
rect 7677 5441 7709 5444
rect 7765 5441 7797 5444
rect 7853 5441 7884 5444
rect 7940 5441 7971 5444
rect 8027 5441 8036 5444
rect 7436 5424 8036 5441
rect 7436 5372 7442 5424
rect 7494 5372 7509 5424
rect 7561 5372 7576 5424
rect 7628 5372 7643 5424
rect 7695 5372 7710 5424
rect 7762 5372 7777 5424
rect 7829 5372 7844 5424
rect 7896 5372 7911 5424
rect 7963 5372 7978 5424
rect 8030 5372 8036 5424
rect 7436 5355 8036 5372
rect 7436 5352 7445 5355
rect 7501 5352 7533 5355
rect 7589 5352 7621 5355
rect 7677 5352 7709 5355
rect 7765 5352 7797 5355
rect 7853 5352 7884 5355
rect 7940 5352 7971 5355
rect 8027 5352 8036 5355
rect 7436 5300 7442 5352
rect 7501 5300 7509 5352
rect 7695 5300 7709 5352
rect 7765 5300 7777 5352
rect 7963 5300 7971 5352
rect 8030 5300 8036 5352
rect 7436 5299 7445 5300
rect 7501 5299 7533 5300
rect 7589 5299 7621 5300
rect 7677 5299 7709 5300
rect 7765 5299 7797 5300
rect 7853 5299 7884 5300
rect 7940 5299 7971 5300
rect 8027 5299 8036 5300
rect 11505 5497 12105 5498
rect 11505 5496 11514 5497
rect 11570 5496 11602 5497
rect 11658 5496 11690 5497
rect 11746 5496 11778 5497
rect 11834 5496 11866 5497
rect 11922 5496 11953 5497
rect 12009 5496 12040 5497
rect 12096 5496 12105 5497
rect 11505 5444 11511 5496
rect 11570 5444 11578 5496
rect 11764 5444 11778 5496
rect 11834 5444 11846 5496
rect 12032 5444 12040 5496
rect 12099 5444 12105 5496
rect 11505 5441 11514 5444
rect 11570 5441 11602 5444
rect 11658 5441 11690 5444
rect 11746 5441 11778 5444
rect 11834 5441 11866 5444
rect 11922 5441 11953 5444
rect 12009 5441 12040 5444
rect 12096 5441 12105 5444
rect 11505 5424 12105 5441
rect 11505 5372 11511 5424
rect 11563 5372 11578 5424
rect 11630 5372 11645 5424
rect 11697 5372 11712 5424
rect 11764 5372 11779 5424
rect 11831 5372 11846 5424
rect 11898 5372 11913 5424
rect 11965 5372 11980 5424
rect 12032 5372 12047 5424
rect 12099 5372 12105 5424
rect 11505 5355 12105 5372
rect 11505 5352 11514 5355
rect 11570 5352 11602 5355
rect 11658 5352 11690 5355
rect 11746 5352 11778 5355
rect 11834 5352 11866 5355
rect 11922 5352 11953 5355
rect 12009 5352 12040 5355
rect 12096 5352 12105 5355
rect 11505 5300 11511 5352
rect 11570 5300 11578 5352
rect 11764 5300 11778 5352
rect 11834 5300 11846 5352
rect 12032 5300 12040 5352
rect 12099 5300 12105 5352
rect 11505 5299 11514 5300
rect 11570 5299 11602 5300
rect 11658 5299 11690 5300
rect 11746 5299 11778 5300
rect 11834 5299 11866 5300
rect 11922 5299 11953 5300
rect 12009 5299 12040 5300
rect 12096 5299 12105 5300
rect 14527 5497 15006 5498
rect 14527 5496 14536 5497
rect 14592 5496 14617 5497
rect 14673 5496 14698 5497
rect 14754 5496 14779 5497
rect 14835 5496 14860 5497
rect 14916 5496 14941 5497
rect 14997 5496 15006 5497
rect 14527 5444 14533 5496
rect 14592 5444 14603 5496
rect 14931 5444 14941 5496
rect 15000 5444 15006 5496
rect 14527 5441 14536 5444
rect 14592 5441 14617 5444
rect 14673 5441 14698 5444
rect 14754 5441 14779 5444
rect 14835 5441 14860 5444
rect 14916 5441 14941 5444
rect 14997 5441 15006 5444
rect 14527 5424 15006 5441
rect 14527 5372 14533 5424
rect 14585 5372 14603 5424
rect 14655 5372 14672 5424
rect 14724 5372 14741 5424
rect 14793 5372 14810 5424
rect 14862 5372 14879 5424
rect 14931 5372 14948 5424
rect 15000 5372 15006 5424
rect 14527 5355 15006 5372
rect 14527 5352 14536 5355
rect 14592 5352 14617 5355
rect 14673 5352 14698 5355
rect 14754 5352 14779 5355
rect 14835 5352 14860 5355
rect 14916 5352 14941 5355
rect 14997 5352 15006 5355
rect 14527 5300 14533 5352
rect 14592 5300 14603 5352
rect 14931 5300 14941 5352
rect 15000 5300 15006 5352
rect 14527 5299 14536 5300
rect 14592 5299 14617 5300
rect 14673 5299 14698 5300
rect 14754 5299 14779 5300
rect 14835 5299 14860 5300
rect 14916 5299 14941 5300
rect 14997 5299 15006 5300
rect 16890 4544 16899 4600
rect 16955 4544 17012 4600
rect 17068 4544 17125 4600
rect 17181 4544 17190 4600
rect 16890 4520 17190 4544
rect 16890 4485 16899 4520
rect 16955 4485 17012 4520
rect 17068 4485 17125 4520
rect 17181 4485 17190 4520
rect 16890 4433 16896 4485
rect 16955 4464 16975 4485
rect 17105 4464 17125 4485
rect 16948 4440 16975 4464
rect 17027 4440 17053 4464
rect 17105 4440 17131 4464
rect 16955 4433 16975 4440
rect 17105 4433 17125 4440
rect 17183 4433 17190 4485
rect 16890 4384 16899 4433
rect 16955 4384 17012 4433
rect 17068 4384 17125 4433
rect 17181 4384 17190 4433
rect 16890 4361 17190 4384
tri 5528 4341 5532 4345 sw
rect 5476 4332 5532 4341
rect 5476 4252 5532 4276
tri 9076 4341 9080 4345 se
tri 9298 4341 9302 4345 sw
rect 9076 4332 9132 4341
rect 9076 4252 9132 4276
rect 5476 4187 5532 4196
tri 5528 4183 5532 4187 nw
rect 7545 4187 7590 4226
tri 7590 4187 7629 4226 sw
rect 9076 4187 9132 4196
rect 9246 4332 9302 4341
rect 9246 4252 9302 4276
rect 9246 4187 9302 4196
tri 13222 4341 13226 4345 se
tri 13444 4341 13448 4345 sw
rect 13222 4332 13278 4341
rect 13222 4252 13278 4276
rect 13222 4187 13278 4196
rect 13392 4332 13448 4341
rect 13392 4252 13448 4276
rect 16890 4309 16896 4361
rect 16948 4360 16975 4361
rect 17027 4360 17053 4361
rect 17105 4360 17131 4361
rect 16955 4309 16975 4360
rect 17105 4309 17125 4360
rect 17183 4309 17190 4361
rect 16890 4304 16899 4309
rect 16955 4304 17012 4309
rect 17068 4304 17125 4309
rect 17181 4304 17190 4309
rect 16890 4280 17190 4304
rect 16890 4224 16899 4280
rect 16955 4224 17012 4280
rect 17068 4224 17125 4280
rect 17181 4224 17190 4280
tri 17368 4341 17372 4345 se
tri 17590 4341 17594 4345 sw
rect 17368 4332 17424 4341
rect 17368 4252 17424 4276
rect 13392 4187 13448 4196
rect 17368 4187 17424 4196
rect 17538 4332 17594 4341
rect 17538 4252 17594 4276
rect 17538 4187 17594 4196
tri 21516 4341 21520 4345 se
tri 25716 4341 25720 4345 sw
rect 21516 4332 21572 4341
rect 21516 4252 21572 4276
rect 21516 4187 21572 4196
rect 21680 4332 21736 4341
rect 21680 4252 21736 4276
rect 25664 4332 25720 4341
rect 25664 4252 25720 4276
rect 21680 4187 21736 4196
rect 25285 4201 25341 4210
rect 7545 4186 7629 4187
tri 7545 4183 7548 4186 ne
rect 7548 4183 7629 4186
tri 7548 4148 7583 4183 ne
rect 7583 4148 7629 4183
tri 7629 4148 7668 4187 sw
tri 7583 4141 7590 4148 ne
rect 7590 4141 7668 4148
tri 7590 4063 7668 4141 ne
tri 7668 4063 7753 4148 sw
tri 7668 4030 7701 4063 ne
tri 4092 3840 4145 3893 sw
rect 4040 3788 4046 3840
rect 4098 3788 4110 3840
rect 4162 3788 4168 3840
rect 2595 3781 2813 3788
tri 2813 3781 2820 3788 nw
rect 2595 3762 2794 3781
tri 2794 3762 2813 3781 nw
rect 2595 3760 2792 3762
tri 2792 3760 2794 3762 nw
rect 2595 3756 2757 3760
rect 2647 3704 2705 3756
tri 2757 3725 2792 3760 nw
rect 7701 3708 7753 4063
tri 7753 3708 7760 3715 sw
rect 2595 3679 2757 3704
tri 3201 3680 3228 3707 se
rect 3228 3680 7313 3707
tri 7313 3680 7340 3707 sw
rect 7701 3680 7760 3708
tri 7760 3680 7788 3708 sw
rect 2647 3627 2705 3679
tri 3173 3652 3201 3680 se
rect 3201 3655 7340 3680
rect 3201 3652 3247 3655
tri 3247 3652 3250 3655 nw
tri 7292 3652 7295 3655 ne
rect 7295 3652 7340 3655
tri 7340 3652 7368 3680 sw
tri 3154 3633 3173 3652 se
rect 3173 3633 3228 3652
tri 3228 3633 3247 3652 nw
tri 7295 3634 7313 3652 ne
rect 7313 3634 7368 3652
tri 7313 3633 7314 3634 ne
rect 7314 3633 7368 3634
tri 3149 3628 3154 3633 se
rect 3154 3628 3223 3633
tri 3223 3628 3228 3633 nw
tri 7314 3628 7319 3633 ne
rect 7319 3628 7368 3633
tri 7368 3628 7392 3652 sw
rect 7701 3628 7707 3680
rect 7759 3628 7771 3680
rect 7823 3628 7829 3680
tri 10478 3628 10485 3635 se
rect 10485 3628 10537 4187
rect 2595 3602 2757 3627
tri 3136 3615 3149 3628 se
rect 3149 3615 3210 3628
tri 3210 3615 3223 3628 nw
tri 7319 3615 7332 3628 ne
rect 7332 3615 7392 3628
tri 7392 3615 7405 3628 sw
tri 10465 3615 10478 3628 se
rect 10478 3615 10537 3628
rect 2647 3550 2705 3602
tri 3121 3600 3136 3615 se
rect 3136 3600 3195 3615
tri 3195 3600 3210 3615 nw
tri 3277 3600 3292 3615 se
rect 3292 3600 7221 3615
tri 7221 3600 7236 3615 sw
tri 7332 3600 7347 3615 ne
rect 7347 3600 7405 3615
tri 7405 3600 7420 3615 sw
tri 10450 3600 10465 3615 se
rect 10465 3600 10537 3615
tri 3081 3560 3121 3600 se
rect 3121 3560 3155 3600
tri 3155 3560 3195 3600 nw
tri 3237 3560 3277 3600 se
rect 3277 3563 7236 3600
rect 3277 3560 3311 3563
tri 3311 3560 3314 3563 nw
tri 7200 3560 7203 3563 ne
rect 7203 3560 7236 3563
tri 7236 3560 7276 3600 sw
tri 7347 3579 7368 3600 ne
rect 7368 3579 7420 3600
tri 7420 3579 7441 3600 sw
tri 7368 3560 7387 3579 ne
rect 7387 3560 8198 3579
tri 3080 3559 3081 3560 se
rect 3081 3559 3154 3560
tri 3154 3559 3155 3560 nw
tri 3236 3559 3237 3560 se
rect 3237 3559 3299 3560
rect 2595 3544 2757 3550
tri 3069 3548 3080 3559 se
rect 3080 3548 3143 3559
tri 3143 3548 3154 3559 nw
tri 3225 3548 3236 3559 se
rect 3236 3548 3299 3559
tri 3299 3548 3311 3560 nw
tri 7203 3548 7215 3560 ne
rect 7215 3548 7276 3560
tri 7276 3548 7288 3560 sw
tri 7387 3548 7399 3560 ne
rect 7399 3548 8198 3560
rect 10409 3548 10415 3600
rect 10467 3548 10479 3600
rect 10531 3548 10537 3600
tri 3065 3544 3069 3548 se
rect 3069 3544 3136 3548
tri 3062 3541 3065 3544 se
rect 3065 3541 3136 3544
tri 3136 3541 3143 3548 nw
tri 3218 3541 3225 3548 se
rect 3225 3541 3292 3548
tri 3292 3541 3299 3548 nw
tri 7215 3542 7221 3548 ne
rect 7221 3542 7288 3548
tri 7221 3541 7222 3542 ne
rect 7222 3541 7288 3542
tri 3053 3532 3062 3541 se
rect 3062 3532 3127 3541
tri 3127 3532 3136 3541 nw
tri 3209 3532 3218 3541 se
rect 3218 3532 3283 3541
tri 3283 3532 3292 3541 nw
tri 7222 3532 7231 3541 ne
rect 7231 3532 7288 3541
tri 7288 3532 7304 3548 sw
tri 7399 3532 7415 3548 ne
rect 7415 3532 8198 3548
tri 3041 3520 3053 3532 se
rect 3053 3520 3115 3532
tri 3115 3520 3127 3532 nw
tri 3197 3520 3209 3532 se
rect 3209 3520 3271 3532
tri 3271 3520 3283 3532 nw
tri 7231 3520 7243 3532 ne
rect 7243 3520 7304 3532
tri 7304 3520 7316 3532 sw
tri 7415 3527 7420 3532 ne
rect 7420 3527 8198 3532
tri 8029 3520 8036 3527 ne
rect 8036 3520 8198 3527
tri 3024 3503 3041 3520 se
rect 3041 3503 3098 3520
tri 3098 3503 3115 3520 nw
tri 3180 3503 3197 3520 se
rect 3197 3503 3254 3520
tri 3254 3503 3271 3520 nw
tri 7243 3503 7260 3520 ne
rect 7260 3503 7316 3520
tri 7316 3503 7333 3520 sw
tri 8036 3503 8053 3520 ne
rect 8053 3503 8198 3520
tri 3018 3497 3024 3503 se
rect 3024 3497 3092 3503
tri 3092 3497 3098 3503 nw
tri 3174 3497 3180 3503 se
rect 3180 3497 3248 3503
tri 3248 3497 3254 3503 nw
rect 3342 3497 3714 3503
tri 3006 3485 3018 3497 se
rect 3018 3485 3080 3497
tri 3080 3485 3092 3497 nw
tri 3162 3485 3174 3497 se
rect 3174 3485 3218 3497
tri 2988 3467 3006 3485 se
rect 3006 3467 3062 3485
tri 3062 3467 3080 3485 nw
tri 3144 3467 3162 3485 se
rect 3162 3467 3218 3485
tri 3218 3467 3248 3497 nw
rect 3342 3494 3351 3497
rect 3403 3494 3415 3497
rect 3467 3494 3479 3497
rect 3531 3494 3543 3497
rect 3595 3494 3714 3497
tri 2982 3461 2988 3467 se
rect 2988 3461 3040 3467
tri 1016 3445 1032 3461 sw
tri 2966 3445 2982 3461 se
rect 2982 3445 3040 3461
tri 3040 3445 3062 3467 nw
tri 3122 3445 3144 3467 se
rect 3144 3445 3196 3467
tri 3196 3445 3218 3467 nw
rect 964 3440 1032 3445
tri 1032 3440 1037 3445 sw
tri 2961 3440 2966 3445 se
rect 2966 3440 3035 3445
tri 3035 3440 3040 3445 nw
tri 3117 3440 3122 3445 se
rect 3122 3440 3191 3445
tri 3191 3440 3196 3445 nw
rect 964 3432 1037 3440
tri 1037 3432 1045 3440 sw
tri 2953 3432 2961 3440 se
rect 2961 3432 3027 3440
tri 3027 3432 3035 3440 nw
tri 3109 3432 3117 3440 se
rect 3117 3432 3183 3440
tri 3183 3432 3191 3440 nw
rect 964 3411 1045 3432
tri 1045 3411 1066 3432 sw
tri 2932 3411 2953 3432 se
rect 2953 3411 3006 3432
tri 3006 3411 3027 3432 nw
tri 3088 3411 3109 3432 se
rect 3109 3411 3144 3432
rect 964 3410 1066 3411
tri 1066 3410 1067 3411 sw
tri 2931 3410 2932 3411 se
rect 2932 3410 3005 3411
tri 3005 3410 3006 3411 nw
tri 3087 3410 3088 3411 se
rect 3088 3410 3144 3411
rect 904 3358 910 3410
rect 962 3358 974 3410
rect 1026 3409 1067 3410
tri 1067 3409 1068 3410 sw
tri 2930 3409 2931 3410 se
rect 2931 3409 2988 3410
rect 1026 3358 1032 3409
tri 2914 3393 2930 3409 se
rect 2930 3393 2988 3409
tri 2988 3393 3005 3410 nw
tri 3070 3393 3087 3410 se
rect 3087 3393 3144 3410
tri 3144 3393 3183 3432 nw
tri 2901 3380 2914 3393 se
rect 2914 3380 2975 3393
tri 2975 3380 2988 3393 nw
tri 3057 3380 3070 3393 se
rect 3070 3380 3131 3393
tri 3131 3380 3144 3393 nw
tri 2888 3367 2901 3380 se
rect 2901 3367 2962 3380
tri 2962 3367 2975 3380 nw
tri 3044 3367 3057 3380 se
rect 3057 3367 3118 3380
tri 3118 3367 3131 3380 nw
tri 2879 3358 2888 3367 se
rect 2888 3358 2953 3367
tri 2953 3358 2962 3367 nw
tri 3035 3358 3044 3367 se
rect 3044 3358 3070 3367
tri 2874 3353 2879 3358 se
rect 2879 3353 2948 3358
tri 2948 3353 2953 3358 nw
tri 3030 3353 3035 3358 se
rect 3035 3353 3070 3358
rect 701 3344 757 3353
tri 2858 3337 2874 3353 se
rect 2874 3337 2932 3353
tri 2932 3337 2948 3353 nw
tri 3014 3337 3030 3353 se
rect 3030 3337 3070 3353
tri 2840 3319 2858 3337 se
rect 2858 3319 2914 3337
tri 2914 3319 2932 3337 nw
tri 2996 3319 3014 3337 se
rect 3014 3319 3070 3337
tri 3070 3319 3118 3367 nw
tri 2836 3315 2840 3319 se
rect 2840 3315 2910 3319
tri 2910 3315 2914 3319 nw
tri 2992 3315 2996 3319 se
rect 2996 3315 3066 3319
tri 3066 3315 3070 3319 nw
tri 2829 3308 2836 3315 se
rect 2836 3308 2903 3315
tri 2903 3308 2910 3315 nw
tri 2985 3308 2992 3315 se
rect 2992 3308 3059 3315
tri 3059 3308 3066 3315 nw
tri 2823 3302 2829 3308 se
rect 2829 3302 2897 3308
tri 2897 3302 2903 3308 nw
tri 2979 3302 2985 3308 se
rect 2985 3302 3053 3308
tri 3053 3302 3059 3308 nw
rect 701 3270 703 3288
rect 755 3270 757 3288
rect 701 3264 757 3270
tri 2784 3263 2823 3302 se
rect 2823 3263 2858 3302
tri 2858 3263 2897 3302 nw
tri 2940 3263 2979 3302 se
rect 2979 3263 3001 3302
tri 2771 3250 2784 3263 se
rect 2784 3250 2845 3263
tri 2845 3250 2858 3263 nw
tri 2927 3250 2940 3263 se
rect 2940 3250 3001 3263
tri 3001 3250 3053 3302 nw
tri 2766 3245 2771 3250 se
rect 2771 3245 2840 3250
tri 2840 3245 2845 3250 nw
tri 2922 3245 2927 3250 se
rect 2927 3245 2996 3250
tri 2996 3245 3001 3250 nw
tri 2758 3237 2766 3245 se
rect 2766 3237 2832 3245
tri 2832 3237 2840 3245 nw
tri 2914 3237 2922 3245 se
rect 2922 3237 2988 3245
tri 2988 3237 2996 3245 nw
rect 701 3206 703 3208
rect 755 3206 757 3208
rect 701 3199 757 3206
tri 2720 3199 2758 3237 se
rect 2758 3199 2794 3237
tri 2794 3199 2832 3237 nw
tri 2876 3199 2914 3237 se
rect 2914 3199 2936 3237
tri 2710 3189 2720 3199 se
rect 2720 3189 2784 3199
tri 2784 3189 2794 3199 nw
tri 2866 3189 2876 3199 se
rect 2876 3189 2936 3199
tri 2706 3185 2710 3189 se
rect 2710 3185 2780 3189
tri 2780 3185 2784 3189 nw
tri 2862 3185 2866 3189 se
rect 2866 3185 2936 3189
tri 2936 3185 2988 3237 nw
rect 3342 3198 3347 3494
rect 3643 3198 3714 3494
tri 7260 3487 7276 3503 ne
rect 7276 3487 7333 3503
tri 7333 3487 7349 3503 sw
tri 8053 3487 8069 3503 ne
rect 8069 3487 8198 3503
tri 7276 3468 7295 3487 ne
rect 7295 3468 7798 3487
tri 8069 3486 8070 3487 ne
tri 7295 3452 7311 3468 ne
rect 7311 3452 7798 3468
tri 7311 3440 7323 3452 ne
rect 7323 3440 7798 3452
tri 7323 3435 7328 3440 ne
rect 7328 3435 7798 3440
tri 7629 3394 7670 3435 ne
rect 7670 3393 7798 3435
rect 7670 3341 7676 3393
rect 7728 3341 7740 3393
rect 7792 3341 7798 3393
rect 8070 3440 8198 3487
tri 10774 3468 10781 3475 se
rect 10781 3468 10833 4187
rect 11192 3468 11198 3520
rect 11250 3468 11262 3520
rect 11314 3468 11320 3520
tri 10758 3452 10774 3468 se
rect 10774 3452 10833 3468
tri 11678 3452 11691 3465 se
rect 11691 3452 11743 4187
tri 11982 3550 11987 3555 se
rect 11987 3550 12039 4187
tri 11964 3532 11982 3550 se
rect 11982 3532 12039 3550
tri 11952 3520 11964 3532 se
rect 11964 3520 12039 3532
rect 11911 3468 11917 3520
rect 11969 3468 11981 3520
rect 12033 3468 12039 3520
rect 14927 3550 14979 4187
tri 14979 3550 14996 3567 sw
rect 14927 3532 14996 3550
tri 14996 3532 15014 3550 sw
rect 14927 3480 14933 3532
rect 14985 3480 14997 3532
rect 15049 3480 15055 3532
rect 15837 3468 15889 4187
tri 19069 3550 19073 3554 se
rect 19073 3550 19125 4187
tri 17022 3498 17074 3550 se
rect 17074 3498 17080 3550
rect 17132 3498 17147 3550
rect 17199 3498 17214 3550
rect 17266 3498 17281 3550
rect 17333 3498 17348 3550
rect 17400 3498 17415 3550
rect 17467 3498 17482 3550
rect 17534 3498 17549 3550
rect 17601 3498 17616 3550
rect 17668 3498 17682 3550
rect 17734 3498 17748 3550
rect 17800 3498 17814 3550
rect 17866 3498 17880 3550
rect 17932 3498 17946 3550
rect 17998 3498 18012 3550
rect 18064 3498 18078 3550
rect 18130 3498 18144 3550
rect 18196 3498 18210 3550
rect 18262 3498 18276 3550
rect 18328 3498 18342 3550
rect 18394 3498 18408 3550
rect 18460 3498 18474 3550
rect 18526 3498 18540 3550
rect 18592 3498 18606 3550
rect 18658 3498 18672 3550
rect 18724 3498 18730 3550
tri 19067 3548 19069 3550 se
rect 19069 3548 19125 3550
rect 20279 3628 20331 4187
rect 22546 3708 22552 3760
rect 22604 3708 22616 3760
rect 22668 3708 22674 3760
tri 22554 3680 22582 3708 ne
rect 22582 3680 22640 3708
tri 20331 3628 20337 3634 sw
rect 20908 3628 20914 3680
rect 20966 3628 20978 3680
rect 21030 3628 21036 3680
tri 22582 3674 22588 3680 ne
rect 20279 3600 20337 3628
tri 20337 3600 20365 3628 sw
tri 20908 3612 20924 3628 ne
rect 20924 3600 20992 3628
tri 20992 3600 21020 3628 nw
rect 20279 3548 20285 3600
rect 20337 3548 20349 3600
rect 20401 3548 20407 3600
tri 19039 3520 19067 3548 se
rect 19067 3520 19125 3548
tri 17011 3487 17022 3498 se
rect 17022 3487 18730 3498
tri 15889 3468 15908 3487 sw
tri 16992 3468 17011 3487 se
rect 17011 3468 18730 3487
rect 18997 3468 19003 3520
rect 19055 3468 19067 3520
rect 19119 3468 19125 3520
tri 10746 3440 10758 3452 se
rect 10758 3440 10833 3452
rect 8070 3388 8076 3440
rect 8128 3388 8140 3440
rect 8192 3388 8198 3440
rect 10705 3388 10711 3440
rect 10763 3388 10775 3440
rect 10827 3388 10833 3440
tri 11656 3430 11678 3452 se
rect 11678 3430 11743 3452
rect 11615 3378 11621 3430
rect 11673 3378 11685 3430
rect 11737 3378 11743 3430
rect 15837 3452 15908 3468
tri 15908 3452 15924 3468 sw
tri 16976 3452 16992 3468 se
rect 16992 3452 18730 3468
rect 15837 3400 15843 3452
rect 15895 3400 15907 3452
rect 15959 3400 15965 3452
tri 16964 3440 16976 3452 se
rect 16976 3440 18730 3452
tri 16924 3400 16964 3440 se
rect 16964 3400 18730 3440
tri 16912 3388 16924 3400 se
rect 16924 3388 18730 3400
tri 16902 3378 16912 3388 se
rect 16912 3378 18730 3388
tri 16884 3360 16902 3378 se
rect 16902 3360 18730 3378
tri 16865 3341 16884 3360 se
rect 16884 3341 18730 3360
tri 16832 3308 16865 3341 se
rect 16865 3308 18730 3341
rect 20924 3360 20976 3600
tri 20976 3584 20992 3600 nw
rect 22408 3548 22414 3600
rect 22466 3548 22478 3600
rect 22530 3548 22536 3600
tri 22450 3520 22478 3548 ne
rect 22478 3520 22536 3548
rect 22304 3468 22310 3520
rect 22362 3468 22374 3520
rect 22426 3468 22432 3520
tri 22478 3514 22484 3520 ne
tri 22346 3440 22374 3468 ne
rect 22374 3440 22432 3468
rect 22198 3388 22204 3440
rect 22256 3388 22268 3440
rect 22320 3428 22326 3440
tri 22326 3428 22338 3440 sw
tri 22374 3434 22380 3440 ne
rect 22320 3388 22338 3428
tri 22252 3378 22262 3388 ne
rect 22262 3378 22338 3388
tri 22262 3364 22276 3378 ne
rect 22276 3364 22338 3378
tri 20976 3360 20980 3364 sw
tri 22276 3360 22280 3364 ne
rect 22280 3360 22338 3364
rect 20924 3330 20980 3360
tri 20924 3308 20946 3330 ne
rect 20946 3308 20980 3330
tri 20980 3308 21032 3360 sw
rect 22090 3308 22096 3360
rect 22148 3308 22160 3360
rect 22212 3308 22218 3360
tri 22280 3354 22286 3360 ne
tri 16808 3284 16832 3308 se
rect 16832 3284 18730 3308
tri 20946 3300 20954 3308 ne
rect 20954 3300 21032 3308
tri 21032 3300 21040 3308 sw
tri 20954 3284 20970 3300 ne
rect 20970 3284 21040 3300
tri 22132 3284 22156 3308 ne
rect 22156 3284 22218 3308
rect 3342 3185 3351 3198
rect 3403 3185 3415 3198
rect 3467 3185 3479 3198
rect 3531 3185 3543 3198
rect 3595 3185 3714 3198
tri 2693 3172 2706 3185 se
rect 2706 3172 2767 3185
tri 2767 3172 2780 3185 nw
tri 2849 3172 2862 3185 se
rect 2862 3172 2923 3185
tri 2923 3172 2936 3185 nw
rect 3342 3173 3714 3185
tri 2692 3171 2693 3172 se
rect 2693 3171 2766 3172
tri 2766 3171 2767 3172 nw
tri 2848 3171 2849 3172 se
rect 2849 3171 2922 3172
tri 2922 3171 2923 3172 nw
rect 1758 3162 1814 3171
rect 1163 3139 1219 3148
rect 1163 3059 1219 3083
tri 2669 3148 2692 3171 se
rect 2692 3148 2743 3171
tri 2743 3148 2766 3171 nw
tri 2825 3148 2848 3171 se
rect 2848 3148 2871 3171
tri 2641 3120 2669 3148 se
rect 2669 3120 2715 3148
tri 2715 3120 2743 3148 nw
tri 2797 3120 2825 3148 se
rect 2825 3120 2871 3148
tri 2871 3120 2922 3171 nw
tri 2636 3115 2641 3120 se
rect 2641 3115 2710 3120
tri 2710 3115 2715 3120 nw
tri 2792 3115 2797 3120 se
rect 2797 3115 2857 3120
tri 2627 3106 2636 3115 se
rect 2636 3106 2701 3115
tri 2701 3106 2710 3115 nw
tri 2783 3106 2792 3115 se
rect 2792 3106 2857 3115
tri 2857 3106 2871 3120 nw
rect 3342 3117 3347 3173
rect 3403 3172 3427 3173
rect 3483 3172 3507 3173
rect 3563 3172 3587 3173
rect 3403 3120 3415 3172
rect 3403 3117 3427 3120
rect 3483 3117 3507 3120
rect 3563 3117 3587 3120
rect 3643 3117 3714 3173
rect 3342 3106 3714 3117
rect 1758 3088 1760 3106
rect 1812 3088 1814 3106
tri 2618 3097 2627 3106 se
rect 2627 3097 2692 3106
tri 2692 3097 2701 3106 nw
tri 2774 3097 2783 3106 se
rect 2783 3097 2848 3106
tri 2848 3097 2857 3106 nw
tri 2611 3090 2618 3097 se
rect 2618 3090 2685 3097
tri 2685 3090 2692 3097 nw
tri 2767 3090 2774 3097 se
rect 2774 3090 2805 3097
rect 1758 3082 1814 3088
rect 1758 3024 1760 3026
rect 1812 3024 1814 3026
rect 1758 3017 1814 3024
rect 2547 3084 2649 3090
rect 2599 3054 2649 3084
tri 2649 3054 2685 3090 nw
tri 2731 3054 2767 3090 se
rect 2767 3054 2805 3090
tri 2805 3054 2848 3097 nw
rect 3342 3092 3351 3106
rect 2599 3040 2635 3054
tri 2635 3040 2649 3054 nw
tri 2717 3040 2731 3054 se
rect 2731 3040 2791 3054
tri 2791 3040 2805 3054 nw
rect 2599 3032 2618 3040
rect 2547 3023 2618 3032
tri 2618 3023 2635 3040 nw
tri 2700 3023 2717 3040 se
rect 2717 3023 2774 3040
tri 2774 3023 2791 3040 nw
rect 3342 3036 3347 3092
rect 3403 3054 3415 3106
rect 3467 3092 3479 3106
rect 3531 3092 3543 3106
rect 3595 3092 3714 3106
rect 3403 3040 3427 3054
rect 3483 3040 3507 3054
rect 3563 3040 3587 3054
rect 2547 3020 2603 3023
rect 1163 2992 1219 3003
rect 1163 2940 1165 2992
rect 1217 2940 1219 2992
rect 2599 3008 2603 3020
tri 2603 3008 2618 3023 nw
tri 2685 3008 2700 3023 se
rect 2700 3008 2739 3023
tri 2599 3004 2603 3008 nw
tri 2681 3004 2685 3008 se
rect 2685 3004 2739 3008
tri 2677 3000 2681 3004 se
rect 2681 3000 2739 3004
tri 2665 2988 2677 3000 se
rect 2677 2988 2739 3000
tri 2739 2988 2774 3023 nw
rect 3342 3011 3351 3036
tri 2651 2974 2665 2988 se
rect 2665 2974 2725 2988
tri 2725 2974 2739 2988 nw
rect 2547 2962 2599 2968
tri 2639 2962 2651 2974 se
rect 2651 2962 2700 2974
tri 2626 2949 2639 2962 se
rect 2639 2949 2700 2962
tri 2700 2949 2725 2974 nw
rect 3342 2955 3347 3011
rect 3403 2988 3415 3040
rect 3643 3036 3714 3092
rect 7436 3228 7445 3284
rect 7501 3228 7533 3284
rect 7589 3228 7621 3284
rect 7677 3228 7709 3284
rect 7765 3228 7797 3284
rect 7853 3228 7884 3284
rect 7940 3228 7971 3284
rect 8027 3228 8036 3284
rect 7436 3144 8036 3228
rect 7436 3088 7445 3144
rect 7501 3088 7533 3144
rect 7589 3088 7621 3144
rect 7677 3088 7709 3144
rect 7765 3088 7797 3144
rect 7853 3088 7884 3144
rect 7940 3088 7971 3144
rect 8027 3088 8036 3144
rect 11505 3228 11514 3284
rect 11570 3228 11602 3284
rect 11658 3228 11690 3284
rect 11746 3228 11778 3284
rect 11834 3228 11866 3284
rect 11922 3228 11953 3284
rect 12009 3228 12040 3284
rect 12096 3228 12105 3284
rect 11505 3144 12105 3228
rect 11505 3088 11514 3144
rect 11570 3088 11602 3144
rect 11658 3088 11690 3144
rect 11746 3088 11778 3144
rect 11834 3088 11866 3144
rect 11922 3088 11953 3144
rect 12009 3088 12040 3144
rect 12096 3088 12105 3144
rect 14527 3228 14536 3284
rect 14592 3228 14624 3284
rect 14680 3228 14712 3284
rect 14768 3228 14800 3284
rect 14856 3228 14888 3284
rect 14944 3228 14975 3284
rect 15031 3228 15062 3284
rect 15118 3228 15127 3284
tri 20970 3279 20975 3284 ne
rect 20975 3280 21040 3284
tri 22156 3280 22160 3284 ne
rect 22160 3280 22218 3284
rect 20975 3279 20988 3280
tri 22160 3279 22161 3280 ne
rect 22161 3279 22218 3280
rect 14527 3144 15127 3228
rect 14527 3088 14536 3144
rect 14592 3088 14624 3144
rect 14680 3088 14712 3144
rect 14768 3088 14800 3144
rect 14856 3088 14888 3144
rect 14944 3088 14975 3144
rect 15031 3088 15062 3144
rect 15118 3088 15127 3144
rect 18260 3223 18269 3279
rect 18325 3223 18368 3279
rect 18424 3223 18466 3279
rect 18522 3223 18531 3279
tri 20975 3278 20976 3279 ne
rect 20976 3278 20988 3279
tri 20976 3274 20980 3278 ne
rect 20980 3274 20988 3278
tri 22161 3274 22166 3279 ne
tri 20980 3266 20988 3274 ne
rect 22166 3265 22218 3279
rect 18260 3149 18531 3223
rect 18260 3093 18269 3149
rect 18325 3093 18368 3149
rect 18424 3093 18466 3149
rect 18522 3093 18531 3149
rect 3467 3011 3479 3036
rect 3531 3011 3543 3036
rect 3595 3011 3714 3036
rect 3403 2974 3427 2988
rect 3483 2974 3507 2988
rect 3563 2974 3587 2988
rect 1163 2934 1219 2940
tri 2611 2934 2626 2949 se
rect 2626 2934 2673 2949
tri 2599 2922 2611 2934 se
rect 2611 2922 2673 2934
tri 2673 2922 2700 2949 nw
rect 3342 2930 3351 2955
tri 2585 2908 2599 2922 se
rect 2599 2908 2659 2922
tri 2659 2908 2673 2922 nw
tri 2572 2895 2585 2908 se
rect 2585 2895 2643 2908
rect 1163 2891 1219 2895
tri 2569 2892 2572 2895 se
rect 2572 2892 2643 2895
tri 2643 2892 2659 2908 nw
rect 2548 2891 2642 2892
tri 2642 2891 2643 2892 nw
rect 1163 2886 1171 2891
rect 1223 2839 1235 2891
rect 1287 2839 1293 2891
rect 2548 2886 2607 2891
rect 1163 2806 1219 2830
rect 2600 2856 2607 2886
tri 2607 2856 2642 2891 nw
rect 3342 2874 3347 2930
rect 3403 2922 3415 2974
rect 3643 2955 3714 3011
rect 3467 2930 3479 2955
rect 3531 2930 3543 2955
rect 3595 2930 3714 2955
rect 3403 2908 3427 2922
rect 3483 2908 3507 2922
rect 3563 2908 3587 2922
rect 3342 2856 3351 2874
rect 3403 2856 3415 2908
rect 3643 2874 3714 2930
rect 3467 2856 3479 2874
rect 3531 2856 3543 2874
rect 3595 2856 3714 2874
tri 2600 2849 2607 2856 nw
rect 3342 2849 3714 2856
rect 2548 2822 2600 2834
rect 3342 2793 3347 2849
rect 3403 2842 3427 2849
rect 3483 2842 3507 2849
rect 3563 2842 3587 2849
rect 3342 2790 3351 2793
rect 3403 2790 3415 2842
rect 3643 2793 3714 2849
rect 3467 2790 3479 2793
rect 3531 2790 3543 2793
rect 3595 2790 3714 2793
rect 3342 2784 3714 2790
rect 4081 3046 4137 3055
rect 4081 2966 4137 2990
rect 4081 2885 4137 2910
rect 4081 2804 4137 2829
rect 2548 2764 2600 2770
rect 1163 2741 1219 2750
rect 4081 2723 4137 2748
rect 4081 2642 4137 2667
rect 1190 2630 1246 2639
rect 1190 2550 1246 2574
rect 1190 2485 1246 2494
tri 22244 2605 22286 2647 se
rect 22286 2605 22338 3360
rect 22380 3280 22432 3440
rect 22484 3280 22536 3520
rect 22588 3278 22640 3680
tri 22917 3548 22923 3554 se
rect 22923 3548 22975 4187
tri 23213 3788 23219 3794 se
rect 23219 3788 23271 4187
tri 23185 3760 23213 3788 se
rect 23213 3760 23271 3788
rect 23143 3708 23149 3760
rect 23201 3708 23213 3760
rect 23265 3708 23271 3760
tri 24123 3708 24129 3714 se
rect 24129 3708 24181 4187
tri 24095 3680 24123 3708 se
rect 24123 3680 24181 3708
rect 24053 3628 24059 3680
rect 24111 3628 24123 3680
rect 24175 3628 24181 3680
tri 22889 3520 22917 3548 se
rect 22917 3520 22975 3548
rect 22847 3468 22853 3520
rect 22905 3468 22917 3520
rect 22969 3468 22975 3520
tri 24419 3468 24425 3474 se
rect 24425 3468 24477 4187
tri 25251 4112 25285 4146 se
rect 25664 4187 25720 4196
tri 25826 4341 25830 4345 se
rect 25826 4332 25882 4341
rect 25826 4252 25882 4276
rect 25826 4187 25882 4196
rect 25285 4121 25341 4145
rect 25281 4065 25285 4112
rect 25281 4060 25341 4065
tri 25281 4056 25285 4060 ne
rect 25285 4056 25341 4060
tri 26133 3840 26164 3871 se
rect 26164 3862 26220 3871
tri 26220 3862 26229 3871 sw
rect 26220 3840 26229 3862
tri 26229 3840 26251 3862 sw
rect 26671 3853 26727 3862
rect 26133 3788 26139 3840
rect 26191 3788 26203 3806
rect 26255 3788 26261 3840
tri 26668 3788 26671 3791 se
rect 26671 3788 26727 3797
tri 26133 3760 26161 3788 ne
rect 26161 3782 26223 3788
rect 26161 3760 26164 3782
tri 26161 3757 26164 3760 ne
rect 26220 3760 26223 3782
tri 26223 3760 26251 3788 nw
tri 26640 3760 26668 3788 se
rect 26668 3773 26727 3788
rect 26668 3760 26671 3773
tri 26220 3757 26223 3760 nw
rect 26164 3717 26220 3726
rect 26599 3708 26605 3760
rect 26657 3708 26669 3760
rect 26721 3708 26727 3717
rect 26797 3773 26853 3782
tri 26794 3708 26797 3711 se
rect 26797 3708 26853 3717
tri 26766 3680 26794 3708 se
rect 26794 3693 26853 3708
rect 26794 3680 26797 3693
rect 26725 3628 26731 3680
rect 26783 3628 26795 3680
rect 26847 3628 26853 3637
rect 26923 3693 26979 3702
tri 26920 3628 26923 3631 se
rect 26923 3628 26979 3637
tri 26914 3622 26920 3628 se
rect 26920 3622 26979 3628
rect 26293 3613 26349 3622
tri 26290 3548 26293 3551 se
rect 26293 3548 26349 3557
tri 26892 3600 26914 3622 se
rect 26914 3613 26979 3622
rect 26914 3600 26923 3613
tri 26979 3600 27010 3631 sw
rect 26892 3548 26898 3600
rect 26950 3548 26962 3557
rect 27014 3548 27020 3600
tri 26262 3520 26290 3548 se
rect 26290 3533 26349 3548
rect 26290 3520 26293 3533
rect 26221 3468 26227 3520
rect 26279 3468 26291 3520
rect 26343 3468 26349 3477
rect 26419 3533 26475 3542
tri 26416 3468 26419 3471 se
rect 26419 3468 26475 3477
tri 24391 3440 24419 3468 se
rect 24419 3440 24477 3468
tri 26388 3440 26416 3468 se
rect 26416 3453 26475 3468
rect 26416 3440 26419 3453
rect 24349 3388 24355 3440
rect 24407 3388 24419 3440
rect 24471 3388 24477 3440
rect 26347 3388 26353 3440
rect 26405 3388 26417 3440
rect 26469 3388 26475 3397
rect 26545 3453 26601 3462
tri 26542 3388 26545 3391 se
rect 26545 3388 26601 3397
tri 27052 3391 27069 3408 se
rect 27069 3391 27121 4187
tri 27331 3600 27365 3634 se
rect 27365 3600 27417 4187
rect 27289 3548 27295 3600
rect 27347 3548 27359 3600
rect 27411 3548 27417 3600
tri 26601 3388 26604 3391 sw
tri 27049 3388 27052 3391 se
rect 27052 3388 27121 3391
rect 27724 3388 27730 3440
rect 27782 3388 27794 3440
rect 27846 3388 27852 3440
tri 26514 3360 26542 3388 se
rect 26542 3373 26604 3388
rect 26542 3360 26545 3373
rect 26601 3360 26604 3373
tri 26604 3360 26632 3388 sw
tri 27021 3360 27049 3388 se
rect 27049 3360 27121 3388
tri 27766 3360 27794 3388 ne
rect 27794 3360 27852 3388
rect 26514 3308 26520 3360
rect 26636 3339 27121 3360
rect 26572 3308 26584 3317
rect 26636 3308 27090 3339
tri 27090 3308 27121 3339 nw
rect 27489 3308 27495 3360
rect 27547 3308 27559 3360
rect 27611 3308 27617 3360
tri 27794 3354 27800 3360 ne
tri 27531 3286 27553 3308 ne
rect 27553 3286 27617 3308
tri 22640 3278 22648 3286 sw
tri 27553 3278 27561 3286 ne
rect 27561 3278 27617 3286
rect 27800 3279 27852 3360
rect 22640 3274 22648 3278
tri 22648 3274 22652 3278 sw
tri 27561 3274 27565 3278 ne
rect 22640 3272 22652 3274
tri 22652 3272 22654 3274 sw
rect 27565 3272 27617 3278
rect 22640 3252 22654 3272
tri 22654 3252 22674 3272 sw
tri 22536 3172 22570 3206 sw
tri 26157 3102 26175 3120 ne
rect 26175 3102 26191 3120
tri 22432 3086 22448 3102 sw
tri 26175 3086 26191 3102 ne
rect 22432 3068 22448 3086
tri 22448 3068 22466 3086 sw
tri 25076 2982 25110 3016 ne
rect 4081 2561 4137 2586
rect 4081 2480 4137 2505
rect 4081 2399 4137 2424
rect 4081 2318 4137 2343
rect 4081 2253 4137 2262
rect 3592 2121 3644 2127
rect 3592 2057 3644 2069
rect 3592 1999 3644 2005
rect 23251 2060 23449 2069
rect 23307 2059 23393 2060
rect 23307 2007 23324 2059
rect 23376 2007 23393 2059
rect 23307 2004 23393 2007
rect 23251 1989 23449 2004
rect 23251 1968 23254 1989
rect 23306 1968 23324 1989
rect 23307 1937 23324 1968
rect 23376 1968 23394 1989
rect 23446 1968 23449 1989
rect 23376 1937 23393 1968
rect 23307 1919 23393 1937
rect 23307 1912 23324 1919
rect 23251 1876 23254 1912
rect 23306 1876 23324 1912
rect 23307 1867 23324 1876
rect 23376 1912 23393 1919
rect 23376 1876 23394 1912
rect 23446 1876 23449 1912
rect 23376 1867 23393 1876
rect 23307 1849 23393 1867
rect 1934 1835 2050 1841
rect 1986 1832 1998 1835
rect 1934 1776 1964 1783
rect 2020 1776 2050 1783
rect 1934 1770 2050 1776
rect 1986 1748 1998 1770
rect 1759 1719 1815 1728
rect 1759 1653 1761 1663
rect 1813 1653 1815 1663
rect 1759 1641 1815 1653
rect 1759 1639 1761 1641
rect 1813 1639 1815 1641
rect 1759 1574 1815 1583
rect 23307 1820 23324 1849
rect 23251 1797 23254 1820
rect 23306 1797 23324 1820
rect 23376 1820 23393 1849
rect 23376 1797 23394 1820
rect 23446 1797 23449 1820
rect 23251 1783 23449 1797
rect 23307 1778 23393 1783
rect 23307 1727 23324 1778
rect 23251 1726 23254 1727
rect 23306 1726 23324 1727
rect 23376 1727 23393 1778
rect 23376 1726 23394 1727
rect 23446 1726 23449 1727
rect 23251 1718 23449 1726
rect 1934 1705 1964 1718
rect 2020 1705 2050 1718
rect 1986 1663 1998 1692
rect 1934 1640 1964 1653
rect 2020 1640 2050 1653
rect 1986 1588 1998 1607
rect 1934 1578 2050 1588
rect 1934 1575 1964 1578
rect 2020 1575 2050 1578
rect 1934 1522 1964 1523
rect 2020 1522 2050 1523
rect 1934 1510 2050 1522
rect 1986 1493 1998 1510
rect 1934 1445 1964 1458
rect 2020 1445 2050 1458
rect 1986 1408 1998 1437
rect 1934 1380 1964 1393
rect 2020 1380 2050 1393
rect 1986 1328 1998 1352
rect 1934 1323 2050 1328
rect 1934 1315 1964 1323
rect 2020 1315 2050 1323
rect 1986 1263 1998 1267
rect 1934 1250 2050 1263
rect 1986 1238 1998 1250
rect 1934 1185 1964 1198
rect 2020 1185 2050 1198
rect 1986 1153 1998 1182
rect 1934 1120 1964 1133
rect 2020 1120 2050 1133
rect 1986 1068 1998 1097
rect 23515 1182 23524 1238
rect 23580 1182 23650 1238
rect 23706 1234 23977 1238
rect 23706 1182 23788 1234
rect 23840 1182 23852 1234
rect 23904 1182 23916 1234
rect 23968 1182 23977 1234
rect 23515 1144 23977 1182
rect 23515 1088 23524 1144
rect 23580 1088 23650 1144
rect 23706 1140 23977 1144
rect 23706 1088 23788 1140
rect 23840 1088 23852 1140
rect 23904 1088 23916 1140
rect 23968 1088 23977 1140
rect 1934 1055 1964 1068
rect 2020 1055 2050 1068
rect 1986 1003 1998 1012
rect 1934 990 2050 1003
rect 1986 983 1998 990
rect 8803 977 8812 1033
rect 8868 977 8892 1033
rect 8948 977 8957 1033
rect 1934 927 1964 938
rect 2020 927 2050 938
rect 1934 925 2050 927
rect 1986 898 1998 925
rect 1934 860 1964 873
rect 2020 860 2050 873
rect 1986 813 1998 842
rect 1934 795 1964 808
rect 2020 795 2050 808
rect 1986 743 1998 757
rect 1934 730 2050 743
rect 1986 728 1998 730
rect 1934 672 1964 678
rect 2020 672 2050 678
rect 1934 664 2050 672
rect 1986 643 1998 664
rect 1934 598 1964 612
rect 2020 598 2050 612
rect 1986 558 1998 587
rect 1934 532 1964 546
rect 2020 532 2050 546
rect 1986 480 1998 502
rect 1934 473 2050 480
rect 1934 466 1964 473
rect 2020 466 2050 473
rect 23515 456 23524 512
rect 23580 456 23650 512
rect 23706 456 23715 512
rect 1986 414 1998 417
rect 1934 408 2050 414
rect 17775 391 18175 427
rect 17775 335 17784 391
rect 17840 335 17866 391
rect 17922 335 17948 391
rect 18004 335 18029 391
rect 18085 335 18110 391
rect 18166 335 18175 391
rect 17775 299 18175 335
rect 18259 410 18535 421
rect 18259 354 18268 410
rect 18324 354 18367 410
rect 18423 354 18465 410
rect 18521 354 18535 410
rect 23515 418 23715 456
rect 23515 362 23524 418
rect 23580 362 23650 418
rect 23706 362 23715 418
rect 18259 230 18535 354
rect 4004 211 4056 217
tri 4056 193 4080 217 sw
rect 4056 183 4080 193
tri 4080 183 4090 193 sw
rect 4056 159 4703 183
rect 4004 147 4703 159
rect 4056 127 4703 147
rect 4759 127 4783 183
rect 4839 127 4848 183
rect 16769 137 16778 193
rect 16834 137 16871 193
rect 16927 137 16964 193
rect 17020 137 17057 193
rect 17113 137 17149 193
rect 17205 137 17241 193
rect 17297 137 17306 193
rect 18259 178 18265 230
rect 18317 178 18336 230
rect 18388 178 18407 230
rect 18459 178 18477 230
rect 18529 178 18535 230
rect 4004 89 4056 95
tri 4056 89 4094 127 nw
rect 16769 63 17306 137
rect 16769 7 16778 63
rect 16834 7 16871 63
rect 16927 7 16964 63
rect 17020 7 17057 63
rect 17113 7 17149 63
rect 17205 7 17241 63
rect 17297 7 17306 63
<< via2 >>
rect 12008 38680 12056 38729
rect 12056 38680 12064 38729
rect 12091 38680 12125 38729
rect 12125 38680 12142 38729
rect 12142 38680 12147 38729
rect 12174 38680 12194 38729
rect 12194 38680 12211 38729
rect 12211 38680 12230 38729
rect 12257 38680 12263 38729
rect 12263 38680 12280 38729
rect 12280 38680 12313 38729
rect 12339 38680 12348 38729
rect 12348 38680 12395 38729
rect 12008 38673 12064 38680
rect 12091 38673 12147 38680
rect 12174 38673 12230 38680
rect 12257 38673 12313 38680
rect 12339 38673 12395 38680
rect 12008 38588 12064 38595
rect 12091 38588 12147 38595
rect 12174 38588 12230 38595
rect 12257 38588 12313 38595
rect 12339 38588 12395 38595
rect 12008 38539 12056 38588
rect 12056 38539 12064 38588
rect 12091 38539 12125 38588
rect 12125 38539 12142 38588
rect 12142 38539 12147 38588
rect 12174 38539 12194 38588
rect 12194 38539 12211 38588
rect 12211 38539 12230 38588
rect 12257 38539 12263 38588
rect 12263 38539 12280 38588
rect 12280 38539 12313 38588
rect 12339 38539 12348 38588
rect 12348 38539 12395 38588
rect 25870 37101 25926 37157
rect 25870 37021 25926 37077
rect 23398 34313 23454 34369
rect 23478 34313 23534 34369
rect 23558 34313 23614 34369
rect 23638 34313 23694 34369
rect 23398 34231 23454 34287
rect 23478 34231 23534 34287
rect 23558 34231 23614 34287
rect 23638 34231 23694 34287
rect 23398 34149 23454 34205
rect 23478 34149 23534 34205
rect 23558 34149 23614 34205
rect 23638 34149 23694 34205
rect 23398 34067 23454 34123
rect 23478 34067 23534 34123
rect 23558 34067 23614 34123
rect 23638 34067 23694 34123
rect 23398 33984 23454 34040
rect 23478 33984 23534 34040
rect 23558 33984 23614 34040
rect 23638 33984 23694 34040
rect 23398 33901 23454 33957
rect 23478 33901 23534 33957
rect 23558 33901 23614 33957
rect 23638 33901 23694 33957
rect 3732 33050 3788 33106
rect 3846 33050 3902 33106
rect 3732 32954 3788 33010
rect 3846 32954 3902 33010
rect 3732 32858 3788 32914
rect 3846 32858 3902 32914
rect 3732 32762 3788 32818
rect 3846 32762 3902 32818
rect 3732 32665 3788 32721
rect 3846 32665 3902 32721
rect 23398 32967 23454 33023
rect 23478 32967 23534 33023
rect 23558 32967 23614 33023
rect 23638 32967 23694 33023
rect 23398 32885 23454 32941
rect 23478 32885 23534 32941
rect 23558 32885 23614 32941
rect 23638 32885 23694 32941
rect 23398 32803 23454 32859
rect 23478 32803 23534 32859
rect 23558 32803 23614 32859
rect 23638 32803 23694 32859
rect 23398 32720 23454 32776
rect 23478 32720 23534 32776
rect 23558 32720 23614 32776
rect 23638 32720 23694 32776
rect 23398 32637 23454 32693
rect 23478 32637 23534 32693
rect 23558 32637 23614 32693
rect 23638 32637 23694 32693
rect 23398 32554 23454 32610
rect 23478 32554 23534 32610
rect 23558 32554 23614 32610
rect 23638 32554 23694 32610
rect 619 32124 675 32180
rect 619 32044 675 32100
rect 619 31964 675 32020
rect 829 31847 885 31903
rect 829 31767 885 31823
rect 829 31687 885 31743
rect 1667 31063 1719 31112
rect 1719 31063 1723 31112
rect 1667 31056 1723 31063
rect 1747 31063 1751 31112
rect 1751 31063 1803 31112
rect 1747 31056 1803 31063
rect 1827 31063 1835 31112
rect 1835 31063 1883 31112
rect 1827 31056 1883 31063
rect 1667 30984 1719 31025
rect 1719 30984 1723 31025
rect 1667 30969 1723 30984
rect 1747 30984 1751 31025
rect 1751 30984 1803 31025
rect 1747 30969 1803 30984
rect 1827 30984 1835 31025
rect 1835 30984 1883 31025
rect 1827 30969 1883 30984
rect 1667 30905 1719 30938
rect 1719 30905 1723 30938
rect 1667 30882 1723 30905
rect 1747 30905 1751 30938
rect 1751 30905 1803 30938
rect 1747 30882 1803 30905
rect 1827 30905 1835 30938
rect 1835 30905 1883 30938
rect 1827 30882 1883 30905
rect 1667 30826 1719 30850
rect 1719 30826 1723 30850
rect 1667 30794 1723 30826
rect 1747 30826 1751 30850
rect 1751 30826 1803 30850
rect 1747 30794 1803 30826
rect 1827 30826 1835 30850
rect 1835 30826 1883 30850
rect 1827 30794 1883 30826
rect 18744 23690 18800 23746
rect 18854 23690 18910 23746
rect 18964 23690 19020 23746
rect 18744 23603 18800 23659
rect 18854 23603 18910 23659
rect 18964 23603 19020 23659
rect 18744 23516 18800 23572
rect 18854 23516 18910 23572
rect 18964 23516 19020 23572
rect 18744 23429 18800 23485
rect 18854 23429 18910 23485
rect 18964 23429 19020 23485
rect 18744 23342 18800 23398
rect 18854 23342 18910 23398
rect 18964 23342 19020 23398
rect 18744 23255 18800 23311
rect 18854 23255 18910 23311
rect 18964 23255 19020 23311
rect 18744 23167 18800 23223
rect 18854 23167 18910 23223
rect 18964 23167 19020 23223
rect 18744 23079 18800 23135
rect 18854 23079 18910 23135
rect 18964 23079 19020 23135
rect 18744 22991 18800 23047
rect 18854 22991 18910 23047
rect 18964 22991 19020 23047
rect 18744 22903 18800 22959
rect 18854 22903 18910 22959
rect 18964 22903 19020 22959
rect 27056 23224 27102 23272
rect 27102 23224 27112 23272
rect 27140 23224 27173 23272
rect 27173 23224 27192 23272
rect 27192 23224 27196 23272
rect 27224 23224 27244 23272
rect 27244 23224 27262 23272
rect 27262 23224 27280 23272
rect 27308 23224 27314 23272
rect 27314 23224 27332 23272
rect 27332 23224 27364 23272
rect 27392 23224 27402 23272
rect 27402 23224 27448 23272
rect 27476 23224 27524 23272
rect 27524 23224 27532 23272
rect 27056 23216 27112 23224
rect 27140 23216 27196 23224
rect 27224 23216 27280 23224
rect 27308 23216 27364 23224
rect 27392 23216 27448 23224
rect 27476 23216 27532 23224
rect 27056 23158 27102 23192
rect 27102 23158 27112 23192
rect 27140 23158 27173 23192
rect 27173 23158 27192 23192
rect 27192 23158 27196 23192
rect 27224 23158 27244 23192
rect 27244 23158 27262 23192
rect 27262 23158 27280 23192
rect 27308 23158 27314 23192
rect 27314 23158 27332 23192
rect 27332 23158 27364 23192
rect 27392 23158 27402 23192
rect 27402 23158 27448 23192
rect 27476 23158 27524 23192
rect 27524 23158 27532 23192
rect 27056 23144 27112 23158
rect 27140 23144 27196 23158
rect 27224 23144 27280 23158
rect 27308 23144 27364 23158
rect 27392 23144 27448 23158
rect 27476 23144 27532 23158
rect 27056 23136 27102 23144
rect 27102 23136 27112 23144
rect 27140 23136 27173 23144
rect 27173 23136 27192 23144
rect 27192 23136 27196 23144
rect 27224 23136 27244 23144
rect 27244 23136 27262 23144
rect 27262 23136 27280 23144
rect 27308 23136 27314 23144
rect 27314 23136 27332 23144
rect 27332 23136 27364 23144
rect 27392 23136 27402 23144
rect 27402 23136 27448 23144
rect 27056 23092 27102 23112
rect 27102 23092 27112 23112
rect 27140 23092 27173 23112
rect 27173 23092 27192 23112
rect 27192 23092 27196 23112
rect 27224 23092 27244 23112
rect 27244 23092 27262 23112
rect 27262 23092 27280 23112
rect 27308 23092 27314 23112
rect 27314 23092 27332 23112
rect 27332 23092 27364 23112
rect 27392 23092 27402 23112
rect 27402 23092 27448 23112
rect 27476 23136 27524 23144
rect 27524 23136 27532 23144
rect 27476 23092 27524 23112
rect 27524 23092 27532 23112
rect 27056 23078 27112 23092
rect 27140 23078 27196 23092
rect 27224 23078 27280 23092
rect 27308 23078 27364 23092
rect 27392 23078 27448 23092
rect 27476 23078 27532 23092
rect 27056 23056 27102 23078
rect 27102 23056 27112 23078
rect 27140 23056 27173 23078
rect 27173 23056 27192 23078
rect 27192 23056 27196 23078
rect 27224 23056 27244 23078
rect 27244 23056 27262 23078
rect 27262 23056 27280 23078
rect 27308 23056 27314 23078
rect 27314 23056 27332 23078
rect 27332 23056 27364 23078
rect 27392 23056 27402 23078
rect 27402 23056 27448 23078
rect 27056 23026 27102 23032
rect 27102 23026 27112 23032
rect 27140 23026 27173 23032
rect 27173 23026 27192 23032
rect 27192 23026 27196 23032
rect 27224 23026 27244 23032
rect 27244 23026 27262 23032
rect 27262 23026 27280 23032
rect 27308 23026 27314 23032
rect 27314 23026 27332 23032
rect 27332 23026 27364 23032
rect 27392 23026 27402 23032
rect 27402 23026 27448 23032
rect 27476 23056 27524 23078
rect 27524 23056 27532 23078
rect 27476 23026 27524 23032
rect 27524 23026 27532 23032
rect 27056 23012 27112 23026
rect 27140 23012 27196 23026
rect 27224 23012 27280 23026
rect 27308 23012 27364 23026
rect 27392 23012 27448 23026
rect 27476 23012 27532 23026
rect 27056 22976 27102 23012
rect 27102 22976 27112 23012
rect 27140 22976 27173 23012
rect 27173 22976 27192 23012
rect 27192 22976 27196 23012
rect 27224 22976 27244 23012
rect 27244 22976 27262 23012
rect 27262 22976 27280 23012
rect 27308 22976 27314 23012
rect 27314 22976 27332 23012
rect 27332 22976 27364 23012
rect 27392 22976 27402 23012
rect 27402 22976 27448 23012
rect 27476 22976 27524 23012
rect 27524 22976 27532 23012
rect 27056 22946 27112 22952
rect 27140 22946 27196 22952
rect 27224 22946 27280 22952
rect 27308 22946 27364 22952
rect 27392 22946 27448 22952
rect 27476 22946 27532 22952
rect 27056 22896 27102 22946
rect 27102 22896 27112 22946
rect 27140 22896 27173 22946
rect 27173 22896 27192 22946
rect 27192 22896 27196 22946
rect 27224 22896 27244 22946
rect 27244 22896 27262 22946
rect 27262 22896 27280 22946
rect 27308 22896 27314 22946
rect 27314 22896 27332 22946
rect 27332 22896 27364 22946
rect 27392 22896 27402 22946
rect 27402 22896 27448 22946
rect 27476 22896 27524 22946
rect 27524 22896 27532 22946
rect 18744 22815 18800 22871
rect 18854 22815 18910 22871
rect 18964 22815 19020 22871
rect 27345 22809 27355 22858
rect 27355 22809 27401 22858
rect 27483 22809 27535 22858
rect 27535 22809 27539 22858
rect 27345 22802 27401 22809
rect 27483 22802 27539 22809
rect 27345 22742 27355 22776
rect 27355 22742 27401 22776
rect 27483 22742 27535 22776
rect 27535 22742 27539 22776
rect 27345 22727 27401 22742
rect 27483 22727 27539 22742
rect 27345 22720 27355 22727
rect 27355 22720 27401 22727
rect 27345 22675 27355 22694
rect 27355 22675 27401 22694
rect 27483 22720 27535 22727
rect 27535 22720 27539 22727
rect 27483 22675 27535 22694
rect 27535 22675 27539 22694
rect 27345 22660 27401 22675
rect 27483 22660 27539 22675
rect 27345 22638 27355 22660
rect 27355 22638 27401 22660
rect 27345 22608 27355 22612
rect 27355 22608 27401 22612
rect 27483 22638 27535 22660
rect 27535 22638 27539 22660
rect 27483 22608 27535 22612
rect 27535 22608 27539 22612
rect 27345 22593 27401 22608
rect 27483 22593 27539 22608
rect 27345 22556 27355 22593
rect 27355 22556 27401 22593
rect 27483 22556 27535 22593
rect 27535 22556 27539 22593
rect 27345 22526 27401 22530
rect 27483 22526 27539 22530
rect 27345 22474 27355 22526
rect 27355 22474 27401 22526
rect 27483 22474 27535 22526
rect 27535 22474 27539 22526
rect 27345 22407 27355 22448
rect 27355 22407 27401 22448
rect 27483 22407 27535 22448
rect 27535 22407 27539 22448
rect 27345 22392 27401 22407
rect 27483 22392 27539 22407
rect 27345 22340 27355 22366
rect 27355 22340 27401 22366
rect 27483 22340 27535 22366
rect 27535 22340 27539 22366
rect 27345 22324 27401 22340
rect 27483 22324 27539 22340
rect 27345 22310 27355 22324
rect 27355 22310 27401 22324
rect 27345 22272 27355 22284
rect 27355 22272 27401 22284
rect 27483 22310 27535 22324
rect 27535 22310 27539 22324
rect 27483 22272 27535 22284
rect 27535 22272 27539 22284
rect 27345 22256 27401 22272
rect 27483 22256 27539 22272
rect 27345 22228 27355 22256
rect 27355 22228 27401 22256
rect 27483 22228 27535 22256
rect 27535 22228 27539 22256
rect 27345 22188 27401 22202
rect 27483 22188 27539 22202
rect 27345 22146 27355 22188
rect 27355 22146 27401 22188
rect 27483 22146 27535 22188
rect 27535 22146 27539 22188
rect 27345 22064 27401 22120
rect 27483 22064 27539 22120
rect 27345 21982 27401 22038
rect 27483 21982 27539 22038
rect 27345 21900 27401 21956
rect 27483 21900 27539 21956
rect 27345 21818 27401 21874
rect 27483 21818 27539 21874
rect 27345 21736 27401 21792
rect 27483 21736 27539 21792
rect 27345 21654 27401 21710
rect 27483 21654 27539 21710
rect 27345 21572 27401 21628
rect 27483 21572 27539 21628
rect 27345 21490 27401 21546
rect 27483 21490 27539 21546
rect 27345 21408 27401 21464
rect 27483 21408 27539 21464
rect 1870 21312 1888 21362
rect 1888 21312 1908 21362
rect 1908 21312 1926 21362
rect 1870 21306 1926 21312
rect 1870 21248 1888 21282
rect 1888 21248 1908 21282
rect 1908 21248 1926 21282
rect 1870 21236 1926 21248
rect 1870 21226 1888 21236
rect 1888 21226 1908 21236
rect 1908 21226 1926 21236
rect 1870 21184 1888 21202
rect 1888 21184 1908 21202
rect 1908 21184 1926 21202
rect 1870 21172 1926 21184
rect 1870 21146 1888 21172
rect 1888 21146 1908 21172
rect 1908 21146 1926 21172
rect 1870 21120 1888 21122
rect 1888 21120 1908 21122
rect 1908 21120 1926 21122
rect 27345 21375 27401 21382
rect 27345 21326 27364 21375
rect 27364 21326 27401 21375
rect 27483 21367 27539 21382
rect 27483 21326 27515 21367
rect 27515 21326 27539 21367
rect 27345 21269 27401 21299
rect 27483 21288 27539 21299
rect 27345 21243 27364 21269
rect 27364 21243 27401 21269
rect 27483 21243 27515 21288
rect 27515 21243 27539 21288
rect 27345 21160 27401 21216
rect 27483 21209 27539 21216
rect 27483 21160 27515 21209
rect 27515 21160 27539 21209
rect 1870 21108 1926 21120
rect 1870 21066 1888 21108
rect 1888 21066 1908 21108
rect 1908 21066 1926 21108
rect 1870 20992 1888 21042
rect 1888 20992 1908 21042
rect 1908 20992 1926 21042
rect 1870 20986 1926 20992
rect 1870 20928 1888 20962
rect 1888 20928 1908 20962
rect 1908 20928 1926 20962
rect 1870 20916 1926 20928
rect 1870 20906 1888 20916
rect 1888 20906 1908 20916
rect 1908 20906 1926 20916
rect 1870 20864 1888 20882
rect 1888 20864 1908 20882
rect 1908 20864 1926 20882
rect 1870 20852 1926 20864
rect 1870 20826 1888 20852
rect 1888 20826 1908 20852
rect 1908 20826 1926 20852
rect 1870 20800 1888 20802
rect 1888 20800 1908 20802
rect 1908 20800 1926 20802
rect 1870 20788 1926 20800
rect 1870 20746 1888 20788
rect 1888 20746 1908 20788
rect 1908 20746 1926 20788
rect 1870 20672 1888 20722
rect 1888 20672 1908 20722
rect 1908 20672 1926 20722
rect 1870 20666 1926 20672
rect 1870 20608 1888 20642
rect 1888 20608 1908 20642
rect 1908 20608 1926 20642
rect 2423 20737 2479 20793
rect 2423 20652 2479 20708
rect 1870 20596 1926 20608
rect 1870 20586 1888 20596
rect 1888 20586 1908 20596
rect 1908 20586 1926 20596
rect 1870 20544 1888 20562
rect 1888 20544 1908 20562
rect 1908 20544 1926 20562
rect 1870 20532 1926 20544
rect 1870 20506 1888 20532
rect 1888 20506 1908 20532
rect 1908 20506 1926 20532
rect 1870 20480 1888 20482
rect 1888 20480 1908 20482
rect 1908 20480 1926 20482
rect 1870 20468 1926 20480
rect 1870 20426 1888 20468
rect 1888 20426 1908 20468
rect 1908 20426 1926 20468
rect 1870 20352 1888 20401
rect 1888 20352 1908 20401
rect 1908 20352 1926 20401
rect 1870 20345 1926 20352
rect 1870 20288 1888 20320
rect 1888 20288 1908 20320
rect 1908 20288 1926 20320
rect 1870 20276 1926 20288
rect 1870 20264 1888 20276
rect 1888 20264 1908 20276
rect 1908 20264 1926 20276
rect 1870 20224 1888 20239
rect 1888 20224 1908 20239
rect 1908 20224 1926 20239
rect 1870 20212 1926 20224
rect 1870 20183 1888 20212
rect 1888 20183 1908 20212
rect 1908 20183 1926 20212
rect 1870 20148 1926 20158
rect 1870 20102 1888 20148
rect 1888 20102 1908 20148
rect 1908 20102 1926 20148
rect 1870 20032 1888 20077
rect 1888 20032 1908 20077
rect 1908 20032 1926 20077
rect 1870 20021 1926 20032
rect 1870 19968 1888 19996
rect 1888 19968 1908 19996
rect 1908 19968 1926 19996
rect 1870 19956 1926 19968
rect 1870 19940 1888 19956
rect 1888 19940 1908 19956
rect 1908 19940 1926 19956
rect 1870 19904 1888 19915
rect 1888 19904 1908 19915
rect 1908 19904 1926 19915
rect 1870 19892 1926 19904
rect 1870 19859 1888 19892
rect 1888 19859 1908 19892
rect 1908 19859 1926 19892
rect 1870 19828 1926 19834
rect 1870 19778 1888 19828
rect 1888 19778 1908 19828
rect 1908 19778 1926 19828
rect 1870 19712 1888 19753
rect 1888 19712 1908 19753
rect 1908 19712 1926 19753
rect 1870 19700 1926 19712
rect 1870 19697 1888 19700
rect 1888 19697 1908 19700
rect 1908 19697 1926 19700
rect 1870 19648 1888 19672
rect 1888 19648 1908 19672
rect 1908 19648 1926 19672
rect 1870 19636 1926 19648
rect 1870 19616 1888 19636
rect 1888 19616 1908 19636
rect 1908 19616 1926 19636
rect 1870 19584 1888 19591
rect 1888 19584 1908 19591
rect 1908 19584 1926 19591
rect 1870 19572 1926 19584
rect 1870 19535 1888 19572
rect 1888 19535 1908 19572
rect 1908 19535 1926 19572
rect 1870 19507 1926 19510
rect 1870 19455 1888 19507
rect 1888 19455 1908 19507
rect 1908 19455 1926 19507
rect 1870 19454 1926 19455
rect 1870 19390 1888 19429
rect 1888 19390 1908 19429
rect 1908 19390 1926 19429
rect 1870 19377 1926 19390
rect 1870 19373 1888 19377
rect 1888 19373 1908 19377
rect 1908 19373 1926 19377
rect 1870 19325 1888 19348
rect 1888 19325 1908 19348
rect 1908 19325 1926 19348
rect 1870 19312 1926 19325
rect 1870 19292 1888 19312
rect 1888 19292 1908 19312
rect 1908 19292 1926 19312
rect 1870 19260 1888 19267
rect 1888 19260 1908 19267
rect 1908 19260 1926 19267
rect 1870 19247 1926 19260
rect 1870 19211 1888 19247
rect 1888 19211 1908 19247
rect 1908 19211 1926 19247
rect 1870 19182 1926 19186
rect 1870 19130 1888 19182
rect 1888 19130 1908 19182
rect 1908 19130 1926 19182
rect 1870 19065 1888 19105
rect 1888 19065 1908 19105
rect 1908 19065 1926 19105
rect 1870 19052 1926 19065
rect 1870 19049 1888 19052
rect 1888 19049 1908 19052
rect 1908 19049 1926 19052
rect 1870 19000 1888 19024
rect 1888 19000 1908 19024
rect 1908 19000 1926 19024
rect 1870 18987 1926 19000
rect 1870 18968 1888 18987
rect 1888 18968 1908 18987
rect 1908 18968 1926 18987
rect 1870 18935 1888 18943
rect 1888 18935 1908 18943
rect 1908 18935 1926 18943
rect 1870 18922 1926 18935
rect 1870 18887 1888 18922
rect 1888 18887 1908 18922
rect 1908 18887 1926 18922
rect 1870 18857 1926 18862
rect 1870 18806 1888 18857
rect 1888 18806 1908 18857
rect 1908 18806 1926 18857
rect 1870 18740 1888 18781
rect 1888 18740 1908 18781
rect 1908 18740 1926 18781
rect 1870 18727 1926 18740
rect 1870 18725 1888 18727
rect 1888 18725 1908 18727
rect 1908 18725 1926 18727
rect 1870 18675 1888 18700
rect 1888 18675 1908 18700
rect 1908 18675 1926 18700
rect 1870 18662 1926 18675
rect 1870 18644 1888 18662
rect 1888 18644 1908 18662
rect 1908 18644 1926 18662
rect 1870 18610 1888 18619
rect 1888 18610 1908 18619
rect 1908 18610 1926 18619
rect 1870 18597 1926 18610
rect 1870 18563 1888 18597
rect 1888 18563 1908 18597
rect 1908 18563 1926 18597
rect 1870 18532 1926 18538
rect 1870 18482 1888 18532
rect 1888 18482 1908 18532
rect 1908 18482 1926 18532
rect 1771 18192 1827 18201
rect 1851 18192 1907 18201
rect 1931 18192 1987 18201
rect 1771 18145 1796 18192
rect 1796 18145 1827 18192
rect 1851 18145 1864 18192
rect 1864 18145 1907 18192
rect 1931 18145 1932 18192
rect 1932 18145 1984 18192
rect 1984 18145 1987 18192
rect 1771 18068 1796 18112
rect 1796 18068 1827 18112
rect 1851 18068 1864 18112
rect 1864 18068 1907 18112
rect 1931 18068 1932 18112
rect 1932 18068 1984 18112
rect 1984 18068 1987 18112
rect 1771 18056 1827 18068
rect 1851 18056 1907 18068
rect 1931 18056 1987 18068
rect 1771 17995 1796 18023
rect 1796 17995 1827 18023
rect 1851 17995 1864 18023
rect 1864 17995 1907 18023
rect 1931 17995 1932 18023
rect 1932 17995 1984 18023
rect 1984 17995 1987 18023
rect 1771 17974 1827 17995
rect 1851 17974 1907 17995
rect 1931 17974 1987 17995
rect 1771 17967 1796 17974
rect 1796 17967 1827 17974
rect 1851 17967 1864 17974
rect 1864 17967 1907 17974
rect 1931 17967 1932 17974
rect 1932 17967 1984 17974
rect 1984 17967 1987 17974
rect 1771 17922 1796 17934
rect 1796 17922 1827 17934
rect 1851 17922 1864 17934
rect 1864 17922 1907 17934
rect 1931 17922 1932 17934
rect 1932 17922 1984 17934
rect 1984 17922 1987 17934
rect 1771 17901 1827 17922
rect 1851 17901 1907 17922
rect 1931 17901 1987 17922
rect 1771 17878 1796 17901
rect 1796 17878 1827 17901
rect 1851 17878 1864 17901
rect 1864 17878 1907 17901
rect 1931 17878 1932 17901
rect 1932 17878 1984 17901
rect 1984 17878 1987 17901
rect 1771 17828 1827 17845
rect 1851 17828 1907 17845
rect 1931 17828 1987 17845
rect 1771 17789 1796 17828
rect 1796 17789 1827 17828
rect 1851 17789 1864 17828
rect 1864 17789 1907 17828
rect 1931 17789 1932 17828
rect 1932 17789 1984 17828
rect 1984 17789 1987 17828
rect 1771 17703 1796 17755
rect 1796 17703 1827 17755
rect 1851 17703 1864 17755
rect 1864 17703 1907 17755
rect 1931 17703 1932 17755
rect 1932 17703 1984 17755
rect 1984 17703 1987 17755
rect 1771 17699 1827 17703
rect 1851 17699 1907 17703
rect 1931 17699 1987 17703
rect 1771 17518 1987 17527
rect 1771 17466 1796 17518
rect 1796 17466 1848 17518
rect 1848 17466 1864 17518
rect 1864 17466 1916 17518
rect 1916 17466 1932 17518
rect 1932 17466 1984 17518
rect 1984 17466 1987 17518
rect 1771 17453 1987 17466
rect 1771 17401 1796 17453
rect 1796 17401 1848 17453
rect 1848 17401 1864 17453
rect 1864 17401 1916 17453
rect 1916 17401 1932 17453
rect 1932 17401 1984 17453
rect 1984 17401 1987 17453
rect 1771 17391 1987 17401
rect 1771 17335 1796 17366
rect 1796 17335 1827 17366
rect 1851 17335 1864 17366
rect 1864 17335 1907 17366
rect 1931 17335 1932 17366
rect 1932 17335 1984 17366
rect 1984 17335 1987 17366
rect 1771 17321 1827 17335
rect 1851 17321 1907 17335
rect 1931 17321 1987 17335
rect 1771 17310 1796 17321
rect 1796 17310 1827 17321
rect 1851 17310 1864 17321
rect 1864 17310 1907 17321
rect 1931 17310 1932 17321
rect 1932 17310 1984 17321
rect 1984 17310 1987 17321
rect 1771 17269 1796 17285
rect 1796 17269 1827 17285
rect 1851 17269 1864 17285
rect 1864 17269 1907 17285
rect 1931 17269 1932 17285
rect 1932 17269 1984 17285
rect 1984 17269 1987 17285
rect 1771 17255 1827 17269
rect 1851 17255 1907 17269
rect 1931 17255 1987 17269
rect 1771 17229 1796 17255
rect 1796 17229 1827 17255
rect 1851 17229 1864 17255
rect 1864 17229 1907 17255
rect 1931 17229 1932 17255
rect 1932 17229 1984 17255
rect 1984 17229 1987 17255
rect 1771 17203 1796 17204
rect 1796 17203 1827 17204
rect 1851 17203 1864 17204
rect 1864 17203 1907 17204
rect 1931 17203 1932 17204
rect 1932 17203 1984 17204
rect 1984 17203 1987 17204
rect 1771 17189 1827 17203
rect 1851 17189 1907 17203
rect 1931 17189 1987 17203
rect 1771 17148 1796 17189
rect 1796 17148 1827 17189
rect 1851 17148 1864 17189
rect 1864 17148 1907 17189
rect 1931 17148 1932 17189
rect 1932 17148 1984 17189
rect 1984 17148 1987 17189
rect 1771 17071 1796 17123
rect 1796 17071 1827 17123
rect 1851 17071 1864 17123
rect 1864 17071 1907 17123
rect 1931 17071 1932 17123
rect 1932 17071 1984 17123
rect 1984 17071 1987 17123
rect 1771 17067 1827 17071
rect 1851 17067 1907 17071
rect 1931 17067 1987 17071
rect 1771 16313 1827 16322
rect 1851 16313 1907 16322
rect 1931 16313 1987 16322
rect 1771 16266 1796 16313
rect 1796 16266 1827 16313
rect 1851 16266 1864 16313
rect 1864 16266 1907 16313
rect 1931 16266 1932 16313
rect 1932 16266 1984 16313
rect 1984 16266 1987 16313
rect 1771 16197 1796 16235
rect 1796 16197 1827 16235
rect 1851 16197 1864 16235
rect 1864 16197 1907 16235
rect 1931 16197 1932 16235
rect 1932 16197 1984 16235
rect 1984 16197 1987 16235
rect 1771 16185 1827 16197
rect 1851 16185 1907 16197
rect 1931 16185 1987 16197
rect 1771 16179 1796 16185
rect 1796 16179 1827 16185
rect 1851 16179 1864 16185
rect 1864 16179 1907 16185
rect 1931 16179 1932 16185
rect 1932 16179 1984 16185
rect 1984 16179 1987 16185
rect 1771 16133 1796 16148
rect 1796 16133 1827 16148
rect 1851 16133 1864 16148
rect 1864 16133 1907 16148
rect 1931 16133 1932 16148
rect 1932 16133 1984 16148
rect 1984 16133 1987 16148
rect 1771 16121 1827 16133
rect 1851 16121 1907 16133
rect 1931 16121 1987 16133
rect 1771 16092 1796 16121
rect 1796 16092 1827 16121
rect 1851 16092 1864 16121
rect 1864 16092 1907 16121
rect 1931 16092 1932 16121
rect 1932 16092 1984 16121
rect 1984 16092 1987 16121
rect 1771 16057 1827 16061
rect 1851 16057 1907 16061
rect 1931 16057 1987 16061
rect 1771 16005 1796 16057
rect 1796 16005 1827 16057
rect 1851 16005 1864 16057
rect 1864 16005 1907 16057
rect 1931 16005 1932 16057
rect 1932 16005 1984 16057
rect 1984 16005 1987 16057
rect 1771 15941 1796 15974
rect 1796 15941 1827 15974
rect 1851 15941 1864 15974
rect 1864 15941 1907 15974
rect 1931 15941 1932 15974
rect 1932 15941 1984 15974
rect 1984 15941 1987 15974
rect 1771 15929 1827 15941
rect 1851 15929 1907 15941
rect 1931 15929 1987 15941
rect 1771 15918 1796 15929
rect 1796 15918 1827 15929
rect 1851 15918 1864 15929
rect 1864 15918 1907 15929
rect 1931 15918 1932 15929
rect 1932 15918 1984 15929
rect 1984 15918 1987 15929
rect 1771 15877 1796 15887
rect 1796 15877 1827 15887
rect 1851 15877 1864 15887
rect 1864 15877 1907 15887
rect 1931 15877 1932 15887
rect 1932 15877 1984 15887
rect 1984 15877 1987 15887
rect 1771 15864 1827 15877
rect 1851 15864 1907 15877
rect 1931 15864 1987 15877
rect 1771 15831 1796 15864
rect 1796 15831 1827 15864
rect 1851 15831 1864 15864
rect 1864 15831 1907 15864
rect 1931 15831 1932 15864
rect 1932 15831 1984 15864
rect 1984 15831 1987 15864
rect 1771 15799 1827 15800
rect 1851 15799 1907 15800
rect 1931 15799 1987 15800
rect 1771 15747 1796 15799
rect 1796 15747 1827 15799
rect 1851 15747 1864 15799
rect 1864 15747 1907 15799
rect 1931 15747 1932 15799
rect 1932 15747 1984 15799
rect 1984 15747 1987 15799
rect 1771 15744 1827 15747
rect 1851 15744 1907 15747
rect 1931 15744 1987 15747
rect 1771 15682 1796 15713
rect 1796 15682 1827 15713
rect 1851 15682 1864 15713
rect 1864 15682 1907 15713
rect 1931 15682 1932 15713
rect 1932 15682 1984 15713
rect 1984 15682 1987 15713
rect 1771 15669 1827 15682
rect 1851 15669 1907 15682
rect 1931 15669 1987 15682
rect 1771 15657 1796 15669
rect 1796 15657 1827 15669
rect 1851 15657 1864 15669
rect 1864 15657 1907 15669
rect 1931 15657 1932 15669
rect 1932 15657 1984 15669
rect 1984 15657 1987 15669
rect 1771 15617 1796 15626
rect 1796 15617 1827 15626
rect 1851 15617 1864 15626
rect 1864 15617 1907 15626
rect 1931 15617 1932 15626
rect 1932 15617 1984 15626
rect 1984 15617 1987 15626
rect 1771 15604 1827 15617
rect 1851 15604 1907 15617
rect 1931 15604 1987 15617
rect 1771 15570 1796 15604
rect 1796 15570 1827 15604
rect 1851 15570 1864 15604
rect 1864 15570 1907 15604
rect 1931 15570 1932 15604
rect 1932 15570 1984 15604
rect 1984 15570 1987 15604
rect 1771 15487 1796 15539
rect 1796 15487 1827 15539
rect 1851 15487 1864 15539
rect 1864 15487 1907 15539
rect 1931 15487 1932 15539
rect 1932 15487 1984 15539
rect 1984 15487 1987 15539
rect 1771 15483 1827 15487
rect 1851 15483 1907 15487
rect 1931 15483 1987 15487
rect 1771 14640 1827 14649
rect 1851 14640 1907 14649
rect 1931 14640 1987 14649
rect 1771 14593 1796 14640
rect 1796 14593 1827 14640
rect 1851 14593 1864 14640
rect 1864 14593 1907 14640
rect 1931 14593 1932 14640
rect 1932 14593 1984 14640
rect 1984 14593 1987 14640
rect 1771 14516 1796 14563
rect 1796 14516 1827 14563
rect 1851 14516 1864 14563
rect 1864 14516 1907 14563
rect 1931 14516 1932 14563
rect 1932 14516 1984 14563
rect 1984 14516 1987 14563
rect 1771 14507 1827 14516
rect 1851 14507 1907 14516
rect 1931 14507 1987 14516
rect 1771 14444 1796 14477
rect 1796 14444 1827 14477
rect 1851 14444 1864 14477
rect 1864 14444 1907 14477
rect 1931 14444 1932 14477
rect 1932 14444 1984 14477
rect 1984 14444 1987 14477
rect 1189 14378 1245 14434
rect 1189 14298 1245 14354
rect 1771 14424 1827 14444
rect 1851 14424 1907 14444
rect 1931 14424 1987 14444
rect 1771 14421 1796 14424
rect 1796 14421 1827 14424
rect 1851 14421 1864 14424
rect 1864 14421 1907 14424
rect 1931 14421 1932 14424
rect 1932 14421 1984 14424
rect 1984 14421 1987 14424
rect 1771 14372 1796 14391
rect 1796 14372 1827 14391
rect 1851 14372 1864 14391
rect 1864 14372 1907 14391
rect 1931 14372 1932 14391
rect 1932 14372 1984 14391
rect 1984 14372 1987 14391
rect 1771 14351 1827 14372
rect 1851 14351 1907 14372
rect 1931 14351 1987 14372
rect 1771 14335 1796 14351
rect 1796 14335 1827 14351
rect 1851 14335 1864 14351
rect 1864 14335 1907 14351
rect 1931 14335 1932 14351
rect 1932 14335 1984 14351
rect 1984 14335 1987 14351
rect 1771 14299 1796 14305
rect 1796 14299 1827 14305
rect 1851 14299 1864 14305
rect 1864 14299 1907 14305
rect 1931 14299 1932 14305
rect 1932 14299 1984 14305
rect 1984 14299 1987 14305
rect 1771 14278 1827 14299
rect 1851 14278 1907 14299
rect 1931 14278 1987 14299
rect 1771 14249 1796 14278
rect 1796 14249 1827 14278
rect 1851 14249 1864 14278
rect 1864 14249 1907 14278
rect 1931 14249 1932 14278
rect 1932 14249 1984 14278
rect 1984 14249 1987 14278
rect 1771 14205 1827 14219
rect 1851 14205 1907 14219
rect 1931 14205 1987 14219
rect 1309 14117 1365 14173
rect 1309 14037 1365 14093
rect 1771 14163 1796 14205
rect 1796 14163 1827 14205
rect 1851 14163 1864 14205
rect 1864 14163 1907 14205
rect 1931 14163 1932 14205
rect 1932 14163 1984 14205
rect 1984 14163 1987 14205
rect 1771 14080 1796 14132
rect 1796 14080 1827 14132
rect 1851 14080 1864 14132
rect 1864 14080 1907 14132
rect 1931 14080 1932 14132
rect 1932 14080 1984 14132
rect 1984 14080 1987 14132
rect 1771 14076 1827 14080
rect 1851 14076 1907 14080
rect 1931 14076 1987 14080
rect 2794 14168 2850 14224
rect 2794 14088 2850 14144
rect 22106 14072 22162 14128
rect 22187 14072 22243 14128
rect 22268 14072 22324 14128
rect 22349 14072 22405 14128
rect 22430 14072 22486 14128
rect 22511 14072 22567 14128
rect 22592 14072 22648 14128
rect 22673 14072 22729 14128
rect 22753 14072 22809 14128
rect 22833 14072 22889 14128
rect 22913 14072 22969 14128
rect 23254 14065 23310 14121
rect 23392 14065 23448 14121
rect 22106 13970 22162 14026
rect 22187 13970 22243 14026
rect 22268 13970 22324 14026
rect 22349 13970 22405 14026
rect 22430 13970 22486 14026
rect 22511 13970 22567 14026
rect 22592 13970 22648 14026
rect 22673 13970 22729 14026
rect 22753 13970 22809 14026
rect 22833 13970 22889 14026
rect 22913 13970 22969 14026
rect 23254 13968 23310 14024
rect 23392 13968 23448 14024
rect 22106 13868 22162 13924
rect 22187 13868 22243 13924
rect 22268 13868 22324 13924
rect 22349 13868 22405 13924
rect 22430 13868 22486 13924
rect 22511 13868 22567 13924
rect 22592 13868 22648 13924
rect 22673 13868 22729 13924
rect 22753 13868 22809 13924
rect 22833 13868 22889 13924
rect 22913 13868 22969 13924
rect 23254 13870 23310 13926
rect 23392 13870 23448 13926
rect 22106 13766 22162 13822
rect 22187 13766 22243 13822
rect 22268 13766 22324 13822
rect 22349 13766 22405 13822
rect 22430 13766 22486 13822
rect 22511 13766 22567 13822
rect 22592 13766 22648 13822
rect 22673 13766 22729 13822
rect 22753 13766 22809 13822
rect 22833 13766 22889 13822
rect 22913 13766 22969 13822
rect 23254 13772 23310 13828
rect 23392 13772 23448 13828
rect 827 12856 883 12865
rect 949 12856 1005 12865
rect 827 12809 878 12856
rect 878 12809 883 12856
rect 949 12809 954 12856
rect 954 12809 1005 12856
rect 827 12781 883 12785
rect 949 12781 1005 12785
rect 827 12729 878 12781
rect 878 12729 883 12781
rect 949 12729 954 12781
rect 954 12729 1005 12781
rect 827 12653 878 12705
rect 878 12653 883 12705
rect 949 12653 954 12705
rect 954 12653 1005 12705
rect 827 12649 883 12653
rect 949 12649 1005 12653
rect 827 12577 878 12625
rect 878 12577 883 12625
rect 949 12577 954 12625
rect 954 12577 1005 12625
rect 23786 12661 23842 12717
rect 23868 12661 23924 12717
rect 23950 12661 24006 12717
rect 24031 12661 24087 12717
rect 24112 12661 24168 12717
rect 827 12569 883 12577
rect 949 12569 1005 12577
rect 15778 11531 15834 11587
rect 15858 11531 15914 11587
rect 3500 11463 3556 11519
rect 3645 11463 3701 11519
rect 3500 11383 3556 11439
rect 3645 11383 3701 11439
rect 20132 11440 20188 11496
rect 20213 11440 20269 11496
rect 20294 11440 20350 11496
rect 20374 11440 20430 11496
rect 20454 11440 20510 11496
rect 14445 11226 14501 11282
rect 14445 11146 14501 11202
rect 700 10920 756 10921
rect 700 10868 707 10920
rect 707 10868 756 10920
rect 700 10865 756 10868
rect 700 10804 707 10841
rect 707 10804 756 10841
rect 700 10785 756 10804
rect 1151 10757 1207 10765
rect 1151 10709 1153 10757
rect 1153 10709 1205 10757
rect 1205 10709 1207 10757
rect 1151 10641 1153 10685
rect 1153 10641 1205 10685
rect 1205 10641 1207 10685
rect 1151 10629 1207 10641
rect 10336 10647 10392 10648
rect 10336 10595 10388 10647
rect 10388 10595 10392 10647
rect 10336 10592 10392 10595
rect 10336 10531 10388 10568
rect 10388 10531 10392 10568
rect 10336 10512 10392 10531
rect 3318 10221 3374 10277
rect 3422 10221 3478 10277
rect 3526 10221 3582 10277
rect 3630 10221 3686 10277
rect 3318 10141 3374 10197
rect 3422 10141 3478 10197
rect 3526 10141 3582 10197
rect 3630 10141 3686 10197
rect 9879 10065 9935 10121
rect 10013 10065 10069 10121
rect 3318 9947 3374 10003
rect 3422 9947 3478 10003
rect 3526 9947 3582 10003
rect 3630 9947 3686 10003
rect 3318 9867 3374 9923
rect 3422 9867 3478 9923
rect 3526 9867 3582 9923
rect 3630 9867 3686 9923
rect 9879 9969 9935 10025
rect 10013 9969 10069 10025
rect 17884 10829 17940 10885
rect 18004 10829 18060 10885
rect 18123 10829 18179 10885
rect 17884 10703 17940 10759
rect 18004 10703 18060 10759
rect 18123 10703 18179 10759
rect 24599 10787 24655 10843
rect 24679 10787 24735 10843
rect 24759 10787 24815 10843
rect 24839 10787 24895 10843
rect 24599 10742 24655 10758
rect 24679 10742 24735 10758
rect 24759 10742 24815 10758
rect 24599 10702 24614 10742
rect 24614 10702 24655 10742
rect 24679 10702 24730 10742
rect 24730 10702 24735 10742
rect 24759 10702 24794 10742
rect 24794 10702 24815 10742
rect 24839 10702 24895 10758
rect 24599 10624 24614 10673
rect 24614 10624 24655 10673
rect 24679 10624 24730 10673
rect 24730 10624 24735 10673
rect 24759 10624 24794 10673
rect 24794 10624 24815 10673
rect 24599 10617 24655 10624
rect 24679 10617 24735 10624
rect 24759 10617 24815 10624
rect 24839 10617 24895 10673
rect 24599 10558 24614 10588
rect 24614 10558 24655 10588
rect 24679 10558 24730 10588
rect 24730 10558 24735 10588
rect 24759 10558 24794 10588
rect 24794 10558 24815 10588
rect 24599 10543 24655 10558
rect 24679 10543 24735 10558
rect 24759 10543 24815 10558
rect 24599 10532 24614 10543
rect 24614 10532 24655 10543
rect 24599 10491 24614 10502
rect 24614 10491 24655 10502
rect 24679 10532 24730 10543
rect 24730 10532 24735 10543
rect 24759 10532 24794 10543
rect 24794 10532 24815 10543
rect 24839 10532 24895 10588
rect 24679 10491 24730 10502
rect 24730 10491 24735 10502
rect 24759 10491 24794 10502
rect 24794 10491 24815 10502
rect 24599 10476 24655 10491
rect 24679 10476 24735 10491
rect 24759 10476 24815 10491
rect 24599 10446 24614 10476
rect 24614 10446 24655 10476
rect 24679 10446 24730 10476
rect 24730 10446 24735 10476
rect 24759 10446 24794 10476
rect 24794 10446 24815 10476
rect 24839 10446 24895 10502
rect 24599 10409 24655 10416
rect 24679 10409 24735 10416
rect 24759 10409 24815 10416
rect 24599 10360 24614 10409
rect 24614 10360 24655 10409
rect 24679 10360 24730 10409
rect 24730 10360 24735 10409
rect 24759 10360 24794 10409
rect 24794 10360 24815 10409
rect 24839 10360 24895 10416
rect 15579 10236 15635 10292
rect 15659 10236 15715 10292
rect 9879 9873 9935 9929
rect 10013 9873 10069 9929
rect 13223 9948 13279 10004
rect 13223 9868 13279 9924
rect 9879 9777 9935 9833
rect 10013 9777 10069 9833
rect 25285 9325 25341 9381
rect 25285 9245 25341 9301
rect 27243 8987 27299 9043
rect 27323 8987 27379 9043
rect 27403 8987 27459 9043
rect 27483 8987 27539 9043
rect 27243 8898 27299 8954
rect 27323 8898 27379 8954
rect 27403 8898 27459 8954
rect 27483 8898 27539 8954
rect 27243 8809 27299 8865
rect 27323 8809 27379 8865
rect 27403 8809 27459 8865
rect 27483 8809 27539 8865
rect 27243 8720 27299 8776
rect 27323 8720 27379 8776
rect 27403 8720 27459 8776
rect 27483 8720 27539 8776
rect 27243 8630 27299 8686
rect 27323 8630 27379 8686
rect 27403 8630 27459 8686
rect 27483 8630 27539 8686
rect 2794 8082 2850 8138
rect 2794 8002 2850 8058
rect 22394 8076 22443 8123
rect 22443 8076 22450 8123
rect 22476 8076 22515 8123
rect 22515 8076 22532 8123
rect 22558 8076 22587 8123
rect 22587 8076 22606 8123
rect 22606 8076 22614 8123
rect 22640 8076 22658 8123
rect 22658 8076 22677 8123
rect 22677 8076 22696 8123
rect 22721 8076 22729 8123
rect 22729 8076 22748 8123
rect 22748 8076 22777 8123
rect 22802 8076 22819 8123
rect 22819 8076 22858 8123
rect 22883 8076 22890 8123
rect 22890 8076 22939 8123
rect 22394 8067 22450 8076
rect 22476 8067 22532 8076
rect 22558 8067 22614 8076
rect 22640 8067 22696 8076
rect 22721 8067 22777 8076
rect 22802 8067 22858 8076
rect 22883 8067 22939 8076
rect 22394 7980 22450 7999
rect 22476 7980 22532 7999
rect 22558 7980 22614 7999
rect 22640 7980 22696 7999
rect 22721 7980 22777 7999
rect 22802 7980 22858 7999
rect 22883 7980 22939 7999
rect 13312 7877 13368 7933
rect 22394 7943 22443 7980
rect 22443 7943 22450 7980
rect 22476 7943 22515 7980
rect 22515 7943 22532 7980
rect 22558 7943 22587 7980
rect 22587 7943 22606 7980
rect 22606 7943 22614 7980
rect 22640 7943 22658 7980
rect 22658 7943 22677 7980
rect 22677 7943 22696 7980
rect 22721 7943 22729 7980
rect 22729 7943 22748 7980
rect 22748 7943 22777 7980
rect 22802 7943 22819 7980
rect 22819 7943 22858 7980
rect 22883 7943 22890 7980
rect 22890 7943 22939 7980
rect 13312 7797 13368 7853
rect 14405 7496 14461 7552
rect 13282 7405 13338 7461
rect 13362 7405 13418 7461
rect 14405 7416 14461 7472
rect 3813 7087 3821 7139
rect 3821 7087 3869 7139
rect 3893 7087 3937 7139
rect 3937 7087 3949 7139
rect 3813 7083 3869 7087
rect 3893 7083 3949 7087
rect 1151 6931 1207 6987
rect 1755 6931 1811 6987
rect 1151 6851 1207 6907
rect 1755 6851 1811 6907
rect 15818 6909 15874 6965
rect 2387 6834 2443 6890
rect 2467 6834 2523 6890
rect 3813 6834 3869 6890
rect 3893 6834 3949 6890
rect 15818 6829 15874 6885
rect 26164 6821 26220 6877
rect 5216 6701 5272 6757
rect 5307 6701 5363 6757
rect 5397 6701 5453 6757
rect 5487 6701 5543 6757
rect 26164 6741 26220 6797
rect 5216 6563 5272 6619
rect 5307 6563 5363 6619
rect 5397 6563 5453 6619
rect 5487 6563 5543 6619
rect 1548 6464 1604 6520
rect 1628 6464 1684 6520
rect 2934 6402 2982 6403
rect 2982 6402 2990 6403
rect 2934 6390 2990 6402
rect 1398 6320 1454 6376
rect 2257 6320 2313 6376
rect 2934 6347 2982 6390
rect 2982 6347 2990 6390
rect 3058 6347 3114 6403
rect 3182 6347 3238 6403
rect 4147 6343 4203 6399
rect 4227 6343 4283 6399
rect 4434 6394 4490 6450
rect 4514 6394 4570 6450
rect 1398 6240 1454 6296
rect 2257 6240 2313 6296
rect 15640 6224 15641 6270
rect 15641 6224 15693 6270
rect 15693 6224 15696 6270
rect 23986 6267 24042 6323
rect 15640 6214 15696 6224
rect 4432 6110 4488 6166
rect 4432 6030 4488 6086
rect 5949 6143 5998 6195
rect 5998 6143 6005 6195
rect 6037 6143 6065 6195
rect 6065 6143 6080 6195
rect 6080 6143 6093 6195
rect 6125 6143 6132 6195
rect 6132 6143 6147 6195
rect 6147 6143 6181 6195
rect 6213 6143 6214 6195
rect 6214 6143 6266 6195
rect 6266 6143 6269 6195
rect 6301 6143 6333 6195
rect 6333 6143 6348 6195
rect 6348 6143 6357 6195
rect 6388 6143 6400 6195
rect 6400 6143 6415 6195
rect 6415 6143 6444 6195
rect 6475 6143 6482 6195
rect 6482 6143 6531 6195
rect 12234 6143 12283 6195
rect 12283 6143 12290 6195
rect 12322 6143 12350 6195
rect 12350 6143 12365 6195
rect 12365 6143 12378 6195
rect 12410 6143 12417 6195
rect 12417 6143 12432 6195
rect 12432 6143 12466 6195
rect 12498 6143 12499 6195
rect 12499 6143 12551 6195
rect 12551 6143 12554 6195
rect 12586 6143 12618 6195
rect 12618 6143 12633 6195
rect 12633 6143 12642 6195
rect 12673 6143 12685 6195
rect 12685 6143 12700 6195
rect 12700 6143 12729 6195
rect 12760 6143 12767 6195
rect 12767 6143 12816 6195
rect 5949 6139 6005 6143
rect 6037 6139 6093 6143
rect 6125 6139 6181 6143
rect 6213 6139 6269 6143
rect 6301 6139 6357 6143
rect 6388 6139 6444 6143
rect 6475 6139 6531 6143
rect 12234 6139 12290 6143
rect 12322 6139 12378 6143
rect 12410 6139 12466 6143
rect 12498 6139 12554 6143
rect 12586 6139 12642 6143
rect 12673 6139 12729 6143
rect 12760 6139 12816 6143
rect 15640 6134 15696 6190
rect 16079 6143 16128 6195
rect 16128 6143 16135 6195
rect 16165 6143 16194 6195
rect 16194 6143 16208 6195
rect 16208 6143 16221 6195
rect 16251 6143 16260 6195
rect 16260 6143 16274 6195
rect 16274 6143 16307 6195
rect 16337 6143 16339 6195
rect 16339 6143 16391 6195
rect 16391 6143 16393 6195
rect 16422 6143 16456 6195
rect 16456 6143 16469 6195
rect 16469 6143 16478 6195
rect 16507 6143 16521 6195
rect 16521 6143 16534 6195
rect 16534 6143 16563 6195
rect 16592 6143 16599 6195
rect 16599 6143 16648 6195
rect 16079 6139 16135 6143
rect 16165 6139 16221 6143
rect 16251 6139 16307 6143
rect 16337 6139 16393 6143
rect 16422 6139 16478 6143
rect 16507 6139 16563 6143
rect 16592 6139 16648 6143
rect 5949 6047 6005 6051
rect 6037 6047 6093 6051
rect 6125 6047 6181 6051
rect 6213 6047 6269 6051
rect 6301 6047 6357 6051
rect 6388 6047 6444 6051
rect 6475 6047 6531 6051
rect 12234 6047 12290 6051
rect 12322 6047 12378 6051
rect 12410 6047 12466 6051
rect 12498 6047 12554 6051
rect 12586 6047 12642 6051
rect 12673 6047 12729 6051
rect 12760 6047 12816 6051
rect 5949 5995 5998 6047
rect 5998 5995 6005 6047
rect 6037 5995 6065 6047
rect 6065 5995 6080 6047
rect 6080 5995 6093 6047
rect 6125 5995 6132 6047
rect 6132 5995 6147 6047
rect 6147 5995 6181 6047
rect 6213 5995 6214 6047
rect 6214 5995 6266 6047
rect 6266 5995 6269 6047
rect 6301 5995 6333 6047
rect 6333 5995 6348 6047
rect 6348 5995 6357 6047
rect 6388 5995 6400 6047
rect 6400 5995 6415 6047
rect 6415 5995 6444 6047
rect 6475 5995 6482 6047
rect 6482 5995 6531 6047
rect 12234 5995 12283 6047
rect 12283 5995 12290 6047
rect 12322 5995 12350 6047
rect 12350 5995 12365 6047
rect 12365 5995 12378 6047
rect 12410 5995 12417 6047
rect 12417 5995 12432 6047
rect 12432 5995 12466 6047
rect 12498 5995 12499 6047
rect 12499 5995 12551 6047
rect 12551 5995 12554 6047
rect 12586 5995 12618 6047
rect 12618 5995 12633 6047
rect 12633 5995 12642 6047
rect 12673 5995 12685 6047
rect 12685 5995 12700 6047
rect 12700 5995 12729 6047
rect 12760 5995 12767 6047
rect 12767 5995 12816 6047
rect 16079 6047 16135 6051
rect 16165 6047 16221 6051
rect 16251 6047 16307 6051
rect 16337 6047 16393 6051
rect 16422 6047 16478 6051
rect 16507 6047 16563 6051
rect 16592 6047 16648 6051
rect 16079 5995 16128 6047
rect 16128 5995 16135 6047
rect 16165 5995 16194 6047
rect 16194 5995 16208 6047
rect 16208 5995 16221 6047
rect 16251 5995 16260 6047
rect 16260 5995 16274 6047
rect 16274 5995 16307 6047
rect 16337 5995 16339 6047
rect 16339 5995 16391 6047
rect 16391 5995 16393 6047
rect 16422 5995 16456 6047
rect 16456 5995 16469 6047
rect 16469 5995 16478 6047
rect 16507 5995 16521 6047
rect 16521 5995 16534 6047
rect 16534 5995 16563 6047
rect 16592 5995 16599 6047
rect 16599 5995 16648 6047
rect 20301 6143 20350 6195
rect 20350 6143 20357 6195
rect 20389 6143 20417 6195
rect 20417 6143 20432 6195
rect 20432 6143 20445 6195
rect 20477 6143 20484 6195
rect 20484 6143 20499 6195
rect 20499 6143 20533 6195
rect 20565 6143 20566 6195
rect 20566 6143 20618 6195
rect 20618 6143 20621 6195
rect 20653 6143 20685 6195
rect 20685 6143 20700 6195
rect 20700 6143 20709 6195
rect 20740 6143 20752 6195
rect 20752 6143 20767 6195
rect 20767 6143 20796 6195
rect 20827 6143 20834 6195
rect 20834 6143 20883 6195
rect 23986 6187 24042 6243
rect 20301 6139 20357 6143
rect 20389 6139 20445 6143
rect 20477 6139 20533 6143
rect 20565 6139 20621 6143
rect 20653 6139 20709 6143
rect 20740 6139 20796 6143
rect 20827 6139 20883 6143
rect 20301 6047 20357 6051
rect 20389 6047 20445 6051
rect 20477 6047 20533 6051
rect 20565 6047 20621 6051
rect 20653 6047 20709 6051
rect 20740 6047 20796 6051
rect 20827 6047 20883 6051
rect 20301 5995 20350 6047
rect 20350 5995 20357 6047
rect 20389 5995 20417 6047
rect 20417 5995 20432 6047
rect 20432 5995 20445 6047
rect 20477 5995 20484 6047
rect 20484 5995 20499 6047
rect 20499 5995 20533 6047
rect 20565 5995 20566 6047
rect 20566 5995 20618 6047
rect 20618 5995 20621 6047
rect 20653 5995 20685 6047
rect 20685 5995 20700 6047
rect 20700 5995 20709 6047
rect 20740 5995 20752 6047
rect 20752 5995 20767 6047
rect 20767 5995 20796 6047
rect 20827 5995 20834 6047
rect 20834 5995 20883 6047
rect 1427 3870 1483 3926
rect 1427 3790 1483 3846
rect 7445 5496 7501 5497
rect 7533 5496 7589 5497
rect 7621 5496 7677 5497
rect 7709 5496 7765 5497
rect 7797 5496 7853 5497
rect 7884 5496 7940 5497
rect 7971 5496 8027 5497
rect 7445 5444 7494 5496
rect 7494 5444 7501 5496
rect 7533 5444 7561 5496
rect 7561 5444 7576 5496
rect 7576 5444 7589 5496
rect 7621 5444 7628 5496
rect 7628 5444 7643 5496
rect 7643 5444 7677 5496
rect 7709 5444 7710 5496
rect 7710 5444 7762 5496
rect 7762 5444 7765 5496
rect 7797 5444 7829 5496
rect 7829 5444 7844 5496
rect 7844 5444 7853 5496
rect 7884 5444 7896 5496
rect 7896 5444 7911 5496
rect 7911 5444 7940 5496
rect 7971 5444 7978 5496
rect 7978 5444 8027 5496
rect 7445 5441 7501 5444
rect 7533 5441 7589 5444
rect 7621 5441 7677 5444
rect 7709 5441 7765 5444
rect 7797 5441 7853 5444
rect 7884 5441 7940 5444
rect 7971 5441 8027 5444
rect 7445 5352 7501 5355
rect 7533 5352 7589 5355
rect 7621 5352 7677 5355
rect 7709 5352 7765 5355
rect 7797 5352 7853 5355
rect 7884 5352 7940 5355
rect 7971 5352 8027 5355
rect 7445 5300 7494 5352
rect 7494 5300 7501 5352
rect 7533 5300 7561 5352
rect 7561 5300 7576 5352
rect 7576 5300 7589 5352
rect 7621 5300 7628 5352
rect 7628 5300 7643 5352
rect 7643 5300 7677 5352
rect 7709 5300 7710 5352
rect 7710 5300 7762 5352
rect 7762 5300 7765 5352
rect 7797 5300 7829 5352
rect 7829 5300 7844 5352
rect 7844 5300 7853 5352
rect 7884 5300 7896 5352
rect 7896 5300 7911 5352
rect 7911 5300 7940 5352
rect 7971 5300 7978 5352
rect 7978 5300 8027 5352
rect 7445 5299 7501 5300
rect 7533 5299 7589 5300
rect 7621 5299 7677 5300
rect 7709 5299 7765 5300
rect 7797 5299 7853 5300
rect 7884 5299 7940 5300
rect 7971 5299 8027 5300
rect 11514 5496 11570 5497
rect 11602 5496 11658 5497
rect 11690 5496 11746 5497
rect 11778 5496 11834 5497
rect 11866 5496 11922 5497
rect 11953 5496 12009 5497
rect 12040 5496 12096 5497
rect 11514 5444 11563 5496
rect 11563 5444 11570 5496
rect 11602 5444 11630 5496
rect 11630 5444 11645 5496
rect 11645 5444 11658 5496
rect 11690 5444 11697 5496
rect 11697 5444 11712 5496
rect 11712 5444 11746 5496
rect 11778 5444 11779 5496
rect 11779 5444 11831 5496
rect 11831 5444 11834 5496
rect 11866 5444 11898 5496
rect 11898 5444 11913 5496
rect 11913 5444 11922 5496
rect 11953 5444 11965 5496
rect 11965 5444 11980 5496
rect 11980 5444 12009 5496
rect 12040 5444 12047 5496
rect 12047 5444 12096 5496
rect 11514 5441 11570 5444
rect 11602 5441 11658 5444
rect 11690 5441 11746 5444
rect 11778 5441 11834 5444
rect 11866 5441 11922 5444
rect 11953 5441 12009 5444
rect 12040 5441 12096 5444
rect 11514 5352 11570 5355
rect 11602 5352 11658 5355
rect 11690 5352 11746 5355
rect 11778 5352 11834 5355
rect 11866 5352 11922 5355
rect 11953 5352 12009 5355
rect 12040 5352 12096 5355
rect 11514 5300 11563 5352
rect 11563 5300 11570 5352
rect 11602 5300 11630 5352
rect 11630 5300 11645 5352
rect 11645 5300 11658 5352
rect 11690 5300 11697 5352
rect 11697 5300 11712 5352
rect 11712 5300 11746 5352
rect 11778 5300 11779 5352
rect 11779 5300 11831 5352
rect 11831 5300 11834 5352
rect 11866 5300 11898 5352
rect 11898 5300 11913 5352
rect 11913 5300 11922 5352
rect 11953 5300 11965 5352
rect 11965 5300 11980 5352
rect 11980 5300 12009 5352
rect 12040 5300 12047 5352
rect 12047 5300 12096 5352
rect 11514 5299 11570 5300
rect 11602 5299 11658 5300
rect 11690 5299 11746 5300
rect 11778 5299 11834 5300
rect 11866 5299 11922 5300
rect 11953 5299 12009 5300
rect 12040 5299 12096 5300
rect 14536 5496 14592 5497
rect 14617 5496 14673 5497
rect 14698 5496 14754 5497
rect 14779 5496 14835 5497
rect 14860 5496 14916 5497
rect 14941 5496 14997 5497
rect 14536 5444 14585 5496
rect 14585 5444 14592 5496
rect 14617 5444 14655 5496
rect 14655 5444 14672 5496
rect 14672 5444 14673 5496
rect 14698 5444 14724 5496
rect 14724 5444 14741 5496
rect 14741 5444 14754 5496
rect 14779 5444 14793 5496
rect 14793 5444 14810 5496
rect 14810 5444 14835 5496
rect 14860 5444 14862 5496
rect 14862 5444 14879 5496
rect 14879 5444 14916 5496
rect 14941 5444 14948 5496
rect 14948 5444 14997 5496
rect 14536 5441 14592 5444
rect 14617 5441 14673 5444
rect 14698 5441 14754 5444
rect 14779 5441 14835 5444
rect 14860 5441 14916 5444
rect 14941 5441 14997 5444
rect 14536 5352 14592 5355
rect 14617 5352 14673 5355
rect 14698 5352 14754 5355
rect 14779 5352 14835 5355
rect 14860 5352 14916 5355
rect 14941 5352 14997 5355
rect 14536 5300 14585 5352
rect 14585 5300 14592 5352
rect 14617 5300 14655 5352
rect 14655 5300 14672 5352
rect 14672 5300 14673 5352
rect 14698 5300 14724 5352
rect 14724 5300 14741 5352
rect 14741 5300 14754 5352
rect 14779 5300 14793 5352
rect 14793 5300 14810 5352
rect 14810 5300 14835 5352
rect 14860 5300 14862 5352
rect 14862 5300 14879 5352
rect 14879 5300 14916 5352
rect 14941 5300 14948 5352
rect 14948 5300 14997 5352
rect 14536 5299 14592 5300
rect 14617 5299 14673 5300
rect 14698 5299 14754 5300
rect 14779 5299 14835 5300
rect 14860 5299 14916 5300
rect 14941 5299 14997 5300
rect 16899 4544 16955 4600
rect 17012 4544 17068 4600
rect 17125 4544 17181 4600
rect 16899 4485 16955 4520
rect 17012 4485 17068 4520
rect 17125 4485 17181 4520
rect 16899 4464 16948 4485
rect 16948 4464 16955 4485
rect 17012 4464 17027 4485
rect 17027 4464 17053 4485
rect 17053 4464 17068 4485
rect 17125 4464 17131 4485
rect 17131 4464 17181 4485
rect 16899 4433 16948 4440
rect 16948 4433 16955 4440
rect 17012 4433 17027 4440
rect 17027 4433 17053 4440
rect 17053 4433 17068 4440
rect 17125 4433 17131 4440
rect 17131 4433 17181 4440
rect 16899 4384 16955 4433
rect 17012 4384 17068 4433
rect 17125 4384 17181 4433
rect 5476 4276 5532 4332
rect 5476 4196 5532 4252
rect 9076 4276 9132 4332
rect 9076 4196 9132 4252
rect 9246 4276 9302 4332
rect 9246 4196 9302 4252
rect 13222 4276 13278 4332
rect 13222 4196 13278 4252
rect 13392 4276 13448 4332
rect 13392 4196 13448 4252
rect 16899 4309 16948 4360
rect 16948 4309 16955 4360
rect 17012 4309 17027 4360
rect 17027 4309 17053 4360
rect 17053 4309 17068 4360
rect 17125 4309 17131 4360
rect 17131 4309 17181 4360
rect 16899 4304 16955 4309
rect 17012 4304 17068 4309
rect 17125 4304 17181 4309
rect 16899 4224 16955 4280
rect 17012 4224 17068 4280
rect 17125 4224 17181 4280
rect 17368 4276 17424 4332
rect 17368 4196 17424 4252
rect 17538 4276 17594 4332
rect 17538 4196 17594 4252
rect 21516 4276 21572 4332
rect 21516 4196 21572 4252
rect 21680 4276 21736 4332
rect 21680 4196 21736 4252
rect 25664 4276 25720 4332
rect 701 3322 757 3344
rect 701 3288 703 3322
rect 703 3288 755 3322
rect 755 3288 757 3322
rect 701 3258 757 3264
rect 701 3208 703 3258
rect 703 3208 755 3258
rect 755 3208 757 3258
rect 3347 3445 3351 3494
rect 3351 3445 3403 3494
rect 3403 3445 3415 3494
rect 3415 3445 3467 3494
rect 3467 3445 3479 3494
rect 3479 3445 3531 3494
rect 3531 3445 3543 3494
rect 3543 3445 3595 3494
rect 3595 3445 3643 3494
rect 3347 3432 3643 3445
rect 3347 3380 3351 3432
rect 3351 3380 3403 3432
rect 3403 3380 3415 3432
rect 3415 3380 3467 3432
rect 3467 3380 3479 3432
rect 3479 3380 3531 3432
rect 3531 3380 3543 3432
rect 3543 3380 3595 3432
rect 3595 3380 3643 3432
rect 3347 3367 3643 3380
rect 3347 3315 3351 3367
rect 3351 3315 3403 3367
rect 3403 3315 3415 3367
rect 3415 3315 3467 3367
rect 3467 3315 3479 3367
rect 3479 3315 3531 3367
rect 3531 3315 3543 3367
rect 3543 3315 3595 3367
rect 3595 3315 3643 3367
rect 3347 3302 3643 3315
rect 3347 3250 3351 3302
rect 3351 3250 3403 3302
rect 3403 3250 3415 3302
rect 3415 3250 3467 3302
rect 3467 3250 3479 3302
rect 3479 3250 3531 3302
rect 3531 3250 3543 3302
rect 3543 3250 3595 3302
rect 3595 3250 3643 3302
rect 3347 3237 3643 3250
rect 3347 3198 3351 3237
rect 3351 3198 3403 3237
rect 3403 3198 3415 3237
rect 3415 3198 3467 3237
rect 3467 3198 3479 3237
rect 3479 3198 3531 3237
rect 3531 3198 3543 3237
rect 3543 3198 3595 3237
rect 3595 3198 3643 3237
rect 1163 3083 1219 3139
rect 1163 3056 1219 3059
rect 1163 3004 1165 3056
rect 1165 3004 1217 3056
rect 1217 3004 1219 3056
rect 1758 3140 1814 3162
rect 1758 3106 1760 3140
rect 1760 3106 1812 3140
rect 1812 3106 1814 3140
rect 3347 3172 3403 3173
rect 3427 3172 3483 3173
rect 3507 3172 3563 3173
rect 3587 3172 3643 3173
rect 3347 3120 3351 3172
rect 3351 3120 3403 3172
rect 3427 3120 3467 3172
rect 3467 3120 3479 3172
rect 3479 3120 3483 3172
rect 3507 3120 3531 3172
rect 3531 3120 3543 3172
rect 3543 3120 3563 3172
rect 3587 3120 3595 3172
rect 3595 3120 3643 3172
rect 3347 3117 3403 3120
rect 3427 3117 3483 3120
rect 3507 3117 3563 3120
rect 3587 3117 3643 3120
rect 1758 3076 1814 3082
rect 1758 3026 1760 3076
rect 1760 3026 1812 3076
rect 1812 3026 1814 3076
rect 3347 3054 3351 3092
rect 3351 3054 3403 3092
rect 3427 3054 3467 3092
rect 3467 3054 3479 3092
rect 3479 3054 3483 3092
rect 3507 3054 3531 3092
rect 3531 3054 3543 3092
rect 3543 3054 3563 3092
rect 3587 3054 3595 3092
rect 3595 3054 3643 3092
rect 3347 3040 3403 3054
rect 3427 3040 3483 3054
rect 3507 3040 3563 3054
rect 3587 3040 3643 3054
rect 3347 3036 3351 3040
rect 3351 3036 3403 3040
rect 1163 3003 1219 3004
rect 3347 2988 3351 3011
rect 3351 2988 3403 3011
rect 3427 3036 3467 3040
rect 3467 3036 3479 3040
rect 3479 3036 3483 3040
rect 3507 3036 3531 3040
rect 3531 3036 3543 3040
rect 3543 3036 3563 3040
rect 3587 3036 3595 3040
rect 3595 3036 3643 3040
rect 7445 3228 7501 3284
rect 7533 3228 7589 3284
rect 7621 3228 7677 3284
rect 7709 3228 7765 3284
rect 7797 3228 7853 3284
rect 7884 3228 7940 3284
rect 7971 3228 8027 3284
rect 7445 3088 7501 3144
rect 7533 3088 7589 3144
rect 7621 3088 7677 3144
rect 7709 3088 7765 3144
rect 7797 3088 7853 3144
rect 7884 3088 7940 3144
rect 7971 3088 8027 3144
rect 11514 3228 11570 3284
rect 11602 3228 11658 3284
rect 11690 3228 11746 3284
rect 11778 3228 11834 3284
rect 11866 3228 11922 3284
rect 11953 3228 12009 3284
rect 12040 3228 12096 3284
rect 11514 3088 11570 3144
rect 11602 3088 11658 3144
rect 11690 3088 11746 3144
rect 11778 3088 11834 3144
rect 11866 3088 11922 3144
rect 11953 3088 12009 3144
rect 12040 3088 12096 3144
rect 14536 3228 14592 3284
rect 14624 3228 14680 3284
rect 14712 3228 14768 3284
rect 14800 3228 14856 3284
rect 14888 3228 14944 3284
rect 14975 3228 15031 3284
rect 15062 3228 15118 3284
rect 14536 3088 14592 3144
rect 14624 3088 14680 3144
rect 14712 3088 14768 3144
rect 14800 3088 14856 3144
rect 14888 3088 14944 3144
rect 14975 3088 15031 3144
rect 15062 3088 15118 3144
rect 18269 3223 18325 3279
rect 18368 3223 18424 3279
rect 18466 3223 18522 3279
rect 18269 3093 18325 3149
rect 18368 3093 18424 3149
rect 18466 3093 18522 3149
rect 3427 2988 3467 3011
rect 3467 2988 3479 3011
rect 3479 2988 3483 3011
rect 3507 2988 3531 3011
rect 3531 2988 3543 3011
rect 3543 2988 3563 3011
rect 3587 2988 3595 3011
rect 3595 2988 3643 3011
rect 3347 2974 3403 2988
rect 3427 2974 3483 2988
rect 3507 2974 3563 2988
rect 3587 2974 3643 2988
rect 3347 2955 3351 2974
rect 3351 2955 3403 2974
rect 1163 2839 1171 2886
rect 1171 2839 1219 2886
rect 1163 2830 1219 2839
rect 1163 2750 1219 2806
rect 3347 2922 3351 2930
rect 3351 2922 3403 2930
rect 3427 2955 3467 2974
rect 3467 2955 3479 2974
rect 3479 2955 3483 2974
rect 3507 2955 3531 2974
rect 3531 2955 3543 2974
rect 3543 2955 3563 2974
rect 3587 2955 3595 2974
rect 3595 2955 3643 2974
rect 3427 2922 3467 2930
rect 3467 2922 3479 2930
rect 3479 2922 3483 2930
rect 3507 2922 3531 2930
rect 3531 2922 3543 2930
rect 3543 2922 3563 2930
rect 3587 2922 3595 2930
rect 3595 2922 3643 2930
rect 3347 2908 3403 2922
rect 3427 2908 3483 2922
rect 3507 2908 3563 2922
rect 3587 2908 3643 2922
rect 3347 2874 3351 2908
rect 3351 2874 3403 2908
rect 3427 2874 3467 2908
rect 3467 2874 3479 2908
rect 3479 2874 3483 2908
rect 3507 2874 3531 2908
rect 3531 2874 3543 2908
rect 3543 2874 3563 2908
rect 3587 2874 3595 2908
rect 3595 2874 3643 2908
rect 3347 2842 3403 2849
rect 3427 2842 3483 2849
rect 3507 2842 3563 2849
rect 3587 2842 3643 2849
rect 3347 2793 3351 2842
rect 3351 2793 3403 2842
rect 3427 2793 3467 2842
rect 3467 2793 3479 2842
rect 3479 2793 3483 2842
rect 3507 2793 3531 2842
rect 3531 2793 3543 2842
rect 3543 2793 3563 2842
rect 3587 2793 3595 2842
rect 3595 2793 3643 2842
rect 4081 2990 4137 3046
rect 4081 2910 4137 2966
rect 4081 2829 4137 2885
rect 4081 2748 4137 2804
rect 4081 2667 4137 2723
rect 1190 2574 1246 2630
rect 1190 2494 1246 2550
rect 4081 2586 4137 2642
rect 25285 4145 25341 4201
rect 25664 4196 25720 4252
rect 25826 4276 25882 4332
rect 25826 4196 25882 4252
rect 25285 4065 25341 4121
rect 26164 3840 26220 3862
rect 26164 3806 26191 3840
rect 26191 3806 26203 3840
rect 26203 3806 26220 3840
rect 26671 3797 26727 3853
rect 26164 3726 26220 3782
rect 26671 3760 26727 3773
rect 26671 3717 26721 3760
rect 26721 3717 26727 3760
rect 26797 3717 26853 3773
rect 26797 3680 26853 3693
rect 26797 3637 26847 3680
rect 26847 3637 26853 3680
rect 26923 3637 26979 3693
rect 26293 3557 26349 3613
rect 26923 3600 26979 3613
rect 26923 3557 26950 3600
rect 26950 3557 26962 3600
rect 26962 3557 26979 3600
rect 26293 3520 26349 3533
rect 26293 3477 26343 3520
rect 26343 3477 26349 3520
rect 26419 3477 26475 3533
rect 26419 3440 26475 3453
rect 26419 3397 26469 3440
rect 26469 3397 26475 3440
rect 26545 3397 26601 3453
rect 26545 3360 26601 3373
rect 26545 3317 26572 3360
rect 26572 3317 26584 3360
rect 26584 3317 26601 3360
rect 4081 2505 4137 2561
rect 4081 2424 4137 2480
rect 4081 2343 4137 2399
rect 4081 2262 4137 2318
rect 23251 2059 23307 2060
rect 23393 2059 23449 2060
rect 23251 2007 23254 2059
rect 23254 2007 23306 2059
rect 23306 2007 23307 2059
rect 23393 2007 23394 2059
rect 23394 2007 23446 2059
rect 23446 2007 23449 2059
rect 23251 2004 23307 2007
rect 23393 2004 23449 2007
rect 23251 1937 23254 1968
rect 23254 1937 23306 1968
rect 23306 1937 23307 1968
rect 23393 1937 23394 1968
rect 23394 1937 23446 1968
rect 23446 1937 23449 1968
rect 23251 1919 23307 1937
rect 23393 1919 23449 1937
rect 23251 1912 23254 1919
rect 23254 1912 23306 1919
rect 23306 1912 23307 1919
rect 23251 1867 23254 1876
rect 23254 1867 23306 1876
rect 23306 1867 23307 1876
rect 23393 1912 23394 1919
rect 23394 1912 23446 1919
rect 23446 1912 23449 1919
rect 23393 1867 23394 1876
rect 23394 1867 23446 1876
rect 23446 1867 23449 1876
rect 23251 1849 23307 1867
rect 23393 1849 23449 1867
rect 1964 1783 1986 1832
rect 1986 1783 1998 1832
rect 1998 1783 2020 1832
rect 1964 1776 2020 1783
rect 1759 1705 1815 1719
rect 1759 1663 1761 1705
rect 1761 1663 1813 1705
rect 1813 1663 1815 1705
rect 1759 1589 1761 1639
rect 1761 1589 1813 1639
rect 1813 1589 1815 1639
rect 1759 1583 1815 1589
rect 1964 1718 1986 1748
rect 1986 1718 1998 1748
rect 1998 1718 2020 1748
rect 23251 1820 23254 1849
rect 23254 1820 23306 1849
rect 23306 1820 23307 1849
rect 23393 1820 23394 1849
rect 23394 1820 23446 1849
rect 23446 1820 23449 1849
rect 23251 1778 23307 1783
rect 23393 1778 23449 1783
rect 23251 1727 23254 1778
rect 23254 1727 23306 1778
rect 23306 1727 23307 1778
rect 23393 1727 23394 1778
rect 23394 1727 23446 1778
rect 23446 1727 23449 1778
rect 1964 1705 2020 1718
rect 1964 1692 1986 1705
rect 1986 1692 1998 1705
rect 1998 1692 2020 1705
rect 1964 1653 1986 1663
rect 1986 1653 1998 1663
rect 1998 1653 2020 1663
rect 1964 1640 2020 1653
rect 1964 1607 1986 1640
rect 1986 1607 1998 1640
rect 1998 1607 2020 1640
rect 1964 1575 2020 1578
rect 1964 1523 1986 1575
rect 1986 1523 1998 1575
rect 1998 1523 2020 1575
rect 1964 1522 2020 1523
rect 1964 1458 1986 1493
rect 1986 1458 1998 1493
rect 1998 1458 2020 1493
rect 1964 1445 2020 1458
rect 1964 1437 1986 1445
rect 1986 1437 1998 1445
rect 1998 1437 2020 1445
rect 1964 1393 1986 1408
rect 1986 1393 1998 1408
rect 1998 1393 2020 1408
rect 1964 1380 2020 1393
rect 1964 1352 1986 1380
rect 1986 1352 1998 1380
rect 1998 1352 2020 1380
rect 1964 1315 2020 1323
rect 1964 1267 1986 1315
rect 1986 1267 1998 1315
rect 1998 1267 2020 1315
rect 1964 1198 1986 1238
rect 1986 1198 1998 1238
rect 1998 1198 2020 1238
rect 1964 1185 2020 1198
rect 1964 1182 1986 1185
rect 1986 1182 1998 1185
rect 1998 1182 2020 1185
rect 1964 1133 1986 1153
rect 1986 1133 1998 1153
rect 1998 1133 2020 1153
rect 1964 1120 2020 1133
rect 1964 1097 1986 1120
rect 1986 1097 1998 1120
rect 1998 1097 2020 1120
rect 23524 1182 23580 1238
rect 23650 1182 23706 1238
rect 23524 1088 23580 1144
rect 23650 1088 23706 1144
rect 1964 1055 2020 1068
rect 1964 1012 1986 1055
rect 1986 1012 1998 1055
rect 1998 1012 2020 1055
rect 1964 938 1986 983
rect 1986 938 1998 983
rect 1998 938 2020 983
rect 8812 977 8868 1033
rect 8892 977 8948 1033
rect 1964 927 2020 938
rect 1964 873 1986 898
rect 1986 873 1998 898
rect 1998 873 2020 898
rect 1964 860 2020 873
rect 1964 842 1986 860
rect 1986 842 1998 860
rect 1998 842 2020 860
rect 1964 808 1986 813
rect 1986 808 1998 813
rect 1998 808 2020 813
rect 1964 795 2020 808
rect 1964 757 1986 795
rect 1986 757 1998 795
rect 1998 757 2020 795
rect 1964 678 1986 728
rect 1986 678 1998 728
rect 1998 678 2020 728
rect 1964 672 2020 678
rect 1964 612 1986 643
rect 1986 612 1998 643
rect 1998 612 2020 643
rect 1964 598 2020 612
rect 1964 587 1986 598
rect 1986 587 1998 598
rect 1998 587 2020 598
rect 1964 546 1986 558
rect 1986 546 1998 558
rect 1998 546 2020 558
rect 1964 532 2020 546
rect 1964 502 1986 532
rect 1986 502 1998 532
rect 1998 502 2020 532
rect 1964 466 2020 473
rect 1964 417 1986 466
rect 1986 417 1998 466
rect 1998 417 2020 466
rect 23524 456 23580 512
rect 23650 456 23706 512
rect 17784 335 17840 391
rect 17866 335 17922 391
rect 17948 335 18004 391
rect 18029 335 18085 391
rect 18110 335 18166 391
rect 18268 354 18324 410
rect 18367 354 18423 410
rect 18465 354 18521 410
rect 23524 362 23580 418
rect 23650 362 23706 418
rect 4703 127 4759 183
rect 4783 127 4839 183
rect 16778 137 16834 193
rect 16871 137 16927 193
rect 16964 137 17020 193
rect 17057 137 17113 193
rect 17149 137 17205 193
rect 17241 137 17297 193
rect 16778 7 16834 63
rect 16871 7 16927 63
rect 16964 7 17020 63
rect 17057 7 17113 63
rect 17149 7 17205 63
rect 17241 7 17297 63
<< metal3 >>
rect 11850 38734 11854 38838
tri 11854 38734 11958 38838 sw
rect 11850 38729 12400 38734
rect 11850 38673 12008 38729
rect 12064 38673 12091 38729
rect 12147 38673 12174 38729
rect 12230 38673 12257 38729
rect 12313 38673 12339 38729
rect 12395 38673 12400 38729
rect 11850 38595 12400 38673
rect 11850 38539 12008 38595
rect 12064 38539 12091 38595
rect 12147 38539 12174 38595
rect 12230 38539 12257 38595
rect 12313 38539 12339 38595
rect 12395 38539 12400 38595
rect 11850 38534 12400 38539
tri 11850 38426 11958 38534 nw
rect 25865 37157 25931 37200
rect 25865 37101 25870 37157
rect 25926 37101 25931 37157
rect 25865 37077 25931 37101
rect 25865 37021 25870 37077
rect 25926 37021 25931 37077
rect 25865 37016 25931 37021
rect 23396 36247 23696 36253
rect 23460 36183 23514 36247
rect 23578 36183 23632 36247
rect 23396 36164 23696 36183
rect 23460 36100 23514 36164
rect 23578 36100 23632 36164
rect 23396 36081 23696 36100
rect 23460 36017 23514 36081
rect 23578 36017 23632 36081
rect 23396 35998 23696 36017
rect 23460 35934 23514 35998
rect 23578 35934 23632 35998
rect 23396 35915 23696 35934
rect 23460 35851 23514 35915
rect 23578 35851 23632 35915
rect 23396 35832 23696 35851
rect 23460 35768 23514 35832
rect 23578 35768 23632 35832
rect 23396 35749 23696 35768
rect 23460 35685 23514 35749
rect 23578 35685 23632 35749
rect 23396 35666 23696 35685
rect 19252 35562 19258 35626
rect 19322 35562 19340 35626
rect 19404 35562 19422 35626
rect 19486 35562 19504 35626
rect 19568 35562 19586 35626
rect 19650 35562 19668 35626
rect 19732 35562 19750 35626
rect 19814 35562 19832 35626
rect 19896 35562 19914 35626
rect 19978 35562 19996 35626
rect 20060 35562 20078 35626
rect 20142 35562 20160 35626
rect 20224 35562 20242 35626
rect 20306 35562 20324 35626
rect 20388 35562 20406 35626
rect 20470 35562 20488 35626
rect 20552 35562 20570 35626
rect 20634 35562 20652 35626
rect 20716 35562 20734 35626
rect 20798 35562 20816 35626
rect 20880 35562 20898 35626
rect 20962 35562 20980 35626
rect 21044 35562 21062 35626
rect 21126 35562 21144 35626
rect 21208 35562 21226 35626
rect 21290 35562 21308 35626
rect 21372 35562 21390 35626
rect 21454 35562 21472 35626
rect 21536 35562 21553 35626
rect 21617 35562 21634 35626
rect 21698 35562 21715 35626
rect 21779 35562 21796 35626
rect 21860 35562 21877 35626
rect 21941 35562 21958 35626
rect 22022 35562 22039 35626
rect 22103 35562 22120 35626
rect 22184 35562 22201 35626
rect 22265 35562 22282 35626
rect 22346 35562 22363 35626
rect 22427 35562 22444 35626
rect 22508 35562 22525 35626
rect 22589 35562 22595 35626
rect 19252 35546 22595 35562
rect 19252 35482 19258 35546
rect 19322 35482 19340 35546
rect 19404 35482 19422 35546
rect 19486 35482 19504 35546
rect 19568 35482 19586 35546
rect 19650 35482 19668 35546
rect 19732 35482 19750 35546
rect 19814 35482 19832 35546
rect 19896 35482 19914 35546
rect 19978 35482 19996 35546
rect 20060 35482 20078 35546
rect 20142 35482 20160 35546
rect 20224 35482 20242 35546
rect 20306 35482 20324 35546
rect 20388 35482 20406 35546
rect 20470 35482 20488 35546
rect 20552 35482 20570 35546
rect 20634 35482 20652 35546
rect 20716 35482 20734 35546
rect 20798 35482 20816 35546
rect 20880 35482 20898 35546
rect 20962 35482 20980 35546
rect 21044 35482 21062 35546
rect 21126 35482 21144 35546
rect 21208 35482 21226 35546
rect 21290 35482 21308 35546
rect 21372 35482 21390 35546
rect 21454 35482 21472 35546
rect 21536 35482 21553 35546
rect 21617 35482 21634 35546
rect 21698 35482 21715 35546
rect 21779 35482 21796 35546
rect 21860 35482 21877 35546
rect 21941 35482 21958 35546
rect 22022 35482 22039 35546
rect 22103 35482 22120 35546
rect 22184 35482 22201 35546
rect 22265 35482 22282 35546
rect 22346 35482 22363 35546
rect 22427 35482 22444 35546
rect 22508 35482 22525 35546
rect 22589 35482 22595 35546
rect 19252 35466 22595 35482
rect 19252 35402 19258 35466
rect 19322 35402 19340 35466
rect 19404 35402 19422 35466
rect 19486 35402 19504 35466
rect 19568 35402 19586 35466
rect 19650 35402 19668 35466
rect 19732 35402 19750 35466
rect 19814 35402 19832 35466
rect 19896 35402 19914 35466
rect 19978 35402 19996 35466
rect 20060 35402 20078 35466
rect 20142 35402 20160 35466
rect 20224 35402 20242 35466
rect 20306 35402 20324 35466
rect 20388 35402 20406 35466
rect 20470 35402 20488 35466
rect 20552 35402 20570 35466
rect 20634 35402 20652 35466
rect 20716 35402 20734 35466
rect 20798 35402 20816 35466
rect 20880 35402 20898 35466
rect 20962 35402 20980 35466
rect 21044 35402 21062 35466
rect 21126 35402 21144 35466
rect 21208 35402 21226 35466
rect 21290 35402 21308 35466
rect 21372 35402 21390 35466
rect 21454 35402 21472 35466
rect 21536 35402 21553 35466
rect 21617 35402 21634 35466
rect 21698 35402 21715 35466
rect 21779 35402 21796 35466
rect 21860 35402 21877 35466
rect 21941 35402 21958 35466
rect 22022 35402 22039 35466
rect 22103 35402 22120 35466
rect 22184 35402 22201 35466
rect 22265 35402 22282 35466
rect 22346 35402 22363 35466
rect 22427 35402 22444 35466
rect 22508 35402 22525 35466
rect 22589 35402 22595 35466
rect 19252 35386 22595 35402
rect 19252 35322 19258 35386
rect 19322 35322 19340 35386
rect 19404 35322 19422 35386
rect 19486 35322 19504 35386
rect 19568 35322 19586 35386
rect 19650 35322 19668 35386
rect 19732 35322 19750 35386
rect 19814 35322 19832 35386
rect 19896 35322 19914 35386
rect 19978 35322 19996 35386
rect 20060 35322 20078 35386
rect 20142 35322 20160 35386
rect 20224 35322 20242 35386
rect 20306 35322 20324 35386
rect 20388 35322 20406 35386
rect 20470 35322 20488 35386
rect 20552 35322 20570 35386
rect 20634 35322 20652 35386
rect 20716 35322 20734 35386
rect 20798 35322 20816 35386
rect 20880 35322 20898 35386
rect 20962 35322 20980 35386
rect 21044 35322 21062 35386
rect 21126 35322 21144 35386
rect 21208 35322 21226 35386
rect 21290 35322 21308 35386
rect 21372 35322 21390 35386
rect 21454 35322 21472 35386
rect 21536 35322 21553 35386
rect 21617 35322 21634 35386
rect 21698 35322 21715 35386
rect 21779 35322 21796 35386
rect 21860 35322 21877 35386
rect 21941 35322 21958 35386
rect 22022 35322 22039 35386
rect 22103 35322 22120 35386
rect 22184 35322 22201 35386
rect 22265 35322 22282 35386
rect 22346 35322 22363 35386
rect 22427 35322 22444 35386
rect 22508 35322 22525 35386
rect 22589 35322 22595 35386
rect 19252 35306 22595 35322
rect 19252 35242 19258 35306
rect 19322 35242 19340 35306
rect 19404 35242 19422 35306
rect 19486 35242 19504 35306
rect 19568 35242 19586 35306
rect 19650 35242 19668 35306
rect 19732 35242 19750 35306
rect 19814 35242 19832 35306
rect 19896 35242 19914 35306
rect 19978 35242 19996 35306
rect 20060 35242 20078 35306
rect 20142 35242 20160 35306
rect 20224 35242 20242 35306
rect 20306 35242 20324 35306
rect 20388 35242 20406 35306
rect 20470 35242 20488 35306
rect 20552 35242 20570 35306
rect 20634 35242 20652 35306
rect 20716 35242 20734 35306
rect 20798 35242 20816 35306
rect 20880 35242 20898 35306
rect 20962 35242 20980 35306
rect 21044 35242 21062 35306
rect 21126 35242 21144 35306
rect 21208 35242 21226 35306
rect 21290 35242 21308 35306
rect 21372 35242 21390 35306
rect 21454 35242 21472 35306
rect 21536 35242 21553 35306
rect 21617 35242 21634 35306
rect 21698 35242 21715 35306
rect 21779 35242 21796 35306
rect 21860 35242 21877 35306
rect 21941 35242 21958 35306
rect 22022 35242 22039 35306
rect 22103 35242 22120 35306
rect 22184 35242 22201 35306
rect 22265 35242 22282 35306
rect 22346 35242 22363 35306
rect 22427 35242 22444 35306
rect 22508 35242 22525 35306
rect 22589 35242 22595 35306
rect 19252 35226 22595 35242
rect 19252 35162 19258 35226
rect 19322 35162 19340 35226
rect 19404 35162 19422 35226
rect 19486 35162 19504 35226
rect 19568 35162 19586 35226
rect 19650 35162 19668 35226
rect 19732 35162 19750 35226
rect 19814 35162 19832 35226
rect 19896 35162 19914 35226
rect 19978 35162 19996 35226
rect 20060 35162 20078 35226
rect 20142 35162 20160 35226
rect 20224 35162 20242 35226
rect 20306 35162 20324 35226
rect 20388 35162 20406 35226
rect 20470 35162 20488 35226
rect 20552 35162 20570 35226
rect 20634 35162 20652 35226
rect 20716 35162 20734 35226
rect 20798 35162 20816 35226
rect 20880 35162 20898 35226
rect 20962 35162 20980 35226
rect 21044 35162 21062 35226
rect 21126 35162 21144 35226
rect 21208 35162 21226 35226
rect 21290 35162 21308 35226
rect 21372 35162 21390 35226
rect 21454 35162 21472 35226
rect 21536 35162 21553 35226
rect 21617 35162 21634 35226
rect 21698 35162 21715 35226
rect 21779 35162 21796 35226
rect 21860 35162 21877 35226
rect 21941 35162 21958 35226
rect 22022 35162 22039 35226
rect 22103 35162 22120 35226
rect 22184 35162 22201 35226
rect 22265 35162 22282 35226
rect 22346 35162 22363 35226
rect 22427 35162 22444 35226
rect 22508 35162 22525 35226
rect 22589 35162 22595 35226
rect 23460 35602 23514 35666
rect 23578 35602 23632 35666
rect 23396 35583 23696 35602
rect 23460 35519 23514 35583
rect 23578 35519 23632 35583
rect 23396 35500 23696 35519
rect 23460 35436 23514 35500
rect 23578 35436 23632 35500
rect 23396 35417 23696 35436
rect 23460 35353 23514 35417
rect 23578 35353 23632 35417
rect 23396 35333 23696 35353
rect 23460 35269 23514 35333
rect 23578 35269 23632 35333
rect 23396 35249 23696 35269
rect 23460 35185 23514 35249
rect 23578 35185 23632 35249
rect 23396 34378 23696 35185
rect 23391 34369 23701 34378
rect 23391 34313 23398 34369
rect 23454 34313 23478 34369
rect 23534 34313 23558 34369
rect 23614 34313 23638 34369
rect 23694 34313 23701 34369
rect 23391 34287 23701 34313
rect 23391 34231 23398 34287
rect 23454 34231 23478 34287
rect 23534 34231 23558 34287
rect 23614 34231 23638 34287
rect 23694 34231 23701 34287
rect 23391 34205 23701 34231
rect 23391 34149 23398 34205
rect 23454 34149 23478 34205
rect 23534 34149 23558 34205
rect 23614 34149 23638 34205
rect 23694 34149 23701 34205
rect 23391 34123 23701 34149
rect 23391 34067 23398 34123
rect 23454 34067 23478 34123
rect 23534 34067 23558 34123
rect 23614 34067 23638 34123
rect 23694 34067 23701 34123
rect 23391 34040 23701 34067
rect 23391 33984 23398 34040
rect 23454 33984 23478 34040
rect 23534 33984 23558 34040
rect 23614 33984 23638 34040
rect 23694 33984 23701 34040
rect 23391 33957 23701 33984
rect 23391 33901 23398 33957
rect 23454 33901 23478 33957
rect 23534 33901 23558 33957
rect 23614 33901 23638 33957
rect 23694 33901 23701 33957
rect 23391 33892 23701 33901
rect 597 32180 717 32189
rect 597 32124 619 32180
rect 675 32124 717 32180
rect 597 32100 717 32124
rect 597 32044 619 32100
rect 675 32044 717 32100
rect 597 32020 717 32044
rect 597 31964 619 32020
rect 675 31964 717 32020
tri 439 14649 597 14807 se
rect 597 14751 717 31964
rect 597 14719 685 14751
tri 685 14719 717 14751 nw
rect 802 31903 923 31912
rect 802 31847 829 31903
rect 885 31847 923 31903
rect 802 31823 923 31847
rect 802 31767 829 31823
rect 885 31767 923 31823
rect 802 31743 923 31767
rect 802 31687 829 31743
rect 885 31687 923 31743
rect 597 14658 624 14719
tri 624 14658 685 14719 nw
tri 741 14658 802 14719 se
rect 802 14662 923 31687
rect 802 14658 910 14662
rect 597 14649 615 14658
tri 615 14649 624 14658 nw
tri 732 14649 741 14658 se
rect 741 14649 910 14658
tri 910 14649 923 14662 nw
rect 993 24578 1113 24584
rect 993 24514 1016 24578
rect 1080 24514 1113 24578
rect 993 24470 1113 24514
rect 993 24406 1016 24470
rect 1080 24406 1113 24470
rect 993 24362 1113 24406
rect 993 24298 1016 24362
rect 1080 24298 1113 24362
tri 426 14636 439 14649 se
rect 439 14636 602 14649
tri 602 14636 615 14649 nw
tri 719 14636 732 14649 se
rect 732 14636 897 14649
tri 897 14636 910 14649 nw
tri 421 14631 426 14636 se
rect 426 14631 597 14636
tri 597 14631 602 14636 nw
tri 714 14631 719 14636 se
rect 719 14631 854 14636
tri 383 14593 421 14631 se
rect 421 14593 559 14631
tri 559 14593 597 14631 nw
tri 676 14593 714 14631 se
rect 714 14593 854 14631
tri 854 14593 897 14636 nw
tri 950 14593 993 14636 se
rect 993 14593 1113 24298
tri 353 14563 383 14593 se
rect 383 14563 529 14593
tri 529 14563 559 14593 nw
tri 646 14563 676 14593 se
rect 676 14566 827 14593
tri 827 14566 854 14593 nw
tri 923 14566 950 14593 se
rect 950 14578 1113 14593
rect 950 14566 1098 14578
rect 676 14563 824 14566
tri 824 14563 827 14566 nw
tri 920 14563 923 14566 se
rect 923 14563 1098 14566
tri 1098 14563 1113 14578 nw
tri 297 14507 353 14563 se
rect 353 14541 507 14563
tri 507 14541 529 14563 nw
tri 624 14541 646 14563 se
rect 646 14541 802 14563
tri 802 14541 824 14563 nw
tri 898 14541 920 14563 se
rect 920 14541 1042 14563
rect 353 14507 473 14541
tri 473 14507 507 14541 nw
tri 590 14507 624 14541 se
rect 624 14507 768 14541
tri 768 14507 802 14541 nw
tri 864 14507 898 14541 se
rect 898 14507 1042 14541
tri 1042 14507 1098 14563 nw
tri 267 14477 297 14507 se
rect 297 14480 446 14507
tri 446 14480 473 14507 nw
tri 563 14480 590 14507 se
rect 590 14480 738 14507
rect 297 14477 443 14480
tri 443 14477 446 14480 nw
tri 560 14477 563 14480 se
rect 563 14477 738 14480
tri 738 14477 768 14507 nw
tri 834 14477 864 14507 se
rect 864 14477 1012 14507
tri 1012 14477 1042 14507 nw
tri 248 14458 267 14477 se
rect 267 14458 424 14477
tri 424 14458 443 14477 nw
tri 541 14458 560 14477 se
rect 560 14458 719 14477
tri 719 14458 738 14477 nw
tri 815 14458 834 14477 se
rect 834 14458 993 14477
tri 993 14458 1012 14477 nw
tri 245 14455 248 14458 se
rect 248 14455 421 14458
tri 421 14455 424 14458 nw
tri 538 14455 541 14458 se
rect 541 14455 706 14458
tri 224 14434 245 14455 se
rect 245 14434 400 14455
tri 400 14434 421 14455 nw
tri 517 14434 538 14455 se
rect 538 14445 706 14455
tri 706 14445 719 14458 nw
tri 802 14445 815 14458 se
rect 815 14445 969 14458
rect 538 14434 695 14445
tri 695 14434 706 14445 nw
tri 791 14434 802 14445 se
rect 802 14434 969 14445
tri 969 14434 993 14458 nw
tri 1184 14439 1190 14445 se
rect 1190 14439 1250 33651
rect 1184 14434 1250 14439
tri 168 14378 224 14434 se
rect 224 14378 344 14434
tri 344 14378 400 14434 nw
tri 461 14378 517 14434 se
rect 517 14378 639 14434
tri 639 14378 695 14434 nw
tri 735 14378 791 14434 se
rect 791 14378 913 14434
tri 913 14378 969 14434 nw
rect 1184 14378 1189 14434
rect 1245 14378 1250 14434
tri 144 14354 168 14378 se
rect 168 14363 329 14378
tri 329 14363 344 14378 nw
tri 446 14363 461 14378 se
rect 461 14363 624 14378
tri 624 14363 639 14378 nw
tri 720 14363 735 14378 se
rect 735 14363 889 14378
rect 168 14354 320 14363
tri 320 14354 329 14363 nw
tri 437 14354 446 14363 se
rect 446 14354 615 14363
tri 615 14354 624 14363 nw
tri 711 14354 720 14363 se
rect 720 14354 889 14363
tri 889 14354 913 14378 nw
rect 1184 14354 1250 14378
tri 88 14298 144 14354 se
rect 144 14302 268 14354
tri 268 14302 320 14354 nw
tri 385 14302 437 14354 se
rect 437 14302 559 14354
rect 144 14298 264 14302
tri 264 14298 268 14302 nw
tri 381 14298 385 14302 se
rect 385 14298 559 14302
tri 559 14298 615 14354 nw
tri 655 14298 711 14354 se
rect 711 14298 833 14354
tri 833 14298 889 14354 nw
rect 1184 14298 1189 14354
rect 1245 14298 1250 14354
tri 70 14280 88 14298 se
rect 88 14280 246 14298
tri 246 14280 264 14298 nw
tri 363 14280 381 14298 se
rect 381 14280 541 14298
tri 541 14280 559 14298 nw
tri 637 14280 655 14298 se
rect 655 14280 815 14298
tri 815 14280 833 14298 nw
rect 1184 14293 1250 14298
tri 69 14279 70 14280 se
rect 70 14279 245 14280
tri 245 14279 246 14280 nw
tri 362 14279 363 14280 se
rect 363 14279 528 14280
tri 66 14276 69 14279 se
rect 69 14276 242 14279
tri 242 14276 245 14279 nw
tri 359 14276 362 14279 se
rect 362 14276 528 14279
rect 66 14249 215 14276
tri 215 14249 242 14276 nw
tri 332 14249 359 14276 se
rect 359 14267 528 14276
tri 528 14267 541 14280 nw
tri 624 14267 637 14280 se
rect 637 14267 784 14280
rect 359 14249 510 14267
tri 510 14249 528 14267 nw
tri 606 14249 624 14267 se
rect 624 14249 784 14267
tri 784 14249 815 14280 nw
rect 66 14224 190 14249
tri 190 14224 215 14249 nw
tri 307 14224 332 14249 se
rect 332 14224 485 14249
tri 485 14224 510 14249 nw
tri 581 14224 606 14249 se
rect 606 14224 759 14249
tri 759 14224 784 14249 nw
rect 66 0 186 14224
tri 186 14220 190 14224 nw
tri 303 14220 307 14224 se
rect 307 14220 480 14224
tri 302 14219 303 14220 se
rect 303 14219 480 14220
tri 480 14219 485 14224 nw
tri 576 14219 581 14224 se
rect 581 14219 754 14224
tri 754 14219 759 14224 nw
tri 268 14185 302 14219 se
rect 302 14185 446 14219
tri 446 14185 480 14219 nw
tri 542 14185 576 14219 se
rect 576 14185 708 14219
tri 256 14173 268 14185 se
rect 268 14173 434 14185
tri 434 14173 446 14185 nw
tri 530 14173 542 14185 se
rect 542 14173 708 14185
tri 708 14173 754 14219 nw
tri 1304 14178 1310 14184 se
rect 1310 14178 1370 33778
rect 1304 14173 1370 14178
tri 248 14165 256 14173 se
rect 256 14165 426 14173
tri 426 14165 434 14173 nw
tri 522 14165 530 14173 se
rect 530 14165 652 14173
rect 248 14117 378 14165
tri 378 14117 426 14165 nw
tri 474 14117 522 14165 se
rect 522 14117 652 14165
tri 652 14117 708 14173 nw
rect 1304 14117 1309 14173
rect 1365 14117 1370 14173
rect 248 1153 368 14117
tri 368 14107 378 14117 nw
tri 464 14107 474 14117 se
rect 474 14107 637 14117
tri 459 14102 464 14107 se
rect 464 14102 637 14107
tri 637 14102 652 14117 nw
tri 450 14093 459 14102 se
rect 459 14093 628 14102
tri 628 14093 637 14102 nw
rect 1304 14093 1370 14117
tri 430 14073 450 14093 se
rect 450 14073 608 14093
tri 608 14073 628 14093 nw
rect 430 14037 572 14073
tri 572 14037 608 14073 nw
rect 1304 14037 1309 14093
rect 1365 14037 1370 14093
rect 430 14026 561 14037
tri 561 14026 572 14037 nw
rect 1304 14032 1370 14037
rect 430 1323 550 14026
tri 550 14015 561 14026 nw
rect 822 12865 1220 12870
rect 822 12809 827 12865
rect 883 12809 949 12865
rect 1005 12809 1220 12865
rect 822 12785 1220 12809
rect 822 12729 827 12785
rect 883 12729 949 12785
rect 1005 12729 1220 12785
rect 822 12705 1220 12729
rect 822 12649 827 12705
rect 883 12649 949 12705
rect 1005 12649 1220 12705
rect 822 12625 1220 12649
rect 822 12569 827 12625
rect 883 12569 949 12625
rect 1005 12569 1220 12625
rect 822 12564 1220 12569
tri 822 12399 987 12564 ne
tri 942 11383 987 11428 se
rect 987 11383 1220 12564
tri 851 11292 942 11383 se
rect 942 11304 1220 11383
rect 942 11292 1208 11304
tri 1208 11292 1220 11304 nw
rect 851 11282 1198 11292
tri 1198 11282 1208 11292 nw
rect 851 11226 1142 11282
tri 1142 11226 1198 11282 nw
rect 851 11202 1118 11226
tri 1118 11202 1142 11226 nw
rect 695 10921 761 10926
rect 695 10865 700 10921
rect 756 10865 761 10921
rect 695 10841 761 10865
rect 695 10785 700 10841
rect 756 10785 761 10841
rect 695 10780 761 10785
tri 695 10775 700 10780 ne
tri 696 3349 700 3353 se
rect 700 3349 761 10780
rect 851 8037 1084 11202
tri 1084 11168 1118 11202 nw
rect 852 8031 1084 8037
rect 916 7967 936 8031
rect 1000 7967 1020 8031
rect 852 7944 1084 7967
rect 916 7880 936 7944
rect 1000 7880 1020 7944
rect 852 7857 1084 7880
rect 916 7793 936 7857
rect 1000 7793 1020 7857
rect 852 7769 1084 7793
rect 916 7705 936 7769
rect 1000 7705 1020 7769
rect 852 7681 1084 7705
rect 916 7617 936 7681
rect 1000 7617 1020 7681
rect 852 7593 1084 7617
rect 916 7529 936 7593
rect 1000 7529 1020 7593
rect 852 7505 1084 7529
rect 916 7441 936 7505
rect 1000 7441 1020 7505
rect 852 7417 1084 7441
rect 916 7353 936 7417
rect 1000 7353 1020 7417
rect 852 7347 1084 7353
rect 1146 10765 1213 10774
rect 1146 10709 1151 10765
rect 1207 10709 1213 10765
rect 1146 10685 1213 10709
rect 1146 10629 1151 10685
rect 1207 10629 1213 10685
rect 1146 10624 1213 10629
rect 1146 6992 1207 10624
tri 1207 10618 1213 10624 nw
tri 1411 10065 1430 10084 se
rect 1430 10065 1490 33646
tri 1371 10025 1411 10065 se
rect 1411 10042 1490 10065
rect 1411 10025 1473 10042
tri 1473 10025 1490 10042 nw
rect 1570 31112 2172 31375
rect 1570 31056 1667 31112
rect 1723 31056 1747 31112
rect 1803 31056 1827 31112
rect 1883 31056 2172 31112
rect 1570 31025 2172 31056
rect 1570 30969 1667 31025
rect 1723 30969 1747 31025
rect 1803 30969 1827 31025
rect 1883 30969 2172 31025
rect 1570 30938 2172 30969
rect 1570 30882 1667 30938
rect 1723 30882 1747 30938
rect 1803 30882 1827 30938
rect 1883 30882 2172 30938
rect 1570 30850 2172 30882
rect 1570 30794 1667 30850
rect 1723 30794 1747 30850
rect 1803 30794 1827 30850
rect 1883 30794 2172 30850
rect 1570 21362 2172 30794
rect 1570 21306 1870 21362
rect 1926 21306 2172 21362
rect 1570 21282 2172 21306
rect 1570 21226 1870 21282
rect 1926 21226 2172 21282
rect 1570 21202 2172 21226
rect 1570 21146 1870 21202
rect 1926 21146 2172 21202
rect 1570 21122 2172 21146
rect 1570 21066 1870 21122
rect 1926 21066 2172 21122
rect 1570 21042 2172 21066
rect 1570 20986 1870 21042
rect 1926 20986 2172 21042
rect 1570 20962 2172 20986
rect 1570 20906 1870 20962
rect 1926 20906 2172 20962
rect 1570 20882 2172 20906
rect 1570 20826 1870 20882
rect 1926 20826 2172 20882
rect 1570 20802 2172 20826
rect 1570 20746 1870 20802
rect 1926 20746 2172 20802
rect 1570 20722 2172 20746
rect 1570 20666 1870 20722
rect 1926 20666 2172 20722
rect 1570 20642 2172 20666
rect 1570 20586 1870 20642
rect 1926 20586 2172 20642
rect 1570 20562 2172 20586
rect 1570 20506 1870 20562
rect 1926 20506 2172 20562
rect 1570 20482 2172 20506
rect 1570 20426 1870 20482
rect 1926 20426 2172 20482
rect 1570 20401 2172 20426
rect 1570 20345 1870 20401
rect 1926 20345 2172 20401
rect 1570 20320 2172 20345
rect 1570 20264 1870 20320
rect 1926 20264 2172 20320
rect 1570 20239 2172 20264
rect 1570 20183 1870 20239
rect 1926 20183 2172 20239
rect 1570 20158 2172 20183
rect 1570 20102 1870 20158
rect 1926 20102 2172 20158
rect 1570 20077 2172 20102
rect 1570 20021 1870 20077
rect 1926 20021 2172 20077
rect 1570 19996 2172 20021
rect 1570 19940 1870 19996
rect 1926 19940 2172 19996
rect 1570 19915 2172 19940
rect 1570 19859 1870 19915
rect 1926 19859 2172 19915
rect 1570 19834 2172 19859
rect 1570 19778 1870 19834
rect 1926 19778 2172 19834
rect 1570 19753 2172 19778
rect 1570 19697 1870 19753
rect 1926 19697 2172 19753
rect 1570 19672 2172 19697
rect 1570 19616 1870 19672
rect 1926 19616 2172 19672
rect 1570 19591 2172 19616
rect 1570 19535 1870 19591
rect 1926 19535 2172 19591
rect 1570 19510 2172 19535
rect 1570 19454 1870 19510
rect 1926 19454 2172 19510
rect 1570 19429 2172 19454
rect 1570 19373 1870 19429
rect 1926 19373 2172 19429
rect 1570 19348 2172 19373
rect 1570 19292 1870 19348
rect 1926 19292 2172 19348
rect 1570 19267 2172 19292
rect 1570 19211 1870 19267
rect 1926 19211 2172 19267
rect 1570 19186 2172 19211
rect 1570 19130 1870 19186
rect 1926 19130 2172 19186
rect 1570 19105 2172 19130
rect 1570 19049 1870 19105
rect 1926 19049 2172 19105
rect 1570 19024 2172 19049
rect 1570 18968 1870 19024
rect 1926 18968 2172 19024
rect 1570 18943 2172 18968
rect 1570 18887 1870 18943
rect 1926 18887 2172 18943
rect 1570 18862 2172 18887
rect 1570 18806 1870 18862
rect 1926 18806 2172 18862
rect 1570 18781 2172 18806
rect 1570 18725 1870 18781
rect 1926 18725 2172 18781
rect 1570 18700 2172 18725
rect 1570 18644 1870 18700
rect 1926 18644 2172 18700
rect 1570 18619 2172 18644
rect 1570 18563 1870 18619
rect 1926 18563 2172 18619
rect 1570 18538 2172 18563
rect 1570 18482 1870 18538
rect 1926 18482 2172 18538
rect 1570 18201 2172 18482
rect 1570 18145 1771 18201
rect 1827 18145 1851 18201
rect 1907 18145 1931 18201
rect 1987 18145 2172 18201
rect 1570 18112 2172 18145
rect 1570 18056 1771 18112
rect 1827 18056 1851 18112
rect 1907 18056 1931 18112
rect 1987 18056 2172 18112
rect 1570 18023 2172 18056
rect 1570 17967 1771 18023
rect 1827 17967 1851 18023
rect 1907 17967 1931 18023
rect 1987 17967 2172 18023
rect 1570 17934 2172 17967
rect 1570 17878 1771 17934
rect 1827 17878 1851 17934
rect 1907 17878 1931 17934
rect 1987 17878 2172 17934
rect 1570 17845 2172 17878
rect 1570 17789 1771 17845
rect 1827 17789 1851 17845
rect 1907 17789 1931 17845
rect 1987 17789 2172 17845
rect 1570 17755 2172 17789
rect 1570 17699 1771 17755
rect 1827 17699 1851 17755
rect 1907 17699 1931 17755
rect 1987 17699 2172 17755
rect 1570 17527 2172 17699
rect 1570 17391 1771 17527
rect 1987 17391 2172 17527
rect 1570 17366 2172 17391
rect 1570 17310 1771 17366
rect 1827 17310 1851 17366
rect 1907 17310 1931 17366
rect 1987 17310 2172 17366
rect 1570 17285 2172 17310
rect 1570 17229 1771 17285
rect 1827 17229 1851 17285
rect 1907 17229 1931 17285
rect 1987 17229 2172 17285
rect 1570 17204 2172 17229
rect 1570 17148 1771 17204
rect 1827 17148 1851 17204
rect 1907 17148 1931 17204
rect 1987 17148 2172 17204
rect 1570 17123 2172 17148
rect 1570 17067 1771 17123
rect 1827 17067 1851 17123
rect 1907 17067 1931 17123
rect 1987 17067 2172 17123
rect 1570 16322 2172 17067
rect 1570 16266 1771 16322
rect 1827 16266 1851 16322
rect 1907 16266 1931 16322
rect 1987 16266 2172 16322
rect 1570 16235 2172 16266
rect 1570 16179 1771 16235
rect 1827 16179 1851 16235
rect 1907 16179 1931 16235
rect 1987 16179 2172 16235
rect 1570 16148 2172 16179
rect 1570 16092 1771 16148
rect 1827 16092 1851 16148
rect 1907 16092 1931 16148
rect 1987 16092 2172 16148
rect 1570 16061 2172 16092
rect 1570 16005 1771 16061
rect 1827 16005 1851 16061
rect 1907 16005 1931 16061
rect 1987 16005 2172 16061
rect 1570 15974 2172 16005
rect 1570 15918 1771 15974
rect 1827 15918 1851 15974
rect 1907 15918 1931 15974
rect 1987 15918 2172 15974
rect 1570 15887 2172 15918
rect 1570 15831 1771 15887
rect 1827 15831 1851 15887
rect 1907 15831 1931 15887
rect 1987 15831 2172 15887
rect 1570 15800 2172 15831
rect 1570 15744 1771 15800
rect 1827 15744 1851 15800
rect 1907 15744 1931 15800
rect 1987 15744 2172 15800
rect 1570 15713 2172 15744
rect 1570 15657 1771 15713
rect 1827 15657 1851 15713
rect 1907 15657 1931 15713
rect 1987 15657 2172 15713
rect 1570 15626 2172 15657
rect 1570 15570 1771 15626
rect 1827 15570 1851 15626
rect 1907 15570 1931 15626
rect 1987 15570 2172 15626
rect 1570 15539 2172 15570
rect 1570 15483 1771 15539
rect 1827 15483 1851 15539
rect 1907 15483 1931 15539
rect 1987 15483 2172 15539
rect 1570 14649 2172 15483
rect 1570 14593 1771 14649
rect 1827 14593 1851 14649
rect 1907 14593 1931 14649
rect 1987 14593 2172 14649
rect 1570 14563 2172 14593
rect 1570 14507 1771 14563
rect 1827 14507 1851 14563
rect 1907 14507 1931 14563
rect 1987 14507 2172 14563
rect 1570 14477 2172 14507
rect 1570 14421 1771 14477
rect 1827 14421 1851 14477
rect 1907 14421 1931 14477
rect 1987 14421 2172 14477
rect 1570 14391 2172 14421
rect 1570 14335 1771 14391
rect 1827 14335 1851 14391
rect 1907 14335 1931 14391
rect 1987 14335 2172 14391
rect 1570 14305 2172 14335
rect 1570 14249 1771 14305
rect 1827 14249 1851 14305
rect 1907 14249 1931 14305
rect 1987 14249 2172 14305
rect 1570 14219 2172 14249
rect 1570 14163 1771 14219
rect 1827 14163 1851 14219
rect 1907 14163 1931 14219
rect 1987 14163 2172 14219
rect 1570 14132 2172 14163
rect 1570 14076 1771 14132
rect 1827 14076 1851 14132
rect 1907 14076 1931 14132
rect 1987 14076 2172 14132
tri 1349 10003 1371 10025 se
rect 1371 10003 1451 10025
tri 1451 10003 1473 10025 nw
tri 1328 9982 1349 10003 se
rect 1349 9982 1430 10003
tri 1430 9982 1451 10003 nw
tri 1293 9947 1328 9982 se
rect 1328 9947 1395 9982
tri 1395 9947 1430 9982 nw
tri 1275 9929 1293 9947 se
rect 1293 9929 1377 9947
tri 1377 9929 1395 9947 nw
tri 1270 9924 1275 9929 se
rect 1275 9924 1372 9929
tri 1372 9924 1377 9929 nw
rect 1270 9923 1371 9924
tri 1371 9923 1372 9924 nw
rect 1270 7126 1331 9923
tri 1331 9883 1371 9923 nw
rect 1570 9240 2172 14076
rect 1570 9176 1595 9240
rect 1659 9176 1675 9240
rect 1739 9176 1755 9240
rect 1819 9176 1835 9240
rect 1899 9176 1915 9240
rect 1979 9176 1995 9240
rect 2059 9176 2075 9240
rect 2139 9176 2172 9240
rect 1570 9155 2172 9176
rect 1570 9091 1595 9155
rect 1659 9091 1675 9155
rect 1739 9091 1755 9155
rect 1819 9091 1835 9155
rect 1899 9091 1915 9155
rect 1979 9091 1995 9155
rect 2059 9091 2075 9155
rect 2139 9091 2172 9155
rect 1570 9070 2172 9091
rect 1570 9006 1595 9070
rect 1659 9006 1675 9070
rect 1739 9006 1755 9070
rect 1819 9006 1835 9070
rect 1899 9006 1915 9070
rect 1979 9006 1995 9070
rect 2059 9006 2075 9070
rect 2139 9006 2172 9070
rect 1570 8985 2172 9006
rect 1570 8921 1595 8985
rect 1659 8921 1675 8985
rect 1739 8921 1755 8985
rect 1819 8921 1835 8985
rect 1899 8921 1915 8985
rect 1979 8921 1995 8985
rect 2059 8921 2075 8985
rect 2139 8921 2172 8985
rect 1570 8900 2172 8921
rect 1570 8836 1595 8900
rect 1659 8836 1675 8900
rect 1739 8836 1755 8900
rect 1819 8836 1835 8900
rect 1899 8836 1915 8900
rect 1979 8836 1995 8900
rect 2059 8836 2075 8900
rect 2139 8836 2172 8900
rect 1570 8815 2172 8836
rect 1570 8751 1595 8815
rect 1659 8751 1675 8815
rect 1739 8751 1755 8815
rect 1819 8751 1835 8815
rect 1899 8751 1915 8815
rect 1979 8751 1995 8815
rect 2059 8751 2075 8815
rect 2139 8751 2172 8815
rect 1570 8730 2172 8751
rect 1570 8666 1595 8730
rect 1659 8666 1675 8730
rect 1739 8666 1755 8730
rect 1819 8666 1835 8730
rect 1899 8666 1915 8730
rect 1979 8666 1995 8730
rect 2059 8666 2075 8730
rect 2139 8666 2172 8730
rect 1570 8645 2172 8666
rect 1570 8581 1595 8645
rect 1659 8581 1675 8645
rect 1739 8581 1755 8645
rect 1819 8581 1835 8645
rect 1899 8581 1915 8645
rect 1979 8581 1995 8645
rect 2059 8581 2075 8645
rect 2139 8581 2172 8645
rect 1570 8560 2172 8581
rect 1570 8496 1595 8560
rect 1659 8496 1675 8560
rect 1739 8496 1755 8560
rect 1819 8496 1835 8560
rect 1899 8496 1915 8560
rect 1979 8496 1995 8560
rect 2059 8496 2075 8560
rect 2139 8496 2172 8560
rect 1570 8474 2172 8496
rect 1570 8410 1595 8474
rect 1659 8410 1675 8474
rect 1739 8410 1755 8474
rect 1819 8410 1835 8474
rect 1899 8410 1915 8474
rect 1979 8410 1995 8474
rect 2059 8410 2075 8474
rect 2139 8410 2172 8474
rect 1570 8388 2172 8410
rect 1570 8324 1595 8388
rect 1659 8324 1675 8388
rect 1739 8324 1755 8388
rect 1819 8324 1835 8388
rect 1899 8324 1915 8388
rect 1979 8324 1995 8388
rect 2059 8324 2075 8388
rect 2139 8324 2172 8388
rect 1570 8317 2172 8324
tri 1331 7126 1336 7131 sw
rect 1270 7094 1336 7126
tri 1270 7089 1275 7094 ne
tri 1207 6992 1212 6997 sw
rect 1146 6987 1212 6992
rect 1146 6931 1151 6987
rect 1207 6931 1212 6987
rect 1146 6907 1212 6931
rect 1146 6851 1151 6907
rect 1207 6851 1212 6907
rect 1146 6846 1212 6851
tri 1270 6702 1275 6707 se
rect 1275 6702 1336 7094
rect 1750 6987 1816 6992
rect 1750 6931 1755 6987
rect 1811 6931 1816 6987
rect 1750 6907 1816 6931
rect 1750 6851 1755 6907
rect 1811 6851 1816 6907
rect 1750 6846 1816 6851
rect 1270 6650 1336 6702
tri 1254 4360 1270 4376 se
rect 1270 4360 1331 6650
tri 1331 6645 1336 6650 nw
rect 1543 6520 1689 6525
rect 1543 6464 1548 6520
rect 1604 6464 1628 6520
rect 1684 6464 1689 6520
rect 1543 6459 1689 6464
tri 1578 6450 1587 6459 ne
rect 1587 6450 1689 6459
tri 1587 6414 1623 6450 ne
tri 1226 4332 1254 4360 se
rect 1254 4345 1331 4360
rect 1254 4332 1318 4345
tri 1318 4332 1331 4345 nw
rect 1393 6376 1459 6381
rect 1393 6320 1398 6376
rect 1454 6320 1459 6376
rect 1393 6296 1459 6320
rect 1393 6240 1398 6296
rect 1454 6240 1459 6296
rect 1393 6235 1459 6240
tri 1178 4284 1226 4332 se
rect 1226 4284 1270 4332
tri 1270 4284 1318 4332 nw
tri 1170 4276 1178 4284 se
rect 1178 4276 1262 4284
tri 1262 4276 1270 4284 nw
tri 1161 4267 1170 4276 se
rect 1170 4267 1253 4276
tri 1253 4267 1262 4276 nw
rect 1161 4252 1238 4267
tri 1238 4252 1253 4267 nw
rect 1161 4249 1235 4252
tri 1235 4249 1238 4252 nw
tri 761 3349 762 3350 sw
rect 696 3344 762 3349
rect 696 3288 701 3344
rect 757 3288 762 3344
rect 696 3264 762 3288
rect 696 3208 701 3264
rect 757 3208 762 3264
rect 696 3203 762 3208
tri 696 3199 700 3203 ne
rect 700 3199 761 3203
tri 761 3202 762 3203 nw
tri 1158 3144 1161 3147 se
rect 1161 3145 1222 4249
tri 1222 4236 1235 4249 nw
tri 1380 4236 1393 4249 se
rect 1393 4236 1454 6235
tri 1454 6230 1459 6235 nw
tri 1539 5058 1623 5142 se
rect 1623 5058 1689 6450
rect 1533 4994 1539 5058
rect 1603 4994 1619 5058
rect 1683 4994 1689 5058
tri 1340 4196 1380 4236 se
rect 1380 4221 1454 4236
rect 1380 4196 1429 4221
tri 1429 4196 1454 4221 nw
tri 1304 4160 1340 4196 se
rect 1340 4160 1393 4196
tri 1393 4160 1429 4196 nw
tri 1289 4145 1304 4160 se
rect 1304 4145 1378 4160
tri 1378 4145 1393 4160 nw
tri 1284 4140 1289 4145 se
rect 1289 4140 1373 4145
tri 1373 4140 1378 4145 nw
rect 1284 4121 1354 4140
tri 1354 4121 1373 4140 nw
tri 1222 3145 1224 3147 sw
rect 1161 3144 1224 3145
rect 1158 3139 1224 3144
rect 1158 3083 1163 3139
rect 1219 3083 1224 3139
rect 1158 3059 1224 3083
rect 1158 3003 1163 3059
rect 1219 3003 1224 3059
rect 1158 2998 1224 3003
tri 1283 2930 1284 2931 se
rect 1284 2930 1345 4121
tri 1345 4112 1354 4121 nw
tri 1244 2891 1283 2930 se
rect 1283 2891 1345 2930
rect 1158 2886 1345 2891
rect 1158 2830 1163 2886
rect 1219 2830 1345 2886
rect 1158 2810 1345 2830
rect 1422 3926 1488 3947
rect 1422 3870 1427 3926
rect 1483 3870 1488 3926
rect 1422 3846 1488 3870
rect 1422 3790 1427 3846
rect 1483 3790 1488 3846
rect 1158 2806 1245 2810
rect 1158 2750 1163 2806
rect 1219 2793 1245 2806
tri 1245 2793 1262 2810 nw
rect 1219 2750 1224 2793
tri 1224 2772 1245 2793 nw
rect 1158 2745 1224 2750
rect 1153 2630 1273 2641
rect 1153 2574 1190 2630
rect 1246 2574 1273 2630
rect 1153 2550 1273 2574
rect 1153 2494 1190 2550
rect 1246 2494 1273 2550
tri 550 1323 554 1327 sw
rect 430 1300 554 1323
tri 554 1300 577 1323 sw
rect 430 1267 577 1300
tri 577 1267 610 1300 sw
rect 430 1252 610 1267
tri 610 1252 625 1267 sw
tri 430 1238 444 1252 ne
rect 444 1238 625 1252
tri 625 1238 639 1252 sw
tri 444 1182 500 1238 ne
rect 500 1182 639 1238
tri 639 1182 695 1238 sw
tri 500 1166 516 1182 ne
rect 516 1180 695 1182
tri 695 1180 697 1182 sw
rect 516 1166 697 1180
tri 368 1153 381 1166 sw
tri 516 1153 529 1166 ne
rect 529 1153 697 1166
rect 248 1105 381 1153
tri 381 1105 429 1153 sw
tri 529 1105 577 1153 ne
rect 248 1097 429 1105
tri 429 1097 437 1105 sw
rect 248 1094 437 1097
tri 437 1094 440 1097 sw
rect 248 1093 440 1094
tri 248 1088 253 1093 ne
rect 253 1088 440 1093
tri 253 1068 273 1088 ne
rect 273 1068 440 1088
tri 273 1021 320 1068 ne
rect 320 0 440 1068
rect 577 0 697 1153
rect 1153 0 1273 2494
rect 1422 0 1488 3790
tri 1753 3167 1755 3169 se
rect 1755 3167 1816 6846
rect 2252 6381 2313 33778
rect 3718 33111 3998 33117
rect 3782 33106 3826 33111
rect 3890 33106 3934 33111
rect 3788 33050 3826 33106
rect 3902 33050 3934 33106
rect 3782 33047 3826 33050
rect 3890 33047 3934 33050
rect 3718 33014 3998 33047
rect 23396 33032 23696 33892
rect 3782 33010 3826 33014
rect 3890 33010 3934 33014
rect 3788 32954 3826 33010
rect 3902 32954 3934 33010
rect 3782 32950 3826 32954
rect 3890 32950 3934 32954
rect 3718 32917 3998 32950
rect 3782 32914 3826 32917
rect 3890 32914 3934 32917
rect 3788 32858 3826 32914
rect 3902 32858 3934 32914
rect 3782 32853 3826 32858
rect 3890 32853 3934 32858
rect 3718 32820 3998 32853
rect 3782 32818 3826 32820
rect 3890 32818 3934 32820
rect 3788 32762 3826 32818
rect 3902 32762 3934 32818
rect 3782 32756 3826 32762
rect 3890 32756 3934 32762
rect 3718 32722 3998 32756
rect 3782 32721 3826 32722
rect 3890 32721 3934 32722
rect 3788 32665 3826 32721
rect 3902 32665 3934 32721
rect 3782 32658 3826 32665
rect 3890 32658 3934 32665
rect 3718 32652 3998 32658
rect 23391 33023 23701 33032
rect 23391 32967 23398 33023
rect 23454 32967 23478 33023
rect 23534 32967 23558 33023
rect 23614 32967 23638 33023
rect 23694 32967 23701 33023
rect 23391 32941 23701 32967
rect 23391 32885 23398 32941
rect 23454 32885 23478 32941
rect 23534 32885 23558 32941
rect 23614 32885 23638 32941
rect 23694 32885 23701 32941
rect 23391 32859 23701 32885
rect 23391 32803 23398 32859
rect 23454 32803 23478 32859
rect 23534 32803 23558 32859
rect 23614 32803 23638 32859
rect 23694 32803 23701 32859
rect 23391 32776 23701 32803
rect 23391 32720 23398 32776
rect 23454 32720 23478 32776
rect 23534 32720 23558 32776
rect 23614 32720 23638 32776
rect 23694 32720 23701 32776
rect 23391 32693 23701 32720
rect 23391 32637 23398 32693
rect 23454 32637 23478 32693
rect 23534 32637 23558 32693
rect 23614 32637 23638 32693
rect 23694 32637 23701 32693
rect 23391 32610 23701 32637
rect 23391 32554 23398 32610
rect 23454 32554 23478 32610
rect 23534 32554 23558 32610
rect 23614 32554 23638 32610
rect 23694 32554 23701 32610
rect 23391 32545 23701 32554
rect 18738 23746 19056 23762
rect 18738 23690 18744 23746
rect 18800 23690 18854 23746
rect 18910 23690 18964 23746
rect 19020 23690 19056 23746
rect 18738 23659 19056 23690
rect 18738 23603 18744 23659
rect 18800 23603 18854 23659
rect 18910 23603 18964 23659
rect 19020 23603 19056 23659
rect 18738 23572 19056 23603
rect 18738 23516 18744 23572
rect 18800 23516 18854 23572
rect 18910 23516 18964 23572
rect 19020 23516 19056 23572
rect 18738 23485 19056 23516
rect 18738 23429 18744 23485
rect 18800 23429 18854 23485
rect 18910 23429 18964 23485
rect 19020 23429 19056 23485
rect 18738 23398 19056 23429
rect 18738 23342 18744 23398
rect 18800 23342 18854 23398
rect 18910 23342 18964 23398
rect 19020 23342 19056 23398
rect 18738 23311 19056 23342
rect 18738 23255 18744 23311
rect 18800 23255 18854 23311
rect 18910 23255 18964 23311
rect 19020 23255 19056 23311
rect 18738 23223 19056 23255
rect 18738 23167 18744 23223
rect 18800 23167 18854 23223
rect 18910 23167 18964 23223
rect 19020 23167 19056 23223
rect 18738 23135 19056 23167
rect 18738 23079 18744 23135
rect 18800 23079 18854 23135
rect 18910 23079 18964 23135
rect 19020 23079 19056 23135
rect 18738 23047 19056 23079
rect 18738 22991 18744 23047
rect 18800 22991 18854 23047
rect 18910 22991 18964 23047
rect 19020 22991 19056 23047
rect 18738 22959 19056 22991
rect 18738 22903 18744 22959
rect 18800 22903 18854 22959
rect 18910 22903 18964 22959
rect 19020 22903 19056 22959
rect 18738 22871 19056 22903
rect 27051 23272 27537 23280
rect 27051 23216 27056 23272
rect 27112 23216 27140 23272
rect 27196 23216 27224 23272
rect 27280 23216 27308 23272
rect 27364 23216 27392 23272
rect 27448 23216 27476 23272
rect 27532 23216 27537 23272
rect 27051 23192 27537 23216
rect 27051 23136 27056 23192
rect 27112 23136 27140 23192
rect 27196 23136 27224 23192
rect 27280 23136 27308 23192
rect 27364 23136 27392 23192
rect 27448 23136 27476 23192
rect 27532 23136 27537 23192
rect 27051 23112 27537 23136
rect 27051 23056 27056 23112
rect 27112 23056 27140 23112
rect 27196 23056 27224 23112
rect 27280 23056 27308 23112
rect 27364 23056 27392 23112
rect 27448 23056 27476 23112
rect 27532 23056 27537 23112
rect 27051 23032 27537 23056
rect 27051 22976 27056 23032
rect 27112 22976 27140 23032
rect 27196 22976 27224 23032
rect 27280 22976 27308 23032
rect 27364 22976 27392 23032
rect 27448 22976 27476 23032
rect 27532 22976 27537 23032
rect 27051 22952 27537 22976
rect 27051 22896 27056 22952
rect 27112 22896 27140 22952
rect 27196 22896 27224 22952
rect 27280 22896 27308 22952
rect 27364 22896 27392 22952
rect 27448 22896 27476 22952
rect 27532 22896 27537 22952
rect 27051 22888 27537 22896
rect 18738 22815 18744 22871
rect 18800 22815 18854 22871
rect 18910 22815 18964 22871
rect 19020 22815 19056 22871
tri 18694 21982 18738 22026 se
rect 18738 21982 19056 22815
rect 27340 22858 27544 22863
rect 27340 22802 27345 22858
rect 27401 22802 27483 22858
rect 27539 22802 27544 22858
rect 27340 22776 27544 22802
rect 27340 22720 27345 22776
rect 27401 22720 27483 22776
rect 27539 22720 27544 22776
rect 27340 22694 27544 22720
rect 27340 22638 27345 22694
rect 27401 22638 27483 22694
rect 27539 22638 27544 22694
rect 27340 22612 27544 22638
rect 27340 22556 27345 22612
rect 27401 22556 27483 22612
rect 27539 22556 27544 22612
rect 27340 22530 27544 22556
rect 27340 22474 27345 22530
rect 27401 22474 27483 22530
rect 27539 22474 27544 22530
rect 27340 22448 27544 22474
rect 27340 22392 27345 22448
rect 27401 22392 27483 22448
rect 27539 22392 27544 22448
rect 27340 22366 27544 22392
rect 27340 22310 27345 22366
rect 27401 22310 27483 22366
rect 27539 22310 27544 22366
tri 23053 22284 23066 22297 sw
rect 27340 22284 27544 22310
rect 23053 22270 23066 22284
tri 23066 22270 23080 22284 sw
rect 22930 22236 23080 22270
tri 22930 22228 22938 22236 ne
rect 22938 22228 23080 22236
tri 23080 22228 23122 22270 sw
rect 27340 22228 27345 22284
rect 27401 22228 27483 22284
rect 27539 22228 27544 22284
tri 22938 22202 22964 22228 ne
rect 22964 22202 23122 22228
tri 23122 22202 23148 22228 sw
rect 27340 22202 27544 22228
tri 22964 22172 22994 22202 ne
rect 22994 22172 23148 22202
tri 23148 22172 23178 22202 sw
tri 22994 22146 23020 22172 ne
rect 23020 22146 23178 22172
tri 23020 22120 23046 22146 ne
rect 23046 22120 23178 22146
tri 23046 22113 23053 22120 ne
rect 23053 22113 23178 22120
tri 23053 22108 23058 22113 ne
tri 18668 21956 18694 21982 se
rect 18694 21956 19056 21982
tri 18612 21900 18668 21956 se
rect 18668 21900 19056 21956
tri 18603 21891 18612 21900 se
rect 18612 21891 19056 21900
rect 2382 20793 2520 20798
rect 2382 20737 2423 20793
rect 2479 20737 2520 20793
rect 2382 20708 2520 20737
rect 2382 20652 2423 20708
rect 2479 20652 2520 20708
rect 2382 6895 2520 20652
rect 8084 18320 8973 18992
rect 12727 18320 13616 18992
rect 14568 18320 15457 18992
rect 19211 18320 20100 18992
rect 21052 18320 21941 18992
rect 2789 14224 2855 14229
rect 2789 14168 2794 14224
rect 2850 14168 2855 14224
rect 2789 14144 2855 14168
rect 2789 14088 2794 14144
rect 2850 14088 2855 14144
rect 22097 14130 22978 14135
rect 2789 8138 2855 14088
rect 22096 14128 22978 14130
rect 22096 14072 22106 14128
rect 22162 14072 22187 14128
rect 22243 14072 22268 14128
rect 22324 14072 22349 14128
rect 22405 14072 22430 14128
rect 22486 14072 22511 14128
rect 22567 14072 22592 14128
rect 22648 14072 22673 14128
rect 22729 14072 22753 14128
rect 22809 14072 22833 14128
rect 22889 14072 22913 14128
rect 22969 14072 22978 14128
rect 22096 14026 22978 14072
tri 2925 13988 2945 14008 se
rect 2945 13988 3607 14008
tri 3607 13988 3627 14008 nw
rect 2789 8082 2794 8138
rect 2850 8082 2855 8138
rect 2789 8058 2855 8082
rect 2789 8002 2794 8058
rect 2850 8002 2855 8058
rect 2789 7997 2855 8002
tri 2920 13983 2925 13988 se
rect 2925 13983 3602 13988
tri 3602 13983 3607 13988 nw
rect 2920 13970 3589 13983
tri 3589 13970 3602 13983 nw
rect 5206 13970 5976 13988
tri 5976 13970 5994 13988 nw
rect 22096 13970 22106 14026
rect 22162 13970 22187 14026
rect 22243 13970 22268 14026
rect 22324 13970 22349 14026
rect 22405 13970 22430 14026
rect 22486 13970 22511 14026
rect 22567 13970 22592 14026
rect 22648 13970 22673 14026
rect 22729 13970 22753 14026
rect 22809 13970 22833 14026
rect 22889 13970 22913 14026
rect 22969 13970 22978 14026
rect 2920 13968 3587 13970
tri 3587 13968 3589 13970 nw
rect 5206 13968 5974 13970
tri 5974 13968 5976 13970 nw
rect 2920 13926 3545 13968
tri 3545 13926 3587 13968 nw
rect 5206 13926 5932 13968
tri 5932 13926 5974 13968 nw
rect 2920 13924 3543 13926
tri 3543 13924 3545 13926 nw
rect 5206 13924 5930 13926
tri 5930 13924 5932 13926 nw
rect 22096 13924 22978 13970
rect 2920 13868 3487 13924
tri 3487 13868 3543 13924 nw
rect 5206 13868 5874 13924
tri 5874 13868 5930 13924 nw
rect 22096 13868 22106 13924
rect 22162 13868 22187 13924
rect 22243 13868 22268 13924
rect 22324 13868 22349 13924
rect 22405 13868 22430 13924
rect 22486 13868 22511 13924
rect 22567 13868 22592 13924
rect 22648 13868 22673 13924
rect 22729 13868 22753 13924
rect 22809 13868 22833 13924
rect 22889 13868 22913 13924
rect 22969 13868 22978 13924
rect 2920 13828 3447 13868
tri 3447 13828 3487 13868 nw
rect 5206 13828 5834 13868
tri 5834 13828 5874 13868 nw
rect 2920 13822 3441 13828
tri 3441 13822 3447 13828 nw
rect 5206 13822 5828 13828
tri 5828 13822 5834 13828 nw
rect 22096 13822 22978 13868
rect 2920 13766 3385 13822
tri 3385 13766 3441 13822 nw
rect 5206 13766 5772 13822
tri 5772 13766 5828 13822 nw
rect 22096 13766 22106 13822
rect 22162 13766 22187 13822
rect 22243 13766 22268 13822
rect 22324 13766 22349 13822
rect 22405 13766 22430 13822
rect 22486 13766 22511 13822
rect 22567 13766 22592 13822
rect 22648 13766 22673 13822
rect 22729 13766 22753 13822
rect 22809 13766 22833 13822
rect 22889 13766 22913 13822
rect 22969 13766 22978 13822
rect 2382 6890 2528 6895
rect 2382 6834 2387 6890
rect 2443 6834 2467 6890
rect 2523 6834 2528 6890
rect 2382 6829 2528 6834
rect 2920 6403 3249 13766
tri 3249 13630 3385 13766 nw
rect 5206 13762 5768 13766
tri 5768 13762 5772 13766 nw
rect 22096 13762 22978 13766
rect 5206 13759 5765 13762
tri 5765 13759 5768 13762 nw
rect 22097 13759 22978 13762
rect 5206 13687 5693 13759
tri 5693 13687 5765 13759 nw
rect 6848 13697 7774 13698
rect 3313 11519 3706 11524
rect 3313 11463 3500 11519
rect 3556 11463 3645 11519
rect 3701 11463 3706 11519
rect 3313 11439 3706 11463
rect 3313 11383 3500 11439
rect 3556 11383 3645 11439
rect 3701 11383 3706 11439
rect 3313 11378 3706 11383
rect 3313 10277 3695 11378
tri 3695 11367 3706 11378 nw
rect 3313 10221 3318 10277
rect 3374 10221 3422 10277
rect 3478 10221 3526 10277
rect 3582 10221 3630 10277
rect 3686 10221 3695 10277
rect 3313 10197 3695 10221
rect 3313 10141 3318 10197
rect 3374 10141 3422 10197
rect 3478 10141 3526 10197
rect 3582 10141 3630 10197
rect 3686 10141 3695 10197
rect 3313 10003 3695 10141
rect 3313 9947 3318 10003
rect 3374 9947 3422 10003
rect 3478 9947 3526 10003
rect 3582 9947 3630 10003
rect 3686 9947 3695 10003
rect 3313 9923 3695 9947
rect 3313 9867 3318 9923
rect 3374 9867 3422 9923
rect 3478 9867 3526 9923
rect 3582 9867 3630 9923
rect 3686 9867 3695 9923
rect 3313 8021 3695 9867
rect 3377 7957 3419 8021
rect 3483 7957 3525 8021
rect 3589 7957 3631 8021
rect 3313 7937 3695 7957
rect 3377 7873 3419 7937
rect 3483 7873 3525 7937
rect 3589 7873 3631 7937
rect 3313 7852 3695 7873
rect 3377 7788 3419 7852
rect 3483 7788 3525 7852
rect 3589 7788 3631 7852
rect 3313 7767 3695 7788
rect 3377 7703 3419 7767
rect 3483 7703 3525 7767
rect 3589 7703 3631 7767
rect 3313 7682 3695 7703
rect 3377 7618 3419 7682
rect 3483 7618 3525 7682
rect 3589 7618 3631 7682
rect 3313 7597 3695 7618
rect 3377 7533 3419 7597
rect 3483 7533 3525 7597
rect 3589 7533 3631 7597
rect 3313 7512 3695 7533
rect 3377 7448 3419 7512
rect 3483 7448 3525 7512
rect 3589 7448 3631 7512
rect 3313 7427 3695 7448
rect 3377 7363 3419 7427
rect 3483 7363 3525 7427
rect 3589 7363 3631 7427
rect 3313 7350 3695 7363
rect 3808 7139 3954 7144
rect 3808 7083 3813 7139
rect 3869 7083 3893 7139
rect 3949 7083 3954 7139
rect 3808 6890 3954 7083
rect 3808 6834 3813 6890
rect 3869 6834 3893 6890
rect 3949 6834 3954 6890
rect 3808 6829 3954 6834
rect 5206 6757 5555 13687
tri 5555 13549 5693 13687 nw
rect 6848 13633 6854 13697
rect 6918 13633 6939 13697
rect 7003 13633 7024 13697
rect 7088 13633 7109 13697
rect 7173 13633 7194 13697
rect 7258 13633 7279 13697
rect 7343 13633 7364 13697
rect 7428 13633 7449 13697
rect 7513 13633 7534 13697
rect 7598 13633 7619 13697
rect 7683 13633 7704 13697
rect 7768 13633 7774 13697
rect 6848 13609 7774 13633
rect 6848 13545 6854 13609
rect 6918 13545 6939 13609
rect 7003 13545 7024 13609
rect 7088 13545 7109 13609
rect 7173 13545 7194 13609
rect 7258 13545 7279 13609
rect 7343 13545 7364 13609
rect 7428 13545 7449 13609
rect 7513 13545 7534 13609
rect 7598 13545 7619 13609
rect 7683 13545 7704 13609
rect 7768 13545 7774 13609
rect 6848 13521 7774 13545
rect 6848 13457 6854 13521
rect 6918 13457 6939 13521
rect 7003 13457 7024 13521
rect 7088 13457 7109 13521
rect 7173 13457 7194 13521
rect 7258 13457 7279 13521
rect 7343 13457 7364 13521
rect 7428 13457 7449 13521
rect 7513 13457 7534 13521
rect 7598 13457 7619 13521
rect 7683 13457 7704 13521
rect 7768 13457 7774 13521
rect 6848 13456 7774 13457
rect 16035 13684 16948 13687
rect 16035 13620 16060 13684
rect 16124 13620 16142 13684
rect 16206 13620 16223 13684
rect 16287 13620 16304 13684
rect 16368 13620 16385 13684
rect 16449 13620 16466 13684
rect 16530 13620 16547 13684
rect 16611 13620 16628 13684
rect 16692 13620 16709 13684
rect 16773 13620 16790 13684
rect 16854 13620 16871 13684
rect 16935 13620 16948 13684
rect 16035 13596 16948 13620
rect 16035 13532 16060 13596
rect 16124 13532 16142 13596
rect 16206 13532 16223 13596
rect 16287 13532 16304 13596
rect 16368 13532 16385 13596
rect 16449 13532 16466 13596
rect 16530 13532 16547 13596
rect 16611 13532 16628 13596
rect 16692 13532 16709 13596
rect 16773 13532 16790 13596
rect 16854 13532 16871 13596
rect 16935 13532 16948 13596
rect 16035 13508 16948 13532
rect 16035 13444 16060 13508
rect 16124 13444 16142 13508
rect 16206 13444 16223 13508
rect 16287 13444 16304 13508
rect 16368 13444 16385 13508
rect 16449 13444 16466 13508
rect 16530 13444 16547 13508
rect 16611 13444 16628 13508
rect 16692 13444 16709 13508
rect 16773 13444 16790 13508
rect 16854 13444 16871 13508
rect 16935 13444 16948 13508
rect 16035 13420 16948 13444
rect 16035 13356 16060 13420
rect 16124 13356 16142 13420
rect 16206 13356 16223 13420
rect 16287 13356 16304 13420
rect 16368 13356 16385 13420
rect 16449 13356 16466 13420
rect 16530 13356 16547 13420
rect 16611 13356 16628 13420
rect 16692 13356 16709 13420
rect 16773 13356 16790 13420
rect 16854 13356 16871 13420
rect 16935 13356 16948 13420
rect 16035 13332 16948 13356
rect 16035 13268 16060 13332
rect 16124 13268 16142 13332
rect 16206 13268 16223 13332
rect 16287 13268 16304 13332
rect 16368 13268 16385 13332
rect 16449 13268 16466 13332
rect 16530 13268 16547 13332
rect 16611 13268 16628 13332
rect 16692 13268 16709 13332
rect 16773 13268 16790 13332
rect 16854 13268 16871 13332
rect 16935 13268 16948 13332
rect 16035 13244 16948 13268
rect 16035 13180 16060 13244
rect 16124 13180 16142 13244
rect 16206 13180 16223 13244
rect 16287 13180 16304 13244
rect 16368 13180 16385 13244
rect 16449 13180 16466 13244
rect 16530 13180 16547 13244
rect 16611 13180 16628 13244
rect 16692 13180 16709 13244
rect 16773 13180 16790 13244
rect 16854 13180 16871 13244
rect 16935 13180 16948 13244
rect 16035 13156 16948 13180
rect 16035 13092 16060 13156
rect 16124 13092 16142 13156
rect 16206 13092 16223 13156
rect 16287 13092 16304 13156
rect 16368 13092 16385 13156
rect 16449 13092 16466 13156
rect 16530 13092 16547 13156
rect 16611 13092 16628 13156
rect 16692 13092 16709 13156
rect 16773 13092 16790 13156
rect 16854 13092 16871 13156
rect 16935 13092 16948 13156
rect 16035 13068 16948 13092
rect 16035 13004 16060 13068
rect 16124 13004 16142 13068
rect 16206 13004 16223 13068
rect 16287 13004 16304 13068
rect 16368 13004 16385 13068
rect 16449 13004 16466 13068
rect 16530 13004 16547 13068
rect 16611 13004 16628 13068
rect 16692 13004 16709 13068
rect 16773 13004 16790 13068
rect 16854 13004 16871 13068
rect 16935 13004 16948 13068
rect 16035 12980 16948 13004
rect 16035 12916 16060 12980
rect 16124 12916 16142 12980
rect 16206 12916 16223 12980
rect 16287 12916 16304 12980
rect 16368 12916 16385 12980
rect 16449 12916 16466 12980
rect 16530 12916 16547 12980
rect 16611 12916 16628 12980
rect 16692 12916 16709 12980
rect 16773 12916 16790 12980
rect 16854 12916 16871 12980
rect 16935 12916 16948 12980
rect 16035 12892 16948 12916
rect 16035 12828 16060 12892
rect 16124 12828 16142 12892
rect 16206 12828 16223 12892
rect 16287 12828 16304 12892
rect 16368 12828 16385 12892
rect 16449 12828 16466 12892
rect 16530 12828 16547 12892
rect 16611 12828 16628 12892
rect 16692 12828 16709 12892
rect 16773 12828 16790 12892
rect 16854 12828 16871 12892
rect 16935 12828 16948 12892
rect 15773 11587 15919 11592
rect 15773 11531 15778 11587
rect 15834 11531 15858 11587
rect 15914 11531 15919 11587
rect 15773 11526 15919 11531
rect 14440 11282 14506 11287
rect 14440 11226 14445 11282
rect 14501 11226 14506 11282
rect 14440 11202 14506 11226
rect 14440 11146 14445 11202
rect 14501 11146 14506 11202
tri 14436 10829 14440 10833 se
rect 14440 10829 14506 11146
tri 14400 10793 14436 10829 se
rect 14436 10793 14506 10829
rect 14400 10787 14500 10793
tri 14500 10787 14506 10793 nw
rect 14400 10759 14472 10787
tri 14472 10759 14500 10787 nw
rect 10331 10648 10397 10653
rect 10331 10592 10336 10648
rect 10392 10592 10397 10648
rect 10331 10568 10397 10592
rect 10331 10512 10336 10568
rect 10392 10512 10397 10568
rect 9874 10121 10074 10130
rect 9874 10065 9879 10121
rect 9935 10065 10013 10121
rect 10069 10065 10074 10121
rect 9874 10025 10074 10065
rect 9874 9969 9879 10025
rect 9935 9969 10013 10025
rect 10069 9969 10074 10025
rect 9874 9929 10074 9969
rect 9874 9873 9879 9929
rect 9935 9873 10013 9929
rect 10069 9873 10074 9929
rect 9874 9833 10074 9873
rect 9874 9777 9879 9833
rect 9935 9777 10013 9833
rect 10069 9777 10074 9833
tri 9873 9772 9874 9773 se
rect 9874 9772 10074 9777
tri 9767 9666 9873 9772 se
rect 9873 9666 10074 9772
rect 5206 6701 5216 6757
rect 5272 6701 5307 6757
rect 5363 6701 5397 6757
rect 5453 6701 5487 6757
rect 5543 6701 5555 6757
rect 5206 6619 5555 6701
rect 5206 6563 5216 6619
rect 5272 6563 5307 6619
rect 5363 6563 5397 6619
rect 5453 6563 5487 6619
rect 5543 6563 5555 6619
rect 5206 6558 5555 6563
rect 7436 9087 8036 9105
rect 7436 9023 7446 9087
rect 7510 9023 7532 9087
rect 7596 9023 7618 9087
rect 7682 9023 7704 9087
rect 7768 9023 7790 9087
rect 7854 9023 7876 9087
rect 7940 9023 7962 9087
rect 8026 9023 8036 9087
rect 7436 9001 8036 9023
rect 7436 8937 7446 9001
rect 7510 8937 7532 9001
rect 7596 8937 7618 9001
rect 7682 8937 7704 9001
rect 7768 8937 7790 9001
rect 7854 8937 7876 9001
rect 7940 8937 7962 9001
rect 8026 8937 8036 9001
rect 7436 8915 8036 8937
rect 7436 8851 7446 8915
rect 7510 8851 7532 8915
rect 7596 8851 7618 8915
rect 7682 8851 7704 8915
rect 7768 8851 7790 8915
rect 7854 8851 7876 8915
rect 7940 8851 7962 8915
rect 8026 8851 8036 8915
rect 7436 8829 8036 8851
rect 7436 8765 7446 8829
rect 7510 8765 7532 8829
rect 7596 8765 7618 8829
rect 7682 8765 7704 8829
rect 7768 8765 7790 8829
rect 7854 8765 7876 8829
rect 7940 8765 7962 8829
rect 8026 8765 8036 8829
rect 7436 8743 8036 8765
rect 7436 8679 7446 8743
rect 7510 8679 7532 8743
rect 7596 8679 7618 8743
rect 7682 8679 7704 8743
rect 7768 8679 7790 8743
rect 7854 8679 7876 8743
rect 7940 8679 7962 8743
rect 8026 8679 8036 8743
rect 7436 8657 8036 8679
rect 7436 8593 7446 8657
rect 7510 8593 7532 8657
rect 7596 8593 7618 8657
rect 7682 8593 7704 8657
rect 7768 8593 7790 8657
rect 7854 8593 7876 8657
rect 7940 8593 7962 8657
rect 8026 8593 8036 8657
rect 7436 8571 8036 8593
rect 7436 8507 7446 8571
rect 7510 8507 7532 8571
rect 7596 8507 7618 8571
rect 7682 8507 7704 8571
rect 7768 8507 7790 8571
rect 7854 8507 7876 8571
rect 7940 8507 7962 8571
rect 8026 8507 8036 8571
rect 7436 8484 8036 8507
rect 7436 8420 7446 8484
rect 7510 8420 7532 8484
rect 7596 8420 7618 8484
rect 7682 8420 7704 8484
rect 7768 8420 7790 8484
rect 7854 8420 7876 8484
rect 7940 8420 7962 8484
rect 8026 8420 8036 8484
rect 7436 8397 8036 8420
rect 7436 8333 7446 8397
rect 7510 8333 7532 8397
rect 7596 8333 7618 8397
rect 7682 8333 7704 8397
rect 7768 8333 7790 8397
rect 7854 8333 7876 8397
rect 7940 8333 7962 8397
rect 8026 8333 8036 8397
rect 4427 6450 4575 6455
tri 2313 6381 2318 6386 sw
rect 2252 6376 2318 6381
rect 2252 6320 2257 6376
rect 2313 6320 2318 6376
rect 2920 6347 2934 6403
rect 2990 6347 3058 6403
rect 3114 6347 3182 6403
rect 3238 6347 3249 6403
rect 2920 6339 3249 6347
rect 4142 6399 4288 6404
rect 4142 6343 4147 6399
rect 4203 6343 4227 6399
rect 4283 6343 4288 6399
rect 4142 6338 4288 6343
rect 4427 6394 4434 6450
rect 4490 6394 4514 6450
rect 4570 6394 4575 6450
rect 4427 6389 4575 6394
rect 2252 6296 2318 6320
rect 2252 6240 2257 6296
rect 2313 6240 2318 6296
rect 2252 6235 2318 6240
rect 4427 6166 4493 6389
tri 4493 6335 4547 6389 nw
rect 4427 6110 4432 6166
rect 4488 6110 4493 6166
rect 4427 6086 4493 6110
rect 4427 6030 4432 6086
rect 4488 6030 4493 6086
rect 2169 4994 2175 5058
rect 2239 4994 2255 5058
rect 2319 4994 2325 5058
tri 2169 4953 2210 4994 ne
rect 2210 4953 2284 4994
tri 2284 4953 2325 4994 nw
tri 2210 4945 2218 4953 ne
rect 1921 3639 2053 3645
rect 1921 3575 1955 3639
rect 2019 3575 2053 3639
rect 1921 3556 2053 3575
rect 1921 3492 1955 3556
rect 2019 3492 2053 3556
rect 1921 3473 2053 3492
rect 1921 3409 1955 3473
rect 2019 3409 2053 3473
rect 1921 3390 2053 3409
rect 1921 3326 1955 3390
rect 2019 3326 2053 3390
rect 1921 3307 2053 3326
rect 1921 3243 1955 3307
rect 2019 3243 2053 3307
rect 1921 3224 2053 3243
tri 1816 3167 1819 3170 sw
rect 1753 3162 1819 3167
rect 1753 3106 1758 3162
rect 1814 3106 1819 3162
rect 1753 3082 1819 3106
rect 1753 3026 1758 3082
rect 1814 3026 1819 3082
rect 1753 3021 1819 3026
rect 1921 3160 1955 3224
rect 2019 3160 2053 3224
rect 1921 3141 2053 3160
rect 1921 3077 1955 3141
rect 2019 3077 2053 3141
rect 1921 3057 2053 3077
rect 1921 2993 1955 3057
rect 2019 2993 2053 3057
rect 1586 2814 1592 2878
rect 1656 2814 1672 2878
rect 1736 2814 1742 2878
tri 1586 2793 1607 2814 ne
rect 1607 2793 1721 2814
tri 1721 2793 1742 2814 nw
tri 1607 2777 1623 2793 ne
rect 1623 2777 1705 2793
tri 1705 2777 1721 2793 nw
rect 1623 0 1689 2777
tri 1689 2761 1705 2777 nw
rect 1921 1832 2053 2993
tri 2210 2919 2218 2927 se
rect 2218 2919 2284 4953
tri 3975 3645 3990 3660 se
rect 3990 3645 4056 4573
tri 3967 3637 3975 3645 se
rect 3975 3637 4056 3645
tri 3943 3613 3967 3637 se
rect 3967 3613 4056 3637
tri 3927 3597 3943 3613 se
rect 3943 3597 4000 3613
rect 3927 3557 4000 3597
tri 4000 3557 4056 3613 nw
rect 3337 3494 3847 3503
rect 3337 3198 3347 3494
rect 3643 3198 3847 3494
rect 3337 3173 3847 3198
rect 3337 3117 3347 3173
rect 3403 3117 3427 3173
rect 3483 3117 3507 3173
rect 3563 3117 3587 3173
rect 3643 3117 3847 3173
rect 3337 3092 3847 3117
rect 3337 3036 3347 3092
rect 3403 3036 3427 3092
rect 3483 3036 3507 3092
rect 3563 3036 3587 3092
rect 3643 3036 3847 3092
rect 3337 3011 3847 3036
rect 3337 2955 3347 3011
rect 3403 2955 3427 3011
rect 3483 2955 3507 3011
rect 3563 2955 3587 3011
rect 3643 2955 3847 3011
rect 3337 2930 3847 2955
tri 2169 2878 2210 2919 se
rect 2210 2878 2284 2919
tri 2284 2878 2325 2919 sw
rect 2169 2814 2175 2878
rect 2239 2814 2255 2878
rect 2319 2814 2325 2878
rect 3337 2874 3347 2930
rect 3403 2874 3427 2930
rect 3483 2874 3507 2930
rect 3563 2874 3587 2930
rect 3643 2874 3847 2930
rect 3337 2849 3847 2874
rect 1921 1776 1964 1832
rect 2020 1776 2053 1832
rect 1921 1748 2053 1776
rect 1754 1719 1820 1724
rect 1754 1663 1759 1719
rect 1815 1663 1820 1719
rect 1754 1639 1820 1663
rect 1754 1583 1759 1639
rect 1815 1583 1820 1639
rect 1754 0 1820 1583
rect 1921 1692 1964 1748
rect 2020 1692 2053 1748
rect 1921 1663 2053 1692
rect 1921 1607 1964 1663
rect 2020 1607 2053 1663
rect 1921 1578 2053 1607
rect 1921 1522 1964 1578
rect 2020 1522 2053 1578
rect 1921 1493 2053 1522
rect 1921 1437 1964 1493
rect 2020 1437 2053 1493
rect 1921 1408 2053 1437
rect 1921 1352 1964 1408
rect 2020 1352 2053 1408
rect 1921 1323 2053 1352
rect 1921 1267 1964 1323
rect 2020 1267 2053 1323
rect 1921 1238 2053 1267
rect 1921 1182 1964 1238
rect 2020 1182 2053 1238
rect 1921 1153 2053 1182
rect 1921 1097 1964 1153
rect 2020 1097 2053 1153
rect 1921 1068 2053 1097
rect 1921 1012 1964 1068
rect 2020 1012 2053 1068
rect 1921 983 2053 1012
rect 1921 927 1964 983
rect 2020 927 2053 983
rect 1921 898 2053 927
rect 1921 842 1964 898
rect 2020 842 2053 898
rect 1921 813 2053 842
rect 1921 757 1964 813
rect 2020 757 2053 813
rect 1921 728 2053 757
rect 1921 672 1964 728
rect 2020 672 2053 728
rect 1921 643 2053 672
rect 1921 587 1964 643
rect 2020 587 2053 643
rect 1921 558 2053 587
rect 1921 502 1964 558
rect 2020 502 2053 558
rect 1921 473 2053 502
rect 1921 417 1964 473
rect 2020 417 2053 473
rect 1921 407 2053 417
rect 3337 2793 3347 2849
rect 3403 2793 3427 2849
rect 3483 2793 3507 2849
rect 3563 2793 3587 2849
rect 3643 2793 3847 2849
rect 3337 1491 3847 2793
rect 3337 1427 3340 1491
rect 3404 1427 3428 1491
rect 3492 1427 3516 1491
rect 3580 1427 3604 1491
rect 3668 1427 3692 1491
rect 3756 1427 3780 1491
rect 3844 1427 3847 1491
rect 3337 1407 3847 1427
rect 3337 1343 3340 1407
rect 3404 1343 3428 1407
rect 3492 1343 3516 1407
rect 3580 1343 3604 1407
rect 3668 1343 3692 1407
rect 3756 1343 3780 1407
rect 3844 1343 3847 1407
rect 3337 1323 3847 1343
rect 3337 1259 3340 1323
rect 3404 1259 3428 1323
rect 3492 1259 3516 1323
rect 3580 1259 3604 1323
rect 3668 1259 3692 1323
rect 3756 1259 3780 1323
rect 3844 1259 3847 1323
rect 3337 1239 3847 1259
rect 3337 1175 3340 1239
rect 3404 1175 3428 1239
rect 3492 1175 3516 1239
rect 3580 1175 3604 1239
rect 3668 1175 3692 1239
rect 3756 1175 3780 1239
rect 3844 1175 3847 1239
rect 3337 1155 3847 1175
rect 3337 1091 3340 1155
rect 3404 1091 3428 1155
rect 3492 1091 3516 1155
rect 3580 1091 3604 1155
rect 3668 1091 3692 1155
rect 3756 1091 3780 1155
rect 3844 1091 3847 1155
rect 3337 1071 3847 1091
rect 3337 1007 3340 1071
rect 3404 1007 3428 1071
rect 3492 1007 3516 1071
rect 3580 1007 3604 1071
rect 3668 1007 3692 1071
rect 3756 1007 3780 1071
rect 3844 1007 3847 1071
rect 3337 987 3847 1007
rect 3337 923 3340 987
rect 3404 923 3428 987
rect 3492 923 3516 987
rect 3580 923 3604 987
rect 3668 923 3692 987
rect 3756 923 3780 987
rect 3844 923 3847 987
rect 3337 902 3847 923
rect 3337 838 3340 902
rect 3404 838 3428 902
rect 3492 838 3516 902
rect 3580 838 3604 902
rect 3668 838 3692 902
rect 3756 838 3780 902
rect 3844 838 3847 902
rect 3337 817 3847 838
rect 3337 753 3340 817
rect 3404 753 3428 817
rect 3492 753 3516 817
rect 3580 753 3604 817
rect 3668 753 3692 817
rect 3756 753 3780 817
rect 3844 753 3847 817
rect 3337 732 3847 753
rect 3337 668 3340 732
rect 3404 668 3428 732
rect 3492 668 3516 732
rect 3580 668 3604 732
rect 3668 668 3692 732
rect 3756 668 3780 732
rect 3844 668 3847 732
rect 3337 647 3847 668
rect 3337 583 3340 647
rect 3404 583 3428 647
rect 3492 583 3516 647
rect 3580 583 3604 647
rect 3668 583 3692 647
rect 3756 583 3780 647
rect 3844 583 3847 647
rect 3337 562 3847 583
rect 3337 498 3340 562
rect 3404 498 3428 562
rect 3492 498 3516 562
rect 3580 498 3604 562
rect 3668 498 3692 562
rect 3756 498 3780 562
rect 3844 498 3847 562
rect 3337 477 3847 498
rect 3337 413 3340 477
rect 3404 413 3428 477
rect 3492 413 3516 477
rect 3580 413 3604 477
rect 3668 413 3692 477
rect 3756 413 3780 477
rect 3844 413 3847 477
rect 3337 407 3847 413
rect 3927 0 3993 3557
tri 3993 3550 4000 3557 nw
rect 4076 3046 4142 3055
rect 4076 2990 4081 3046
rect 4137 2990 4142 3046
rect 4076 2966 4142 2990
rect 4076 2910 4081 2966
rect 4137 2910 4142 2966
rect 4076 2885 4142 2910
rect 4076 2829 4081 2885
rect 4137 2829 4142 2885
rect 4076 2804 4142 2829
rect 4076 2748 4081 2804
rect 4137 2748 4142 2804
rect 4076 2723 4142 2748
rect 4076 2667 4081 2723
rect 4137 2667 4142 2723
rect 4076 2642 4142 2667
rect 4076 2586 4081 2642
rect 4137 2586 4142 2642
rect 4076 2561 4142 2586
rect 4076 2505 4081 2561
rect 4137 2505 4142 2561
rect 4076 2480 4142 2505
rect 4076 2424 4081 2480
rect 4137 2424 4142 2480
rect 4076 2399 4142 2424
rect 4076 2343 4081 2399
rect 4137 2343 4142 2399
rect 4076 2318 4142 2343
rect 4076 2262 4081 2318
rect 4137 2262 4142 2318
rect 4076 0 4142 2262
rect 4427 0 4493 6030
rect 5940 6195 6540 6200
rect 5940 6139 5949 6195
rect 6005 6139 6037 6195
rect 6093 6139 6125 6195
rect 6181 6139 6213 6195
rect 6269 6139 6301 6195
rect 6357 6139 6388 6195
rect 6444 6139 6475 6195
rect 6531 6139 6540 6195
rect 5940 6051 6540 6139
rect 5940 5995 5949 6051
rect 6005 5995 6037 6051
rect 6093 5995 6125 6051
rect 6181 5995 6213 6051
rect 6269 5995 6301 6051
rect 6357 5995 6388 6051
rect 6444 5995 6475 6051
rect 6531 5995 6540 6051
rect 5471 4332 5537 4337
rect 5471 4276 5476 4332
rect 5532 4276 5537 4332
rect 5471 4252 5537 4276
rect 5471 4196 5476 4252
rect 5532 4196 5537 4252
tri 5433 3477 5471 3515 se
rect 5471 3487 5537 4196
rect 5471 3477 5527 3487
tri 5527 3477 5537 3487 nw
tri 5409 3453 5433 3477 se
rect 5433 3453 5503 3477
tri 5503 3453 5527 3477 nw
tri 5377 3421 5409 3453 se
rect 5409 3421 5471 3453
tri 5471 3421 5503 3453 nw
tri 5353 3397 5377 3421 se
rect 5377 3397 5447 3421
tri 5447 3397 5471 3421 nw
tri 5329 3373 5353 3397 se
rect 5353 3373 5423 3397
tri 5423 3373 5447 3397 nw
tri 5283 3327 5329 3373 se
rect 5329 3327 5377 3373
tri 5377 3327 5423 3373 nw
tri 5273 3317 5283 3327 se
rect 5283 3317 5367 3327
tri 5367 3317 5377 3327 nw
tri 5240 3284 5273 3317 se
rect 5273 3284 5334 3317
tri 5334 3284 5367 3317 nw
tri 5189 3233 5240 3284 se
rect 5240 3233 5283 3284
tri 5283 3233 5334 3284 nw
tri 5184 3228 5189 3233 se
rect 5189 3228 5278 3233
tri 5278 3228 5283 3233 nw
tri 5179 3223 5184 3228 se
rect 5184 3223 5273 3228
tri 5273 3223 5278 3228 nw
tri 5105 3149 5179 3223 se
rect 5179 3149 5245 3223
tri 5245 3195 5273 3223 nw
tri 5100 3144 5105 3149 se
rect 5105 3144 5245 3149
tri 5089 3133 5100 3144 se
rect 5100 3133 5245 3144
rect 5089 2875 5245 3133
rect 5089 2811 5095 2875
rect 5159 2811 5175 2875
rect 5239 2811 5245 2875
rect 5380 2811 5386 2875
rect 5450 2811 5466 2875
rect 5530 2811 5536 2875
tri 5380 2720 5471 2811 ne
rect 4698 183 4942 188
rect 4698 127 4703 183
rect 4759 127 4783 183
rect 4839 127 4942 183
rect 4698 122 4942 127
tri 4819 65 4876 122 ne
rect 4876 0 4942 122
rect 5471 0 5537 2811
rect 5940 2701 6540 5995
rect 7436 5497 8036 8333
rect 7436 5441 7445 5497
rect 7501 5441 7533 5497
rect 7589 5441 7621 5497
rect 7677 5441 7709 5497
rect 7765 5441 7797 5497
rect 7853 5441 7884 5497
rect 7940 5441 7971 5497
rect 8027 5441 8036 5497
rect 7436 5355 8036 5441
rect 7436 5299 7445 5355
rect 7501 5299 7533 5355
rect 7589 5299 7621 5355
rect 7677 5299 7709 5355
rect 7765 5299 7797 5355
rect 7853 5299 7884 5355
rect 7940 5299 7971 5355
rect 8027 5299 8036 5355
rect 7436 3284 8036 5299
rect 7436 3228 7445 3284
rect 7501 3228 7533 3284
rect 7589 3228 7621 3284
rect 7677 3228 7709 3284
rect 7765 3228 7797 3284
rect 7853 3228 7884 3284
rect 7940 3228 7971 3284
rect 8027 3228 8036 3284
rect 7436 3144 8036 3228
rect 7436 3088 7445 3144
rect 7501 3088 7533 3144
rect 7589 3088 7621 3144
rect 7677 3088 7709 3144
rect 7765 3088 7797 3144
rect 7853 3088 7884 3144
rect 7940 3088 7971 3144
rect 8027 3088 8036 3144
rect 7436 3083 8036 3088
rect 9071 4332 9137 4337
rect 9071 4276 9076 4332
rect 9132 4276 9137 4332
rect 9071 4252 9137 4276
rect 9071 4196 9076 4252
rect 9132 4196 9137 4252
rect 5940 2637 5944 2701
rect 6008 2637 6032 2701
rect 6096 2637 6120 2701
rect 6184 2637 6208 2701
rect 6272 2637 6296 2701
rect 6360 2637 6384 2701
rect 6448 2637 6472 2701
rect 6536 2637 6540 2701
rect 5940 2616 6540 2637
rect 5940 2552 5944 2616
rect 6008 2552 6032 2616
rect 6096 2552 6120 2616
rect 6184 2552 6208 2616
rect 6272 2552 6296 2616
rect 6360 2552 6384 2616
rect 6448 2552 6472 2616
rect 6536 2552 6540 2616
rect 5940 2531 6540 2552
rect 5940 2467 5944 2531
rect 6008 2467 6032 2531
rect 6096 2467 6120 2531
rect 6184 2467 6208 2531
rect 6272 2467 6296 2531
rect 6360 2467 6384 2531
rect 6448 2467 6472 2531
rect 6536 2467 6540 2531
rect 5940 2446 6540 2467
rect 5940 2382 5944 2446
rect 6008 2382 6032 2446
rect 6096 2382 6120 2446
rect 6184 2382 6208 2446
rect 6272 2382 6296 2446
rect 6360 2382 6384 2446
rect 6448 2382 6472 2446
rect 6536 2382 6540 2446
rect 5940 2361 6540 2382
rect 5940 2297 5944 2361
rect 6008 2297 6032 2361
rect 6096 2297 6120 2361
rect 6184 2297 6208 2361
rect 6272 2297 6296 2361
rect 6360 2297 6384 2361
rect 6448 2297 6472 2361
rect 6536 2297 6540 2361
rect 5940 2276 6540 2297
rect 5940 2212 5944 2276
rect 6008 2212 6032 2276
rect 6096 2212 6120 2276
rect 6184 2212 6208 2276
rect 6272 2212 6296 2276
rect 6360 2212 6384 2276
rect 6448 2212 6472 2276
rect 6536 2212 6540 2276
rect 5940 2191 6540 2212
tri 8977 2198 9071 2292 se
rect 9071 2264 9137 4196
tri 9071 2198 9137 2264 nw
rect 9241 4332 9307 4337
rect 9241 4276 9246 4332
rect 9302 4276 9307 4332
rect 9241 4252 9307 4276
rect 9241 4196 9246 4252
rect 9302 4196 9307 4252
rect 5940 2127 5944 2191
rect 6008 2127 6032 2191
rect 6096 2127 6120 2191
rect 6184 2127 6208 2191
rect 6272 2127 6296 2191
rect 6360 2127 6384 2191
rect 6448 2127 6472 2191
rect 6536 2127 6540 2191
rect 5940 2105 6540 2127
rect 5940 2041 5944 2105
rect 6008 2041 6032 2105
rect 6096 2041 6120 2105
rect 6184 2041 6208 2105
rect 6272 2041 6296 2105
rect 6360 2041 6384 2105
rect 6448 2041 6472 2105
rect 6536 2041 6540 2105
tri 8883 2104 8977 2198 se
tri 8977 2104 9071 2198 nw
tri 8839 2060 8883 2104 se
rect 8883 2060 8933 2104
tri 8933 2060 8977 2104 nw
rect 5940 2019 6540 2041
rect 5940 1955 5944 2019
rect 6008 1955 6032 2019
rect 6096 1955 6120 2019
rect 6184 1955 6208 2019
rect 6272 1955 6296 2019
rect 6360 1955 6384 2019
rect 6448 1955 6472 2019
rect 6536 1955 6540 2019
tri 8789 2010 8839 2060 se
rect 8839 2010 8883 2060
tri 8883 2010 8933 2060 nw
tri 8783 2004 8789 2010 se
rect 8789 2004 8877 2010
tri 8877 2004 8883 2010 nw
tri 8747 1968 8783 2004 se
rect 8783 1968 8846 2004
tri 8846 1973 8877 2004 nw
rect 5940 1933 6540 1955
rect 5940 1869 5944 1933
rect 6008 1869 6032 1933
rect 6096 1869 6120 1933
rect 6184 1869 6208 1933
rect 6272 1869 6296 1933
rect 6360 1869 6384 1933
rect 6448 1869 6472 1933
rect 6536 1869 6540 1933
tri 8691 1912 8747 1968 se
rect 8747 1912 8846 1968
rect 5940 1847 6540 1869
rect 5940 1783 5944 1847
rect 6008 1783 6032 1847
rect 6096 1783 6120 1847
rect 6184 1783 6208 1847
rect 6272 1783 6296 1847
rect 6360 1783 6384 1847
rect 6448 1783 6472 1847
rect 6536 1783 6540 1847
rect 5940 1777 6540 1783
tri 8690 1911 8691 1912 se
rect 8691 1911 8846 1912
rect 8690 1676 8846 1911
rect 8690 1612 8696 1676
rect 8760 1612 8776 1676
rect 8840 1612 8846 1676
rect 8981 1612 8987 1676
rect 9051 1612 9067 1676
rect 9131 1612 9137 1676
tri 8981 1522 9071 1612 ne
rect 8807 1033 8953 1038
rect 8807 977 8812 1033
rect 8868 977 8892 1033
rect 8948 977 8953 1033
rect 8807 972 8953 977
rect 8807 0 8873 972
tri 8873 892 8953 972 nw
rect 9071 0 9137 1612
rect 9241 0 9307 4196
rect 9767 3664 10074 9666
rect 9767 3600 9768 3664
rect 9832 3600 9848 3664
rect 9912 3600 9928 3664
rect 9992 3600 10008 3664
rect 10072 3600 10074 3664
rect 9767 3579 10074 3600
rect 9767 3515 9768 3579
rect 9832 3515 9848 3579
rect 9912 3515 9928 3579
rect 9992 3515 10008 3579
rect 10072 3515 10074 3579
rect 9767 3494 10074 3515
rect 9767 3430 9768 3494
rect 9832 3430 9848 3494
rect 9912 3430 9928 3494
rect 9992 3430 10008 3494
rect 10072 3430 10074 3494
rect 9767 3409 10074 3430
rect 9767 3345 9768 3409
rect 9832 3345 9848 3409
rect 9912 3345 9928 3409
rect 9992 3345 10008 3409
rect 10072 3345 10074 3409
rect 9767 3323 10074 3345
rect 9767 3259 9768 3323
rect 9832 3259 9848 3323
rect 9912 3259 9928 3323
rect 9992 3259 10008 3323
rect 10072 3259 10074 3323
rect 9767 3237 10074 3259
rect 9767 3173 9768 3237
rect 9832 3173 9848 3237
rect 9912 3173 9928 3237
rect 9992 3173 10008 3237
rect 10072 3173 10074 3237
rect 9767 3151 10074 3173
rect 9767 3087 9768 3151
rect 9832 3087 9848 3151
rect 9912 3087 9928 3151
rect 9992 3087 10008 3151
rect 10072 3087 10074 3151
rect 9767 3065 10074 3087
rect 9767 3001 9768 3065
rect 9832 3001 9848 3065
rect 9912 3001 9928 3065
rect 9992 3001 10008 3065
rect 10072 3001 10074 3065
rect 9767 2989 10074 3001
rect 10331 2071 10397 10512
rect 11505 9228 12105 9246
rect 11505 9164 11516 9228
rect 11580 9164 11602 9228
rect 11666 9164 11688 9228
rect 11752 9164 11774 9228
rect 11838 9164 11860 9228
rect 11924 9164 11946 9228
rect 12010 9164 12032 9228
rect 12096 9164 12105 9228
rect 11505 9145 12105 9164
rect 11505 9081 11516 9145
rect 11580 9081 11602 9145
rect 11666 9081 11688 9145
rect 11752 9081 11774 9145
rect 11838 9081 11860 9145
rect 11924 9081 11946 9145
rect 12010 9081 12032 9145
rect 12096 9081 12105 9145
rect 11505 9062 12105 9081
rect 11505 8998 11516 9062
rect 11580 8998 11602 9062
rect 11666 8998 11688 9062
rect 11752 8998 11774 9062
rect 11838 8998 11860 9062
rect 11924 8998 11946 9062
rect 12010 8998 12032 9062
rect 12096 8998 12105 9062
rect 11505 8979 12105 8998
rect 11505 8915 11516 8979
rect 11580 8915 11602 8979
rect 11666 8915 11688 8979
rect 11752 8915 11774 8979
rect 11838 8915 11860 8979
rect 11924 8915 11946 8979
rect 12010 8915 12032 8979
rect 12096 8915 12105 8979
rect 11505 8896 12105 8915
rect 11505 8832 11516 8896
rect 11580 8832 11602 8896
rect 11666 8832 11688 8896
rect 11752 8832 11774 8896
rect 11838 8832 11860 8896
rect 11924 8832 11946 8896
rect 12010 8832 12032 8896
rect 12096 8832 12105 8896
rect 11505 8813 12105 8832
rect 11505 8749 11516 8813
rect 11580 8749 11602 8813
rect 11666 8749 11688 8813
rect 11752 8749 11774 8813
rect 11838 8749 11860 8813
rect 11924 8749 11946 8813
rect 12010 8749 12032 8813
rect 12096 8749 12105 8813
rect 11505 8730 12105 8749
rect 11505 8666 11516 8730
rect 11580 8666 11602 8730
rect 11666 8666 11688 8730
rect 11752 8666 11774 8730
rect 11838 8666 11860 8730
rect 11924 8666 11946 8730
rect 12010 8666 12032 8730
rect 12096 8666 12105 8730
rect 11505 8647 12105 8666
rect 11505 8583 11516 8647
rect 11580 8583 11602 8647
rect 11666 8583 11688 8647
rect 11752 8583 11774 8647
rect 11838 8583 11860 8647
rect 11924 8583 11946 8647
rect 12010 8583 12032 8647
rect 12096 8583 12105 8647
rect 11505 8564 12105 8583
rect 11505 8500 11516 8564
rect 11580 8500 11602 8564
rect 11666 8500 11688 8564
rect 11752 8500 11774 8564
rect 11838 8500 11860 8564
rect 11924 8500 11946 8564
rect 12010 8500 12032 8564
rect 12096 8500 12105 8564
rect 11505 8480 12105 8500
rect 11505 8416 11516 8480
rect 11580 8416 11602 8480
rect 11666 8416 11688 8480
rect 11752 8416 11774 8480
rect 11838 8416 11860 8480
rect 11924 8416 11946 8480
rect 12010 8416 12032 8480
rect 12096 8416 12105 8480
rect 11505 8396 12105 8416
rect 11505 8332 11516 8396
rect 11580 8332 11602 8396
rect 11666 8332 11688 8396
rect 11752 8332 11774 8396
rect 11838 8332 11860 8396
rect 11924 8332 11946 8396
rect 12010 8332 12032 8396
rect 12096 8332 12105 8396
rect 11505 5497 12105 8332
rect 11505 5441 11514 5497
rect 11570 5441 11602 5497
rect 11658 5441 11690 5497
rect 11746 5441 11778 5497
rect 11834 5441 11866 5497
rect 11922 5441 11953 5497
rect 12009 5441 12040 5497
rect 12096 5441 12105 5497
rect 11505 5355 12105 5441
rect 11505 5299 11514 5355
rect 11570 5299 11602 5355
rect 11658 5299 11690 5355
rect 11746 5299 11778 5355
rect 11834 5299 11866 5355
rect 11922 5299 11953 5355
rect 12009 5299 12040 5355
rect 12096 5299 12105 5355
rect 11505 3284 12105 5299
rect 11505 3228 11514 3284
rect 11570 3228 11602 3284
rect 11658 3228 11690 3284
rect 11746 3228 11778 3284
rect 11834 3228 11866 3284
rect 11922 3228 11953 3284
rect 12009 3228 12040 3284
rect 12096 3228 12105 3284
rect 11505 3144 12105 3228
rect 11505 3088 11514 3144
rect 11570 3088 11602 3144
rect 11658 3088 11690 3144
rect 11746 3088 11778 3144
rect 11834 3088 11866 3144
rect 11922 3088 11953 3144
rect 12009 3088 12040 3144
rect 12096 3088 12105 3144
rect 11505 3083 12105 3088
rect 12225 6200 12817 10356
rect 13218 10004 13284 10013
rect 13218 9948 13223 10004
rect 13279 9948 13284 10004
rect 13218 9924 13284 9948
rect 13218 9868 13223 9924
rect 13279 9868 13284 9924
tri 13112 9649 13218 9755 se
rect 13218 9715 13284 9868
tri 13218 9649 13284 9715 nw
tri 13047 9584 13112 9649 se
rect 13112 9584 13153 9649
tri 13153 9584 13218 9649 nw
tri 12817 6200 12825 6208 sw
rect 12225 6195 12825 6200
rect 12225 6139 12234 6195
rect 12290 6139 12322 6195
rect 12378 6139 12410 6195
rect 12466 6139 12498 6195
rect 12554 6139 12586 6195
rect 12642 6139 12673 6195
rect 12729 6139 12760 6195
rect 12816 6139 12825 6195
rect 12225 6051 12825 6139
rect 12225 5995 12234 6051
rect 12290 5995 12322 6051
rect 12378 5995 12410 6051
rect 12466 5995 12498 6051
rect 12554 5995 12586 6051
rect 12642 5995 12673 6051
rect 12729 5995 12760 6051
rect 12816 5995 12825 6051
rect 12225 2701 12825 5995
rect 12225 2637 12229 2701
rect 12293 2637 12317 2701
rect 12381 2637 12405 2701
rect 12469 2637 12493 2701
rect 12557 2637 12581 2701
rect 12645 2637 12669 2701
rect 12733 2637 12757 2701
rect 12821 2637 12825 2701
rect 12225 2616 12825 2637
rect 12225 2552 12229 2616
rect 12293 2552 12317 2616
rect 12381 2552 12405 2616
rect 12469 2552 12493 2616
rect 12557 2552 12581 2616
rect 12645 2552 12669 2616
rect 12733 2552 12757 2616
rect 12821 2552 12825 2616
rect 12225 2531 12825 2552
rect 12225 2467 12229 2531
rect 12293 2467 12317 2531
rect 12381 2467 12405 2531
rect 12469 2467 12493 2531
rect 12557 2467 12581 2531
rect 12645 2467 12669 2531
rect 12733 2467 12757 2531
rect 12821 2467 12825 2531
rect 12225 2446 12825 2467
rect 12225 2382 12229 2446
rect 12293 2382 12317 2446
rect 12381 2382 12405 2446
rect 12469 2382 12493 2446
rect 12557 2382 12581 2446
rect 12645 2382 12669 2446
rect 12733 2382 12757 2446
rect 12821 2382 12825 2446
rect 12225 2361 12825 2382
rect 12225 2297 12229 2361
rect 12293 2297 12317 2361
rect 12381 2297 12405 2361
rect 12469 2297 12493 2361
rect 12557 2297 12581 2361
rect 12645 2297 12669 2361
rect 12733 2297 12757 2361
rect 12821 2297 12825 2361
rect 12225 2276 12825 2297
rect 12225 2212 12229 2276
rect 12293 2212 12317 2276
rect 12381 2212 12405 2276
rect 12469 2212 12493 2276
rect 12557 2212 12581 2276
rect 12645 2212 12669 2276
rect 12733 2212 12757 2276
rect 12821 2212 12825 2276
rect 12225 2191 12825 2212
rect 12225 2127 12229 2191
rect 12293 2127 12317 2191
rect 12381 2127 12405 2191
rect 12469 2127 12493 2191
rect 12557 2127 12581 2191
rect 12645 2127 12669 2191
rect 12733 2127 12757 2191
rect 12821 2127 12825 2191
rect 12225 2105 12825 2127
tri 10331 2062 10340 2071 ne
rect 10340 2062 10397 2071
tri 10397 2062 10434 2099 sw
tri 10340 2060 10342 2062 ne
rect 10342 2060 10434 2062
tri 10434 2060 10436 2062 sw
tri 10342 2005 10397 2060 ne
rect 10397 2005 10436 2060
tri 10397 2004 10398 2005 ne
rect 10398 2004 10436 2005
tri 10436 2004 10492 2060 sw
rect 12225 2041 12229 2105
rect 12293 2041 12317 2105
rect 12381 2041 12405 2105
rect 12469 2041 12493 2105
rect 12557 2041 12581 2105
rect 12645 2041 12669 2105
rect 12733 2041 12757 2105
rect 12821 2041 12825 2105
rect 12225 2019 12825 2041
tri 10398 1968 10434 2004 ne
rect 10434 1968 10492 2004
tri 10492 1968 10528 2004 sw
tri 10434 1912 10490 1968 ne
rect 10490 1912 10528 1968
tri 10528 1912 10584 1968 sw
rect 12225 1955 12229 2019
rect 12293 1955 12317 2019
rect 12381 1955 12405 2019
rect 12469 1955 12493 2019
rect 12557 1955 12581 2019
rect 12645 1955 12669 2019
rect 12733 1955 12757 2019
rect 12821 1955 12825 2019
rect 12225 1933 12825 1955
tri 10490 1876 10526 1912 ne
rect 10526 1876 10584 1912
tri 10584 1876 10620 1912 sw
tri 10526 1874 10528 1876 ne
rect 10528 1874 10620 1876
tri 10620 1874 10622 1876 sw
tri 10528 1820 10582 1874 ne
rect 10582 1820 10622 1874
tri 10622 1820 10676 1874 sw
rect 12225 1869 12229 1933
rect 12293 1869 12317 1933
rect 12381 1869 12405 1933
rect 12469 1869 12493 1933
rect 12557 1869 12581 1933
rect 12645 1869 12669 1933
rect 12733 1869 12757 1933
rect 12821 1869 12825 1933
rect 12225 1847 12825 1869
tri 10582 1783 10619 1820 ne
rect 10619 1783 10676 1820
tri 10676 1783 10713 1820 sw
rect 12225 1783 12229 1847
rect 12293 1783 12317 1847
rect 12381 1783 12405 1847
rect 12469 1783 12493 1847
rect 12557 1783 12581 1847
rect 12645 1783 12669 1847
rect 12733 1783 12757 1847
rect 12821 1783 12825 1847
tri 10619 1780 10622 1783 ne
rect 10622 1780 10713 1783
tri 10713 1780 10716 1783 sw
rect 10622 1777 10716 1780
tri 10716 1777 10719 1780 sw
rect 12225 1777 12825 1783
rect 10622 1727 10719 1777
tri 10719 1727 10769 1777 sw
rect 10622 1718 10769 1727
tri 10769 1718 10778 1727 sw
rect 10622 1676 10778 1718
rect 10331 1612 10337 1676
rect 10401 1612 10417 1676
rect 10481 1612 10487 1676
rect 10622 1612 10628 1676
rect 10692 1612 10708 1676
rect 10772 1612 10778 1676
rect 10331 0 10397 1612
tri 10397 1552 10457 1612 nw
tri 12953 626 13047 720 se
rect 13047 692 13113 9584
tri 13113 9544 13153 9584 nw
rect 13307 7933 13373 7938
rect 13307 7877 13312 7933
rect 13368 7877 13373 7933
rect 13307 7853 13373 7877
rect 13307 7797 13312 7853
rect 13368 7797 13373 7853
rect 13307 7792 13373 7797
tri 13283 7472 13307 7496 se
rect 13307 7472 13367 7792
tri 13367 7786 13373 7792 nw
rect 14400 7552 14466 10759
tri 14466 10753 14472 10759 nw
rect 15574 10292 15720 10297
rect 15574 10236 15579 10292
rect 15635 10236 15659 10292
rect 15715 10236 15720 10292
rect 15574 10231 15720 10236
rect 14400 7496 14405 7552
rect 14461 7496 14466 7552
tri 13367 7472 13391 7496 sw
rect 14400 7472 14466 7496
tri 13277 7466 13283 7472 se
rect 13283 7466 13391 7472
tri 13391 7466 13397 7472 sw
rect 13277 7461 13423 7466
rect 13277 7405 13282 7461
rect 13338 7405 13362 7461
rect 13418 7405 13423 7461
rect 14400 7416 14405 7472
rect 14461 7416 14466 7472
rect 14400 7411 14466 7416
rect 14527 9235 15127 9247
rect 14527 9171 14540 9235
rect 14604 9171 14626 9235
rect 14690 9171 14712 9235
rect 14776 9171 14798 9235
rect 14862 9171 14884 9235
rect 14948 9171 14970 9235
rect 15034 9171 15056 9235
rect 15120 9171 15127 9235
rect 14527 9152 15127 9171
rect 14527 9088 14540 9152
rect 14604 9088 14626 9152
rect 14690 9088 14712 9152
rect 14776 9088 14798 9152
rect 14862 9088 14884 9152
rect 14948 9088 14970 9152
rect 15034 9088 15056 9152
rect 15120 9088 15127 9152
rect 14527 9068 15127 9088
rect 14527 9004 14540 9068
rect 14604 9004 14626 9068
rect 14690 9004 14712 9068
rect 14776 9004 14798 9068
rect 14862 9004 14884 9068
rect 14948 9004 14970 9068
rect 15034 9004 15056 9068
rect 15120 9004 15127 9068
rect 14527 8984 15127 9004
rect 14527 8920 14540 8984
rect 14604 8920 14626 8984
rect 14690 8920 14712 8984
rect 14776 8920 14798 8984
rect 14862 8920 14884 8984
rect 14948 8920 14970 8984
rect 15034 8920 15056 8984
rect 15120 8920 15127 8984
rect 14527 8900 15127 8920
rect 14527 8836 14540 8900
rect 14604 8836 14626 8900
rect 14690 8836 14712 8900
rect 14776 8836 14798 8900
rect 14862 8836 14884 8900
rect 14948 8836 14970 8900
rect 15034 8836 15056 8900
rect 15120 8836 15127 8900
rect 14527 8816 15127 8836
rect 14527 8752 14540 8816
rect 14604 8752 14626 8816
rect 14690 8752 14712 8816
rect 14776 8752 14798 8816
rect 14862 8752 14884 8816
rect 14948 8752 14970 8816
rect 15034 8752 15056 8816
rect 15120 8752 15127 8816
rect 14527 8732 15127 8752
rect 14527 8668 14540 8732
rect 14604 8668 14626 8732
rect 14690 8668 14712 8732
rect 14776 8668 14798 8732
rect 14862 8668 14884 8732
rect 14948 8668 14970 8732
rect 15034 8668 15056 8732
rect 15120 8668 15127 8732
rect 14527 8648 15127 8668
rect 14527 8584 14540 8648
rect 14604 8584 14626 8648
rect 14690 8584 14712 8648
rect 14776 8584 14798 8648
rect 14862 8584 14884 8648
rect 14948 8584 14970 8648
rect 15034 8584 15056 8648
rect 15120 8584 15127 8648
rect 14527 8564 15127 8584
rect 14527 8500 14540 8564
rect 14604 8500 14626 8564
rect 14690 8500 14712 8564
rect 14776 8500 14798 8564
rect 14862 8500 14884 8564
rect 14948 8500 14970 8564
rect 15034 8500 15056 8564
rect 15120 8500 15127 8564
rect 14527 8480 15127 8500
rect 14527 8416 14540 8480
rect 14604 8416 14626 8480
rect 14690 8416 14712 8480
rect 14776 8416 14798 8480
rect 14862 8416 14884 8480
rect 14948 8416 14970 8480
rect 15034 8416 15056 8480
rect 15120 8416 15127 8480
rect 14527 8396 15127 8416
rect 14527 8332 14540 8396
rect 14604 8332 14626 8396
rect 14690 8332 14712 8396
rect 14776 8332 14798 8396
rect 14862 8332 14884 8396
rect 14948 8332 14970 8396
rect 15034 8332 15056 8396
rect 15120 8332 15127 8396
rect 13277 7400 13423 7405
rect 14527 5497 15127 8332
tri 15623 6829 15635 6841 se
rect 15635 6829 15701 10231
tri 15615 6821 15623 6829 se
rect 15623 6821 15701 6829
rect 15813 6965 15879 11526
rect 16035 11235 16948 12828
tri 16035 10996 16274 11235 ne
rect 15813 6909 15818 6965
rect 15874 6909 15879 6965
rect 15813 6885 15879 6909
rect 15813 6829 15818 6885
rect 15874 6829 15879 6885
rect 15813 6824 15879 6829
rect 16274 7061 16948 11235
rect 20127 11496 20515 11529
rect 20127 11440 20132 11496
rect 20188 11440 20213 11496
rect 20269 11440 20294 11496
rect 20350 11440 20374 11496
rect 20430 11440 20454 11496
rect 20510 11440 20515 11496
rect 17879 10885 18184 10890
rect 17879 10829 17884 10885
rect 17940 10829 18004 10885
rect 18060 10829 18123 10885
rect 18179 10829 18184 10885
rect 17879 10759 18184 10829
rect 17879 10703 17884 10759
rect 17940 10703 18004 10759
rect 18060 10703 18123 10759
rect 18179 10703 18184 10759
rect 17879 9239 18184 10703
rect 17879 9175 17880 9239
rect 17944 9175 17960 9239
rect 18024 9175 18040 9239
rect 18104 9175 18120 9239
rect 17879 9154 18184 9175
rect 17879 9090 17880 9154
rect 17944 9090 17960 9154
rect 18024 9090 18040 9154
rect 18104 9090 18120 9154
rect 17879 9069 18184 9090
rect 17879 9005 17880 9069
rect 17944 9005 17960 9069
rect 18024 9005 18040 9069
rect 18104 9005 18120 9069
rect 17879 8984 18184 9005
rect 17879 8920 17880 8984
rect 17944 8920 17960 8984
rect 18024 8920 18040 8984
rect 18104 8920 18120 8984
rect 17879 8899 18184 8920
rect 17879 8835 17880 8899
rect 17944 8835 17960 8899
rect 18024 8835 18040 8899
rect 18104 8835 18120 8899
rect 17879 8814 18184 8835
rect 17879 8750 17880 8814
rect 17944 8750 17960 8814
rect 18024 8750 18040 8814
rect 18104 8750 18120 8814
rect 17879 8729 18184 8750
rect 17879 8665 17880 8729
rect 17944 8665 17960 8729
rect 18024 8665 18040 8729
rect 18104 8665 18120 8729
rect 17879 8644 18184 8665
rect 17879 8580 17880 8644
rect 17944 8580 17960 8644
rect 18024 8580 18040 8644
rect 18104 8580 18120 8644
rect 17879 8559 18184 8580
rect 17879 8495 17880 8559
rect 17944 8495 17960 8559
rect 18024 8495 18040 8559
rect 18104 8495 18120 8559
rect 17879 8474 18184 8495
rect 17879 8410 17880 8474
rect 17944 8410 17960 8474
rect 18024 8410 18040 8474
rect 18104 8410 18120 8474
rect 17879 8388 18184 8410
rect 17879 8324 17880 8388
rect 17944 8324 17960 8388
rect 18024 8324 18040 8388
rect 18104 8324 18120 8388
rect 17879 8317 18184 8324
rect 20127 9239 20515 11440
rect 20127 9175 20130 9239
rect 20194 9175 20210 9239
rect 20274 9175 20290 9239
rect 20354 9175 20370 9239
rect 20434 9175 20450 9239
rect 20514 9175 20515 9239
rect 20127 9154 20515 9175
rect 20127 9090 20130 9154
rect 20194 9090 20210 9154
rect 20274 9090 20290 9154
rect 20354 9090 20370 9154
rect 20434 9090 20450 9154
rect 20514 9090 20515 9154
rect 20127 9069 20515 9090
rect 20127 9005 20130 9069
rect 20194 9005 20210 9069
rect 20274 9005 20290 9069
rect 20354 9005 20370 9069
rect 20434 9005 20450 9069
rect 20514 9005 20515 9069
rect 20127 8984 20515 9005
rect 20127 8920 20130 8984
rect 20194 8920 20210 8984
rect 20274 8920 20290 8984
rect 20354 8920 20370 8984
rect 20434 8920 20450 8984
rect 20514 8920 20515 8984
rect 20127 8899 20515 8920
rect 20127 8835 20130 8899
rect 20194 8835 20210 8899
rect 20274 8835 20290 8899
rect 20354 8835 20370 8899
rect 20434 8835 20450 8899
rect 20514 8835 20515 8899
rect 20127 8814 20515 8835
rect 20127 8750 20130 8814
rect 20194 8750 20210 8814
rect 20274 8750 20290 8814
rect 20354 8750 20370 8814
rect 20434 8750 20450 8814
rect 20514 8750 20515 8814
rect 20127 8729 20515 8750
rect 20127 8665 20130 8729
rect 20194 8665 20210 8729
rect 20274 8665 20290 8729
rect 20354 8665 20370 8729
rect 20434 8665 20450 8729
rect 20514 8665 20515 8729
rect 20127 8644 20515 8665
rect 20127 8580 20130 8644
rect 20194 8580 20210 8644
rect 20274 8580 20290 8644
rect 20354 8580 20370 8644
rect 20434 8580 20450 8644
rect 20514 8580 20515 8644
rect 20127 8559 20515 8580
rect 20127 8495 20130 8559
rect 20194 8495 20210 8559
rect 20274 8495 20290 8559
rect 20354 8495 20370 8559
rect 20434 8495 20450 8559
rect 20514 8495 20515 8559
rect 20127 8474 20515 8495
rect 20127 8410 20130 8474
rect 20194 8410 20210 8474
rect 20274 8410 20290 8474
rect 20354 8410 20370 8474
rect 20434 8410 20450 8474
rect 20514 8410 20515 8474
rect 20127 8388 20515 8410
rect 20127 8324 20130 8388
rect 20194 8324 20210 8388
rect 20274 8324 20290 8388
rect 20354 8324 20370 8388
rect 20434 8324 20450 8388
rect 20514 8324 20515 8388
rect 20127 8317 20515 8324
rect 22389 8123 22944 8128
rect 22389 8067 22394 8123
rect 22450 8067 22476 8123
rect 22532 8067 22558 8123
rect 22614 8067 22640 8123
rect 22696 8067 22721 8123
rect 22777 8067 22802 8123
rect 22858 8067 22883 8123
rect 22939 8067 22944 8123
rect 22389 7999 22944 8067
rect 22389 7943 22394 7999
rect 22450 7943 22476 7999
rect 22532 7943 22558 7999
rect 22614 7943 22640 7999
rect 22696 7943 22721 7999
rect 22777 7943 22802 7999
rect 22858 7943 22883 7999
rect 22939 7943 22944 7999
tri 16948 7061 17053 7166 sw
rect 16274 6877 17053 7061
tri 17053 6877 17237 7061 sw
rect 21869 7055 22305 7061
rect 21869 6991 21871 7055
rect 21935 6991 21963 7055
rect 22027 6991 22055 7055
rect 22119 6991 22147 7055
rect 22211 6991 22239 7055
rect 22303 6991 22305 7055
rect 21869 6969 22305 6991
rect 21869 6905 21871 6969
rect 21935 6905 21963 6969
rect 22027 6905 22055 6969
rect 22119 6905 22147 6969
rect 22211 6905 22239 6969
rect 22303 6905 22305 6969
rect 21869 6883 22305 6905
tri 15606 6812 15615 6821 se
rect 15615 6812 15701 6821
tri 15591 6797 15606 6812 se
rect 15606 6797 15686 6812
tri 15686 6797 15701 6812 nw
rect 16274 6821 17237 6877
tri 17237 6821 17293 6877 sw
rect 16274 6812 17293 6821
tri 17293 6812 17302 6821 sw
tri 15590 6796 15591 6797 se
rect 15591 6796 15656 6797
rect 15590 6293 15656 6796
tri 15656 6767 15686 6797 nw
rect 16274 6756 17302 6812
tri 16274 6741 16289 6756 ne
rect 16289 6741 17302 6756
tri 16289 6381 16649 6741 ne
rect 16649 6381 17302 6741
rect 21869 6819 21871 6883
rect 21935 6819 21963 6883
rect 22027 6819 22055 6883
rect 22119 6819 22147 6883
rect 22211 6819 22239 6883
rect 22303 6819 22305 6883
rect 21869 6797 22305 6819
rect 21869 6733 21871 6797
rect 21935 6733 21963 6797
rect 22027 6733 22055 6797
rect 22119 6733 22147 6797
rect 22211 6733 22239 6797
rect 22303 6733 22305 6797
rect 21869 6711 22305 6733
rect 21869 6647 21871 6711
rect 21935 6647 21963 6711
rect 22027 6647 22055 6711
rect 22119 6647 22147 6711
rect 22211 6647 22239 6711
rect 22303 6647 22305 6711
rect 21869 6625 22305 6647
rect 21869 6561 21871 6625
rect 21935 6561 21963 6625
rect 22027 6561 22055 6625
rect 22119 6561 22147 6625
rect 22211 6561 22239 6625
rect 22303 6561 22305 6625
rect 21869 6538 22305 6561
rect 21869 6474 21871 6538
rect 21935 6474 21963 6538
rect 22027 6474 22055 6538
rect 22119 6474 22147 6538
rect 22211 6474 22239 6538
rect 22303 6474 22305 6538
rect 21869 6451 22305 6474
rect 21869 6387 21871 6451
rect 21935 6387 21963 6451
rect 22027 6387 22055 6451
rect 22119 6387 22147 6451
rect 22211 6387 22239 6451
rect 22303 6387 22305 6451
rect 21869 6381 22305 6387
tri 16649 6323 16707 6381 ne
rect 16707 6323 17302 6381
tri 16707 6322 16708 6323 ne
rect 16708 6322 17302 6323
tri 15590 6277 15606 6293 ne
rect 15606 6277 15656 6293
tri 15656 6277 15701 6322 sw
tri 16708 6277 16753 6322 ne
rect 16753 6277 17302 6322
tri 15606 6270 15613 6277 ne
rect 15613 6270 15701 6277
tri 15613 6248 15635 6270 ne
rect 14527 5441 14536 5497
rect 14592 5441 14617 5497
rect 14673 5441 14698 5497
rect 14754 5441 14779 5497
rect 14835 5441 14860 5497
rect 14916 5441 14941 5497
rect 14997 5441 15127 5497
rect 14527 5355 15127 5441
rect 14527 5299 14536 5355
rect 14592 5299 14617 5355
rect 14673 5299 14698 5355
rect 14754 5299 14779 5355
rect 14835 5299 14860 5355
rect 14916 5299 14941 5355
rect 14997 5299 15127 5355
tri 13047 626 13113 692 nw
rect 13217 4332 13283 4337
rect 13217 4276 13222 4332
rect 13278 4276 13283 4332
rect 13217 4252 13283 4276
rect 13217 4196 13222 4252
rect 13278 4196 13283 4252
tri 12859 532 12953 626 se
tri 12953 532 13047 626 nw
tri 12839 512 12859 532 se
rect 12859 512 12933 532
tri 12933 512 12953 532 nw
tri 12783 456 12839 512 se
rect 12839 456 12877 512
tri 12877 456 12933 512 nw
tri 12765 438 12783 456 se
rect 12783 438 12859 456
tri 12859 438 12877 456 nw
tri 12745 418 12765 438 se
rect 12765 418 12839 438
tri 12839 418 12859 438 nw
tri 12737 410 12745 418 se
rect 12745 410 12831 418
tri 12831 410 12839 418 nw
tri 12718 391 12737 410 se
rect 12737 391 12822 410
tri 12822 401 12831 410 nw
tri 12666 339 12718 391 se
rect 12718 339 12822 391
rect 12666 297 12822 339
rect 12666 233 12672 297
rect 12736 233 12752 297
rect 12816 233 12822 297
rect 12957 233 12963 297
rect 13027 233 13043 297
rect 13107 233 13113 297
tri 12997 193 13037 233 ne
rect 13037 193 13113 233
tri 13037 183 13047 193 ne
rect 13047 0 13113 193
rect 13217 0 13283 4196
rect 13387 4332 13453 4337
rect 13387 4276 13392 4332
rect 13448 4276 13453 4332
rect 13387 4252 13453 4276
rect 13387 4196 13392 4252
rect 13448 4196 13453 4252
rect 13387 0 13453 4196
rect 14527 3284 15127 5299
rect 14527 3228 14536 3284
rect 14592 3228 14624 3284
rect 14680 3228 14712 3284
rect 14768 3228 14800 3284
rect 14856 3228 14888 3284
rect 14944 3228 14975 3284
rect 15031 3228 15062 3284
rect 15118 3228 15127 3284
rect 14527 3144 15127 3228
rect 14527 3088 14536 3144
rect 14592 3088 14624 3144
rect 14680 3088 14712 3144
rect 14768 3088 14800 3144
rect 14856 3088 14888 3144
rect 14944 3088 14975 3144
rect 15031 3088 15062 3144
rect 15118 3088 15127 3144
rect 14527 3083 15127 3088
rect 15635 6214 15640 6270
rect 15696 6214 15701 6270
tri 16753 6267 16763 6277 ne
rect 16763 6267 17302 6277
tri 16763 6264 16766 6267 ne
rect 15635 6190 15701 6214
rect 15635 6134 15640 6190
rect 15696 6134 15701 6190
tri 15556 2973 15635 3052 se
rect 15635 2973 15701 6134
rect 14825 2907 15701 2973
rect 16057 6195 16657 6200
rect 16057 6139 16079 6195
rect 16135 6139 16165 6195
rect 16221 6139 16251 6195
rect 16307 6139 16337 6195
rect 16393 6139 16422 6195
rect 16478 6139 16507 6195
rect 16563 6139 16592 6195
rect 16648 6139 16657 6195
rect 16057 6051 16657 6139
rect 16057 5995 16079 6051
rect 16135 5995 16165 6051
rect 16221 5995 16251 6051
rect 16307 5995 16337 6051
rect 16393 5995 16422 6051
rect 16478 5995 16507 6051
rect 16563 5995 16592 6051
rect 16648 5995 16657 6051
rect 14825 0 14891 2907
tri 14891 2828 14970 2907 nw
rect 16057 2701 16657 5995
rect 16057 2637 16061 2701
rect 16125 2637 16149 2701
rect 16213 2637 16237 2701
rect 16301 2637 16325 2701
rect 16389 2637 16413 2701
rect 16477 2637 16501 2701
rect 16565 2637 16589 2701
rect 16653 2637 16657 2701
rect 16057 2616 16657 2637
rect 16057 2552 16061 2616
rect 16125 2552 16149 2616
rect 16213 2552 16237 2616
rect 16301 2552 16325 2616
rect 16389 2552 16413 2616
rect 16477 2552 16501 2616
rect 16565 2552 16589 2616
rect 16653 2552 16657 2616
rect 16057 2531 16657 2552
rect 16057 2467 16061 2531
rect 16125 2467 16149 2531
rect 16213 2467 16237 2531
rect 16301 2467 16325 2531
rect 16389 2467 16413 2531
rect 16477 2467 16501 2531
rect 16565 2467 16589 2531
rect 16653 2467 16657 2531
rect 16057 2446 16657 2467
rect 16057 2382 16061 2446
rect 16125 2382 16149 2446
rect 16213 2382 16237 2446
rect 16301 2382 16325 2446
rect 16389 2382 16413 2446
rect 16477 2382 16501 2446
rect 16565 2382 16589 2446
rect 16653 2382 16657 2446
rect 16057 2361 16657 2382
rect 16057 2297 16061 2361
rect 16125 2297 16149 2361
rect 16213 2297 16237 2361
rect 16301 2297 16325 2361
rect 16389 2297 16413 2361
rect 16477 2297 16501 2361
rect 16565 2297 16589 2361
rect 16653 2297 16657 2361
rect 16057 2276 16657 2297
rect 16057 2212 16061 2276
rect 16125 2212 16149 2276
rect 16213 2212 16237 2276
rect 16301 2212 16325 2276
rect 16389 2212 16413 2276
rect 16477 2212 16501 2276
rect 16565 2212 16589 2276
rect 16653 2212 16657 2276
rect 16057 2191 16657 2212
rect 16057 2127 16061 2191
rect 16125 2127 16149 2191
rect 16213 2127 16237 2191
rect 16301 2127 16325 2191
rect 16389 2127 16413 2191
rect 16477 2127 16501 2191
rect 16565 2127 16589 2191
rect 16653 2127 16657 2191
rect 16057 2105 16657 2127
rect 16057 2041 16061 2105
rect 16125 2041 16149 2105
rect 16213 2041 16237 2105
rect 16301 2041 16325 2105
rect 16389 2041 16413 2105
rect 16477 2041 16501 2105
rect 16565 2041 16589 2105
rect 16653 2041 16657 2105
rect 16057 2019 16657 2041
rect 16057 1955 16061 2019
rect 16125 1955 16149 2019
rect 16213 1955 16237 2019
rect 16301 1955 16325 2019
rect 16389 1955 16413 2019
rect 16477 1955 16501 2019
rect 16565 1955 16589 2019
rect 16653 1955 16657 2019
rect 16057 1933 16657 1955
rect 16057 1869 16061 1933
rect 16125 1869 16149 1933
rect 16213 1869 16237 1933
rect 16301 1869 16325 1933
rect 16389 1869 16413 1933
rect 16477 1869 16501 1933
rect 16565 1869 16589 1933
rect 16653 1869 16657 1933
rect 16057 1847 16657 1869
rect 16057 1783 16061 1847
rect 16125 1783 16149 1847
rect 16213 1783 16237 1847
rect 16301 1783 16325 1847
rect 16389 1783 16413 1847
rect 16477 1783 16501 1847
rect 16565 1783 16589 1847
rect 16653 1783 16657 1847
rect 16057 1777 16657 1783
rect 16766 4600 17302 6267
rect 16766 4544 16899 4600
rect 16955 4544 17012 4600
rect 17068 4544 17125 4600
rect 17181 4544 17302 4600
rect 16766 4520 17302 4544
rect 16766 4464 16899 4520
rect 16955 4464 17012 4520
rect 17068 4464 17125 4520
rect 17181 4464 17302 4520
rect 16766 4440 17302 4464
rect 16766 4384 16899 4440
rect 16955 4384 17012 4440
rect 17068 4384 17125 4440
rect 17181 4384 17302 4440
rect 16766 4360 17302 4384
rect 16766 4304 16899 4360
rect 16955 4304 17012 4360
rect 17068 4304 17125 4360
rect 17181 4304 17302 4360
rect 20292 6195 20892 6200
rect 20292 6139 20301 6195
rect 20357 6139 20389 6195
rect 20445 6139 20477 6195
rect 20533 6139 20565 6195
rect 20621 6139 20653 6195
rect 20709 6139 20740 6195
rect 20796 6139 20827 6195
rect 20883 6139 20892 6195
rect 20292 6051 20892 6139
rect 20292 5995 20301 6051
rect 20357 5995 20389 6051
rect 20445 5995 20477 6051
rect 20533 5995 20565 6051
rect 20621 5995 20653 6051
rect 20709 5995 20740 6051
rect 20796 5995 20827 6051
rect 20883 5995 20892 6051
rect 16766 4280 17302 4304
rect 16766 4224 16899 4280
rect 16955 4224 17012 4280
rect 17068 4224 17125 4280
rect 17181 4224 17302 4280
rect 16766 193 17302 4224
rect 16766 137 16778 193
rect 16834 137 16871 193
rect 16927 137 16964 193
rect 17020 137 17057 193
rect 17113 137 17149 193
rect 17205 137 17241 193
rect 17297 137 17302 193
rect 16766 63 17302 137
rect 16766 7 16778 63
rect 16834 7 16871 63
rect 16927 7 16964 63
rect 17020 7 17057 63
rect 17113 7 17149 63
rect 17205 7 17241 63
rect 17297 7 17302 63
rect 16766 0 17302 7
rect 17363 4332 17429 4337
rect 17363 4276 17368 4332
rect 17424 4276 17429 4332
rect 17363 4252 17429 4276
rect 17363 4196 17368 4252
rect 17424 4196 17429 4252
rect 17363 0 17429 4196
rect 17533 4332 17599 4337
rect 17533 4276 17538 4332
rect 17594 4276 17599 4332
rect 17533 4252 17599 4276
rect 17533 4196 17538 4252
rect 17594 4196 17599 4252
rect 17533 0 17599 4196
rect 18259 3279 18535 3284
rect 18259 3223 18269 3279
rect 18325 3223 18368 3279
rect 18424 3223 18466 3279
rect 18522 3223 18535 3279
rect 18259 3149 18535 3223
rect 18259 3093 18269 3149
rect 18325 3093 18368 3149
rect 18424 3093 18466 3149
rect 18522 3093 18535 3149
rect 17775 1491 18175 1497
rect 17839 1427 17859 1491
rect 17923 1427 17943 1491
rect 18007 1427 18027 1491
rect 18091 1427 18111 1491
rect 17775 1407 18175 1427
rect 17839 1343 17859 1407
rect 17923 1343 17943 1407
rect 18007 1343 18027 1407
rect 18091 1343 18111 1407
rect 17775 1323 18175 1343
rect 17839 1259 17859 1323
rect 17923 1259 17943 1323
rect 18007 1259 18027 1323
rect 18091 1259 18111 1323
rect 17775 1239 18175 1259
rect 17839 1175 17859 1239
rect 17923 1175 17943 1239
rect 18007 1175 18027 1239
rect 18091 1175 18111 1239
rect 17775 1155 18175 1175
rect 17839 1091 17859 1155
rect 17923 1091 17943 1155
rect 18007 1091 18027 1155
rect 18091 1091 18111 1155
rect 17775 1071 18175 1091
rect 17839 1007 17859 1071
rect 17923 1007 17943 1071
rect 18007 1007 18027 1071
rect 18091 1007 18111 1071
rect 17775 987 18175 1007
rect 17839 923 17859 987
rect 17923 923 17943 987
rect 18007 923 18027 987
rect 18091 923 18111 987
rect 17775 902 18175 923
rect 17839 838 17859 902
rect 17923 838 17943 902
rect 18007 838 18027 902
rect 18091 838 18111 902
rect 17775 817 18175 838
rect 17839 753 17859 817
rect 17923 753 17943 817
rect 18007 753 18027 817
rect 18091 753 18111 817
rect 17775 732 18175 753
rect 17839 668 17859 732
rect 17923 668 17943 732
rect 18007 668 18027 732
rect 18091 668 18111 732
rect 17775 647 18175 668
rect 17839 583 17859 647
rect 17923 583 17943 647
rect 18007 583 18027 647
rect 18091 583 18111 647
rect 17775 562 18175 583
rect 17839 498 17859 562
rect 17923 498 17943 562
rect 18007 498 18027 562
rect 18091 498 18111 562
rect 17775 477 18175 498
rect 17839 413 17859 477
rect 17923 413 17943 477
rect 18007 413 18027 477
rect 18091 413 18111 477
rect 17775 391 18175 413
rect 17775 335 17784 391
rect 17840 335 17866 391
rect 17922 335 17948 391
rect 18004 335 18029 391
rect 18085 335 18110 391
rect 18166 335 18175 391
rect 18259 410 18535 3093
rect 20292 2701 20892 5995
rect 21511 4332 21577 4337
rect 21511 4276 21516 4332
rect 21572 4276 21577 4332
rect 21511 4252 21577 4276
rect 21511 4196 21516 4252
rect 21572 4196 21577 4252
rect 21511 4191 21577 4196
rect 21675 4332 21741 4337
rect 21675 4276 21680 4332
rect 21736 4276 21741 4332
rect 21675 4252 21741 4276
rect 21675 4196 21680 4252
rect 21736 4196 21741 4252
rect 20292 2637 20296 2701
rect 20360 2637 20384 2701
rect 20448 2637 20472 2701
rect 20536 2637 20560 2701
rect 20624 2637 20648 2701
rect 20712 2637 20736 2701
rect 20800 2637 20824 2701
rect 20888 2637 20892 2701
rect 20292 2616 20892 2637
rect 20292 2552 20296 2616
rect 20360 2552 20384 2616
rect 20448 2552 20472 2616
rect 20536 2552 20560 2616
rect 20624 2552 20648 2616
rect 20712 2552 20736 2616
rect 20800 2552 20824 2616
rect 20888 2552 20892 2616
rect 20292 2531 20892 2552
rect 20292 2467 20296 2531
rect 20360 2467 20384 2531
rect 20448 2467 20472 2531
rect 20536 2467 20560 2531
rect 20624 2467 20648 2531
rect 20712 2467 20736 2531
rect 20800 2467 20824 2531
rect 20888 2467 20892 2531
rect 20292 2446 20892 2467
rect 20292 2382 20296 2446
rect 20360 2382 20384 2446
rect 20448 2382 20472 2446
rect 20536 2382 20560 2446
rect 20624 2382 20648 2446
rect 20712 2382 20736 2446
rect 20800 2382 20824 2446
rect 20888 2382 20892 2446
rect 20292 2361 20892 2382
rect 20292 2297 20296 2361
rect 20360 2297 20384 2361
rect 20448 2297 20472 2361
rect 20536 2297 20560 2361
rect 20624 2297 20648 2361
rect 20712 2297 20736 2361
rect 20800 2297 20824 2361
rect 20888 2297 20892 2361
rect 20292 2276 20892 2297
rect 20292 2212 20296 2276
rect 20360 2212 20384 2276
rect 20448 2212 20472 2276
rect 20536 2212 20560 2276
rect 20624 2212 20648 2276
rect 20712 2212 20736 2276
rect 20800 2212 20824 2276
rect 20888 2212 20892 2276
rect 20292 2191 20892 2212
rect 20292 2127 20296 2191
rect 20360 2127 20384 2191
rect 20448 2127 20472 2191
rect 20536 2127 20560 2191
rect 20624 2127 20648 2191
rect 20712 2127 20736 2191
rect 20800 2127 20824 2191
rect 20888 2127 20892 2191
rect 20292 2105 20892 2127
rect 20292 2041 20296 2105
rect 20360 2041 20384 2105
rect 20448 2041 20472 2105
rect 20536 2041 20560 2105
rect 20624 2041 20648 2105
rect 20712 2041 20736 2105
rect 20800 2041 20824 2105
rect 20888 2041 20892 2105
tri 21470 2060 21509 2099 se
rect 21509 2071 21575 4191
rect 21675 4128 21741 4196
rect 21675 4056 21745 4128
rect 21509 2060 21564 2071
tri 21564 2060 21575 2071 nw
rect 20292 2019 20892 2041
rect 20292 1955 20296 2019
rect 20360 1955 20384 2019
rect 20448 1955 20472 2019
rect 20536 1955 20560 2019
rect 20624 1955 20648 2019
rect 20712 1955 20736 2019
rect 20800 1955 20824 2019
rect 20888 1955 20892 2019
tri 21415 2005 21470 2060 se
rect 21470 2005 21509 2060
tri 21509 2005 21564 2060 nw
tri 21414 2004 21415 2005 se
rect 21415 2004 21508 2005
tri 21508 2004 21509 2005 nw
tri 21378 1968 21414 2004 se
rect 21414 1968 21472 2004
tri 21472 1968 21508 2004 nw
rect 20292 1933 20892 1955
rect 20292 1869 20296 1933
rect 20360 1869 20384 1933
rect 20448 1869 20472 1933
rect 20536 1869 20560 1933
rect 20624 1869 20648 1933
rect 20712 1869 20736 1933
rect 20800 1869 20824 1933
rect 20888 1869 20892 1933
tri 21322 1912 21378 1968 se
rect 21378 1912 21416 1968
tri 21416 1912 21472 1968 nw
tri 21321 1911 21322 1912 se
rect 21322 1911 21415 1912
tri 21415 1911 21416 1912 nw
tri 21286 1876 21321 1911 se
rect 21321 1876 21380 1911
tri 21380 1876 21415 1911 nw
rect 20292 1847 20892 1869
rect 20292 1783 20296 1847
rect 20360 1783 20384 1847
rect 20448 1783 20472 1847
rect 20536 1783 20560 1847
rect 20624 1783 20648 1847
rect 20712 1783 20736 1847
rect 20800 1783 20824 1847
rect 20888 1783 20892 1847
tri 21230 1820 21286 1876 se
rect 21286 1820 21324 1876
tri 21324 1820 21380 1876 nw
tri 21227 1817 21230 1820 se
rect 21230 1817 21321 1820
tri 21321 1817 21324 1820 nw
tri 21193 1783 21227 1817 se
rect 21227 1783 21287 1817
tri 21287 1783 21321 1817 nw
rect 20292 1777 20892 1783
tri 21187 1777 21193 1783 se
rect 21193 1777 21284 1783
tri 21284 1780 21287 1783 nw
tri 21137 1727 21187 1777 se
rect 21187 1727 21284 1777
tri 21128 1718 21137 1727 se
rect 21137 1718 21284 1727
rect 21128 1676 21284 1718
rect 21128 1612 21134 1676
rect 21198 1612 21214 1676
rect 21278 1612 21284 1676
rect 21419 1612 21425 1676
rect 21489 1612 21505 1676
rect 21569 1612 21575 1676
tri 21456 1559 21509 1612 ne
rect 18259 354 18268 410
rect 18324 354 18367 410
rect 18423 354 18465 410
rect 18521 354 18535 410
rect 18259 338 18535 354
rect 17775 294 18175 335
rect 19169 0 19243 348
rect 21509 0 21575 1612
rect 21679 0 21745 4056
tri 22276 1494 22389 1607 se
rect 22389 1494 22944 7943
rect 22276 1488 22944 1494
rect 22276 1424 22281 1488
rect 22345 1424 22365 1488
rect 22429 1424 22449 1488
rect 22513 1424 22533 1488
rect 22597 1424 22617 1488
rect 22681 1424 22701 1488
rect 22765 1424 22785 1488
rect 22849 1424 22869 1488
rect 22933 1424 22944 1488
rect 22276 1405 22944 1424
rect 22276 1341 22281 1405
rect 22345 1341 22365 1405
rect 22429 1341 22449 1405
rect 22513 1341 22533 1405
rect 22597 1341 22617 1405
rect 22681 1341 22701 1405
rect 22765 1341 22785 1405
rect 22849 1341 22869 1405
rect 22933 1341 22944 1405
rect 22276 1322 22944 1341
rect 22276 1258 22281 1322
rect 22345 1258 22365 1322
rect 22429 1258 22449 1322
rect 22513 1258 22533 1322
rect 22597 1258 22617 1322
rect 22681 1258 22701 1322
rect 22765 1258 22785 1322
rect 22849 1258 22869 1322
rect 22933 1258 22944 1322
rect 22276 1238 22944 1258
rect 22276 1174 22281 1238
rect 22345 1174 22365 1238
rect 22429 1174 22449 1238
rect 22513 1174 22533 1238
rect 22597 1174 22617 1238
rect 22681 1174 22701 1238
rect 22765 1174 22785 1238
rect 22849 1174 22869 1238
rect 22933 1174 22944 1238
rect 22276 1154 22944 1174
rect 22276 1090 22281 1154
rect 22345 1090 22365 1154
rect 22429 1090 22449 1154
rect 22513 1090 22533 1154
rect 22597 1090 22617 1154
rect 22681 1090 22701 1154
rect 22765 1090 22785 1154
rect 22849 1090 22869 1154
rect 22933 1090 22944 1154
rect 22276 1070 22944 1090
rect 22276 1006 22281 1070
rect 22345 1006 22365 1070
rect 22429 1006 22449 1070
rect 22513 1006 22533 1070
rect 22597 1006 22617 1070
rect 22681 1006 22701 1070
rect 22765 1006 22785 1070
rect 22849 1006 22869 1070
rect 22933 1006 22944 1070
rect 22276 986 22944 1006
rect 22276 922 22281 986
rect 22345 922 22365 986
rect 22429 922 22449 986
rect 22513 922 22533 986
rect 22597 922 22617 986
rect 22681 922 22701 986
rect 22765 922 22785 986
rect 22849 922 22869 986
rect 22933 922 22944 986
rect 22276 902 22944 922
rect 22276 838 22281 902
rect 22345 838 22365 902
rect 22429 838 22449 902
rect 22513 838 22533 902
rect 22597 838 22617 902
rect 22681 838 22701 902
rect 22765 838 22785 902
rect 22849 838 22869 902
rect 22933 838 22944 902
rect 22276 818 22944 838
rect 22276 754 22281 818
rect 22345 754 22365 818
rect 22429 754 22449 818
rect 22513 754 22533 818
rect 22597 754 22617 818
rect 22681 754 22701 818
rect 22765 754 22785 818
rect 22849 754 22869 818
rect 22933 754 22944 818
rect 22276 734 22944 754
rect 22276 670 22281 734
rect 22345 670 22365 734
rect 22429 670 22449 734
rect 22513 670 22533 734
rect 22597 670 22617 734
rect 22681 670 22701 734
rect 22765 670 22785 734
rect 22849 670 22869 734
rect 22933 670 22944 734
rect 22276 650 22944 670
rect 22276 586 22281 650
rect 22345 586 22365 650
rect 22429 586 22449 650
rect 22513 586 22533 650
rect 22597 586 22617 650
rect 22681 586 22701 650
rect 22765 586 22785 650
rect 22849 586 22869 650
rect 22933 586 22944 650
rect 22276 566 22944 586
rect 22276 502 22281 566
rect 22345 502 22365 566
rect 22429 502 22449 566
rect 22513 502 22533 566
rect 22597 502 22617 566
rect 22681 502 22701 566
rect 22765 502 22785 566
rect 22849 502 22869 566
rect 22933 502 22944 566
rect 22276 482 22944 502
rect 22276 418 22281 482
rect 22345 418 22365 482
rect 22429 418 22449 482
rect 22513 418 22533 482
rect 22597 418 22617 482
rect 22681 418 22701 482
rect 22765 418 22785 482
rect 22849 418 22869 482
rect 22933 418 22944 482
rect 22276 412 22944 418
rect 23058 0 23178 22113
rect 26092 22041 26228 22187
tri 26130 22038 26133 22041 ne
rect 26133 22038 26228 22041
tri 26133 22009 26162 22038 ne
rect 23849 18991 23987 18997
rect 23849 18927 23886 18991
rect 23950 18927 23987 18991
rect 23849 18910 23987 18927
rect 23849 18846 23886 18910
rect 23950 18846 23987 18910
rect 23849 18829 23987 18846
rect 23849 18765 23886 18829
rect 23950 18765 23987 18829
rect 23849 18748 23987 18765
rect 23849 18684 23886 18748
rect 23950 18684 23987 18748
rect 23849 18666 23987 18684
rect 23849 18602 23886 18666
rect 23950 18602 23987 18666
rect 23849 18584 23987 18602
rect 23849 18520 23886 18584
rect 23950 18520 23987 18584
rect 23849 18502 23987 18520
rect 23849 18438 23886 18502
rect 23950 18438 23987 18502
rect 23849 18420 23987 18438
rect 23849 18356 23886 18420
rect 23950 18356 23987 18420
rect 23849 18338 23987 18356
rect 23849 18274 23886 18338
rect 23950 18274 23987 18338
rect 23849 18256 23987 18274
rect 23849 18192 23886 18256
rect 23950 18192 23987 18256
rect 23849 18174 23987 18192
rect 23849 18110 23886 18174
rect 23950 18110 23987 18174
rect 23849 18092 23987 18110
rect 23849 18028 23886 18092
rect 23950 18028 23987 18092
rect 23849 18010 23987 18028
rect 23849 17946 23886 18010
rect 23950 17946 23987 18010
rect 23849 17928 23987 17946
rect 23849 17864 23886 17928
rect 23950 17864 23987 17928
rect 23849 17846 23987 17864
rect 23849 17782 23886 17846
rect 23950 17782 23987 17846
rect 23849 17764 23987 17782
rect 23849 17700 23886 17764
rect 23950 17700 23987 17764
rect 23849 17682 23987 17700
rect 23849 17618 23886 17682
rect 23950 17618 23987 17682
rect 23849 17600 23987 17618
rect 23849 17536 23886 17600
rect 23950 17536 23987 17600
rect 23849 17518 23987 17536
rect 23849 17454 23886 17518
rect 23950 17454 23987 17518
rect 23849 17436 23987 17454
rect 23849 17372 23886 17436
rect 23950 17372 23987 17436
rect 23849 17354 23987 17372
rect 23849 17290 23886 17354
rect 23950 17290 23987 17354
rect 23849 17272 23987 17290
rect 23849 17208 23886 17272
rect 23950 17208 23987 17272
rect 23849 17190 23987 17208
rect 23849 17126 23886 17190
rect 23950 17126 23987 17190
rect 23849 17108 23987 17126
rect 23849 17044 23886 17108
rect 23950 17044 23987 17108
rect 23849 17026 23987 17044
rect 23849 16962 23886 17026
rect 23950 16962 23987 17026
rect 23849 16944 23987 16962
rect 23849 16880 23886 16944
rect 23950 16880 23987 16944
rect 23849 16862 23987 16880
rect 23849 16798 23886 16862
rect 23950 16798 23987 16862
rect 23849 16780 23987 16798
rect 23849 16716 23886 16780
rect 23950 16716 23987 16780
rect 23849 16698 23987 16716
rect 23849 16634 23886 16698
rect 23950 16634 23987 16698
rect 23849 16616 23987 16634
rect 23849 16552 23886 16616
rect 23950 16552 23987 16616
rect 23849 16546 23987 16552
rect 23246 14121 23454 14135
rect 23246 14065 23254 14121
rect 23310 14065 23392 14121
rect 23448 14065 23454 14121
rect 23246 14024 23454 14065
rect 23246 13968 23254 14024
rect 23310 13968 23392 14024
rect 23448 13968 23454 14024
rect 23246 13926 23454 13968
rect 23246 13870 23254 13926
rect 23310 13870 23392 13926
rect 23448 13870 23454 13926
rect 23246 13828 23454 13870
rect 23246 13772 23254 13828
rect 23310 13772 23392 13828
rect 23448 13772 23454 13828
rect 23246 2060 23454 13772
rect 24550 13698 24945 13707
rect 24550 13634 24565 13698
rect 24629 13634 24667 13698
rect 24731 13634 24769 13698
rect 24833 13634 24871 13698
rect 24935 13634 24945 13698
rect 24550 13618 24945 13634
rect 24550 13554 24565 13618
rect 24629 13554 24667 13618
rect 24731 13554 24769 13618
rect 24833 13554 24871 13618
rect 24935 13554 24945 13618
rect 24550 13538 24945 13554
rect 24550 13474 24565 13538
rect 24629 13474 24667 13538
rect 24731 13474 24769 13538
rect 24833 13474 24871 13538
rect 24935 13474 24945 13538
rect 24550 13458 24945 13474
rect 24550 13394 24565 13458
rect 24629 13394 24667 13458
rect 24731 13394 24769 13458
rect 24833 13394 24871 13458
rect 24935 13394 24945 13458
rect 24550 13378 24945 13394
rect 24550 13314 24565 13378
rect 24629 13314 24667 13378
rect 24731 13314 24769 13378
rect 24833 13314 24871 13378
rect 24935 13314 24945 13378
rect 24550 13298 24945 13314
rect 24550 13234 24565 13298
rect 24629 13234 24667 13298
rect 24731 13234 24769 13298
rect 24833 13234 24871 13298
rect 24935 13234 24945 13298
rect 24550 13218 24945 13234
rect 24550 13154 24565 13218
rect 24629 13154 24667 13218
rect 24731 13154 24769 13218
rect 24833 13154 24871 13218
rect 24935 13154 24945 13218
rect 24550 13138 24945 13154
rect 24550 13074 24565 13138
rect 24629 13074 24667 13138
rect 24731 13074 24769 13138
rect 24833 13074 24871 13138
rect 24935 13074 24945 13138
rect 24550 13058 24945 13074
rect 24550 12994 24565 13058
rect 24629 12994 24667 13058
rect 24731 12994 24769 13058
rect 24833 12994 24871 13058
rect 24935 12994 24945 13058
rect 24550 12978 24945 12994
rect 24550 12914 24565 12978
rect 24629 12914 24667 12978
rect 24731 12914 24769 12978
rect 24833 12914 24871 12978
rect 24935 12914 24945 12978
rect 24550 12898 24945 12914
rect 23777 12717 24177 12869
rect 23777 12661 23786 12717
rect 23842 12661 23868 12717
rect 23924 12661 23950 12717
rect 24006 12661 24031 12717
rect 24087 12661 24112 12717
rect 24168 12661 24177 12717
rect 23246 2004 23251 2060
rect 23307 2004 23393 2060
rect 23449 2004 23454 2060
rect 23246 1968 23454 2004
rect 23246 1912 23251 1968
rect 23307 1912 23393 1968
rect 23449 1912 23454 1968
rect 23246 1876 23454 1912
rect 23246 1820 23251 1876
rect 23307 1820 23393 1876
rect 23449 1820 23454 1876
rect 23246 1783 23454 1820
rect 23246 1727 23251 1783
rect 23307 1727 23393 1783
rect 23449 1727 23454 1783
rect 23246 1715 23454 1727
rect 23514 1238 23717 9248
rect 23777 8023 24177 12661
rect 24550 12834 24565 12898
rect 24629 12834 24667 12898
rect 24731 12834 24769 12898
rect 24833 12834 24871 12898
rect 24935 12834 24945 12898
rect 24550 10843 24945 12834
tri 26058 12394 26162 12498 se
rect 26162 12460 26228 22038
rect 27340 22146 27345 22202
rect 27401 22146 27483 22202
rect 27539 22146 27544 22202
rect 27340 22120 27544 22146
rect 27340 22064 27345 22120
rect 27401 22064 27483 22120
rect 27539 22064 27544 22120
rect 27340 22038 27544 22064
rect 27340 21982 27345 22038
rect 27401 21982 27483 22038
rect 27539 21982 27544 22038
rect 27340 21956 27544 21982
rect 27340 21900 27345 21956
rect 27401 21900 27483 21956
rect 27539 21900 27544 21956
rect 27340 21874 27544 21900
rect 27340 21818 27345 21874
rect 27401 21818 27483 21874
rect 27539 21818 27544 21874
rect 27340 21792 27544 21818
rect 27340 21736 27345 21792
rect 27401 21736 27483 21792
rect 27539 21736 27544 21792
rect 27340 21710 27544 21736
rect 27340 21654 27345 21710
rect 27401 21654 27483 21710
rect 27539 21654 27544 21710
rect 27340 21628 27544 21654
rect 27340 21572 27345 21628
rect 27401 21572 27483 21628
rect 27539 21572 27544 21628
rect 27340 21546 27544 21572
rect 27340 21490 27345 21546
rect 27401 21490 27483 21546
rect 27539 21490 27544 21546
rect 27340 21464 27544 21490
rect 27340 21408 27345 21464
rect 27401 21408 27483 21464
rect 27539 21408 27544 21464
rect 27340 21382 27544 21408
rect 27340 21326 27345 21382
rect 27401 21326 27483 21382
rect 27539 21326 27544 21382
rect 27340 21299 27544 21326
rect 27340 21243 27345 21299
rect 27401 21243 27483 21299
rect 27539 21243 27544 21299
rect 27340 21216 27544 21243
rect 27340 21160 27345 21216
rect 27401 21160 27483 21216
rect 27539 21160 27544 21216
rect 27340 21155 27544 21160
tri 26162 12394 26228 12460 nw
rect 24550 10787 24599 10843
rect 24655 10787 24679 10843
rect 24735 10787 24759 10843
rect 24815 10787 24839 10843
rect 24895 10787 24945 10843
rect 24550 10758 24945 10787
rect 24550 10702 24599 10758
rect 24655 10702 24679 10758
rect 24735 10702 24759 10758
rect 24815 10702 24839 10758
rect 24895 10702 24945 10758
rect 24550 10673 24945 10702
rect 24550 10617 24599 10673
rect 24655 10617 24679 10673
rect 24735 10617 24759 10673
rect 24815 10617 24839 10673
rect 24895 10617 24945 10673
rect 24550 10588 24945 10617
rect 24550 10532 24599 10588
rect 24655 10532 24679 10588
rect 24735 10532 24759 10588
rect 24815 10532 24839 10588
rect 24895 10532 24945 10588
rect 24550 10502 24945 10532
rect 24550 10446 24599 10502
rect 24655 10446 24679 10502
rect 24735 10446 24759 10502
rect 24815 10446 24839 10502
rect 24895 10446 24945 10502
rect 24550 10416 24945 10446
rect 24550 10360 24599 10416
rect 24655 10360 24679 10416
rect 24735 10360 24759 10416
rect 24815 10360 24839 10416
rect 24895 10360 24945 10416
rect 24550 10350 24945 10360
tri 25995 12331 26058 12394 se
rect 26058 12331 26099 12394
tri 26099 12331 26162 12394 nw
rect 25280 9381 25346 9386
rect 25280 9325 25285 9381
rect 25341 9325 25346 9381
rect 25280 9301 25346 9325
rect 25280 9245 25285 9301
rect 25341 9245 25346 9301
rect 25280 9240 25346 9245
rect 23777 7959 23784 8023
rect 23848 7959 23890 8023
rect 23954 7959 23996 8023
rect 24060 7959 24102 8023
rect 24166 7959 24177 8023
rect 23777 7939 24177 7959
rect 23777 7875 23784 7939
rect 23848 7875 23890 7939
rect 23954 7875 23996 7939
rect 24060 7875 24102 7939
rect 24166 7875 24177 7939
rect 23777 7854 24177 7875
rect 23777 7790 23784 7854
rect 23848 7790 23890 7854
rect 23954 7790 23996 7854
rect 24060 7790 24102 7854
rect 24166 7790 24177 7854
rect 23777 7769 24177 7790
rect 23777 7705 23784 7769
rect 23848 7705 23890 7769
rect 23954 7705 23996 7769
rect 24060 7705 24102 7769
rect 24166 7705 24177 7769
rect 23777 7684 24177 7705
rect 23777 7620 23784 7684
rect 23848 7620 23890 7684
rect 23954 7620 23996 7684
rect 24060 7620 24102 7684
rect 24166 7620 24177 7684
rect 23777 7599 24177 7620
rect 23777 7535 23784 7599
rect 23848 7535 23890 7599
rect 23954 7535 23996 7599
rect 24060 7535 24102 7599
rect 24166 7535 24177 7599
rect 23777 7514 24177 7535
rect 23777 7450 23784 7514
rect 23848 7450 23890 7514
rect 23954 7450 23996 7514
rect 24060 7450 24102 7514
rect 24166 7450 24177 7514
rect 23777 7443 24177 7450
rect 23981 6323 24047 6328
rect 23981 6267 23986 6323
rect 24042 6284 24047 6323
tri 24047 6284 24079 6316 sw
tri 24744 6284 24776 6316 se
rect 24776 6284 24842 6316
rect 24042 6267 24842 6284
rect 23981 6243 24842 6267
rect 23981 6187 23986 6243
rect 24042 6224 24842 6243
rect 24042 6187 24047 6224
tri 24047 6189 24082 6224 nw
rect 23981 6182 24047 6187
tri 24889 6102 24902 6115 se
rect 24902 6102 24968 6284
rect 24889 6080 24968 6102
tri 24777 3892 24889 4004 se
rect 24889 3939 24955 6080
tri 24955 6067 24968 6080 nw
rect 24889 3892 24908 3939
tri 24908 3892 24955 3939 nw
rect 24777 3865 24881 3892
tri 24881 3865 24908 3892 nw
rect 24777 3862 24878 3865
tri 24878 3862 24881 3865 nw
tri 25025 3862 25028 3865 se
rect 25028 3862 25094 6278
rect 25154 5966 25220 6261
rect 25280 4201 25346 6261
rect 25280 4145 25285 4201
rect 25341 4145 25346 4201
rect 25280 4121 25346 4145
rect 25280 4065 25285 4121
rect 25341 4065 25346 4121
rect 25280 4060 25346 4065
rect 25659 4332 25725 4337
rect 25659 4276 25664 4332
rect 25720 4276 25725 4332
rect 25659 4252 25725 4276
rect 25659 4196 25664 4252
rect 25720 4196 25725 4252
rect 24777 2364 24843 3862
tri 24843 3827 24878 3862 nw
tri 24990 3827 25025 3862 se
rect 25025 3827 25094 3862
tri 24969 3806 24990 3827 se
rect 24990 3806 25094 3827
tri 24960 3797 24969 3806 se
rect 24969 3797 25085 3806
tri 25085 3797 25094 3806 nw
tri 25655 4036 25659 4040 se
rect 25659 4036 25725 4196
rect 25821 4332 25887 4337
rect 25821 4276 25826 4332
rect 25882 4276 25887 4332
rect 25821 4252 25887 4276
rect 25821 4196 25826 4252
rect 25882 4196 25887 4252
rect 25821 4191 25887 4196
rect 25655 3979 25725 4036
tri 24945 3782 24960 3797 se
rect 24960 3782 25070 3797
tri 25070 3782 25085 3797 nw
tri 24916 3753 24945 3782 se
rect 24945 3753 25014 3782
rect 24916 3726 25014 3753
tri 25014 3726 25070 3782 nw
rect 24916 3717 25005 3726
tri 25005 3717 25014 3726 nw
rect 24916 2430 24982 3717
tri 24982 3694 25005 3717 nw
tri 24916 2393 24953 2430 ne
rect 24953 2393 24982 2430
tri 24982 2393 25094 2505 sw
tri 24953 2366 24980 2393 ne
rect 24980 2366 25094 2393
tri 24843 2364 24845 2366 sw
tri 24980 2364 24982 2366 ne
rect 24982 2364 25094 2366
rect 24777 2320 24845 2364
tri 24845 2320 24889 2364 sw
tri 24982 2320 25026 2364 ne
rect 25026 2320 25094 2364
rect 24777 2318 24889 2320
tri 24889 2318 24891 2320 sw
tri 25026 2318 25028 2320 ne
rect 24777 2298 24891 2318
tri 24891 2298 24911 2318 sw
tri 24777 2186 24889 2298 ne
rect 24889 2254 24911 2298
tri 24911 2254 24955 2298 sw
tri 24795 2005 24889 2099 se
rect 24889 2071 24955 2254
tri 24889 2005 24955 2071 nw
tri 24701 1911 24795 2005 se
tri 24795 1911 24889 2005 nw
tri 24607 1817 24701 1911 se
tri 24701 1817 24795 1911 nw
tri 24508 1718 24607 1817 se
rect 24607 1718 24664 1817
tri 24664 1780 24701 1817 nw
rect 24508 1676 24664 1718
rect 24508 1612 24514 1676
rect 24578 1612 24594 1676
rect 24658 1612 24664 1676
rect 24799 1612 24805 1676
rect 24869 1612 24885 1676
rect 24949 1612 24955 1676
tri 24841 1564 24889 1612 ne
rect 23514 1182 23524 1238
rect 23580 1182 23650 1238
rect 23706 1182 23717 1238
rect 23514 1144 23717 1182
rect 23514 1088 23524 1144
rect 23580 1088 23650 1144
rect 23706 1088 23717 1144
rect 23514 512 23717 1088
rect 23514 456 23524 512
rect 23580 456 23650 512
rect 23706 456 23717 512
rect 23514 418 23717 456
rect 23514 362 23524 418
rect 23580 362 23650 418
rect 23706 362 23717 418
rect 23514 358 23717 362
rect 23519 357 23711 358
rect 24889 0 24955 1612
rect 25028 0 25094 2320
rect 25655 0 25721 3979
tri 25721 3975 25725 3979 nw
rect 25825 0 25891 4191
rect 25995 0 26061 12331
tri 26061 12293 26099 12331 nw
rect 27238 9043 27544 9048
rect 27238 8987 27243 9043
rect 27299 8987 27323 9043
rect 27379 8987 27403 9043
rect 27459 8987 27483 9043
rect 27539 8987 27544 9043
rect 27238 8954 27544 8987
rect 27238 8898 27243 8954
rect 27299 8898 27323 8954
rect 27379 8898 27403 8954
rect 27459 8898 27483 8954
rect 27539 8898 27544 8954
rect 27238 8865 27544 8898
rect 27238 8809 27243 8865
rect 27299 8809 27323 8865
rect 27379 8809 27403 8865
rect 27459 8809 27483 8865
rect 27539 8809 27544 8865
rect 27238 8776 27544 8809
rect 27238 8720 27243 8776
rect 27299 8720 27323 8776
rect 27379 8720 27403 8776
rect 27459 8720 27483 8776
rect 27539 8720 27544 8776
rect 27238 8686 27544 8720
rect 27238 8630 27243 8686
rect 27299 8630 27323 8686
rect 27379 8630 27403 8686
rect 27459 8630 27483 8686
rect 27539 8630 27544 8686
rect 27238 8625 27544 8630
rect 26159 6877 26225 6882
rect 26159 6821 26164 6877
rect 26220 6821 26225 6877
rect 26159 6797 26225 6821
rect 26159 6741 26164 6797
rect 26220 6741 26225 6797
rect 26159 3862 26225 6741
rect 26159 3806 26164 3862
rect 26220 3806 26225 3862
rect 26159 3782 26225 3806
rect 26159 3726 26164 3782
rect 26220 3726 26225 3782
rect 26159 3721 26225 3726
rect 26288 3613 26354 6216
rect 26288 3557 26293 3613
rect 26349 3557 26354 3613
rect 26288 3533 26354 3557
rect 26288 3477 26293 3533
rect 26349 3477 26354 3533
rect 26288 3468 26354 3477
rect 26414 3533 26480 6216
rect 26414 3477 26419 3533
rect 26475 3477 26480 3533
rect 26414 3453 26480 3477
rect 26414 3397 26419 3453
rect 26475 3397 26480 3453
rect 26414 3388 26480 3397
rect 26540 3453 26606 6216
rect 26666 3853 26732 6216
rect 26666 3797 26671 3853
rect 26727 3797 26732 3853
rect 26666 3773 26732 3797
rect 26666 3717 26671 3773
rect 26727 3717 26732 3773
rect 26666 3707 26732 3717
rect 26792 3773 26858 6216
rect 26792 3717 26797 3773
rect 26853 3717 26858 3773
rect 26792 3693 26858 3717
rect 26792 3637 26797 3693
rect 26853 3637 26858 3693
rect 26792 3632 26858 3637
rect 26918 3693 26984 6216
rect 26918 3637 26923 3693
rect 26979 3637 26984 3693
rect 26918 3613 26984 3637
rect 26918 3557 26923 3613
rect 26979 3557 26984 3613
rect 26918 3548 26984 3557
rect 26540 3397 26545 3453
rect 26601 3397 26606 3453
rect 26540 3373 26606 3397
rect 26540 3317 26545 3373
rect 26601 3317 26606 3373
rect 26540 3308 26606 3317
rect 27652 2692 27988 2698
rect 27652 2628 27653 2692
rect 27717 2628 27743 2692
rect 27807 2628 27833 2692
rect 27897 2628 27923 2692
rect 27987 2628 27988 2692
rect 27652 2608 27988 2628
rect 27652 2544 27653 2608
rect 27717 2544 27743 2608
rect 27807 2544 27833 2608
rect 27897 2544 27923 2608
rect 27987 2544 27988 2608
rect 27652 2524 27988 2544
rect 27652 2460 27653 2524
rect 27717 2460 27743 2524
rect 27807 2460 27833 2524
rect 27897 2460 27923 2524
rect 27987 2460 27988 2524
rect 27652 2440 27988 2460
rect 27652 2376 27653 2440
rect 27717 2376 27743 2440
rect 27807 2376 27833 2440
rect 27897 2376 27923 2440
rect 27987 2376 27988 2440
rect 27652 2356 27988 2376
rect 27652 2292 27653 2356
rect 27717 2292 27743 2356
rect 27807 2292 27833 2356
rect 27897 2292 27923 2356
rect 27987 2292 27988 2356
rect 27652 2272 27988 2292
rect 27652 2208 27653 2272
rect 27717 2208 27743 2272
rect 27807 2208 27833 2272
rect 27897 2208 27923 2272
rect 27987 2208 27988 2272
rect 27652 2188 27988 2208
rect 27652 2124 27653 2188
rect 27717 2124 27743 2188
rect 27807 2124 27833 2188
rect 27897 2124 27923 2188
rect 27987 2124 27988 2188
rect 27652 2104 27988 2124
rect 27652 2040 27653 2104
rect 27717 2040 27743 2104
rect 27807 2040 27833 2104
rect 27897 2040 27923 2104
rect 27987 2040 27988 2104
rect 27652 2020 27988 2040
rect 27652 1956 27653 2020
rect 27717 1956 27743 2020
rect 27807 1956 27833 2020
rect 27897 1956 27923 2020
rect 27987 1956 27988 2020
rect 27652 1936 27988 1956
rect 27652 1872 27653 1936
rect 27717 1872 27743 1936
rect 27807 1872 27833 1936
rect 27897 1872 27923 1936
rect 27987 1872 27988 1936
rect 27652 1851 27988 1872
rect 27652 1787 27653 1851
rect 27717 1787 27743 1851
rect 27807 1787 27833 1851
rect 27897 1787 27923 1851
rect 27987 1787 27988 1851
rect 27652 1781 27988 1787
<< via3 >>
rect 23396 36183 23460 36247
rect 23514 36183 23578 36247
rect 23632 36183 23696 36247
rect 23396 36100 23460 36164
rect 23514 36100 23578 36164
rect 23632 36100 23696 36164
rect 23396 36017 23460 36081
rect 23514 36017 23578 36081
rect 23632 36017 23696 36081
rect 23396 35934 23460 35998
rect 23514 35934 23578 35998
rect 23632 35934 23696 35998
rect 23396 35851 23460 35915
rect 23514 35851 23578 35915
rect 23632 35851 23696 35915
rect 23396 35768 23460 35832
rect 23514 35768 23578 35832
rect 23632 35768 23696 35832
rect 23396 35685 23460 35749
rect 23514 35685 23578 35749
rect 23632 35685 23696 35749
rect 19258 35562 19322 35626
rect 19340 35562 19404 35626
rect 19422 35562 19486 35626
rect 19504 35562 19568 35626
rect 19586 35562 19650 35626
rect 19668 35562 19732 35626
rect 19750 35562 19814 35626
rect 19832 35562 19896 35626
rect 19914 35562 19978 35626
rect 19996 35562 20060 35626
rect 20078 35562 20142 35626
rect 20160 35562 20224 35626
rect 20242 35562 20306 35626
rect 20324 35562 20388 35626
rect 20406 35562 20470 35626
rect 20488 35562 20552 35626
rect 20570 35562 20634 35626
rect 20652 35562 20716 35626
rect 20734 35562 20798 35626
rect 20816 35562 20880 35626
rect 20898 35562 20962 35626
rect 20980 35562 21044 35626
rect 21062 35562 21126 35626
rect 21144 35562 21208 35626
rect 21226 35562 21290 35626
rect 21308 35562 21372 35626
rect 21390 35562 21454 35626
rect 21472 35562 21536 35626
rect 21553 35562 21617 35626
rect 21634 35562 21698 35626
rect 21715 35562 21779 35626
rect 21796 35562 21860 35626
rect 21877 35562 21941 35626
rect 21958 35562 22022 35626
rect 22039 35562 22103 35626
rect 22120 35562 22184 35626
rect 22201 35562 22265 35626
rect 22282 35562 22346 35626
rect 22363 35562 22427 35626
rect 22444 35562 22508 35626
rect 22525 35562 22589 35626
rect 19258 35482 19322 35546
rect 19340 35482 19404 35546
rect 19422 35482 19486 35546
rect 19504 35482 19568 35546
rect 19586 35482 19650 35546
rect 19668 35482 19732 35546
rect 19750 35482 19814 35546
rect 19832 35482 19896 35546
rect 19914 35482 19978 35546
rect 19996 35482 20060 35546
rect 20078 35482 20142 35546
rect 20160 35482 20224 35546
rect 20242 35482 20306 35546
rect 20324 35482 20388 35546
rect 20406 35482 20470 35546
rect 20488 35482 20552 35546
rect 20570 35482 20634 35546
rect 20652 35482 20716 35546
rect 20734 35482 20798 35546
rect 20816 35482 20880 35546
rect 20898 35482 20962 35546
rect 20980 35482 21044 35546
rect 21062 35482 21126 35546
rect 21144 35482 21208 35546
rect 21226 35482 21290 35546
rect 21308 35482 21372 35546
rect 21390 35482 21454 35546
rect 21472 35482 21536 35546
rect 21553 35482 21617 35546
rect 21634 35482 21698 35546
rect 21715 35482 21779 35546
rect 21796 35482 21860 35546
rect 21877 35482 21941 35546
rect 21958 35482 22022 35546
rect 22039 35482 22103 35546
rect 22120 35482 22184 35546
rect 22201 35482 22265 35546
rect 22282 35482 22346 35546
rect 22363 35482 22427 35546
rect 22444 35482 22508 35546
rect 22525 35482 22589 35546
rect 19258 35402 19322 35466
rect 19340 35402 19404 35466
rect 19422 35402 19486 35466
rect 19504 35402 19568 35466
rect 19586 35402 19650 35466
rect 19668 35402 19732 35466
rect 19750 35402 19814 35466
rect 19832 35402 19896 35466
rect 19914 35402 19978 35466
rect 19996 35402 20060 35466
rect 20078 35402 20142 35466
rect 20160 35402 20224 35466
rect 20242 35402 20306 35466
rect 20324 35402 20388 35466
rect 20406 35402 20470 35466
rect 20488 35402 20552 35466
rect 20570 35402 20634 35466
rect 20652 35402 20716 35466
rect 20734 35402 20798 35466
rect 20816 35402 20880 35466
rect 20898 35402 20962 35466
rect 20980 35402 21044 35466
rect 21062 35402 21126 35466
rect 21144 35402 21208 35466
rect 21226 35402 21290 35466
rect 21308 35402 21372 35466
rect 21390 35402 21454 35466
rect 21472 35402 21536 35466
rect 21553 35402 21617 35466
rect 21634 35402 21698 35466
rect 21715 35402 21779 35466
rect 21796 35402 21860 35466
rect 21877 35402 21941 35466
rect 21958 35402 22022 35466
rect 22039 35402 22103 35466
rect 22120 35402 22184 35466
rect 22201 35402 22265 35466
rect 22282 35402 22346 35466
rect 22363 35402 22427 35466
rect 22444 35402 22508 35466
rect 22525 35402 22589 35466
rect 19258 35322 19322 35386
rect 19340 35322 19404 35386
rect 19422 35322 19486 35386
rect 19504 35322 19568 35386
rect 19586 35322 19650 35386
rect 19668 35322 19732 35386
rect 19750 35322 19814 35386
rect 19832 35322 19896 35386
rect 19914 35322 19978 35386
rect 19996 35322 20060 35386
rect 20078 35322 20142 35386
rect 20160 35322 20224 35386
rect 20242 35322 20306 35386
rect 20324 35322 20388 35386
rect 20406 35322 20470 35386
rect 20488 35322 20552 35386
rect 20570 35322 20634 35386
rect 20652 35322 20716 35386
rect 20734 35322 20798 35386
rect 20816 35322 20880 35386
rect 20898 35322 20962 35386
rect 20980 35322 21044 35386
rect 21062 35322 21126 35386
rect 21144 35322 21208 35386
rect 21226 35322 21290 35386
rect 21308 35322 21372 35386
rect 21390 35322 21454 35386
rect 21472 35322 21536 35386
rect 21553 35322 21617 35386
rect 21634 35322 21698 35386
rect 21715 35322 21779 35386
rect 21796 35322 21860 35386
rect 21877 35322 21941 35386
rect 21958 35322 22022 35386
rect 22039 35322 22103 35386
rect 22120 35322 22184 35386
rect 22201 35322 22265 35386
rect 22282 35322 22346 35386
rect 22363 35322 22427 35386
rect 22444 35322 22508 35386
rect 22525 35322 22589 35386
rect 19258 35242 19322 35306
rect 19340 35242 19404 35306
rect 19422 35242 19486 35306
rect 19504 35242 19568 35306
rect 19586 35242 19650 35306
rect 19668 35242 19732 35306
rect 19750 35242 19814 35306
rect 19832 35242 19896 35306
rect 19914 35242 19978 35306
rect 19996 35242 20060 35306
rect 20078 35242 20142 35306
rect 20160 35242 20224 35306
rect 20242 35242 20306 35306
rect 20324 35242 20388 35306
rect 20406 35242 20470 35306
rect 20488 35242 20552 35306
rect 20570 35242 20634 35306
rect 20652 35242 20716 35306
rect 20734 35242 20798 35306
rect 20816 35242 20880 35306
rect 20898 35242 20962 35306
rect 20980 35242 21044 35306
rect 21062 35242 21126 35306
rect 21144 35242 21208 35306
rect 21226 35242 21290 35306
rect 21308 35242 21372 35306
rect 21390 35242 21454 35306
rect 21472 35242 21536 35306
rect 21553 35242 21617 35306
rect 21634 35242 21698 35306
rect 21715 35242 21779 35306
rect 21796 35242 21860 35306
rect 21877 35242 21941 35306
rect 21958 35242 22022 35306
rect 22039 35242 22103 35306
rect 22120 35242 22184 35306
rect 22201 35242 22265 35306
rect 22282 35242 22346 35306
rect 22363 35242 22427 35306
rect 22444 35242 22508 35306
rect 22525 35242 22589 35306
rect 19258 35162 19322 35226
rect 19340 35162 19404 35226
rect 19422 35162 19486 35226
rect 19504 35162 19568 35226
rect 19586 35162 19650 35226
rect 19668 35162 19732 35226
rect 19750 35162 19814 35226
rect 19832 35162 19896 35226
rect 19914 35162 19978 35226
rect 19996 35162 20060 35226
rect 20078 35162 20142 35226
rect 20160 35162 20224 35226
rect 20242 35162 20306 35226
rect 20324 35162 20388 35226
rect 20406 35162 20470 35226
rect 20488 35162 20552 35226
rect 20570 35162 20634 35226
rect 20652 35162 20716 35226
rect 20734 35162 20798 35226
rect 20816 35162 20880 35226
rect 20898 35162 20962 35226
rect 20980 35162 21044 35226
rect 21062 35162 21126 35226
rect 21144 35162 21208 35226
rect 21226 35162 21290 35226
rect 21308 35162 21372 35226
rect 21390 35162 21454 35226
rect 21472 35162 21536 35226
rect 21553 35162 21617 35226
rect 21634 35162 21698 35226
rect 21715 35162 21779 35226
rect 21796 35162 21860 35226
rect 21877 35162 21941 35226
rect 21958 35162 22022 35226
rect 22039 35162 22103 35226
rect 22120 35162 22184 35226
rect 22201 35162 22265 35226
rect 22282 35162 22346 35226
rect 22363 35162 22427 35226
rect 22444 35162 22508 35226
rect 22525 35162 22589 35226
rect 23396 35602 23460 35666
rect 23514 35602 23578 35666
rect 23632 35602 23696 35666
rect 23396 35519 23460 35583
rect 23514 35519 23578 35583
rect 23632 35519 23696 35583
rect 23396 35436 23460 35500
rect 23514 35436 23578 35500
rect 23632 35436 23696 35500
rect 23396 35353 23460 35417
rect 23514 35353 23578 35417
rect 23632 35353 23696 35417
rect 23396 35269 23460 35333
rect 23514 35269 23578 35333
rect 23632 35269 23696 35333
rect 23396 35185 23460 35249
rect 23514 35185 23578 35249
rect 23632 35185 23696 35249
rect 1016 24514 1080 24578
rect 1016 24406 1080 24470
rect 1016 24298 1080 24362
rect 852 7967 916 8031
rect 936 7967 1000 8031
rect 1020 7967 1084 8031
rect 852 7880 916 7944
rect 936 7880 1000 7944
rect 1020 7880 1084 7944
rect 852 7793 916 7857
rect 936 7793 1000 7857
rect 1020 7793 1084 7857
rect 852 7705 916 7769
rect 936 7705 1000 7769
rect 1020 7705 1084 7769
rect 852 7617 916 7681
rect 936 7617 1000 7681
rect 1020 7617 1084 7681
rect 852 7529 916 7593
rect 936 7529 1000 7593
rect 1020 7529 1084 7593
rect 852 7441 916 7505
rect 936 7441 1000 7505
rect 1020 7441 1084 7505
rect 852 7353 916 7417
rect 936 7353 1000 7417
rect 1020 7353 1084 7417
rect 1595 9176 1659 9240
rect 1675 9176 1739 9240
rect 1755 9176 1819 9240
rect 1835 9176 1899 9240
rect 1915 9176 1979 9240
rect 1995 9176 2059 9240
rect 2075 9176 2139 9240
rect 1595 9091 1659 9155
rect 1675 9091 1739 9155
rect 1755 9091 1819 9155
rect 1835 9091 1899 9155
rect 1915 9091 1979 9155
rect 1995 9091 2059 9155
rect 2075 9091 2139 9155
rect 1595 9006 1659 9070
rect 1675 9006 1739 9070
rect 1755 9006 1819 9070
rect 1835 9006 1899 9070
rect 1915 9006 1979 9070
rect 1995 9006 2059 9070
rect 2075 9006 2139 9070
rect 1595 8921 1659 8985
rect 1675 8921 1739 8985
rect 1755 8921 1819 8985
rect 1835 8921 1899 8985
rect 1915 8921 1979 8985
rect 1995 8921 2059 8985
rect 2075 8921 2139 8985
rect 1595 8836 1659 8900
rect 1675 8836 1739 8900
rect 1755 8836 1819 8900
rect 1835 8836 1899 8900
rect 1915 8836 1979 8900
rect 1995 8836 2059 8900
rect 2075 8836 2139 8900
rect 1595 8751 1659 8815
rect 1675 8751 1739 8815
rect 1755 8751 1819 8815
rect 1835 8751 1899 8815
rect 1915 8751 1979 8815
rect 1995 8751 2059 8815
rect 2075 8751 2139 8815
rect 1595 8666 1659 8730
rect 1675 8666 1739 8730
rect 1755 8666 1819 8730
rect 1835 8666 1899 8730
rect 1915 8666 1979 8730
rect 1995 8666 2059 8730
rect 2075 8666 2139 8730
rect 1595 8581 1659 8645
rect 1675 8581 1739 8645
rect 1755 8581 1819 8645
rect 1835 8581 1899 8645
rect 1915 8581 1979 8645
rect 1995 8581 2059 8645
rect 2075 8581 2139 8645
rect 1595 8496 1659 8560
rect 1675 8496 1739 8560
rect 1755 8496 1819 8560
rect 1835 8496 1899 8560
rect 1915 8496 1979 8560
rect 1995 8496 2059 8560
rect 2075 8496 2139 8560
rect 1595 8410 1659 8474
rect 1675 8410 1739 8474
rect 1755 8410 1819 8474
rect 1835 8410 1899 8474
rect 1915 8410 1979 8474
rect 1995 8410 2059 8474
rect 2075 8410 2139 8474
rect 1595 8324 1659 8388
rect 1675 8324 1739 8388
rect 1755 8324 1819 8388
rect 1835 8324 1899 8388
rect 1915 8324 1979 8388
rect 1995 8324 2059 8388
rect 2075 8324 2139 8388
rect 1539 4994 1603 5058
rect 1619 4994 1683 5058
rect 3718 33106 3782 33111
rect 3826 33106 3890 33111
rect 3718 33050 3732 33106
rect 3732 33050 3782 33106
rect 3826 33050 3846 33106
rect 3846 33050 3890 33106
rect 3718 33047 3782 33050
rect 3826 33047 3890 33050
rect 3934 33047 3998 33111
rect 3718 33010 3782 33014
rect 3826 33010 3890 33014
rect 3718 32954 3732 33010
rect 3732 32954 3782 33010
rect 3826 32954 3846 33010
rect 3846 32954 3890 33010
rect 3718 32950 3782 32954
rect 3826 32950 3890 32954
rect 3934 32950 3998 33014
rect 3718 32914 3782 32917
rect 3826 32914 3890 32917
rect 3718 32858 3732 32914
rect 3732 32858 3782 32914
rect 3826 32858 3846 32914
rect 3846 32858 3890 32914
rect 3718 32853 3782 32858
rect 3826 32853 3890 32858
rect 3934 32853 3998 32917
rect 3718 32818 3782 32820
rect 3826 32818 3890 32820
rect 3718 32762 3732 32818
rect 3732 32762 3782 32818
rect 3826 32762 3846 32818
rect 3846 32762 3890 32818
rect 3718 32756 3782 32762
rect 3826 32756 3890 32762
rect 3934 32756 3998 32820
rect 3718 32721 3782 32722
rect 3826 32721 3890 32722
rect 3718 32665 3732 32721
rect 3732 32665 3782 32721
rect 3826 32665 3846 32721
rect 3846 32665 3890 32721
rect 3718 32658 3782 32665
rect 3826 32658 3890 32665
rect 3934 32658 3998 32722
rect 3313 7957 3377 8021
rect 3419 7957 3483 8021
rect 3525 7957 3589 8021
rect 3631 7957 3695 8021
rect 3313 7873 3377 7937
rect 3419 7873 3483 7937
rect 3525 7873 3589 7937
rect 3631 7873 3695 7937
rect 3313 7788 3377 7852
rect 3419 7788 3483 7852
rect 3525 7788 3589 7852
rect 3631 7788 3695 7852
rect 3313 7703 3377 7767
rect 3419 7703 3483 7767
rect 3525 7703 3589 7767
rect 3631 7703 3695 7767
rect 3313 7618 3377 7682
rect 3419 7618 3483 7682
rect 3525 7618 3589 7682
rect 3631 7618 3695 7682
rect 3313 7533 3377 7597
rect 3419 7533 3483 7597
rect 3525 7533 3589 7597
rect 3631 7533 3695 7597
rect 3313 7448 3377 7512
rect 3419 7448 3483 7512
rect 3525 7448 3589 7512
rect 3631 7448 3695 7512
rect 3313 7363 3377 7427
rect 3419 7363 3483 7427
rect 3525 7363 3589 7427
rect 3631 7363 3695 7427
rect 6854 13633 6918 13697
rect 6939 13633 7003 13697
rect 7024 13633 7088 13697
rect 7109 13633 7173 13697
rect 7194 13633 7258 13697
rect 7279 13633 7343 13697
rect 7364 13633 7428 13697
rect 7449 13633 7513 13697
rect 7534 13633 7598 13697
rect 7619 13633 7683 13697
rect 7704 13633 7768 13697
rect 6854 13545 6918 13609
rect 6939 13545 7003 13609
rect 7024 13545 7088 13609
rect 7109 13545 7173 13609
rect 7194 13545 7258 13609
rect 7279 13545 7343 13609
rect 7364 13545 7428 13609
rect 7449 13545 7513 13609
rect 7534 13545 7598 13609
rect 7619 13545 7683 13609
rect 7704 13545 7768 13609
rect 6854 13457 6918 13521
rect 6939 13457 7003 13521
rect 7024 13457 7088 13521
rect 7109 13457 7173 13521
rect 7194 13457 7258 13521
rect 7279 13457 7343 13521
rect 7364 13457 7428 13521
rect 7449 13457 7513 13521
rect 7534 13457 7598 13521
rect 7619 13457 7683 13521
rect 7704 13457 7768 13521
rect 16060 13620 16124 13684
rect 16142 13620 16206 13684
rect 16223 13620 16287 13684
rect 16304 13620 16368 13684
rect 16385 13620 16449 13684
rect 16466 13620 16530 13684
rect 16547 13620 16611 13684
rect 16628 13620 16692 13684
rect 16709 13620 16773 13684
rect 16790 13620 16854 13684
rect 16871 13620 16935 13684
rect 16060 13532 16124 13596
rect 16142 13532 16206 13596
rect 16223 13532 16287 13596
rect 16304 13532 16368 13596
rect 16385 13532 16449 13596
rect 16466 13532 16530 13596
rect 16547 13532 16611 13596
rect 16628 13532 16692 13596
rect 16709 13532 16773 13596
rect 16790 13532 16854 13596
rect 16871 13532 16935 13596
rect 16060 13444 16124 13508
rect 16142 13444 16206 13508
rect 16223 13444 16287 13508
rect 16304 13444 16368 13508
rect 16385 13444 16449 13508
rect 16466 13444 16530 13508
rect 16547 13444 16611 13508
rect 16628 13444 16692 13508
rect 16709 13444 16773 13508
rect 16790 13444 16854 13508
rect 16871 13444 16935 13508
rect 16060 13356 16124 13420
rect 16142 13356 16206 13420
rect 16223 13356 16287 13420
rect 16304 13356 16368 13420
rect 16385 13356 16449 13420
rect 16466 13356 16530 13420
rect 16547 13356 16611 13420
rect 16628 13356 16692 13420
rect 16709 13356 16773 13420
rect 16790 13356 16854 13420
rect 16871 13356 16935 13420
rect 16060 13268 16124 13332
rect 16142 13268 16206 13332
rect 16223 13268 16287 13332
rect 16304 13268 16368 13332
rect 16385 13268 16449 13332
rect 16466 13268 16530 13332
rect 16547 13268 16611 13332
rect 16628 13268 16692 13332
rect 16709 13268 16773 13332
rect 16790 13268 16854 13332
rect 16871 13268 16935 13332
rect 16060 13180 16124 13244
rect 16142 13180 16206 13244
rect 16223 13180 16287 13244
rect 16304 13180 16368 13244
rect 16385 13180 16449 13244
rect 16466 13180 16530 13244
rect 16547 13180 16611 13244
rect 16628 13180 16692 13244
rect 16709 13180 16773 13244
rect 16790 13180 16854 13244
rect 16871 13180 16935 13244
rect 16060 13092 16124 13156
rect 16142 13092 16206 13156
rect 16223 13092 16287 13156
rect 16304 13092 16368 13156
rect 16385 13092 16449 13156
rect 16466 13092 16530 13156
rect 16547 13092 16611 13156
rect 16628 13092 16692 13156
rect 16709 13092 16773 13156
rect 16790 13092 16854 13156
rect 16871 13092 16935 13156
rect 16060 13004 16124 13068
rect 16142 13004 16206 13068
rect 16223 13004 16287 13068
rect 16304 13004 16368 13068
rect 16385 13004 16449 13068
rect 16466 13004 16530 13068
rect 16547 13004 16611 13068
rect 16628 13004 16692 13068
rect 16709 13004 16773 13068
rect 16790 13004 16854 13068
rect 16871 13004 16935 13068
rect 16060 12916 16124 12980
rect 16142 12916 16206 12980
rect 16223 12916 16287 12980
rect 16304 12916 16368 12980
rect 16385 12916 16449 12980
rect 16466 12916 16530 12980
rect 16547 12916 16611 12980
rect 16628 12916 16692 12980
rect 16709 12916 16773 12980
rect 16790 12916 16854 12980
rect 16871 12916 16935 12980
rect 16060 12828 16124 12892
rect 16142 12828 16206 12892
rect 16223 12828 16287 12892
rect 16304 12828 16368 12892
rect 16385 12828 16449 12892
rect 16466 12828 16530 12892
rect 16547 12828 16611 12892
rect 16628 12828 16692 12892
rect 16709 12828 16773 12892
rect 16790 12828 16854 12892
rect 16871 12828 16935 12892
rect 7446 9023 7510 9087
rect 7532 9023 7596 9087
rect 7618 9023 7682 9087
rect 7704 9023 7768 9087
rect 7790 9023 7854 9087
rect 7876 9023 7940 9087
rect 7962 9023 8026 9087
rect 7446 8937 7510 9001
rect 7532 8937 7596 9001
rect 7618 8937 7682 9001
rect 7704 8937 7768 9001
rect 7790 8937 7854 9001
rect 7876 8937 7940 9001
rect 7962 8937 8026 9001
rect 7446 8851 7510 8915
rect 7532 8851 7596 8915
rect 7618 8851 7682 8915
rect 7704 8851 7768 8915
rect 7790 8851 7854 8915
rect 7876 8851 7940 8915
rect 7962 8851 8026 8915
rect 7446 8765 7510 8829
rect 7532 8765 7596 8829
rect 7618 8765 7682 8829
rect 7704 8765 7768 8829
rect 7790 8765 7854 8829
rect 7876 8765 7940 8829
rect 7962 8765 8026 8829
rect 7446 8679 7510 8743
rect 7532 8679 7596 8743
rect 7618 8679 7682 8743
rect 7704 8679 7768 8743
rect 7790 8679 7854 8743
rect 7876 8679 7940 8743
rect 7962 8679 8026 8743
rect 7446 8593 7510 8657
rect 7532 8593 7596 8657
rect 7618 8593 7682 8657
rect 7704 8593 7768 8657
rect 7790 8593 7854 8657
rect 7876 8593 7940 8657
rect 7962 8593 8026 8657
rect 7446 8507 7510 8571
rect 7532 8507 7596 8571
rect 7618 8507 7682 8571
rect 7704 8507 7768 8571
rect 7790 8507 7854 8571
rect 7876 8507 7940 8571
rect 7962 8507 8026 8571
rect 7446 8420 7510 8484
rect 7532 8420 7596 8484
rect 7618 8420 7682 8484
rect 7704 8420 7768 8484
rect 7790 8420 7854 8484
rect 7876 8420 7940 8484
rect 7962 8420 8026 8484
rect 7446 8333 7510 8397
rect 7532 8333 7596 8397
rect 7618 8333 7682 8397
rect 7704 8333 7768 8397
rect 7790 8333 7854 8397
rect 7876 8333 7940 8397
rect 7962 8333 8026 8397
rect 2175 4994 2239 5058
rect 2255 4994 2319 5058
rect 1955 3575 2019 3639
rect 1955 3492 2019 3556
rect 1955 3409 2019 3473
rect 1955 3326 2019 3390
rect 1955 3243 2019 3307
rect 1955 3160 2019 3224
rect 1955 3077 2019 3141
rect 1955 2993 2019 3057
rect 1592 2814 1656 2878
rect 1672 2814 1736 2878
rect 2175 2814 2239 2878
rect 2255 2814 2319 2878
rect 3340 1427 3404 1491
rect 3428 1427 3492 1491
rect 3516 1427 3580 1491
rect 3604 1427 3668 1491
rect 3692 1427 3756 1491
rect 3780 1427 3844 1491
rect 3340 1343 3404 1407
rect 3428 1343 3492 1407
rect 3516 1343 3580 1407
rect 3604 1343 3668 1407
rect 3692 1343 3756 1407
rect 3780 1343 3844 1407
rect 3340 1259 3404 1323
rect 3428 1259 3492 1323
rect 3516 1259 3580 1323
rect 3604 1259 3668 1323
rect 3692 1259 3756 1323
rect 3780 1259 3844 1323
rect 3340 1175 3404 1239
rect 3428 1175 3492 1239
rect 3516 1175 3580 1239
rect 3604 1175 3668 1239
rect 3692 1175 3756 1239
rect 3780 1175 3844 1239
rect 3340 1091 3404 1155
rect 3428 1091 3492 1155
rect 3516 1091 3580 1155
rect 3604 1091 3668 1155
rect 3692 1091 3756 1155
rect 3780 1091 3844 1155
rect 3340 1007 3404 1071
rect 3428 1007 3492 1071
rect 3516 1007 3580 1071
rect 3604 1007 3668 1071
rect 3692 1007 3756 1071
rect 3780 1007 3844 1071
rect 3340 923 3404 987
rect 3428 923 3492 987
rect 3516 923 3580 987
rect 3604 923 3668 987
rect 3692 923 3756 987
rect 3780 923 3844 987
rect 3340 838 3404 902
rect 3428 838 3492 902
rect 3516 838 3580 902
rect 3604 838 3668 902
rect 3692 838 3756 902
rect 3780 838 3844 902
rect 3340 753 3404 817
rect 3428 753 3492 817
rect 3516 753 3580 817
rect 3604 753 3668 817
rect 3692 753 3756 817
rect 3780 753 3844 817
rect 3340 668 3404 732
rect 3428 668 3492 732
rect 3516 668 3580 732
rect 3604 668 3668 732
rect 3692 668 3756 732
rect 3780 668 3844 732
rect 3340 583 3404 647
rect 3428 583 3492 647
rect 3516 583 3580 647
rect 3604 583 3668 647
rect 3692 583 3756 647
rect 3780 583 3844 647
rect 3340 498 3404 562
rect 3428 498 3492 562
rect 3516 498 3580 562
rect 3604 498 3668 562
rect 3692 498 3756 562
rect 3780 498 3844 562
rect 3340 413 3404 477
rect 3428 413 3492 477
rect 3516 413 3580 477
rect 3604 413 3668 477
rect 3692 413 3756 477
rect 3780 413 3844 477
rect 5095 2811 5159 2875
rect 5175 2811 5239 2875
rect 5386 2811 5450 2875
rect 5466 2811 5530 2875
rect 5944 2637 6008 2701
rect 6032 2637 6096 2701
rect 6120 2637 6184 2701
rect 6208 2637 6272 2701
rect 6296 2637 6360 2701
rect 6384 2637 6448 2701
rect 6472 2637 6536 2701
rect 5944 2552 6008 2616
rect 6032 2552 6096 2616
rect 6120 2552 6184 2616
rect 6208 2552 6272 2616
rect 6296 2552 6360 2616
rect 6384 2552 6448 2616
rect 6472 2552 6536 2616
rect 5944 2467 6008 2531
rect 6032 2467 6096 2531
rect 6120 2467 6184 2531
rect 6208 2467 6272 2531
rect 6296 2467 6360 2531
rect 6384 2467 6448 2531
rect 6472 2467 6536 2531
rect 5944 2382 6008 2446
rect 6032 2382 6096 2446
rect 6120 2382 6184 2446
rect 6208 2382 6272 2446
rect 6296 2382 6360 2446
rect 6384 2382 6448 2446
rect 6472 2382 6536 2446
rect 5944 2297 6008 2361
rect 6032 2297 6096 2361
rect 6120 2297 6184 2361
rect 6208 2297 6272 2361
rect 6296 2297 6360 2361
rect 6384 2297 6448 2361
rect 6472 2297 6536 2361
rect 5944 2212 6008 2276
rect 6032 2212 6096 2276
rect 6120 2212 6184 2276
rect 6208 2212 6272 2276
rect 6296 2212 6360 2276
rect 6384 2212 6448 2276
rect 6472 2212 6536 2276
rect 5944 2127 6008 2191
rect 6032 2127 6096 2191
rect 6120 2127 6184 2191
rect 6208 2127 6272 2191
rect 6296 2127 6360 2191
rect 6384 2127 6448 2191
rect 6472 2127 6536 2191
rect 5944 2041 6008 2105
rect 6032 2041 6096 2105
rect 6120 2041 6184 2105
rect 6208 2041 6272 2105
rect 6296 2041 6360 2105
rect 6384 2041 6448 2105
rect 6472 2041 6536 2105
rect 5944 1955 6008 2019
rect 6032 1955 6096 2019
rect 6120 1955 6184 2019
rect 6208 1955 6272 2019
rect 6296 1955 6360 2019
rect 6384 1955 6448 2019
rect 6472 1955 6536 2019
rect 5944 1869 6008 1933
rect 6032 1869 6096 1933
rect 6120 1869 6184 1933
rect 6208 1869 6272 1933
rect 6296 1869 6360 1933
rect 6384 1869 6448 1933
rect 6472 1869 6536 1933
rect 5944 1783 6008 1847
rect 6032 1783 6096 1847
rect 6120 1783 6184 1847
rect 6208 1783 6272 1847
rect 6296 1783 6360 1847
rect 6384 1783 6448 1847
rect 6472 1783 6536 1847
rect 8696 1612 8760 1676
rect 8776 1612 8840 1676
rect 8987 1612 9051 1676
rect 9067 1612 9131 1676
rect 9768 3600 9832 3664
rect 9848 3600 9912 3664
rect 9928 3600 9992 3664
rect 10008 3600 10072 3664
rect 9768 3515 9832 3579
rect 9848 3515 9912 3579
rect 9928 3515 9992 3579
rect 10008 3515 10072 3579
rect 9768 3430 9832 3494
rect 9848 3430 9912 3494
rect 9928 3430 9992 3494
rect 10008 3430 10072 3494
rect 9768 3345 9832 3409
rect 9848 3345 9912 3409
rect 9928 3345 9992 3409
rect 10008 3345 10072 3409
rect 9768 3259 9832 3323
rect 9848 3259 9912 3323
rect 9928 3259 9992 3323
rect 10008 3259 10072 3323
rect 9768 3173 9832 3237
rect 9848 3173 9912 3237
rect 9928 3173 9992 3237
rect 10008 3173 10072 3237
rect 9768 3087 9832 3151
rect 9848 3087 9912 3151
rect 9928 3087 9992 3151
rect 10008 3087 10072 3151
rect 9768 3001 9832 3065
rect 9848 3001 9912 3065
rect 9928 3001 9992 3065
rect 10008 3001 10072 3065
rect 11516 9164 11580 9228
rect 11602 9164 11666 9228
rect 11688 9164 11752 9228
rect 11774 9164 11838 9228
rect 11860 9164 11924 9228
rect 11946 9164 12010 9228
rect 12032 9164 12096 9228
rect 11516 9081 11580 9145
rect 11602 9081 11666 9145
rect 11688 9081 11752 9145
rect 11774 9081 11838 9145
rect 11860 9081 11924 9145
rect 11946 9081 12010 9145
rect 12032 9081 12096 9145
rect 11516 8998 11580 9062
rect 11602 8998 11666 9062
rect 11688 8998 11752 9062
rect 11774 8998 11838 9062
rect 11860 8998 11924 9062
rect 11946 8998 12010 9062
rect 12032 8998 12096 9062
rect 11516 8915 11580 8979
rect 11602 8915 11666 8979
rect 11688 8915 11752 8979
rect 11774 8915 11838 8979
rect 11860 8915 11924 8979
rect 11946 8915 12010 8979
rect 12032 8915 12096 8979
rect 11516 8832 11580 8896
rect 11602 8832 11666 8896
rect 11688 8832 11752 8896
rect 11774 8832 11838 8896
rect 11860 8832 11924 8896
rect 11946 8832 12010 8896
rect 12032 8832 12096 8896
rect 11516 8749 11580 8813
rect 11602 8749 11666 8813
rect 11688 8749 11752 8813
rect 11774 8749 11838 8813
rect 11860 8749 11924 8813
rect 11946 8749 12010 8813
rect 12032 8749 12096 8813
rect 11516 8666 11580 8730
rect 11602 8666 11666 8730
rect 11688 8666 11752 8730
rect 11774 8666 11838 8730
rect 11860 8666 11924 8730
rect 11946 8666 12010 8730
rect 12032 8666 12096 8730
rect 11516 8583 11580 8647
rect 11602 8583 11666 8647
rect 11688 8583 11752 8647
rect 11774 8583 11838 8647
rect 11860 8583 11924 8647
rect 11946 8583 12010 8647
rect 12032 8583 12096 8647
rect 11516 8500 11580 8564
rect 11602 8500 11666 8564
rect 11688 8500 11752 8564
rect 11774 8500 11838 8564
rect 11860 8500 11924 8564
rect 11946 8500 12010 8564
rect 12032 8500 12096 8564
rect 11516 8416 11580 8480
rect 11602 8416 11666 8480
rect 11688 8416 11752 8480
rect 11774 8416 11838 8480
rect 11860 8416 11924 8480
rect 11946 8416 12010 8480
rect 12032 8416 12096 8480
rect 11516 8332 11580 8396
rect 11602 8332 11666 8396
rect 11688 8332 11752 8396
rect 11774 8332 11838 8396
rect 11860 8332 11924 8396
rect 11946 8332 12010 8396
rect 12032 8332 12096 8396
rect 12229 2637 12293 2701
rect 12317 2637 12381 2701
rect 12405 2637 12469 2701
rect 12493 2637 12557 2701
rect 12581 2637 12645 2701
rect 12669 2637 12733 2701
rect 12757 2637 12821 2701
rect 12229 2552 12293 2616
rect 12317 2552 12381 2616
rect 12405 2552 12469 2616
rect 12493 2552 12557 2616
rect 12581 2552 12645 2616
rect 12669 2552 12733 2616
rect 12757 2552 12821 2616
rect 12229 2467 12293 2531
rect 12317 2467 12381 2531
rect 12405 2467 12469 2531
rect 12493 2467 12557 2531
rect 12581 2467 12645 2531
rect 12669 2467 12733 2531
rect 12757 2467 12821 2531
rect 12229 2382 12293 2446
rect 12317 2382 12381 2446
rect 12405 2382 12469 2446
rect 12493 2382 12557 2446
rect 12581 2382 12645 2446
rect 12669 2382 12733 2446
rect 12757 2382 12821 2446
rect 12229 2297 12293 2361
rect 12317 2297 12381 2361
rect 12405 2297 12469 2361
rect 12493 2297 12557 2361
rect 12581 2297 12645 2361
rect 12669 2297 12733 2361
rect 12757 2297 12821 2361
rect 12229 2212 12293 2276
rect 12317 2212 12381 2276
rect 12405 2212 12469 2276
rect 12493 2212 12557 2276
rect 12581 2212 12645 2276
rect 12669 2212 12733 2276
rect 12757 2212 12821 2276
rect 12229 2127 12293 2191
rect 12317 2127 12381 2191
rect 12405 2127 12469 2191
rect 12493 2127 12557 2191
rect 12581 2127 12645 2191
rect 12669 2127 12733 2191
rect 12757 2127 12821 2191
rect 12229 2041 12293 2105
rect 12317 2041 12381 2105
rect 12405 2041 12469 2105
rect 12493 2041 12557 2105
rect 12581 2041 12645 2105
rect 12669 2041 12733 2105
rect 12757 2041 12821 2105
rect 12229 1955 12293 2019
rect 12317 1955 12381 2019
rect 12405 1955 12469 2019
rect 12493 1955 12557 2019
rect 12581 1955 12645 2019
rect 12669 1955 12733 2019
rect 12757 1955 12821 2019
rect 12229 1869 12293 1933
rect 12317 1869 12381 1933
rect 12405 1869 12469 1933
rect 12493 1869 12557 1933
rect 12581 1869 12645 1933
rect 12669 1869 12733 1933
rect 12757 1869 12821 1933
rect 12229 1783 12293 1847
rect 12317 1783 12381 1847
rect 12405 1783 12469 1847
rect 12493 1783 12557 1847
rect 12581 1783 12645 1847
rect 12669 1783 12733 1847
rect 12757 1783 12821 1847
rect 10337 1612 10401 1676
rect 10417 1612 10481 1676
rect 10628 1612 10692 1676
rect 10708 1612 10772 1676
rect 14540 9171 14604 9235
rect 14626 9171 14690 9235
rect 14712 9171 14776 9235
rect 14798 9171 14862 9235
rect 14884 9171 14948 9235
rect 14970 9171 15034 9235
rect 15056 9171 15120 9235
rect 14540 9088 14604 9152
rect 14626 9088 14690 9152
rect 14712 9088 14776 9152
rect 14798 9088 14862 9152
rect 14884 9088 14948 9152
rect 14970 9088 15034 9152
rect 15056 9088 15120 9152
rect 14540 9004 14604 9068
rect 14626 9004 14690 9068
rect 14712 9004 14776 9068
rect 14798 9004 14862 9068
rect 14884 9004 14948 9068
rect 14970 9004 15034 9068
rect 15056 9004 15120 9068
rect 14540 8920 14604 8984
rect 14626 8920 14690 8984
rect 14712 8920 14776 8984
rect 14798 8920 14862 8984
rect 14884 8920 14948 8984
rect 14970 8920 15034 8984
rect 15056 8920 15120 8984
rect 14540 8836 14604 8900
rect 14626 8836 14690 8900
rect 14712 8836 14776 8900
rect 14798 8836 14862 8900
rect 14884 8836 14948 8900
rect 14970 8836 15034 8900
rect 15056 8836 15120 8900
rect 14540 8752 14604 8816
rect 14626 8752 14690 8816
rect 14712 8752 14776 8816
rect 14798 8752 14862 8816
rect 14884 8752 14948 8816
rect 14970 8752 15034 8816
rect 15056 8752 15120 8816
rect 14540 8668 14604 8732
rect 14626 8668 14690 8732
rect 14712 8668 14776 8732
rect 14798 8668 14862 8732
rect 14884 8668 14948 8732
rect 14970 8668 15034 8732
rect 15056 8668 15120 8732
rect 14540 8584 14604 8648
rect 14626 8584 14690 8648
rect 14712 8584 14776 8648
rect 14798 8584 14862 8648
rect 14884 8584 14948 8648
rect 14970 8584 15034 8648
rect 15056 8584 15120 8648
rect 14540 8500 14604 8564
rect 14626 8500 14690 8564
rect 14712 8500 14776 8564
rect 14798 8500 14862 8564
rect 14884 8500 14948 8564
rect 14970 8500 15034 8564
rect 15056 8500 15120 8564
rect 14540 8416 14604 8480
rect 14626 8416 14690 8480
rect 14712 8416 14776 8480
rect 14798 8416 14862 8480
rect 14884 8416 14948 8480
rect 14970 8416 15034 8480
rect 15056 8416 15120 8480
rect 14540 8332 14604 8396
rect 14626 8332 14690 8396
rect 14712 8332 14776 8396
rect 14798 8332 14862 8396
rect 14884 8332 14948 8396
rect 14970 8332 15034 8396
rect 15056 8332 15120 8396
rect 17880 9175 17944 9239
rect 17960 9175 18024 9239
rect 18040 9175 18104 9239
rect 18120 9175 18184 9239
rect 17880 9090 17944 9154
rect 17960 9090 18024 9154
rect 18040 9090 18104 9154
rect 18120 9090 18184 9154
rect 17880 9005 17944 9069
rect 17960 9005 18024 9069
rect 18040 9005 18104 9069
rect 18120 9005 18184 9069
rect 17880 8920 17944 8984
rect 17960 8920 18024 8984
rect 18040 8920 18104 8984
rect 18120 8920 18184 8984
rect 17880 8835 17944 8899
rect 17960 8835 18024 8899
rect 18040 8835 18104 8899
rect 18120 8835 18184 8899
rect 17880 8750 17944 8814
rect 17960 8750 18024 8814
rect 18040 8750 18104 8814
rect 18120 8750 18184 8814
rect 17880 8665 17944 8729
rect 17960 8665 18024 8729
rect 18040 8665 18104 8729
rect 18120 8665 18184 8729
rect 17880 8580 17944 8644
rect 17960 8580 18024 8644
rect 18040 8580 18104 8644
rect 18120 8580 18184 8644
rect 17880 8495 17944 8559
rect 17960 8495 18024 8559
rect 18040 8495 18104 8559
rect 18120 8495 18184 8559
rect 17880 8410 17944 8474
rect 17960 8410 18024 8474
rect 18040 8410 18104 8474
rect 18120 8410 18184 8474
rect 17880 8324 17944 8388
rect 17960 8324 18024 8388
rect 18040 8324 18104 8388
rect 18120 8324 18184 8388
rect 20130 9175 20194 9239
rect 20210 9175 20274 9239
rect 20290 9175 20354 9239
rect 20370 9175 20434 9239
rect 20450 9175 20514 9239
rect 20130 9090 20194 9154
rect 20210 9090 20274 9154
rect 20290 9090 20354 9154
rect 20370 9090 20434 9154
rect 20450 9090 20514 9154
rect 20130 9005 20194 9069
rect 20210 9005 20274 9069
rect 20290 9005 20354 9069
rect 20370 9005 20434 9069
rect 20450 9005 20514 9069
rect 20130 8920 20194 8984
rect 20210 8920 20274 8984
rect 20290 8920 20354 8984
rect 20370 8920 20434 8984
rect 20450 8920 20514 8984
rect 20130 8835 20194 8899
rect 20210 8835 20274 8899
rect 20290 8835 20354 8899
rect 20370 8835 20434 8899
rect 20450 8835 20514 8899
rect 20130 8750 20194 8814
rect 20210 8750 20274 8814
rect 20290 8750 20354 8814
rect 20370 8750 20434 8814
rect 20450 8750 20514 8814
rect 20130 8665 20194 8729
rect 20210 8665 20274 8729
rect 20290 8665 20354 8729
rect 20370 8665 20434 8729
rect 20450 8665 20514 8729
rect 20130 8580 20194 8644
rect 20210 8580 20274 8644
rect 20290 8580 20354 8644
rect 20370 8580 20434 8644
rect 20450 8580 20514 8644
rect 20130 8495 20194 8559
rect 20210 8495 20274 8559
rect 20290 8495 20354 8559
rect 20370 8495 20434 8559
rect 20450 8495 20514 8559
rect 20130 8410 20194 8474
rect 20210 8410 20274 8474
rect 20290 8410 20354 8474
rect 20370 8410 20434 8474
rect 20450 8410 20514 8474
rect 20130 8324 20194 8388
rect 20210 8324 20274 8388
rect 20290 8324 20354 8388
rect 20370 8324 20434 8388
rect 20450 8324 20514 8388
rect 21871 6991 21935 7055
rect 21963 6991 22027 7055
rect 22055 6991 22119 7055
rect 22147 6991 22211 7055
rect 22239 6991 22303 7055
rect 21871 6905 21935 6969
rect 21963 6905 22027 6969
rect 22055 6905 22119 6969
rect 22147 6905 22211 6969
rect 22239 6905 22303 6969
rect 21871 6819 21935 6883
rect 21963 6819 22027 6883
rect 22055 6819 22119 6883
rect 22147 6819 22211 6883
rect 22239 6819 22303 6883
rect 21871 6733 21935 6797
rect 21963 6733 22027 6797
rect 22055 6733 22119 6797
rect 22147 6733 22211 6797
rect 22239 6733 22303 6797
rect 21871 6647 21935 6711
rect 21963 6647 22027 6711
rect 22055 6647 22119 6711
rect 22147 6647 22211 6711
rect 22239 6647 22303 6711
rect 21871 6561 21935 6625
rect 21963 6561 22027 6625
rect 22055 6561 22119 6625
rect 22147 6561 22211 6625
rect 22239 6561 22303 6625
rect 21871 6474 21935 6538
rect 21963 6474 22027 6538
rect 22055 6474 22119 6538
rect 22147 6474 22211 6538
rect 22239 6474 22303 6538
rect 21871 6387 21935 6451
rect 21963 6387 22027 6451
rect 22055 6387 22119 6451
rect 22147 6387 22211 6451
rect 22239 6387 22303 6451
rect 12672 233 12736 297
rect 12752 233 12816 297
rect 12963 233 13027 297
rect 13043 233 13107 297
rect 16061 2637 16125 2701
rect 16149 2637 16213 2701
rect 16237 2637 16301 2701
rect 16325 2637 16389 2701
rect 16413 2637 16477 2701
rect 16501 2637 16565 2701
rect 16589 2637 16653 2701
rect 16061 2552 16125 2616
rect 16149 2552 16213 2616
rect 16237 2552 16301 2616
rect 16325 2552 16389 2616
rect 16413 2552 16477 2616
rect 16501 2552 16565 2616
rect 16589 2552 16653 2616
rect 16061 2467 16125 2531
rect 16149 2467 16213 2531
rect 16237 2467 16301 2531
rect 16325 2467 16389 2531
rect 16413 2467 16477 2531
rect 16501 2467 16565 2531
rect 16589 2467 16653 2531
rect 16061 2382 16125 2446
rect 16149 2382 16213 2446
rect 16237 2382 16301 2446
rect 16325 2382 16389 2446
rect 16413 2382 16477 2446
rect 16501 2382 16565 2446
rect 16589 2382 16653 2446
rect 16061 2297 16125 2361
rect 16149 2297 16213 2361
rect 16237 2297 16301 2361
rect 16325 2297 16389 2361
rect 16413 2297 16477 2361
rect 16501 2297 16565 2361
rect 16589 2297 16653 2361
rect 16061 2212 16125 2276
rect 16149 2212 16213 2276
rect 16237 2212 16301 2276
rect 16325 2212 16389 2276
rect 16413 2212 16477 2276
rect 16501 2212 16565 2276
rect 16589 2212 16653 2276
rect 16061 2127 16125 2191
rect 16149 2127 16213 2191
rect 16237 2127 16301 2191
rect 16325 2127 16389 2191
rect 16413 2127 16477 2191
rect 16501 2127 16565 2191
rect 16589 2127 16653 2191
rect 16061 2041 16125 2105
rect 16149 2041 16213 2105
rect 16237 2041 16301 2105
rect 16325 2041 16389 2105
rect 16413 2041 16477 2105
rect 16501 2041 16565 2105
rect 16589 2041 16653 2105
rect 16061 1955 16125 2019
rect 16149 1955 16213 2019
rect 16237 1955 16301 2019
rect 16325 1955 16389 2019
rect 16413 1955 16477 2019
rect 16501 1955 16565 2019
rect 16589 1955 16653 2019
rect 16061 1869 16125 1933
rect 16149 1869 16213 1933
rect 16237 1869 16301 1933
rect 16325 1869 16389 1933
rect 16413 1869 16477 1933
rect 16501 1869 16565 1933
rect 16589 1869 16653 1933
rect 16061 1783 16125 1847
rect 16149 1783 16213 1847
rect 16237 1783 16301 1847
rect 16325 1783 16389 1847
rect 16413 1783 16477 1847
rect 16501 1783 16565 1847
rect 16589 1783 16653 1847
rect 17775 1427 17839 1491
rect 17859 1427 17923 1491
rect 17943 1427 18007 1491
rect 18027 1427 18091 1491
rect 18111 1427 18175 1491
rect 17775 1343 17839 1407
rect 17859 1343 17923 1407
rect 17943 1343 18007 1407
rect 18027 1343 18091 1407
rect 18111 1343 18175 1407
rect 17775 1259 17839 1323
rect 17859 1259 17923 1323
rect 17943 1259 18007 1323
rect 18027 1259 18091 1323
rect 18111 1259 18175 1323
rect 17775 1175 17839 1239
rect 17859 1175 17923 1239
rect 17943 1175 18007 1239
rect 18027 1175 18091 1239
rect 18111 1175 18175 1239
rect 17775 1091 17839 1155
rect 17859 1091 17923 1155
rect 17943 1091 18007 1155
rect 18027 1091 18091 1155
rect 18111 1091 18175 1155
rect 17775 1007 17839 1071
rect 17859 1007 17923 1071
rect 17943 1007 18007 1071
rect 18027 1007 18091 1071
rect 18111 1007 18175 1071
rect 17775 923 17839 987
rect 17859 923 17923 987
rect 17943 923 18007 987
rect 18027 923 18091 987
rect 18111 923 18175 987
rect 17775 838 17839 902
rect 17859 838 17923 902
rect 17943 838 18007 902
rect 18027 838 18091 902
rect 18111 838 18175 902
rect 17775 753 17839 817
rect 17859 753 17923 817
rect 17943 753 18007 817
rect 18027 753 18091 817
rect 18111 753 18175 817
rect 17775 668 17839 732
rect 17859 668 17923 732
rect 17943 668 18007 732
rect 18027 668 18091 732
rect 18111 668 18175 732
rect 17775 583 17839 647
rect 17859 583 17923 647
rect 17943 583 18007 647
rect 18027 583 18091 647
rect 18111 583 18175 647
rect 17775 498 17839 562
rect 17859 498 17923 562
rect 17943 498 18007 562
rect 18027 498 18091 562
rect 18111 498 18175 562
rect 17775 413 17839 477
rect 17859 413 17923 477
rect 17943 413 18007 477
rect 18027 413 18091 477
rect 18111 413 18175 477
rect 20296 2637 20360 2701
rect 20384 2637 20448 2701
rect 20472 2637 20536 2701
rect 20560 2637 20624 2701
rect 20648 2637 20712 2701
rect 20736 2637 20800 2701
rect 20824 2637 20888 2701
rect 20296 2552 20360 2616
rect 20384 2552 20448 2616
rect 20472 2552 20536 2616
rect 20560 2552 20624 2616
rect 20648 2552 20712 2616
rect 20736 2552 20800 2616
rect 20824 2552 20888 2616
rect 20296 2467 20360 2531
rect 20384 2467 20448 2531
rect 20472 2467 20536 2531
rect 20560 2467 20624 2531
rect 20648 2467 20712 2531
rect 20736 2467 20800 2531
rect 20824 2467 20888 2531
rect 20296 2382 20360 2446
rect 20384 2382 20448 2446
rect 20472 2382 20536 2446
rect 20560 2382 20624 2446
rect 20648 2382 20712 2446
rect 20736 2382 20800 2446
rect 20824 2382 20888 2446
rect 20296 2297 20360 2361
rect 20384 2297 20448 2361
rect 20472 2297 20536 2361
rect 20560 2297 20624 2361
rect 20648 2297 20712 2361
rect 20736 2297 20800 2361
rect 20824 2297 20888 2361
rect 20296 2212 20360 2276
rect 20384 2212 20448 2276
rect 20472 2212 20536 2276
rect 20560 2212 20624 2276
rect 20648 2212 20712 2276
rect 20736 2212 20800 2276
rect 20824 2212 20888 2276
rect 20296 2127 20360 2191
rect 20384 2127 20448 2191
rect 20472 2127 20536 2191
rect 20560 2127 20624 2191
rect 20648 2127 20712 2191
rect 20736 2127 20800 2191
rect 20824 2127 20888 2191
rect 20296 2041 20360 2105
rect 20384 2041 20448 2105
rect 20472 2041 20536 2105
rect 20560 2041 20624 2105
rect 20648 2041 20712 2105
rect 20736 2041 20800 2105
rect 20824 2041 20888 2105
rect 20296 1955 20360 2019
rect 20384 1955 20448 2019
rect 20472 1955 20536 2019
rect 20560 1955 20624 2019
rect 20648 1955 20712 2019
rect 20736 1955 20800 2019
rect 20824 1955 20888 2019
rect 20296 1869 20360 1933
rect 20384 1869 20448 1933
rect 20472 1869 20536 1933
rect 20560 1869 20624 1933
rect 20648 1869 20712 1933
rect 20736 1869 20800 1933
rect 20824 1869 20888 1933
rect 20296 1783 20360 1847
rect 20384 1783 20448 1847
rect 20472 1783 20536 1847
rect 20560 1783 20624 1847
rect 20648 1783 20712 1847
rect 20736 1783 20800 1847
rect 20824 1783 20888 1847
rect 21134 1612 21198 1676
rect 21214 1612 21278 1676
rect 21425 1612 21489 1676
rect 21505 1612 21569 1676
rect 22281 1424 22345 1488
rect 22365 1424 22429 1488
rect 22449 1424 22513 1488
rect 22533 1424 22597 1488
rect 22617 1424 22681 1488
rect 22701 1424 22765 1488
rect 22785 1424 22849 1488
rect 22869 1424 22933 1488
rect 22281 1341 22345 1405
rect 22365 1341 22429 1405
rect 22449 1341 22513 1405
rect 22533 1341 22597 1405
rect 22617 1341 22681 1405
rect 22701 1341 22765 1405
rect 22785 1341 22849 1405
rect 22869 1341 22933 1405
rect 22281 1258 22345 1322
rect 22365 1258 22429 1322
rect 22449 1258 22513 1322
rect 22533 1258 22597 1322
rect 22617 1258 22681 1322
rect 22701 1258 22765 1322
rect 22785 1258 22849 1322
rect 22869 1258 22933 1322
rect 22281 1174 22345 1238
rect 22365 1174 22429 1238
rect 22449 1174 22513 1238
rect 22533 1174 22597 1238
rect 22617 1174 22681 1238
rect 22701 1174 22765 1238
rect 22785 1174 22849 1238
rect 22869 1174 22933 1238
rect 22281 1090 22345 1154
rect 22365 1090 22429 1154
rect 22449 1090 22513 1154
rect 22533 1090 22597 1154
rect 22617 1090 22681 1154
rect 22701 1090 22765 1154
rect 22785 1090 22849 1154
rect 22869 1090 22933 1154
rect 22281 1006 22345 1070
rect 22365 1006 22429 1070
rect 22449 1006 22513 1070
rect 22533 1006 22597 1070
rect 22617 1006 22681 1070
rect 22701 1006 22765 1070
rect 22785 1006 22849 1070
rect 22869 1006 22933 1070
rect 22281 922 22345 986
rect 22365 922 22429 986
rect 22449 922 22513 986
rect 22533 922 22597 986
rect 22617 922 22681 986
rect 22701 922 22765 986
rect 22785 922 22849 986
rect 22869 922 22933 986
rect 22281 838 22345 902
rect 22365 838 22429 902
rect 22449 838 22513 902
rect 22533 838 22597 902
rect 22617 838 22681 902
rect 22701 838 22765 902
rect 22785 838 22849 902
rect 22869 838 22933 902
rect 22281 754 22345 818
rect 22365 754 22429 818
rect 22449 754 22513 818
rect 22533 754 22597 818
rect 22617 754 22681 818
rect 22701 754 22765 818
rect 22785 754 22849 818
rect 22869 754 22933 818
rect 22281 670 22345 734
rect 22365 670 22429 734
rect 22449 670 22513 734
rect 22533 670 22597 734
rect 22617 670 22681 734
rect 22701 670 22765 734
rect 22785 670 22849 734
rect 22869 670 22933 734
rect 22281 586 22345 650
rect 22365 586 22429 650
rect 22449 586 22513 650
rect 22533 586 22597 650
rect 22617 586 22681 650
rect 22701 586 22765 650
rect 22785 586 22849 650
rect 22869 586 22933 650
rect 22281 502 22345 566
rect 22365 502 22429 566
rect 22449 502 22513 566
rect 22533 502 22597 566
rect 22617 502 22681 566
rect 22701 502 22765 566
rect 22785 502 22849 566
rect 22869 502 22933 566
rect 22281 418 22345 482
rect 22365 418 22429 482
rect 22449 418 22513 482
rect 22533 418 22597 482
rect 22617 418 22681 482
rect 22701 418 22765 482
rect 22785 418 22849 482
rect 22869 418 22933 482
rect 23886 18927 23950 18991
rect 23886 18846 23950 18910
rect 23886 18765 23950 18829
rect 23886 18684 23950 18748
rect 23886 18602 23950 18666
rect 23886 18520 23950 18584
rect 23886 18438 23950 18502
rect 23886 18356 23950 18420
rect 23886 18274 23950 18338
rect 23886 18192 23950 18256
rect 23886 18110 23950 18174
rect 23886 18028 23950 18092
rect 23886 17946 23950 18010
rect 23886 17864 23950 17928
rect 23886 17782 23950 17846
rect 23886 17700 23950 17764
rect 23886 17618 23950 17682
rect 23886 17536 23950 17600
rect 23886 17454 23950 17518
rect 23886 17372 23950 17436
rect 23886 17290 23950 17354
rect 23886 17208 23950 17272
rect 23886 17126 23950 17190
rect 23886 17044 23950 17108
rect 23886 16962 23950 17026
rect 23886 16880 23950 16944
rect 23886 16798 23950 16862
rect 23886 16716 23950 16780
rect 23886 16634 23950 16698
rect 23886 16552 23950 16616
rect 24565 13634 24629 13698
rect 24667 13634 24731 13698
rect 24769 13634 24833 13698
rect 24871 13634 24935 13698
rect 24565 13554 24629 13618
rect 24667 13554 24731 13618
rect 24769 13554 24833 13618
rect 24871 13554 24935 13618
rect 24565 13474 24629 13538
rect 24667 13474 24731 13538
rect 24769 13474 24833 13538
rect 24871 13474 24935 13538
rect 24565 13394 24629 13458
rect 24667 13394 24731 13458
rect 24769 13394 24833 13458
rect 24871 13394 24935 13458
rect 24565 13314 24629 13378
rect 24667 13314 24731 13378
rect 24769 13314 24833 13378
rect 24871 13314 24935 13378
rect 24565 13234 24629 13298
rect 24667 13234 24731 13298
rect 24769 13234 24833 13298
rect 24871 13234 24935 13298
rect 24565 13154 24629 13218
rect 24667 13154 24731 13218
rect 24769 13154 24833 13218
rect 24871 13154 24935 13218
rect 24565 13074 24629 13138
rect 24667 13074 24731 13138
rect 24769 13074 24833 13138
rect 24871 13074 24935 13138
rect 24565 12994 24629 13058
rect 24667 12994 24731 13058
rect 24769 12994 24833 13058
rect 24871 12994 24935 13058
rect 24565 12914 24629 12978
rect 24667 12914 24731 12978
rect 24769 12914 24833 12978
rect 24871 12914 24935 12978
rect 24565 12834 24629 12898
rect 24667 12834 24731 12898
rect 24769 12834 24833 12898
rect 24871 12834 24935 12898
rect 23784 7959 23848 8023
rect 23890 7959 23954 8023
rect 23996 7959 24060 8023
rect 24102 7959 24166 8023
rect 23784 7875 23848 7939
rect 23890 7875 23954 7939
rect 23996 7875 24060 7939
rect 24102 7875 24166 7939
rect 23784 7790 23848 7854
rect 23890 7790 23954 7854
rect 23996 7790 24060 7854
rect 24102 7790 24166 7854
rect 23784 7705 23848 7769
rect 23890 7705 23954 7769
rect 23996 7705 24060 7769
rect 24102 7705 24166 7769
rect 23784 7620 23848 7684
rect 23890 7620 23954 7684
rect 23996 7620 24060 7684
rect 24102 7620 24166 7684
rect 23784 7535 23848 7599
rect 23890 7535 23954 7599
rect 23996 7535 24060 7599
rect 24102 7535 24166 7599
rect 23784 7450 23848 7514
rect 23890 7450 23954 7514
rect 23996 7450 24060 7514
rect 24102 7450 24166 7514
rect 24514 1612 24578 1676
rect 24594 1612 24658 1676
rect 24805 1612 24869 1676
rect 24885 1612 24949 1676
rect 27653 2628 27717 2692
rect 27743 2628 27807 2692
rect 27833 2628 27897 2692
rect 27923 2628 27987 2692
rect 27653 2544 27717 2608
rect 27743 2544 27807 2608
rect 27833 2544 27897 2608
rect 27923 2544 27987 2608
rect 27653 2460 27717 2524
rect 27743 2460 27807 2524
rect 27833 2460 27897 2524
rect 27923 2460 27987 2524
rect 27653 2376 27717 2440
rect 27743 2376 27807 2440
rect 27833 2376 27897 2440
rect 27923 2376 27987 2440
rect 27653 2292 27717 2356
rect 27743 2292 27807 2356
rect 27833 2292 27897 2356
rect 27923 2292 27987 2356
rect 27653 2208 27717 2272
rect 27743 2208 27807 2272
rect 27833 2208 27897 2272
rect 27923 2208 27987 2272
rect 27653 2124 27717 2188
rect 27743 2124 27807 2188
rect 27833 2124 27897 2188
rect 27923 2124 27987 2188
rect 27653 2040 27717 2104
rect 27743 2040 27807 2104
rect 27833 2040 27897 2104
rect 27923 2040 27987 2104
rect 27653 1956 27717 2020
rect 27743 1956 27807 2020
rect 27833 1956 27897 2020
rect 27923 1956 27987 2020
rect 27653 1872 27717 1936
rect 27743 1872 27807 1936
rect 27833 1872 27897 1936
rect 27923 1872 27987 1936
rect 27653 1787 27717 1851
rect 27743 1787 27807 1851
rect 27833 1787 27897 1851
rect 27923 1787 27987 1851
<< metal4 >>
rect 0 35157 254 40000
rect 23395 36247 23697 36248
rect 23395 36183 23396 36247
rect 23460 36183 23514 36247
rect 23578 36183 23632 36247
rect 23696 36183 23697 36247
rect 23395 36164 23697 36183
rect 23395 36100 23396 36164
rect 23460 36100 23514 36164
rect 23578 36100 23632 36164
rect 23696 36100 23697 36164
rect 23395 36081 23697 36100
rect 23395 36017 23396 36081
rect 23460 36017 23514 36081
rect 23578 36017 23632 36081
rect 23696 36017 23697 36081
rect 23395 35998 23697 36017
rect 23395 35934 23396 35998
rect 23460 35934 23514 35998
rect 23578 35934 23632 35998
rect 23696 35934 23697 35998
rect 23395 35915 23697 35934
rect 23395 35851 23396 35915
rect 23460 35851 23514 35915
rect 23578 35851 23632 35915
rect 23696 35851 23697 35915
rect 23395 35832 23697 35851
rect 23395 35768 23396 35832
rect 23460 35768 23514 35832
rect 23578 35768 23632 35832
rect 23696 35768 23697 35832
rect 23395 35749 23697 35768
rect 23395 35685 23396 35749
rect 23460 35685 23514 35749
rect 23578 35685 23632 35749
rect 23696 35685 23697 35749
rect 23395 35666 23697 35685
rect 19257 35626 22590 35627
rect 19257 35562 19258 35626
rect 19322 35562 19340 35626
rect 19404 35562 19422 35626
rect 19486 35562 19504 35626
rect 19568 35562 19586 35626
rect 19650 35562 19668 35626
rect 19732 35562 19750 35626
rect 19814 35562 19832 35626
rect 19896 35562 19914 35626
rect 19978 35562 19996 35626
rect 20060 35562 20078 35626
rect 20142 35562 20160 35626
rect 20224 35562 20242 35626
rect 20306 35562 20324 35626
rect 20388 35562 20406 35626
rect 20470 35562 20488 35626
rect 20552 35562 20570 35626
rect 20634 35562 20652 35626
rect 20716 35562 20734 35626
rect 20798 35562 20816 35626
rect 20880 35562 20898 35626
rect 20962 35562 20980 35626
rect 21044 35562 21062 35626
rect 21126 35562 21144 35626
rect 21208 35562 21226 35626
rect 21290 35562 21308 35626
rect 21372 35562 21390 35626
rect 21454 35562 21472 35626
rect 21536 35562 21553 35626
rect 21617 35562 21634 35626
rect 21698 35562 21715 35626
rect 21779 35562 21796 35626
rect 21860 35562 21877 35626
rect 21941 35562 21958 35626
rect 22022 35562 22039 35626
rect 22103 35562 22120 35626
rect 22184 35562 22201 35626
rect 22265 35562 22282 35626
rect 22346 35562 22363 35626
rect 22427 35562 22444 35626
rect 22508 35562 22525 35626
rect 22589 35562 22590 35626
rect 19257 35546 22590 35562
rect 19257 35482 19258 35546
rect 19322 35482 19340 35546
rect 19404 35482 19422 35546
rect 19486 35482 19504 35546
rect 19568 35482 19586 35546
rect 19650 35482 19668 35546
rect 19732 35482 19750 35546
rect 19814 35482 19832 35546
rect 19896 35482 19914 35546
rect 19978 35482 19996 35546
rect 20060 35482 20078 35546
rect 20142 35482 20160 35546
rect 20224 35482 20242 35546
rect 20306 35482 20324 35546
rect 20388 35482 20406 35546
rect 20470 35482 20488 35546
rect 20552 35482 20570 35546
rect 20634 35482 20652 35546
rect 20716 35482 20734 35546
rect 20798 35482 20816 35546
rect 20880 35482 20898 35546
rect 20962 35482 20980 35546
rect 21044 35482 21062 35546
rect 21126 35482 21144 35546
rect 21208 35482 21226 35546
rect 21290 35482 21308 35546
rect 21372 35482 21390 35546
rect 21454 35482 21472 35546
rect 21536 35482 21553 35546
rect 21617 35482 21634 35546
rect 21698 35482 21715 35546
rect 21779 35482 21796 35546
rect 21860 35482 21877 35546
rect 21941 35482 21958 35546
rect 22022 35482 22039 35546
rect 22103 35482 22120 35546
rect 22184 35482 22201 35546
rect 22265 35482 22282 35546
rect 22346 35482 22363 35546
rect 22427 35482 22444 35546
rect 22508 35482 22525 35546
rect 22589 35482 22590 35546
rect 19257 35466 22590 35482
rect 19257 35402 19258 35466
rect 19322 35402 19340 35466
rect 19404 35402 19422 35466
rect 19486 35402 19504 35466
rect 19568 35402 19586 35466
rect 19650 35402 19668 35466
rect 19732 35402 19750 35466
rect 19814 35402 19832 35466
rect 19896 35402 19914 35466
rect 19978 35402 19996 35466
rect 20060 35402 20078 35466
rect 20142 35402 20160 35466
rect 20224 35402 20242 35466
rect 20306 35402 20324 35466
rect 20388 35402 20406 35466
rect 20470 35402 20488 35466
rect 20552 35402 20570 35466
rect 20634 35402 20652 35466
rect 20716 35402 20734 35466
rect 20798 35402 20816 35466
rect 20880 35402 20898 35466
rect 20962 35402 20980 35466
rect 21044 35402 21062 35466
rect 21126 35402 21144 35466
rect 21208 35402 21226 35466
rect 21290 35402 21308 35466
rect 21372 35402 21390 35466
rect 21454 35402 21472 35466
rect 21536 35402 21553 35466
rect 21617 35402 21634 35466
rect 21698 35402 21715 35466
rect 21779 35402 21796 35466
rect 21860 35402 21877 35466
rect 21941 35402 21958 35466
rect 22022 35402 22039 35466
rect 22103 35402 22120 35466
rect 22184 35402 22201 35466
rect 22265 35402 22282 35466
rect 22346 35402 22363 35466
rect 22427 35402 22444 35466
rect 22508 35402 22525 35466
rect 22589 35402 22590 35466
rect 19257 35386 22590 35402
rect 19257 35322 19258 35386
rect 19322 35322 19340 35386
rect 19404 35322 19422 35386
rect 19486 35322 19504 35386
rect 19568 35322 19586 35386
rect 19650 35322 19668 35386
rect 19732 35322 19750 35386
rect 19814 35322 19832 35386
rect 19896 35322 19914 35386
rect 19978 35322 19996 35386
rect 20060 35322 20078 35386
rect 20142 35322 20160 35386
rect 20224 35322 20242 35386
rect 20306 35322 20324 35386
rect 20388 35322 20406 35386
rect 20470 35322 20488 35386
rect 20552 35322 20570 35386
rect 20634 35322 20652 35386
rect 20716 35322 20734 35386
rect 20798 35322 20816 35386
rect 20880 35322 20898 35386
rect 20962 35322 20980 35386
rect 21044 35322 21062 35386
rect 21126 35322 21144 35386
rect 21208 35322 21226 35386
rect 21290 35322 21308 35386
rect 21372 35322 21390 35386
rect 21454 35322 21472 35386
rect 21536 35322 21553 35386
rect 21617 35322 21634 35386
rect 21698 35322 21715 35386
rect 21779 35322 21796 35386
rect 21860 35322 21877 35386
rect 21941 35322 21958 35386
rect 22022 35322 22039 35386
rect 22103 35322 22120 35386
rect 22184 35322 22201 35386
rect 22265 35322 22282 35386
rect 22346 35322 22363 35386
rect 22427 35322 22444 35386
rect 22508 35322 22525 35386
rect 22589 35322 22590 35386
rect 19257 35306 22590 35322
rect 19257 35242 19258 35306
rect 19322 35242 19340 35306
rect 19404 35242 19422 35306
rect 19486 35242 19504 35306
rect 19568 35242 19586 35306
rect 19650 35242 19668 35306
rect 19732 35242 19750 35306
rect 19814 35242 19832 35306
rect 19896 35242 19914 35306
rect 19978 35242 19996 35306
rect 20060 35242 20078 35306
rect 20142 35242 20160 35306
rect 20224 35242 20242 35306
rect 20306 35242 20324 35306
rect 20388 35242 20406 35306
rect 20470 35242 20488 35306
rect 20552 35242 20570 35306
rect 20634 35242 20652 35306
rect 20716 35242 20734 35306
rect 20798 35242 20816 35306
rect 20880 35242 20898 35306
rect 20962 35242 20980 35306
rect 21044 35242 21062 35306
rect 21126 35242 21144 35306
rect 21208 35242 21226 35306
rect 21290 35242 21308 35306
rect 21372 35242 21390 35306
rect 21454 35242 21472 35306
rect 21536 35242 21553 35306
rect 21617 35242 21634 35306
rect 21698 35242 21715 35306
rect 21779 35242 21796 35306
rect 21860 35242 21877 35306
rect 21941 35242 21958 35306
rect 22022 35242 22039 35306
rect 22103 35242 22120 35306
rect 22184 35242 22201 35306
rect 22265 35242 22282 35306
rect 22346 35242 22363 35306
rect 22427 35242 22444 35306
rect 22508 35242 22525 35306
rect 22589 35242 22590 35306
rect 19257 35226 22590 35242
rect 19257 35162 19258 35226
rect 19322 35162 19340 35226
rect 19404 35162 19422 35226
rect 19486 35162 19504 35226
rect 19568 35162 19586 35226
rect 19650 35162 19668 35226
rect 19732 35162 19750 35226
rect 19814 35162 19832 35226
rect 19896 35162 19914 35226
rect 19978 35162 19996 35226
rect 20060 35162 20078 35226
rect 20142 35162 20160 35226
rect 20224 35162 20242 35226
rect 20306 35162 20324 35226
rect 20388 35162 20406 35226
rect 20470 35162 20488 35226
rect 20552 35162 20570 35226
rect 20634 35162 20652 35226
rect 20716 35162 20734 35226
rect 20798 35162 20816 35226
rect 20880 35162 20898 35226
rect 20962 35162 20980 35226
rect 21044 35162 21062 35226
rect 21126 35162 21144 35226
rect 21208 35162 21226 35226
rect 21290 35162 21308 35226
rect 21372 35162 21390 35226
rect 21454 35162 21472 35226
rect 21536 35162 21553 35226
rect 21617 35162 21634 35226
rect 21698 35162 21715 35226
rect 21779 35162 21796 35226
rect 21860 35162 21877 35226
rect 21941 35162 21958 35226
rect 22022 35162 22039 35226
rect 22103 35162 22120 35226
rect 22184 35162 22201 35226
rect 22265 35162 22282 35226
rect 22346 35162 22363 35226
rect 22427 35162 22444 35226
rect 22508 35162 22525 35226
rect 22589 35162 22590 35226
rect 23395 35602 23396 35666
rect 23460 35602 23514 35666
rect 23578 35602 23632 35666
rect 23696 35602 23697 35666
rect 23395 35583 23697 35602
rect 23395 35519 23396 35583
rect 23460 35519 23514 35583
rect 23578 35519 23632 35583
rect 23696 35519 23697 35583
rect 23395 35500 23697 35519
rect 23395 35436 23396 35500
rect 23460 35436 23514 35500
rect 23578 35436 23632 35500
rect 23696 35436 23697 35500
rect 23395 35417 23697 35436
rect 23395 35353 23396 35417
rect 23460 35353 23514 35417
rect 23578 35353 23632 35417
rect 23696 35353 23697 35417
rect 23395 35333 23697 35353
rect 23395 35269 23396 35333
rect 23460 35269 23514 35333
rect 23578 35269 23632 35333
rect 23696 35269 23697 35333
rect 23395 35249 23697 35269
rect 23395 35185 23396 35249
rect 23460 35185 23514 35249
rect 23578 35185 23632 35249
rect 23696 35185 23697 35249
rect 23395 35184 23697 35185
rect 19257 35161 22590 35162
rect 27746 35157 28000 40000
rect 3717 33111 3999 33112
rect 3717 33047 3718 33111
rect 3782 33047 3826 33111
rect 3890 33047 3934 33111
rect 3998 33047 3999 33111
rect 3717 33014 3999 33047
rect 3717 32950 3718 33014
rect 3782 32950 3826 33014
rect 3890 32950 3934 33014
rect 3998 32950 3999 33014
rect 3717 32917 3999 32950
rect 3717 32853 3718 32917
rect 3782 32853 3826 32917
rect 3890 32853 3934 32917
rect 3998 32853 3999 32917
rect 3717 32820 3999 32853
rect 3717 32756 3718 32820
rect 3782 32756 3826 32820
rect 3890 32756 3934 32820
rect 3998 32756 3999 32820
rect 3717 32722 3999 32756
rect 3717 32658 3718 32722
rect 3782 32658 3826 32722
rect 3890 32658 3934 32722
rect 3998 32658 3999 32722
rect 3717 32657 3999 32658
rect 1015 24578 1109 24579
rect 1015 24514 1016 24578
rect 1080 24522 1109 24578
tri 1109 24522 1166 24579 sw
rect 1080 24514 2257 24522
rect 1015 24470 2257 24514
rect 1015 24406 1016 24470
rect 1080 24406 2257 24470
rect 1015 24362 2257 24406
rect 1015 24298 1016 24362
rect 1080 24346 2257 24362
rect 2259 24346 2504 24522
rect 1080 24298 1092 24346
rect 1015 24297 1092 24298
tri 1092 24297 1141 24346 nw
rect 0 14007 254 19000
rect 23848 18991 23988 18992
rect 23848 18927 23886 18991
rect 23950 18927 23988 18991
rect 23848 18910 23988 18927
rect 23848 18846 23886 18910
rect 23950 18846 23988 18910
rect 23848 18829 23988 18846
rect 23848 18765 23886 18829
rect 23950 18765 23988 18829
rect 23848 18748 23988 18765
rect 23848 18684 23886 18748
rect 23950 18684 23988 18748
rect 23848 18666 23988 18684
rect 23848 18602 23886 18666
rect 23950 18602 23988 18666
rect 23848 18584 23988 18602
rect 23848 18520 23886 18584
rect 23950 18520 23988 18584
rect 23848 18502 23988 18520
rect 23848 18438 23886 18502
rect 23950 18438 23988 18502
rect 23848 18420 23988 18438
rect 23848 18356 23886 18420
rect 23950 18356 23988 18420
rect 23848 18338 23988 18356
rect 23848 18274 23886 18338
rect 23950 18274 23988 18338
rect 23848 18256 23988 18274
rect 23848 18192 23886 18256
rect 23950 18192 23988 18256
rect 23848 18174 23988 18192
rect 23848 18110 23886 18174
rect 23950 18110 23988 18174
rect 23848 18092 23988 18110
rect 23848 18028 23886 18092
rect 23950 18028 23988 18092
rect 23848 18010 23988 18028
rect 23848 17946 23886 18010
rect 23950 17946 23988 18010
rect 23848 17928 23988 17946
rect 23848 17864 23886 17928
rect 23950 17864 23988 17928
rect 23848 17846 23988 17864
rect 23848 17782 23886 17846
rect 23950 17782 23988 17846
rect 23848 17764 23988 17782
rect 23848 17700 23886 17764
rect 23950 17700 23988 17764
rect 23848 17682 23988 17700
rect 23848 17618 23886 17682
rect 23950 17618 23988 17682
rect 23848 17600 23988 17618
rect 23848 17536 23886 17600
rect 23950 17536 23988 17600
rect 23848 17518 23988 17536
rect 23848 17454 23886 17518
rect 23950 17454 23988 17518
rect 23848 17436 23988 17454
rect 23848 17372 23886 17436
rect 23950 17372 23988 17436
rect 23848 17354 23988 17372
rect 23848 17290 23886 17354
rect 23950 17290 23988 17354
rect 23848 17272 23988 17290
rect 23848 17208 23886 17272
rect 23950 17208 23988 17272
rect 23848 17190 23988 17208
rect 23848 17126 23886 17190
rect 23950 17126 23988 17190
rect 23848 17108 23988 17126
rect 23848 17044 23886 17108
rect 23950 17044 23988 17108
rect 23848 17026 23988 17044
rect 23848 16962 23886 17026
rect 23950 16962 23988 17026
rect 23848 16944 23988 16962
rect 23848 16880 23886 16944
rect 23950 16880 23988 16944
rect 23848 16862 23988 16880
rect 23848 16798 23886 16862
rect 23950 16798 23988 16862
rect 23848 16780 23988 16798
rect 23848 16716 23886 16780
rect 23950 16716 23988 16780
rect 23848 16698 23988 16716
rect 23848 16634 23886 16698
rect 23950 16634 23988 16698
rect 23848 16616 23988 16634
rect 23848 16552 23886 16616
rect 23950 16552 23988 16616
rect 23848 16551 23988 16552
rect 27746 14007 28000 19000
rect 0 12817 254 13707
rect 6853 13697 7769 13699
rect 6853 13633 6854 13697
rect 6918 13633 6939 13697
rect 7003 13633 7024 13697
rect 7088 13633 7109 13697
rect 7173 13633 7194 13697
rect 7258 13633 7279 13697
rect 7343 13633 7364 13697
rect 7428 13633 7449 13697
rect 7513 13633 7534 13697
rect 7598 13633 7619 13697
rect 7683 13633 7704 13697
rect 7768 13633 7769 13697
rect 24564 13698 24936 13699
rect 6853 13609 7769 13633
rect 6853 13545 6854 13609
rect 6918 13545 6939 13609
rect 7003 13545 7024 13609
rect 7088 13545 7109 13609
rect 7173 13545 7194 13609
rect 7258 13545 7279 13609
rect 7343 13545 7364 13609
rect 7428 13545 7449 13609
rect 7513 13545 7534 13609
rect 7598 13545 7619 13609
rect 7683 13545 7704 13609
rect 7768 13545 7769 13609
rect 6853 13521 7769 13545
rect 6853 13457 6854 13521
rect 6918 13457 6939 13521
rect 7003 13457 7024 13521
rect 7088 13457 7109 13521
rect 7173 13457 7194 13521
rect 7258 13457 7279 13521
rect 7343 13457 7364 13521
rect 7428 13457 7449 13521
rect 7513 13457 7534 13521
rect 7598 13457 7619 13521
rect 7683 13457 7704 13521
rect 7768 13457 7769 13521
rect 6853 13455 7769 13457
rect 16059 13684 16936 13688
rect 16059 13620 16060 13684
rect 16124 13620 16142 13684
rect 16206 13620 16223 13684
rect 16287 13620 16304 13684
rect 16368 13620 16385 13684
rect 16449 13620 16466 13684
rect 16530 13620 16547 13684
rect 16611 13620 16628 13684
rect 16692 13620 16709 13684
rect 16773 13620 16790 13684
rect 16854 13620 16871 13684
rect 16935 13620 16936 13684
rect 16059 13596 16936 13620
rect 16059 13532 16060 13596
rect 16124 13532 16142 13596
rect 16206 13532 16223 13596
rect 16287 13532 16304 13596
rect 16368 13532 16385 13596
rect 16449 13532 16466 13596
rect 16530 13532 16547 13596
rect 16611 13532 16628 13596
rect 16692 13532 16709 13596
rect 16773 13532 16790 13596
rect 16854 13532 16871 13596
rect 16935 13532 16936 13596
rect 16059 13508 16936 13532
rect 16059 13444 16060 13508
rect 16124 13444 16142 13508
rect 16206 13444 16223 13508
rect 16287 13444 16304 13508
rect 16368 13444 16385 13508
rect 16449 13444 16466 13508
rect 16530 13444 16547 13508
rect 16611 13444 16628 13508
rect 16692 13444 16709 13508
rect 16773 13444 16790 13508
rect 16854 13444 16871 13508
rect 16935 13444 16936 13508
rect 16059 13420 16936 13444
rect 16059 13356 16060 13420
rect 16124 13356 16142 13420
rect 16206 13356 16223 13420
rect 16287 13356 16304 13420
rect 16368 13356 16385 13420
rect 16449 13356 16466 13420
rect 16530 13356 16547 13420
rect 16611 13356 16628 13420
rect 16692 13356 16709 13420
rect 16773 13356 16790 13420
rect 16854 13356 16871 13420
rect 16935 13356 16936 13420
rect 16059 13332 16936 13356
rect 16059 13268 16060 13332
rect 16124 13268 16142 13332
rect 16206 13268 16223 13332
rect 16287 13268 16304 13332
rect 16368 13268 16385 13332
rect 16449 13268 16466 13332
rect 16530 13268 16547 13332
rect 16611 13268 16628 13332
rect 16692 13268 16709 13332
rect 16773 13268 16790 13332
rect 16854 13268 16871 13332
rect 16935 13268 16936 13332
rect 16059 13244 16936 13268
rect 16059 13180 16060 13244
rect 16124 13180 16142 13244
rect 16206 13180 16223 13244
rect 16287 13180 16304 13244
rect 16368 13180 16385 13244
rect 16449 13180 16466 13244
rect 16530 13180 16547 13244
rect 16611 13180 16628 13244
rect 16692 13180 16709 13244
rect 16773 13180 16790 13244
rect 16854 13180 16871 13244
rect 16935 13180 16936 13244
rect 16059 13156 16936 13180
rect 16059 13092 16060 13156
rect 16124 13092 16142 13156
rect 16206 13092 16223 13156
rect 16287 13092 16304 13156
rect 16368 13092 16385 13156
rect 16449 13092 16466 13156
rect 16530 13092 16547 13156
rect 16611 13092 16628 13156
rect 16692 13092 16709 13156
rect 16773 13092 16790 13156
rect 16854 13092 16871 13156
rect 16935 13092 16936 13156
rect 16059 13068 16936 13092
rect 16059 13004 16060 13068
rect 16124 13004 16142 13068
rect 16206 13004 16223 13068
rect 16287 13004 16304 13068
rect 16368 13004 16385 13068
rect 16449 13004 16466 13068
rect 16530 13004 16547 13068
rect 16611 13004 16628 13068
rect 16692 13004 16709 13068
rect 16773 13004 16790 13068
rect 16854 13004 16871 13068
rect 16935 13004 16936 13068
rect 16059 12980 16936 13004
rect 16059 12916 16060 12980
rect 16124 12916 16142 12980
rect 16206 12916 16223 12980
rect 16287 12916 16304 12980
rect 16368 12916 16385 12980
rect 16449 12916 16466 12980
rect 16530 12916 16547 12980
rect 16611 12916 16628 12980
rect 16692 12916 16709 12980
rect 16773 12916 16790 12980
rect 16854 12916 16871 12980
rect 16935 12916 16936 12980
rect 16059 12892 16936 12916
rect 16059 12828 16060 12892
rect 16124 12828 16142 12892
rect 16206 12828 16223 12892
rect 16287 12828 16304 12892
rect 16368 12828 16385 12892
rect 16449 12828 16466 12892
rect 16530 12828 16547 12892
rect 16611 12828 16628 12892
rect 16692 12828 16709 12892
rect 16773 12828 16790 12892
rect 16854 12828 16871 12892
rect 16935 12828 16936 12892
rect 24564 13634 24565 13698
rect 24629 13634 24667 13698
rect 24731 13634 24769 13698
rect 24833 13634 24871 13698
rect 24935 13634 24936 13698
rect 24564 13618 24936 13634
rect 24564 13554 24565 13618
rect 24629 13554 24667 13618
rect 24731 13554 24769 13618
rect 24833 13554 24871 13618
rect 24935 13554 24936 13618
rect 24564 13538 24936 13554
rect 24564 13474 24565 13538
rect 24629 13474 24667 13538
rect 24731 13474 24769 13538
rect 24833 13474 24871 13538
rect 24935 13474 24936 13538
rect 24564 13458 24936 13474
rect 24564 13394 24565 13458
rect 24629 13394 24667 13458
rect 24731 13394 24769 13458
rect 24833 13394 24871 13458
rect 24935 13394 24936 13458
rect 24564 13378 24936 13394
rect 24564 13314 24565 13378
rect 24629 13314 24667 13378
rect 24731 13314 24769 13378
rect 24833 13314 24871 13378
rect 24935 13314 24936 13378
rect 24564 13298 24936 13314
rect 24564 13234 24565 13298
rect 24629 13234 24667 13298
rect 24731 13234 24769 13298
rect 24833 13234 24871 13298
rect 24935 13234 24936 13298
rect 24564 13218 24936 13234
rect 24564 13154 24565 13218
rect 24629 13154 24667 13218
rect 24731 13154 24769 13218
rect 24833 13154 24871 13218
rect 24935 13154 24936 13218
rect 24564 13138 24936 13154
rect 24564 13074 24565 13138
rect 24629 13074 24667 13138
rect 24731 13074 24769 13138
rect 24833 13074 24871 13138
rect 24935 13074 24936 13138
rect 24564 13058 24936 13074
rect 24564 12994 24565 13058
rect 24629 12994 24667 13058
rect 24731 12994 24769 13058
rect 24833 12994 24871 13058
rect 24935 12994 24936 13058
rect 24564 12978 24936 12994
rect 24564 12914 24565 12978
rect 24629 12914 24667 12978
rect 24731 12914 24769 12978
rect 24833 12914 24871 12978
rect 24935 12914 24936 12978
rect 24564 12898 24936 12914
rect 24564 12834 24565 12898
rect 24629 12834 24667 12898
rect 24731 12834 24769 12898
rect 24833 12834 24871 12898
rect 24935 12834 24936 12898
rect 24564 12833 24936 12834
rect 16059 12824 16936 12828
rect 27746 12817 28000 13707
rect 0 11647 254 12537
rect 27746 11647 28000 12537
rect 0 11281 254 11347
rect 27746 11281 28000 11347
rect 0 10625 254 11221
rect 27746 10625 28000 11221
rect 0 10329 254 10565
rect 27746 10329 28000 10565
rect 0 9673 254 10269
rect 27746 9673 28000 10269
rect 0 9547 254 9613
rect 27746 9547 28000 9613
rect 0 8317 254 9247
rect 1594 9240 2140 9241
rect 1594 9176 1595 9240
rect 1659 9176 1675 9240
rect 1739 9176 1755 9240
rect 1819 9176 1835 9240
rect 1899 9176 1915 9240
rect 1979 9176 1995 9240
rect 2059 9176 2075 9240
rect 2139 9176 2140 9240
rect 17879 9239 18185 9240
rect 14538 9235 15122 9236
rect 1594 9155 2140 9176
rect 1594 9091 1595 9155
rect 1659 9091 1675 9155
rect 1739 9091 1755 9155
rect 1819 9091 1835 9155
rect 1899 9091 1915 9155
rect 1979 9091 1995 9155
rect 2059 9091 2075 9155
rect 2139 9091 2140 9155
rect 1594 9070 2140 9091
rect 11514 9228 12098 9229
rect 11514 9164 11516 9228
rect 11580 9164 11602 9228
rect 11666 9164 11688 9228
rect 11752 9164 11774 9228
rect 11838 9164 11860 9228
rect 11924 9164 11946 9228
rect 12010 9164 12032 9228
rect 12096 9164 12098 9228
rect 11514 9145 12098 9164
rect 1594 9006 1595 9070
rect 1659 9006 1675 9070
rect 1739 9006 1755 9070
rect 1819 9006 1835 9070
rect 1899 9006 1915 9070
rect 1979 9006 1995 9070
rect 2059 9006 2075 9070
rect 2139 9006 2140 9070
rect 1594 8985 2140 9006
rect 1594 8921 1595 8985
rect 1659 8921 1675 8985
rect 1739 8921 1755 8985
rect 1819 8921 1835 8985
rect 1899 8921 1915 8985
rect 1979 8921 1995 8985
rect 2059 8921 2075 8985
rect 2139 8921 2140 8985
rect 1594 8900 2140 8921
rect 1594 8836 1595 8900
rect 1659 8836 1675 8900
rect 1739 8836 1755 8900
rect 1819 8836 1835 8900
rect 1899 8836 1915 8900
rect 1979 8836 1995 8900
rect 2059 8836 2075 8900
rect 2139 8836 2140 8900
rect 1594 8815 2140 8836
rect 1594 8751 1595 8815
rect 1659 8751 1675 8815
rect 1739 8751 1755 8815
rect 1819 8751 1835 8815
rect 1899 8751 1915 8815
rect 1979 8751 1995 8815
rect 2059 8751 2075 8815
rect 2139 8751 2140 8815
rect 1594 8730 2140 8751
rect 1594 8666 1595 8730
rect 1659 8666 1675 8730
rect 1739 8666 1755 8730
rect 1819 8666 1835 8730
rect 1899 8666 1915 8730
rect 1979 8666 1995 8730
rect 2059 8666 2075 8730
rect 2139 8666 2140 8730
rect 1594 8645 2140 8666
rect 1594 8581 1595 8645
rect 1659 8581 1675 8645
rect 1739 8581 1755 8645
rect 1819 8581 1835 8645
rect 1899 8581 1915 8645
rect 1979 8581 1995 8645
rect 2059 8581 2075 8645
rect 2139 8581 2140 8645
rect 1594 8560 2140 8581
rect 1594 8496 1595 8560
rect 1659 8496 1675 8560
rect 1739 8496 1755 8560
rect 1819 8496 1835 8560
rect 1899 8496 1915 8560
rect 1979 8496 1995 8560
rect 2059 8496 2075 8560
rect 2139 8496 2140 8560
rect 1594 8474 2140 8496
rect 1594 8410 1595 8474
rect 1659 8410 1675 8474
rect 1739 8410 1755 8474
rect 1819 8410 1835 8474
rect 1899 8410 1915 8474
rect 1979 8410 1995 8474
rect 2059 8410 2075 8474
rect 2139 8410 2140 8474
rect 1594 8388 2140 8410
rect 1594 8324 1595 8388
rect 1659 8324 1675 8388
rect 1739 8324 1755 8388
rect 1819 8324 1835 8388
rect 1899 8324 1915 8388
rect 1979 8324 1995 8388
rect 2059 8324 2075 8388
rect 2139 8324 2140 8388
rect 7445 9087 8027 9088
rect 7445 9023 7446 9087
rect 7510 9023 7532 9087
rect 7596 9023 7618 9087
rect 7682 9023 7704 9087
rect 7768 9023 7790 9087
rect 7854 9023 7876 9087
rect 7940 9023 7962 9087
rect 8026 9023 8027 9087
rect 7445 9001 8027 9023
rect 7445 8937 7446 9001
rect 7510 8937 7532 9001
rect 7596 8937 7618 9001
rect 7682 8937 7704 9001
rect 7768 8937 7790 9001
rect 7854 8937 7876 9001
rect 7940 8937 7962 9001
rect 8026 8937 8027 9001
rect 7445 8915 8027 8937
rect 7445 8851 7446 8915
rect 7510 8851 7532 8915
rect 7596 8851 7618 8915
rect 7682 8851 7704 8915
rect 7768 8851 7790 8915
rect 7854 8851 7876 8915
rect 7940 8851 7962 8915
rect 8026 8851 8027 8915
rect 7445 8829 8027 8851
rect 7445 8765 7446 8829
rect 7510 8765 7532 8829
rect 7596 8765 7618 8829
rect 7682 8765 7704 8829
rect 7768 8765 7790 8829
rect 7854 8765 7876 8829
rect 7940 8765 7962 8829
rect 8026 8765 8027 8829
rect 7445 8743 8027 8765
rect 7445 8679 7446 8743
rect 7510 8679 7532 8743
rect 7596 8679 7618 8743
rect 7682 8679 7704 8743
rect 7768 8679 7790 8743
rect 7854 8679 7876 8743
rect 7940 8679 7962 8743
rect 8026 8679 8027 8743
rect 7445 8657 8027 8679
rect 7445 8593 7446 8657
rect 7510 8593 7532 8657
rect 7596 8593 7618 8657
rect 7682 8593 7704 8657
rect 7768 8593 7790 8657
rect 7854 8593 7876 8657
rect 7940 8593 7962 8657
rect 8026 8593 8027 8657
rect 7445 8571 8027 8593
rect 7445 8507 7446 8571
rect 7510 8507 7532 8571
rect 7596 8507 7618 8571
rect 7682 8507 7704 8571
rect 7768 8507 7790 8571
rect 7854 8507 7876 8571
rect 7940 8507 7962 8571
rect 8026 8507 8027 8571
rect 7445 8484 8027 8507
rect 7445 8420 7446 8484
rect 7510 8420 7532 8484
rect 7596 8420 7618 8484
rect 7682 8420 7704 8484
rect 7768 8420 7790 8484
rect 7854 8420 7876 8484
rect 7940 8420 7962 8484
rect 8026 8420 8027 8484
rect 7445 8397 8027 8420
rect 7445 8333 7446 8397
rect 7510 8333 7532 8397
rect 7596 8333 7618 8397
rect 7682 8333 7704 8397
rect 7768 8333 7790 8397
rect 7854 8333 7876 8397
rect 7940 8333 7962 8397
rect 8026 8333 8027 8397
rect 7445 8332 8027 8333
rect 11514 9081 11516 9145
rect 11580 9081 11602 9145
rect 11666 9081 11688 9145
rect 11752 9081 11774 9145
rect 11838 9081 11860 9145
rect 11924 9081 11946 9145
rect 12010 9081 12032 9145
rect 12096 9081 12098 9145
rect 11514 9062 12098 9081
rect 11514 8998 11516 9062
rect 11580 8998 11602 9062
rect 11666 8998 11688 9062
rect 11752 8998 11774 9062
rect 11838 8998 11860 9062
rect 11924 8998 11946 9062
rect 12010 8998 12032 9062
rect 12096 8998 12098 9062
rect 11514 8979 12098 8998
rect 11514 8915 11516 8979
rect 11580 8915 11602 8979
rect 11666 8915 11688 8979
rect 11752 8915 11774 8979
rect 11838 8915 11860 8979
rect 11924 8915 11946 8979
rect 12010 8915 12032 8979
rect 12096 8915 12098 8979
rect 11514 8896 12098 8915
rect 11514 8832 11516 8896
rect 11580 8832 11602 8896
rect 11666 8832 11688 8896
rect 11752 8832 11774 8896
rect 11838 8832 11860 8896
rect 11924 8832 11946 8896
rect 12010 8832 12032 8896
rect 12096 8832 12098 8896
rect 11514 8813 12098 8832
rect 11514 8749 11516 8813
rect 11580 8749 11602 8813
rect 11666 8749 11688 8813
rect 11752 8749 11774 8813
rect 11838 8749 11860 8813
rect 11924 8749 11946 8813
rect 12010 8749 12032 8813
rect 12096 8749 12098 8813
rect 11514 8730 12098 8749
rect 11514 8666 11516 8730
rect 11580 8666 11602 8730
rect 11666 8666 11688 8730
rect 11752 8666 11774 8730
rect 11838 8666 11860 8730
rect 11924 8666 11946 8730
rect 12010 8666 12032 8730
rect 12096 8666 12098 8730
rect 11514 8647 12098 8666
rect 11514 8583 11516 8647
rect 11580 8583 11602 8647
rect 11666 8583 11688 8647
rect 11752 8583 11774 8647
rect 11838 8583 11860 8647
rect 11924 8583 11946 8647
rect 12010 8583 12032 8647
rect 12096 8583 12098 8647
rect 11514 8564 12098 8583
rect 11514 8500 11516 8564
rect 11580 8500 11602 8564
rect 11666 8500 11688 8564
rect 11752 8500 11774 8564
rect 11838 8500 11860 8564
rect 11924 8500 11946 8564
rect 12010 8500 12032 8564
rect 12096 8500 12098 8564
rect 11514 8480 12098 8500
rect 11514 8416 11516 8480
rect 11580 8416 11602 8480
rect 11666 8416 11688 8480
rect 11752 8416 11774 8480
rect 11838 8416 11860 8480
rect 11924 8416 11946 8480
rect 12010 8416 12032 8480
rect 12096 8416 12098 8480
rect 11514 8396 12098 8416
rect 11514 8332 11516 8396
rect 11580 8332 11602 8396
rect 11666 8332 11688 8396
rect 11752 8332 11774 8396
rect 11838 8332 11860 8396
rect 11924 8332 11946 8396
rect 12010 8332 12032 8396
rect 12096 8332 12098 8396
rect 11514 8331 12098 8332
rect 14538 9171 14540 9235
rect 14604 9171 14626 9235
rect 14690 9171 14712 9235
rect 14776 9171 14798 9235
rect 14862 9171 14884 9235
rect 14948 9171 14970 9235
rect 15034 9171 15056 9235
rect 15120 9171 15122 9235
rect 14538 9152 15122 9171
rect 14538 9088 14540 9152
rect 14604 9088 14626 9152
rect 14690 9088 14712 9152
rect 14776 9088 14798 9152
rect 14862 9088 14884 9152
rect 14948 9088 14970 9152
rect 15034 9088 15056 9152
rect 15120 9088 15122 9152
rect 14538 9068 15122 9088
rect 14538 9004 14540 9068
rect 14604 9004 14626 9068
rect 14690 9004 14712 9068
rect 14776 9004 14798 9068
rect 14862 9004 14884 9068
rect 14948 9004 14970 9068
rect 15034 9004 15056 9068
rect 15120 9004 15122 9068
rect 14538 8984 15122 9004
rect 14538 8920 14540 8984
rect 14604 8920 14626 8984
rect 14690 8920 14712 8984
rect 14776 8920 14798 8984
rect 14862 8920 14884 8984
rect 14948 8920 14970 8984
rect 15034 8920 15056 8984
rect 15120 8920 15122 8984
rect 14538 8900 15122 8920
rect 14538 8836 14540 8900
rect 14604 8836 14626 8900
rect 14690 8836 14712 8900
rect 14776 8836 14798 8900
rect 14862 8836 14884 8900
rect 14948 8836 14970 8900
rect 15034 8836 15056 8900
rect 15120 8836 15122 8900
rect 14538 8816 15122 8836
rect 14538 8752 14540 8816
rect 14604 8752 14626 8816
rect 14690 8752 14712 8816
rect 14776 8752 14798 8816
rect 14862 8752 14884 8816
rect 14948 8752 14970 8816
rect 15034 8752 15056 8816
rect 15120 8752 15122 8816
rect 14538 8732 15122 8752
rect 14538 8668 14540 8732
rect 14604 8668 14626 8732
rect 14690 8668 14712 8732
rect 14776 8668 14798 8732
rect 14862 8668 14884 8732
rect 14948 8668 14970 8732
rect 15034 8668 15056 8732
rect 15120 8668 15122 8732
rect 14538 8648 15122 8668
rect 14538 8584 14540 8648
rect 14604 8584 14626 8648
rect 14690 8584 14712 8648
rect 14776 8584 14798 8648
rect 14862 8584 14884 8648
rect 14948 8584 14970 8648
rect 15034 8584 15056 8648
rect 15120 8584 15122 8648
rect 14538 8564 15122 8584
rect 14538 8500 14540 8564
rect 14604 8500 14626 8564
rect 14690 8500 14712 8564
rect 14776 8500 14798 8564
rect 14862 8500 14884 8564
rect 14948 8500 14970 8564
rect 15034 8500 15056 8564
rect 15120 8500 15122 8564
rect 14538 8480 15122 8500
rect 14538 8416 14540 8480
rect 14604 8416 14626 8480
rect 14690 8416 14712 8480
rect 14776 8416 14798 8480
rect 14862 8416 14884 8480
rect 14948 8416 14970 8480
rect 15034 8416 15056 8480
rect 15120 8416 15122 8480
rect 14538 8396 15122 8416
rect 14538 8332 14540 8396
rect 14604 8332 14626 8396
rect 14690 8332 14712 8396
rect 14776 8332 14798 8396
rect 14862 8332 14884 8396
rect 14948 8332 14970 8396
rect 15034 8332 15056 8396
rect 15120 8332 15122 8396
rect 14538 8331 15122 8332
rect 17879 9175 17880 9239
rect 17944 9175 17960 9239
rect 18024 9175 18040 9239
rect 18104 9175 18120 9239
rect 18184 9175 18185 9239
rect 17879 9154 18185 9175
rect 17879 9090 17880 9154
rect 17944 9090 17960 9154
rect 18024 9090 18040 9154
rect 18104 9090 18120 9154
rect 18184 9090 18185 9154
rect 17879 9069 18185 9090
rect 17879 9005 17880 9069
rect 17944 9005 17960 9069
rect 18024 9005 18040 9069
rect 18104 9005 18120 9069
rect 18184 9005 18185 9069
rect 17879 8984 18185 9005
rect 17879 8920 17880 8984
rect 17944 8920 17960 8984
rect 18024 8920 18040 8984
rect 18104 8920 18120 8984
rect 18184 8920 18185 8984
rect 17879 8899 18185 8920
rect 17879 8835 17880 8899
rect 17944 8835 17960 8899
rect 18024 8835 18040 8899
rect 18104 8835 18120 8899
rect 18184 8835 18185 8899
rect 17879 8814 18185 8835
rect 17879 8750 17880 8814
rect 17944 8750 17960 8814
rect 18024 8750 18040 8814
rect 18104 8750 18120 8814
rect 18184 8750 18185 8814
rect 17879 8729 18185 8750
rect 17879 8665 17880 8729
rect 17944 8665 17960 8729
rect 18024 8665 18040 8729
rect 18104 8665 18120 8729
rect 18184 8665 18185 8729
rect 17879 8644 18185 8665
rect 17879 8580 17880 8644
rect 17944 8580 17960 8644
rect 18024 8580 18040 8644
rect 18104 8580 18120 8644
rect 18184 8580 18185 8644
rect 17879 8559 18185 8580
rect 17879 8495 17880 8559
rect 17944 8495 17960 8559
rect 18024 8495 18040 8559
rect 18104 8495 18120 8559
rect 18184 8495 18185 8559
rect 17879 8474 18185 8495
rect 17879 8410 17880 8474
rect 17944 8410 17960 8474
rect 18024 8410 18040 8474
rect 18104 8410 18120 8474
rect 18184 8410 18185 8474
rect 17879 8388 18185 8410
rect 1594 8323 2140 8324
rect 17879 8324 17880 8388
rect 17944 8324 17960 8388
rect 18024 8324 18040 8388
rect 18104 8324 18120 8388
rect 18184 8324 18185 8388
rect 17879 8323 18185 8324
rect 20129 9239 20515 9240
rect 20129 9175 20130 9239
rect 20194 9175 20210 9239
rect 20274 9175 20290 9239
rect 20354 9175 20370 9239
rect 20434 9175 20450 9239
rect 20514 9175 20515 9239
rect 20129 9154 20515 9175
rect 20129 9090 20130 9154
rect 20194 9090 20210 9154
rect 20274 9090 20290 9154
rect 20354 9090 20370 9154
rect 20434 9090 20450 9154
rect 20514 9090 20515 9154
rect 20129 9069 20515 9090
rect 20129 9005 20130 9069
rect 20194 9005 20210 9069
rect 20274 9005 20290 9069
rect 20354 9005 20370 9069
rect 20434 9005 20450 9069
rect 20514 9005 20515 9069
rect 20129 8984 20515 9005
rect 20129 8920 20130 8984
rect 20194 8920 20210 8984
rect 20274 8920 20290 8984
rect 20354 8920 20370 8984
rect 20434 8920 20450 8984
rect 20514 8920 20515 8984
rect 20129 8899 20515 8920
rect 20129 8835 20130 8899
rect 20194 8835 20210 8899
rect 20274 8835 20290 8899
rect 20354 8835 20370 8899
rect 20434 8835 20450 8899
rect 20514 8835 20515 8899
rect 20129 8814 20515 8835
rect 20129 8750 20130 8814
rect 20194 8750 20210 8814
rect 20274 8750 20290 8814
rect 20354 8750 20370 8814
rect 20434 8750 20450 8814
rect 20514 8750 20515 8814
rect 20129 8729 20515 8750
rect 20129 8665 20130 8729
rect 20194 8665 20210 8729
rect 20274 8665 20290 8729
rect 20354 8665 20370 8729
rect 20434 8665 20450 8729
rect 20514 8665 20515 8729
rect 20129 8644 20515 8665
rect 20129 8580 20130 8644
rect 20194 8580 20210 8644
rect 20274 8580 20290 8644
rect 20354 8580 20370 8644
rect 20434 8580 20450 8644
rect 20514 8580 20515 8644
rect 20129 8559 20515 8580
rect 20129 8495 20130 8559
rect 20194 8495 20210 8559
rect 20274 8495 20290 8559
rect 20354 8495 20370 8559
rect 20434 8495 20450 8559
rect 20514 8495 20515 8559
rect 20129 8474 20515 8495
rect 20129 8410 20130 8474
rect 20194 8410 20210 8474
rect 20274 8410 20290 8474
rect 20354 8410 20370 8474
rect 20434 8410 20450 8474
rect 20514 8410 20515 8474
rect 20129 8388 20515 8410
rect 20129 8324 20130 8388
rect 20194 8324 20210 8388
rect 20274 8324 20290 8388
rect 20354 8324 20370 8388
rect 20434 8324 20450 8388
rect 20514 8324 20515 8388
rect 20129 8323 20515 8324
rect 27746 8317 28000 9247
rect 0 7347 254 8037
rect 851 8031 1084 8037
rect 851 7967 852 8031
rect 916 7967 936 8031
rect 1000 7967 1020 8031
rect 23783 8023 24167 8024
rect 851 7944 1084 7967
rect 851 7880 852 7944
rect 916 7880 936 7944
rect 1000 7880 1020 7944
rect 851 7857 1084 7880
rect 851 7793 852 7857
rect 916 7793 936 7857
rect 1000 7793 1020 7857
rect 851 7769 1084 7793
rect 851 7705 852 7769
rect 916 7705 936 7769
rect 1000 7705 1020 7769
rect 851 7681 1084 7705
rect 851 7617 852 7681
rect 916 7617 936 7681
rect 1000 7617 1020 7681
rect 851 7593 1084 7617
rect 851 7529 852 7593
rect 916 7529 936 7593
rect 1000 7529 1020 7593
rect 851 7505 1084 7529
rect 851 7441 852 7505
rect 916 7441 936 7505
rect 1000 7441 1020 7505
rect 851 7417 1084 7441
rect 851 7353 852 7417
rect 916 7353 936 7417
rect 1000 7353 1020 7417
rect 3312 8021 3696 8022
rect 3312 7957 3313 8021
rect 3377 7957 3419 8021
rect 3483 7957 3525 8021
rect 3589 7957 3631 8021
rect 3695 7957 3696 8021
rect 3312 7937 3696 7957
rect 3312 7873 3313 7937
rect 3377 7873 3419 7937
rect 3483 7873 3525 7937
rect 3589 7873 3631 7937
rect 3695 7873 3696 7937
rect 3312 7852 3696 7873
rect 3312 7788 3313 7852
rect 3377 7788 3419 7852
rect 3483 7788 3525 7852
rect 3589 7788 3631 7852
rect 3695 7788 3696 7852
rect 3312 7767 3696 7788
rect 3312 7703 3313 7767
rect 3377 7703 3419 7767
rect 3483 7703 3525 7767
rect 3589 7703 3631 7767
rect 3695 7703 3696 7767
rect 3312 7682 3696 7703
rect 3312 7618 3313 7682
rect 3377 7618 3419 7682
rect 3483 7618 3525 7682
rect 3589 7618 3631 7682
rect 3695 7618 3696 7682
rect 3312 7597 3696 7618
rect 3312 7533 3313 7597
rect 3377 7533 3419 7597
rect 3483 7533 3525 7597
rect 3589 7533 3631 7597
rect 3695 7533 3696 7597
rect 3312 7512 3696 7533
rect 3312 7448 3313 7512
rect 3377 7448 3419 7512
rect 3483 7448 3525 7512
rect 3589 7448 3631 7512
rect 3695 7448 3696 7512
rect 23783 7959 23784 8023
rect 23848 7959 23890 8023
rect 23954 7959 23996 8023
rect 24060 7959 24102 8023
rect 24166 7959 24167 8023
rect 23783 7939 24167 7959
rect 23783 7875 23784 7939
rect 23848 7875 23890 7939
rect 23954 7875 23996 7939
rect 24060 7875 24102 7939
rect 24166 7875 24167 7939
rect 23783 7854 24167 7875
rect 23783 7790 23784 7854
rect 23848 7790 23890 7854
rect 23954 7790 23996 7854
rect 24060 7790 24102 7854
rect 24166 7790 24167 7854
rect 23783 7769 24167 7790
rect 23783 7705 23784 7769
rect 23848 7705 23890 7769
rect 23954 7705 23996 7769
rect 24060 7705 24102 7769
rect 24166 7705 24167 7769
rect 23783 7684 24167 7705
rect 23783 7620 23784 7684
rect 23848 7620 23890 7684
rect 23954 7620 23996 7684
rect 24060 7620 24102 7684
rect 24166 7620 24167 7684
rect 23783 7599 24167 7620
rect 23783 7535 23784 7599
rect 23848 7535 23890 7599
rect 23954 7535 23996 7599
rect 24060 7535 24102 7599
rect 24166 7535 24167 7599
rect 23783 7514 24167 7535
rect 23783 7450 23784 7514
rect 23848 7450 23890 7514
rect 23954 7450 23996 7514
rect 24060 7450 24102 7514
rect 24166 7450 24167 7514
rect 23783 7449 24167 7450
rect 3312 7427 3696 7448
rect 3312 7363 3313 7427
rect 3377 7363 3419 7427
rect 3483 7363 3525 7427
rect 3589 7363 3631 7427
rect 3695 7363 3696 7427
rect 3312 7362 3696 7363
rect 851 7347 1084 7353
rect 27746 7347 28000 8037
rect 0 6377 254 7067
rect 21868 7055 22306 7056
rect 21868 6991 21871 7055
rect 21935 6991 21963 7055
rect 22027 6991 22055 7055
rect 22119 6991 22147 7055
rect 22211 6991 22239 7055
rect 22303 6991 22306 7055
rect 21868 6969 22306 6991
rect 21868 6905 21871 6969
rect 21935 6905 21963 6969
rect 22027 6905 22055 6969
rect 22119 6905 22147 6969
rect 22211 6905 22239 6969
rect 22303 6905 22306 6969
rect 21868 6883 22306 6905
rect 21868 6819 21871 6883
rect 21935 6819 21963 6883
rect 22027 6819 22055 6883
rect 22119 6819 22147 6883
rect 22211 6819 22239 6883
rect 22303 6819 22306 6883
rect 21868 6797 22306 6819
rect 21868 6733 21871 6797
rect 21935 6733 21963 6797
rect 22027 6733 22055 6797
rect 22119 6733 22147 6797
rect 22211 6733 22239 6797
rect 22303 6733 22306 6797
rect 21868 6711 22306 6733
rect 21868 6647 21871 6711
rect 21935 6647 21963 6711
rect 22027 6647 22055 6711
rect 22119 6647 22147 6711
rect 22211 6647 22239 6711
rect 22303 6647 22306 6711
rect 21868 6625 22306 6647
rect 21868 6561 21871 6625
rect 21935 6561 21963 6625
rect 22027 6561 22055 6625
rect 22119 6561 22147 6625
rect 22211 6561 22239 6625
rect 22303 6561 22306 6625
rect 21868 6538 22306 6561
rect 21868 6474 21871 6538
rect 21935 6474 21963 6538
rect 22027 6474 22055 6538
rect 22119 6474 22147 6538
rect 22211 6474 22239 6538
rect 22303 6474 22306 6538
rect 21868 6451 22306 6474
rect 21868 6387 21871 6451
rect 21935 6387 21963 6451
rect 22027 6387 22055 6451
rect 22119 6387 22147 6451
rect 22211 6387 22239 6451
rect 22303 6387 22306 6451
rect 21868 6386 22306 6387
rect 27746 6377 28000 7067
rect 0 5167 254 6097
rect 27746 5167 28000 6097
rect 1538 5058 2320 5059
rect 1538 4994 1539 5058
rect 1603 4994 1619 5058
rect 1683 4994 2175 5058
rect 2239 4994 2255 5058
rect 2319 4994 2320 5058
rect 1538 4993 2320 4994
rect 0 3957 254 4887
rect 27746 3957 28000 4887
rect 0 2987 193 3677
rect 1921 3639 2053 3677
rect 1921 3575 1955 3639
rect 2019 3575 2053 3639
rect 1921 3556 2053 3575
rect 1921 3492 1955 3556
rect 2019 3492 2053 3556
rect 1921 3473 2053 3492
rect 1921 3409 1955 3473
rect 2019 3409 2053 3473
rect 1921 3390 2053 3409
rect 1921 3326 1955 3390
rect 2019 3326 2053 3390
rect 1921 3307 2053 3326
rect 1921 3243 1955 3307
rect 2019 3243 2053 3307
rect 1921 3224 2053 3243
rect 1921 3160 1955 3224
rect 2019 3160 2053 3224
rect 1921 3141 2053 3160
rect 1921 3077 1955 3141
rect 2019 3077 2053 3141
rect 1921 3057 2053 3077
rect 1921 2993 1955 3057
rect 2019 2993 2053 3057
rect 9767 3664 10073 3665
rect 9767 3600 9768 3664
rect 9832 3600 9848 3664
rect 9912 3600 9928 3664
rect 9992 3600 10008 3664
rect 10072 3600 10073 3664
rect 9767 3579 10073 3600
rect 9767 3515 9768 3579
rect 9832 3515 9848 3579
rect 9912 3515 9928 3579
rect 9992 3515 10008 3579
rect 10072 3515 10073 3579
rect 9767 3494 10073 3515
rect 9767 3430 9768 3494
rect 9832 3430 9848 3494
rect 9912 3430 9928 3494
rect 9992 3430 10008 3494
rect 10072 3430 10073 3494
rect 9767 3409 10073 3430
rect 9767 3345 9768 3409
rect 9832 3345 9848 3409
rect 9912 3345 9928 3409
rect 9992 3345 10008 3409
rect 10072 3345 10073 3409
rect 9767 3323 10073 3345
rect 9767 3259 9768 3323
rect 9832 3259 9848 3323
rect 9912 3259 9928 3323
rect 9992 3259 10008 3323
rect 10072 3259 10073 3323
rect 9767 3237 10073 3259
rect 9767 3173 9768 3237
rect 9832 3173 9848 3237
rect 9912 3173 9928 3237
rect 9992 3173 10008 3237
rect 10072 3173 10073 3237
rect 9767 3151 10073 3173
rect 9767 3087 9768 3151
rect 9832 3087 9848 3151
rect 9912 3087 9928 3151
rect 9992 3087 10008 3151
rect 10072 3087 10073 3151
rect 9767 3065 10073 3087
rect 9767 3001 9768 3065
rect 9832 3001 9848 3065
rect 9912 3001 9928 3065
rect 9992 3001 10008 3065
rect 10072 3001 10073 3065
rect 9767 3000 10073 3001
rect 1921 2987 2053 2993
rect 27807 2987 28000 3677
rect 1591 2878 2320 2879
rect 1591 2814 1592 2878
rect 1656 2814 1672 2878
rect 1736 2814 2175 2878
rect 2239 2814 2255 2878
rect 2319 2814 2320 2878
rect 1591 2813 2320 2814
rect 5094 2875 5531 2876
rect 5094 2811 5095 2875
rect 5159 2811 5175 2875
rect 5239 2811 5386 2875
rect 5450 2811 5466 2875
rect 5530 2811 5531 2875
rect 5094 2810 5531 2811
rect 0 1777 254 2707
rect 5940 2701 6540 2707
rect 5940 2637 5944 2701
rect 6008 2637 6032 2701
rect 6096 2637 6120 2701
rect 6184 2637 6208 2701
rect 6272 2637 6296 2701
rect 6360 2637 6384 2701
rect 6448 2637 6472 2701
rect 6536 2637 6540 2701
rect 5940 2616 6540 2637
rect 5940 2552 5944 2616
rect 6008 2552 6032 2616
rect 6096 2552 6120 2616
rect 6184 2552 6208 2616
rect 6272 2552 6296 2616
rect 6360 2552 6384 2616
rect 6448 2552 6472 2616
rect 6536 2552 6540 2616
rect 5940 2531 6540 2552
rect 5940 2467 5944 2531
rect 6008 2467 6032 2531
rect 6096 2467 6120 2531
rect 6184 2467 6208 2531
rect 6272 2467 6296 2531
rect 6360 2467 6384 2531
rect 6448 2467 6472 2531
rect 6536 2467 6540 2531
rect 5940 2446 6540 2467
rect 5940 2382 5944 2446
rect 6008 2382 6032 2446
rect 6096 2382 6120 2446
rect 6184 2382 6208 2446
rect 6272 2382 6296 2446
rect 6360 2382 6384 2446
rect 6448 2382 6472 2446
rect 6536 2382 6540 2446
rect 5940 2361 6540 2382
rect 5940 2297 5944 2361
rect 6008 2297 6032 2361
rect 6096 2297 6120 2361
rect 6184 2297 6208 2361
rect 6272 2297 6296 2361
rect 6360 2297 6384 2361
rect 6448 2297 6472 2361
rect 6536 2297 6540 2361
rect 5940 2276 6540 2297
rect 5940 2212 5944 2276
rect 6008 2212 6032 2276
rect 6096 2212 6120 2276
rect 6184 2212 6208 2276
rect 6272 2212 6296 2276
rect 6360 2212 6384 2276
rect 6448 2212 6472 2276
rect 6536 2212 6540 2276
rect 5940 2191 6540 2212
rect 5940 2127 5944 2191
rect 6008 2127 6032 2191
rect 6096 2127 6120 2191
rect 6184 2127 6208 2191
rect 6272 2127 6296 2191
rect 6360 2127 6384 2191
rect 6448 2127 6472 2191
rect 6536 2127 6540 2191
rect 5940 2105 6540 2127
rect 5940 2041 5944 2105
rect 6008 2041 6032 2105
rect 6096 2041 6120 2105
rect 6184 2041 6208 2105
rect 6272 2041 6296 2105
rect 6360 2041 6384 2105
rect 6448 2041 6472 2105
rect 6536 2041 6540 2105
rect 5940 2019 6540 2041
rect 5940 1955 5944 2019
rect 6008 1955 6032 2019
rect 6096 1955 6120 2019
rect 6184 1955 6208 2019
rect 6272 1955 6296 2019
rect 6360 1955 6384 2019
rect 6448 1955 6472 2019
rect 6536 1955 6540 2019
rect 5940 1933 6540 1955
rect 5940 1869 5944 1933
rect 6008 1869 6032 1933
rect 6096 1869 6120 1933
rect 6184 1869 6208 1933
rect 6272 1869 6296 1933
rect 6360 1869 6384 1933
rect 6448 1869 6472 1933
rect 6536 1869 6540 1933
rect 5940 1847 6540 1869
rect 5940 1783 5944 1847
rect 6008 1783 6032 1847
rect 6096 1783 6120 1847
rect 6184 1783 6208 1847
rect 6272 1783 6296 1847
rect 6360 1783 6384 1847
rect 6448 1783 6472 1847
rect 6536 1783 6540 1847
rect 5940 1777 6540 1783
rect 12225 2701 12825 2707
rect 12225 2637 12229 2701
rect 12293 2637 12317 2701
rect 12381 2637 12405 2701
rect 12469 2637 12493 2701
rect 12557 2637 12581 2701
rect 12645 2637 12669 2701
rect 12733 2637 12757 2701
rect 12821 2637 12825 2701
rect 12225 2616 12825 2637
rect 12225 2552 12229 2616
rect 12293 2552 12317 2616
rect 12381 2552 12405 2616
rect 12469 2552 12493 2616
rect 12557 2552 12581 2616
rect 12645 2552 12669 2616
rect 12733 2552 12757 2616
rect 12821 2552 12825 2616
rect 12225 2531 12825 2552
rect 12225 2467 12229 2531
rect 12293 2467 12317 2531
rect 12381 2467 12405 2531
rect 12469 2467 12493 2531
rect 12557 2467 12581 2531
rect 12645 2467 12669 2531
rect 12733 2467 12757 2531
rect 12821 2467 12825 2531
rect 12225 2446 12825 2467
rect 12225 2382 12229 2446
rect 12293 2382 12317 2446
rect 12381 2382 12405 2446
rect 12469 2382 12493 2446
rect 12557 2382 12581 2446
rect 12645 2382 12669 2446
rect 12733 2382 12757 2446
rect 12821 2382 12825 2446
rect 12225 2361 12825 2382
rect 12225 2297 12229 2361
rect 12293 2297 12317 2361
rect 12381 2297 12405 2361
rect 12469 2297 12493 2361
rect 12557 2297 12581 2361
rect 12645 2297 12669 2361
rect 12733 2297 12757 2361
rect 12821 2297 12825 2361
rect 12225 2276 12825 2297
rect 12225 2212 12229 2276
rect 12293 2212 12317 2276
rect 12381 2212 12405 2276
rect 12469 2212 12493 2276
rect 12557 2212 12581 2276
rect 12645 2212 12669 2276
rect 12733 2212 12757 2276
rect 12821 2212 12825 2276
rect 12225 2191 12825 2212
rect 12225 2127 12229 2191
rect 12293 2127 12317 2191
rect 12381 2127 12405 2191
rect 12469 2127 12493 2191
rect 12557 2127 12581 2191
rect 12645 2127 12669 2191
rect 12733 2127 12757 2191
rect 12821 2127 12825 2191
rect 12225 2105 12825 2127
rect 12225 2041 12229 2105
rect 12293 2041 12317 2105
rect 12381 2041 12405 2105
rect 12469 2041 12493 2105
rect 12557 2041 12581 2105
rect 12645 2041 12669 2105
rect 12733 2041 12757 2105
rect 12821 2041 12825 2105
rect 12225 2019 12825 2041
rect 12225 1955 12229 2019
rect 12293 1955 12317 2019
rect 12381 1955 12405 2019
rect 12469 1955 12493 2019
rect 12557 1955 12581 2019
rect 12645 1955 12669 2019
rect 12733 1955 12757 2019
rect 12821 1955 12825 2019
rect 12225 1933 12825 1955
rect 12225 1869 12229 1933
rect 12293 1869 12317 1933
rect 12381 1869 12405 1933
rect 12469 1869 12493 1933
rect 12557 1869 12581 1933
rect 12645 1869 12669 1933
rect 12733 1869 12757 1933
rect 12821 1869 12825 1933
rect 12225 1847 12825 1869
rect 12225 1783 12229 1847
rect 12293 1783 12317 1847
rect 12381 1783 12405 1847
rect 12469 1783 12493 1847
rect 12557 1783 12581 1847
rect 12645 1783 12669 1847
rect 12733 1783 12757 1847
rect 12821 1783 12825 1847
rect 12225 1777 12825 1783
rect 16057 2701 16657 2707
rect 16057 2637 16061 2701
rect 16125 2637 16149 2701
rect 16213 2637 16237 2701
rect 16301 2637 16325 2701
rect 16389 2637 16413 2701
rect 16477 2637 16501 2701
rect 16565 2637 16589 2701
rect 16653 2637 16657 2701
rect 16057 2616 16657 2637
rect 16057 2552 16061 2616
rect 16125 2552 16149 2616
rect 16213 2552 16237 2616
rect 16301 2552 16325 2616
rect 16389 2552 16413 2616
rect 16477 2552 16501 2616
rect 16565 2552 16589 2616
rect 16653 2552 16657 2616
rect 16057 2531 16657 2552
rect 16057 2467 16061 2531
rect 16125 2467 16149 2531
rect 16213 2467 16237 2531
rect 16301 2467 16325 2531
rect 16389 2467 16413 2531
rect 16477 2467 16501 2531
rect 16565 2467 16589 2531
rect 16653 2467 16657 2531
rect 16057 2446 16657 2467
rect 16057 2382 16061 2446
rect 16125 2382 16149 2446
rect 16213 2382 16237 2446
rect 16301 2382 16325 2446
rect 16389 2382 16413 2446
rect 16477 2382 16501 2446
rect 16565 2382 16589 2446
rect 16653 2382 16657 2446
rect 16057 2361 16657 2382
rect 16057 2297 16061 2361
rect 16125 2297 16149 2361
rect 16213 2297 16237 2361
rect 16301 2297 16325 2361
rect 16389 2297 16413 2361
rect 16477 2297 16501 2361
rect 16565 2297 16589 2361
rect 16653 2297 16657 2361
rect 16057 2276 16657 2297
rect 16057 2212 16061 2276
rect 16125 2212 16149 2276
rect 16213 2212 16237 2276
rect 16301 2212 16325 2276
rect 16389 2212 16413 2276
rect 16477 2212 16501 2276
rect 16565 2212 16589 2276
rect 16653 2212 16657 2276
rect 16057 2191 16657 2212
rect 16057 2127 16061 2191
rect 16125 2127 16149 2191
rect 16213 2127 16237 2191
rect 16301 2127 16325 2191
rect 16389 2127 16413 2191
rect 16477 2127 16501 2191
rect 16565 2127 16589 2191
rect 16653 2127 16657 2191
rect 16057 2105 16657 2127
rect 16057 2041 16061 2105
rect 16125 2041 16149 2105
rect 16213 2041 16237 2105
rect 16301 2041 16325 2105
rect 16389 2041 16413 2105
rect 16477 2041 16501 2105
rect 16565 2041 16589 2105
rect 16653 2041 16657 2105
rect 16057 2019 16657 2041
rect 16057 1955 16061 2019
rect 16125 1955 16149 2019
rect 16213 1955 16237 2019
rect 16301 1955 16325 2019
rect 16389 1955 16413 2019
rect 16477 1955 16501 2019
rect 16565 1955 16589 2019
rect 16653 1955 16657 2019
rect 16057 1933 16657 1955
rect 16057 1869 16061 1933
rect 16125 1869 16149 1933
rect 16213 1869 16237 1933
rect 16301 1869 16325 1933
rect 16389 1869 16413 1933
rect 16477 1869 16501 1933
rect 16565 1869 16589 1933
rect 16653 1869 16657 1933
rect 16057 1847 16657 1869
rect 16057 1783 16061 1847
rect 16125 1783 16149 1847
rect 16213 1783 16237 1847
rect 16301 1783 16325 1847
rect 16389 1783 16413 1847
rect 16477 1783 16501 1847
rect 16565 1783 16589 1847
rect 16653 1783 16657 1847
rect 16057 1777 16657 1783
rect 20292 2701 20892 2707
rect 20292 2637 20296 2701
rect 20360 2637 20384 2701
rect 20448 2637 20472 2701
rect 20536 2637 20560 2701
rect 20624 2637 20648 2701
rect 20712 2637 20736 2701
rect 20800 2637 20824 2701
rect 20888 2637 20892 2701
rect 27746 2693 28000 2707
rect 20292 2616 20892 2637
rect 20292 2552 20296 2616
rect 20360 2552 20384 2616
rect 20448 2552 20472 2616
rect 20536 2552 20560 2616
rect 20624 2552 20648 2616
rect 20712 2552 20736 2616
rect 20800 2552 20824 2616
rect 20888 2552 20892 2616
rect 20292 2531 20892 2552
rect 20292 2467 20296 2531
rect 20360 2467 20384 2531
rect 20448 2467 20472 2531
rect 20536 2467 20560 2531
rect 20624 2467 20648 2531
rect 20712 2467 20736 2531
rect 20800 2467 20824 2531
rect 20888 2467 20892 2531
rect 20292 2446 20892 2467
rect 20292 2382 20296 2446
rect 20360 2382 20384 2446
rect 20448 2382 20472 2446
rect 20536 2382 20560 2446
rect 20624 2382 20648 2446
rect 20712 2382 20736 2446
rect 20800 2382 20824 2446
rect 20888 2382 20892 2446
rect 20292 2361 20892 2382
rect 20292 2297 20296 2361
rect 20360 2297 20384 2361
rect 20448 2297 20472 2361
rect 20536 2297 20560 2361
rect 20624 2297 20648 2361
rect 20712 2297 20736 2361
rect 20800 2297 20824 2361
rect 20888 2297 20892 2361
rect 20292 2276 20892 2297
rect 20292 2212 20296 2276
rect 20360 2212 20384 2276
rect 20448 2212 20472 2276
rect 20536 2212 20560 2276
rect 20624 2212 20648 2276
rect 20712 2212 20736 2276
rect 20800 2212 20824 2276
rect 20888 2212 20892 2276
rect 20292 2191 20892 2212
rect 20292 2127 20296 2191
rect 20360 2127 20384 2191
rect 20448 2127 20472 2191
rect 20536 2127 20560 2191
rect 20624 2127 20648 2191
rect 20712 2127 20736 2191
rect 20800 2127 20824 2191
rect 20888 2127 20892 2191
rect 20292 2105 20892 2127
rect 20292 2041 20296 2105
rect 20360 2041 20384 2105
rect 20448 2041 20472 2105
rect 20536 2041 20560 2105
rect 20624 2041 20648 2105
rect 20712 2041 20736 2105
rect 20800 2041 20824 2105
rect 20888 2041 20892 2105
rect 20292 2019 20892 2041
rect 20292 1955 20296 2019
rect 20360 1955 20384 2019
rect 20448 1955 20472 2019
rect 20536 1955 20560 2019
rect 20624 1955 20648 2019
rect 20712 1955 20736 2019
rect 20800 1955 20824 2019
rect 20888 1955 20892 2019
rect 20292 1933 20892 1955
rect 20292 1869 20296 1933
rect 20360 1869 20384 1933
rect 20448 1869 20472 1933
rect 20536 1869 20560 1933
rect 20624 1869 20648 1933
rect 20712 1869 20736 1933
rect 20800 1869 20824 1933
rect 20888 1869 20892 1933
rect 20292 1847 20892 1869
rect 20292 1783 20296 1847
rect 20360 1783 20384 1847
rect 20448 1783 20472 1847
rect 20536 1783 20560 1847
rect 20624 1783 20648 1847
rect 20712 1783 20736 1847
rect 20800 1783 20824 1847
rect 20888 1783 20892 1847
rect 27651 2692 28000 2693
rect 27651 2628 27653 2692
rect 27717 2628 27743 2692
rect 27807 2628 27833 2692
rect 27897 2628 27923 2692
rect 27987 2628 28000 2692
rect 27651 2608 28000 2628
rect 27651 2544 27653 2608
rect 27717 2544 27743 2608
rect 27807 2544 27833 2608
rect 27897 2544 27923 2608
rect 27987 2544 28000 2608
rect 27651 2524 28000 2544
rect 27651 2460 27653 2524
rect 27717 2460 27743 2524
rect 27807 2460 27833 2524
rect 27897 2460 27923 2524
rect 27987 2460 28000 2524
rect 27651 2440 28000 2460
rect 27651 2376 27653 2440
rect 27717 2376 27743 2440
rect 27807 2376 27833 2440
rect 27897 2376 27923 2440
rect 27987 2376 28000 2440
rect 27651 2356 28000 2376
rect 27651 2292 27653 2356
rect 27717 2292 27743 2356
rect 27807 2292 27833 2356
rect 27897 2292 27923 2356
rect 27987 2292 28000 2356
rect 27651 2272 28000 2292
rect 27651 2208 27653 2272
rect 27717 2208 27743 2272
rect 27807 2208 27833 2272
rect 27897 2208 27923 2272
rect 27987 2208 28000 2272
rect 27651 2188 28000 2208
rect 27651 2124 27653 2188
rect 27717 2124 27743 2188
rect 27807 2124 27833 2188
rect 27897 2124 27923 2188
rect 27987 2124 28000 2188
rect 27651 2104 28000 2124
rect 27651 2040 27653 2104
rect 27717 2040 27743 2104
rect 27807 2040 27833 2104
rect 27897 2040 27923 2104
rect 27987 2040 28000 2104
rect 27651 2020 28000 2040
rect 27651 1956 27653 2020
rect 27717 1956 27743 2020
rect 27807 1956 27833 2020
rect 27897 1956 27923 2020
rect 27987 1956 28000 2020
rect 27651 1936 28000 1956
rect 27651 1872 27653 1936
rect 27717 1872 27743 1936
rect 27807 1872 27833 1936
rect 27897 1872 27923 1936
rect 27987 1872 28000 1936
rect 27651 1851 28000 1872
rect 27651 1787 27653 1851
rect 27717 1787 27743 1851
rect 27807 1787 27833 1851
rect 27897 1787 27923 1851
rect 27987 1787 28000 1851
rect 27651 1786 28000 1787
rect 20292 1777 20892 1783
rect 27746 1777 28000 1786
rect 8695 1676 9132 1677
rect 8695 1612 8696 1676
rect 8760 1612 8776 1676
rect 8840 1612 8987 1676
rect 9051 1612 9067 1676
rect 9131 1612 9132 1676
rect 8695 1611 9132 1612
rect 10336 1676 10773 1677
rect 10336 1612 10337 1676
rect 10401 1612 10417 1676
rect 10481 1612 10628 1676
rect 10692 1612 10708 1676
rect 10772 1612 10773 1676
rect 10336 1611 10773 1612
rect 21133 1676 21570 1677
rect 21133 1612 21134 1676
rect 21198 1612 21214 1676
rect 21278 1612 21425 1676
rect 21489 1612 21505 1676
rect 21569 1612 21570 1676
rect 21133 1611 21570 1612
rect 24513 1676 24950 1677
rect 24513 1612 24514 1676
rect 24578 1612 24594 1676
rect 24658 1612 24805 1676
rect 24869 1612 24885 1676
rect 24949 1612 24950 1676
rect 24513 1611 24950 1612
rect 0 407 254 1497
rect 3337 1491 3847 1497
rect 3337 1427 3340 1491
rect 3404 1427 3428 1491
rect 3492 1427 3516 1491
rect 3580 1427 3604 1491
rect 3668 1427 3692 1491
rect 3756 1427 3780 1491
rect 3844 1427 3847 1491
rect 3337 1407 3847 1427
rect 3337 1343 3340 1407
rect 3404 1343 3428 1407
rect 3492 1343 3516 1407
rect 3580 1343 3604 1407
rect 3668 1343 3692 1407
rect 3756 1343 3780 1407
rect 3844 1343 3847 1407
rect 3337 1323 3847 1343
rect 3337 1259 3340 1323
rect 3404 1259 3428 1323
rect 3492 1259 3516 1323
rect 3580 1259 3604 1323
rect 3668 1259 3692 1323
rect 3756 1259 3780 1323
rect 3844 1259 3847 1323
rect 3337 1239 3847 1259
rect 3337 1175 3340 1239
rect 3404 1175 3428 1239
rect 3492 1175 3516 1239
rect 3580 1175 3604 1239
rect 3668 1175 3692 1239
rect 3756 1175 3780 1239
rect 3844 1175 3847 1239
rect 3337 1155 3847 1175
rect 3337 1091 3340 1155
rect 3404 1091 3428 1155
rect 3492 1091 3516 1155
rect 3580 1091 3604 1155
rect 3668 1091 3692 1155
rect 3756 1091 3780 1155
rect 3844 1091 3847 1155
rect 3337 1071 3847 1091
rect 3337 1007 3340 1071
rect 3404 1007 3428 1071
rect 3492 1007 3516 1071
rect 3580 1007 3604 1071
rect 3668 1007 3692 1071
rect 3756 1007 3780 1071
rect 3844 1007 3847 1071
rect 3337 987 3847 1007
rect 3337 923 3340 987
rect 3404 923 3428 987
rect 3492 923 3516 987
rect 3580 923 3604 987
rect 3668 923 3692 987
rect 3756 923 3780 987
rect 3844 923 3847 987
rect 3337 902 3847 923
rect 3337 838 3340 902
rect 3404 838 3428 902
rect 3492 838 3516 902
rect 3580 838 3604 902
rect 3668 838 3692 902
rect 3756 838 3780 902
rect 3844 838 3847 902
rect 3337 817 3847 838
rect 3337 753 3340 817
rect 3404 753 3428 817
rect 3492 753 3516 817
rect 3580 753 3604 817
rect 3668 753 3692 817
rect 3756 753 3780 817
rect 3844 753 3847 817
rect 3337 732 3847 753
rect 3337 668 3340 732
rect 3404 668 3428 732
rect 3492 668 3516 732
rect 3580 668 3604 732
rect 3668 668 3692 732
rect 3756 668 3780 732
rect 3844 668 3847 732
rect 3337 647 3847 668
rect 3337 583 3340 647
rect 3404 583 3428 647
rect 3492 583 3516 647
rect 3580 583 3604 647
rect 3668 583 3692 647
rect 3756 583 3780 647
rect 3844 583 3847 647
rect 3337 562 3847 583
rect 3337 498 3340 562
rect 3404 498 3428 562
rect 3492 498 3516 562
rect 3580 498 3604 562
rect 3668 498 3692 562
rect 3756 498 3780 562
rect 3844 498 3847 562
rect 3337 477 3847 498
rect 3337 413 3340 477
rect 3404 413 3428 477
rect 3492 413 3516 477
rect 3580 413 3604 477
rect 3668 413 3692 477
rect 3756 413 3780 477
rect 3844 413 3847 477
rect 3337 407 3847 413
rect 17775 1491 18175 1497
rect 17839 1427 17859 1491
rect 17923 1427 17943 1491
rect 18007 1427 18027 1491
rect 18091 1427 18111 1491
rect 17775 1407 18175 1427
rect 17839 1343 17859 1407
rect 17923 1343 17943 1407
rect 18007 1343 18027 1407
rect 18091 1343 18111 1407
rect 17775 1323 18175 1343
rect 17839 1259 17859 1323
rect 17923 1259 17943 1323
rect 18007 1259 18027 1323
rect 18091 1259 18111 1323
rect 17775 1239 18175 1259
rect 17839 1175 17859 1239
rect 17923 1175 17943 1239
rect 18007 1175 18027 1239
rect 18091 1175 18111 1239
rect 17775 1155 18175 1175
rect 17839 1091 17859 1155
rect 17923 1091 17943 1155
rect 18007 1091 18027 1155
rect 18091 1091 18111 1155
rect 17775 1071 18175 1091
rect 17839 1007 17859 1071
rect 17923 1007 17943 1071
rect 18007 1007 18027 1071
rect 18091 1007 18111 1071
rect 17775 987 18175 1007
rect 17839 923 17859 987
rect 17923 923 17943 987
rect 18007 923 18027 987
rect 18091 923 18111 987
rect 17775 902 18175 923
rect 17839 838 17859 902
rect 17923 838 17943 902
rect 18007 838 18027 902
rect 18091 838 18111 902
rect 17775 817 18175 838
rect 17839 753 17859 817
rect 17923 753 17943 817
rect 18007 753 18027 817
rect 18091 753 18111 817
rect 17775 732 18175 753
rect 17839 668 17859 732
rect 17923 668 17943 732
rect 18007 668 18027 732
rect 18091 668 18111 732
rect 17775 647 18175 668
rect 17839 583 17859 647
rect 17923 583 17943 647
rect 18007 583 18027 647
rect 18091 583 18111 647
rect 17775 562 18175 583
rect 17839 498 17859 562
rect 17923 498 17943 562
rect 18007 498 18027 562
rect 18091 498 18111 562
rect 17775 477 18175 498
rect 17839 413 17859 477
rect 17923 413 17943 477
rect 18007 413 18027 477
rect 18091 413 18111 477
rect 22275 1488 22939 1489
rect 22275 1424 22281 1488
rect 22345 1424 22365 1488
rect 22429 1424 22449 1488
rect 22513 1424 22533 1488
rect 22597 1424 22617 1488
rect 22681 1424 22701 1488
rect 22765 1424 22785 1488
rect 22849 1424 22869 1488
rect 22933 1424 22939 1488
rect 22275 1405 22939 1424
rect 22275 1341 22281 1405
rect 22345 1341 22365 1405
rect 22429 1341 22449 1405
rect 22513 1341 22533 1405
rect 22597 1341 22617 1405
rect 22681 1341 22701 1405
rect 22765 1341 22785 1405
rect 22849 1341 22869 1405
rect 22933 1341 22939 1405
rect 22275 1322 22939 1341
rect 22275 1258 22281 1322
rect 22345 1258 22365 1322
rect 22429 1258 22449 1322
rect 22513 1258 22533 1322
rect 22597 1258 22617 1322
rect 22681 1258 22701 1322
rect 22765 1258 22785 1322
rect 22849 1258 22869 1322
rect 22933 1258 22939 1322
rect 22275 1238 22939 1258
rect 22275 1174 22281 1238
rect 22345 1174 22365 1238
rect 22429 1174 22449 1238
rect 22513 1174 22533 1238
rect 22597 1174 22617 1238
rect 22681 1174 22701 1238
rect 22765 1174 22785 1238
rect 22849 1174 22869 1238
rect 22933 1174 22939 1238
rect 22275 1154 22939 1174
rect 22275 1090 22281 1154
rect 22345 1090 22365 1154
rect 22429 1090 22449 1154
rect 22513 1090 22533 1154
rect 22597 1090 22617 1154
rect 22681 1090 22701 1154
rect 22765 1090 22785 1154
rect 22849 1090 22869 1154
rect 22933 1090 22939 1154
rect 22275 1070 22939 1090
rect 22275 1006 22281 1070
rect 22345 1006 22365 1070
rect 22429 1006 22449 1070
rect 22513 1006 22533 1070
rect 22597 1006 22617 1070
rect 22681 1006 22701 1070
rect 22765 1006 22785 1070
rect 22849 1006 22869 1070
rect 22933 1006 22939 1070
rect 22275 986 22939 1006
rect 22275 922 22281 986
rect 22345 922 22365 986
rect 22429 922 22449 986
rect 22513 922 22533 986
rect 22597 922 22617 986
rect 22681 922 22701 986
rect 22765 922 22785 986
rect 22849 922 22869 986
rect 22933 922 22939 986
rect 22275 902 22939 922
rect 22275 838 22281 902
rect 22345 838 22365 902
rect 22429 838 22449 902
rect 22513 838 22533 902
rect 22597 838 22617 902
rect 22681 838 22701 902
rect 22765 838 22785 902
rect 22849 838 22869 902
rect 22933 838 22939 902
rect 22275 818 22939 838
rect 22275 754 22281 818
rect 22345 754 22365 818
rect 22429 754 22449 818
rect 22513 754 22533 818
rect 22597 754 22617 818
rect 22681 754 22701 818
rect 22765 754 22785 818
rect 22849 754 22869 818
rect 22933 754 22939 818
rect 22275 734 22939 754
rect 22275 670 22281 734
rect 22345 670 22365 734
rect 22429 670 22449 734
rect 22513 670 22533 734
rect 22597 670 22617 734
rect 22681 670 22701 734
rect 22765 670 22785 734
rect 22849 670 22869 734
rect 22933 670 22939 734
rect 22275 650 22939 670
rect 22275 586 22281 650
rect 22345 586 22365 650
rect 22429 586 22449 650
rect 22513 586 22533 650
rect 22597 586 22617 650
rect 22681 586 22701 650
rect 22765 586 22785 650
rect 22849 586 22869 650
rect 22933 586 22939 650
rect 22275 566 22939 586
rect 22275 502 22281 566
rect 22345 502 22365 566
rect 22429 502 22449 566
rect 22513 502 22533 566
rect 22597 502 22617 566
rect 22681 502 22701 566
rect 22765 502 22785 566
rect 22849 502 22869 566
rect 22933 502 22939 566
rect 22275 482 22939 502
rect 22275 418 22281 482
rect 22345 418 22365 482
rect 22429 418 22449 482
rect 22513 418 22533 482
rect 22597 418 22617 482
rect 22681 418 22701 482
rect 22765 418 22785 482
rect 22849 418 22869 482
rect 22933 418 22939 482
rect 22275 417 22939 418
rect 17775 407 18175 413
rect 27746 407 28000 1497
rect 12671 297 13108 298
rect 12671 233 12672 297
rect 12736 233 12752 297
rect 12816 233 12963 297
rect 13027 233 13043 297
rect 13107 233 13108 297
rect 12671 232 13108 233
<< rmetal4 >>
rect 2257 24346 2259 24522
<< metal5 >>
rect 0 35157 254 40000
rect 27746 35157 28000 40000
rect 8019 26541 12627 29546
rect 0 14007 254 18997
rect 27746 14007 28000 18997
rect 0 12837 254 13687
rect 27746 12837 28000 13687
rect 0 11667 254 12517
rect 27746 11667 28000 12517
rect 0 9547 254 11347
rect 27746 9547 28000 11347
rect 0 8337 254 9227
rect 27746 8337 28000 9227
rect 0 7368 254 8017
rect 27746 7368 28000 8017
rect 0 6397 254 7047
rect 27746 6397 28000 7047
rect 0 5187 254 6077
rect 27746 5187 28000 6077
rect 0 3977 254 4867
rect 27746 3977 28000 4867
rect 0 3007 193 3657
rect 27807 3007 28000 3657
rect 0 1797 254 2687
rect 27746 1797 28000 2687
rect 0 427 254 1477
rect 27746 427 28000 1477
use sky130_fd_io__gpio_ctlv2_i2c_fix  sky130_fd_io__gpio_ctlv2_i2c_fix_0
timestamp 1666464484
transform 1 0 421 0 1 4115
box 173 -4115 27579 2717
use sky130_fd_io__gpio_ovtv2_amux_i2c_fix  sky130_fd_io__gpio_ovtv2_amux_i2c_fix_0
timestamp 1666464484
transform 1 0 1288 0 1 8163
box -1368 -8163 26923 25429
use sky130_fd_io__gpio_ovtv2_busses  sky130_fd_io__gpio_ovtv2_busses_0
timestamp 1666464484
transform 1 0 3360 0 1 549
box -3360 -142 24640 39451
use sky130_fd_io__gpio_ovtv2_ipath  sky130_fd_io__gpio_ovtv2_ipath_0
timestamp 1666464484
transform -1 0 28000 0 -1 3318
box 0 -5000 25393 3465
use sky130_fd_io__gpio_ovtv2_opath_i2c_fix_leak_fix  sky130_fd_io__gpio_ovtv2_opath_i2c_fix_leak_fix_0
timestamp 1666464484
transform 1 0 1 0 1 6235
box 136 -5849 28210 33916
use sky130_fd_io__gpio_ovtv2_tap_i2c_fix  sky130_fd_io__gpio_ovtv2_tap_i2c_fix_0
timestamp 1666464484
transform 1 0 26 0 1 26
box 50 1591 27974 39950
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_0
timestamp 1666464484
transform 0 -1 2648 -1 0 34282
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_1
timestamp 1666464484
transform 0 -1 2648 -1 0 33400
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_2
timestamp 1666464484
transform 0 -1 3152 -1 0 34282
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_3
timestamp 1666464484
transform 0 -1 3152 -1 0 33400
box 0 0 882 404
use sky130_fd_pr__antenna_diode_pw2nd_05v5__example_55959141808556  sky130_fd_pr__antenna_diode_pw2nd_05v5__example_55959141808556_0
timestamp 1666464484
transform 1 0 27419 0 1 37419
box 0 0 1 1
use sky130_fd_pr__m4short__example_55959141808557  sky130_fd_pr__m4short__example_55959141808557_0
timestamp 1666464484
transform 1 0 2198 0 1 24346
box 0 0 1 1
<< labels >>
flabel metal5 s 27746 11667 28000 12517 3 FreeSans 520 180 0 0 VSSIO_Q
port 1 nsew ground bidirectional
flabel metal5 s 27746 6397 28000 7047 3 FreeSans 520 180 0 0 VSWITCH
port 2 nsew power bidirectional
flabel metal5 s 27746 5187 28000 6077 3 FreeSans 520 180 0 0 VSSIO
port 3 nsew ground bidirectional
flabel metal5 s 27746 8337 28000 9227 3 FreeSans 520 180 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal5 s 27746 7368 28000 8017 3 FreeSans 520 180 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal5 s 27746 12837 28000 13687 3 FreeSans 520 180 0 0 VDDIO_Q
port 6 nsew power bidirectional
flabel metal5 s 27746 14007 28000 18997 3 FreeSans 520 180 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal5 s 27807 3007 28000 3657 3 FreeSans 520 180 0 0 VDDA
port 8 nsew power bidirectional
flabel metal5 s 27746 427 28000 1477 3 FreeSans 520 180 0 0 VCCHIB
port 9 nsew power bidirectional
flabel metal5 s 27746 1797 28000 2687 3 FreeSans 520 180 0 0 VCCD
port 10 nsew power bidirectional
flabel metal5 s 27746 3977 28000 4867 3 FreeSans 520 180 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal5 s 27746 9547 28000 11347 3 FreeSans 520 180 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal5 s 27746 35157 28000 40000 3 FreeSans 520 180 0 0 VSSIO
port 3 nsew ground bidirectional
flabel metal5 s 0 11667 254 12517 3 FreeSans 520 0 0 0 VSSIO_Q
port 1 nsew ground bidirectional
flabel metal5 s 0 6397 254 7047 3 FreeSans 520 0 0 0 VSWITCH
port 2 nsew power bidirectional
flabel metal5 s 0 5187 254 6077 3 FreeSans 520 0 0 0 VSSIO
port 3 nsew ground bidirectional
flabel metal5 s 0 8337 254 9227 3 FreeSans 520 0 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal5 s 0 7368 254 8017 3 FreeSans 520 0 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal5 s 0 12837 254 13687 3 FreeSans 520 0 0 0 VDDIO_Q
port 6 nsew power bidirectional
flabel metal5 s 0 14007 254 18997 3 FreeSans 520 0 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal5 s 0 3007 193 3657 3 FreeSans 520 0 0 0 VDDA
port 8 nsew power bidirectional
flabel metal5 s 0 427 254 1477 3 FreeSans 520 0 0 0 VCCHIB
port 9 nsew power bidirectional
flabel metal5 s 0 1797 254 2687 3 FreeSans 520 0 0 0 VCCD
port 10 nsew power bidirectional
flabel metal5 s 0 3977 254 4867 3 FreeSans 520 0 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal5 s 0 9547 254 11347 3 FreeSans 520 0 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal5 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 3 nsew ground bidirectional
flabel metal5 s 8019 26541 12627 29546 3 FreeSans 8000 0 0 0 PAD
port 11 nsew signal bidirectional
flabel metal4 s 27746 10329 28000 10565 3 FreeSans 520 180 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 27746 9547 28000 9613 3 FreeSans 520 180 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 27746 11647 28000 12537 3 FreeSans 520 180 0 0 VSSIO_Q
port 1 nsew ground bidirectional
flabel metal4 s 27746 11281 28000 11347 3 FreeSans 520 180 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 27746 35157 28000 40000 3 FreeSans 520 180 0 0 VSSIO
port 3 nsew ground bidirectional
flabel metal4 s 27746 407 28000 1497 3 FreeSans 520 180 0 0 VCCHIB
port 9 nsew power bidirectional
flabel metal4 s 27746 1777 28000 2707 3 FreeSans 520 180 0 0 VCCD
port 10 nsew power bidirectional
flabel metal4 s 27807 2987 28000 3677 3 FreeSans 520 180 0 0 VDDA
port 8 nsew power bidirectional
flabel metal4 s 27746 3957 28000 4887 3 FreeSans 520 180 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal4 s 27746 5167 28000 6097 3 FreeSans 520 180 0 0 VSSIO
port 3 nsew ground bidirectional
flabel metal4 s 27746 6377 28000 7067 3 FreeSans 520 180 0 0 VSWITCH
port 2 nsew power bidirectional
flabel metal4 s 27746 14007 28000 19000 3 FreeSans 520 180 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal4 s 27746 12817 28000 13707 3 FreeSans 520 180 0 0 VDDIO_Q
port 6 nsew power bidirectional
flabel metal4 s 27746 10625 28000 11221 3 FreeSans 520 180 0 0 AMUXBUS_A
port 12 nsew signal bidirectional
flabel metal4 s 27746 9673 28000 10269 3 FreeSans 520 180 0 0 AMUXBUS_B
port 13 nsew signal bidirectional
flabel metal4 s 27746 8317 28000 9247 3 FreeSans 520 180 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal4 s 27746 7347 28000 8037 3 FreeSans 520 180 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 0 10329 254 10565 3 FreeSans 520 0 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 0 9547 254 9613 3 FreeSans 520 0 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 0 11647 254 12537 3 FreeSans 520 0 0 0 VSSIO_Q
port 1 nsew ground bidirectional
flabel metal4 s 0 11281 254 11347 3 FreeSans 520 0 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 3 nsew ground bidirectional
flabel metal4 s 0 407 254 1497 3 FreeSans 520 0 0 0 VCCHIB
port 9 nsew power bidirectional
flabel metal4 s 0 1777 254 2707 3 FreeSans 520 0 0 0 VCCD
port 10 nsew power bidirectional
flabel metal4 s 0 2987 193 3677 3 FreeSans 520 0 0 0 VDDA
port 8 nsew power bidirectional
flabel metal4 s 0 3957 254 4887 3 FreeSans 520 0 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal4 s 0 5167 254 6097 3 FreeSans 520 0 0 0 VSSIO
port 3 nsew ground bidirectional
flabel metal4 s 0 6377 254 7067 3 FreeSans 520 0 0 0 VSWITCH
port 2 nsew power bidirectional
flabel metal4 s 0 14007 254 19000 3 FreeSans 520 0 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal4 s 0 12817 254 13707 3 FreeSans 520 0 0 0 VDDIO_Q
port 6 nsew power bidirectional
flabel metal4 s 0 10625 254 11221 3 FreeSans 520 0 0 0 AMUXBUS_A
port 12 nsew signal bidirectional
flabel metal4 s 0 9673 254 10269 3 FreeSans 520 0 0 0 AMUXBUS_B
port 13 nsew signal bidirectional
flabel metal4 s 0 8317 254 9247 3 FreeSans 520 0 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal4 s 0 7347 254 8037 3 FreeSans 520 0 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal3 s 25825 0 25891 134 3 FreeSans 200 0 0 0 DM[0]
port 14 nsew signal input
flabel metal3 s 25655 0 25721 134 3 FreeSans 200 0 0 0 DM[1]
port 15 nsew signal input
flabel metal3 s 21679 0 21745 134 3 FreeSans 200 0 0 0 DM[2]
port 16 nsew signal input
flabel metal3 s 21509 0 21575 134 3 FreeSans 200 0 0 0 INP_DIS
port 17 nsew signal input
flabel metal3 s 17533 0 17599 134 3 FreeSans 200 0 0 0 VTRIP_SEL
port 18 nsew signal input
flabel metal3 s 17363 0 17429 134 3 FreeSans 200 180 0 0 IB_MODE_SEL[0]
port 19 nsew signal input
flabel metal3 s 13387 0 13453 134 3 FreeSans 200 0 0 0 IB_MODE_SEL[1]
port 20 nsew signal input
flabel metal3 s 13217 0 13283 134 3 FreeSans 200 0 0 0 SLEW_CTL[0]
port 21 nsew signal input
flabel metal3 s 9241 0 9307 134 3 FreeSans 200 0 0 0 SLEW_CTL[1]
port 22 nsew signal input
flabel metal3 s 9071 0 9137 134 3 FreeSans 200 0 0 0 HYS_TRIM
port 23 nsew signal input
flabel metal3 s 5471 0 5537 134 3 FreeSans 200 0 0 0 HLD_OVR
port 24 nsew signal input
flabel metal3 s 4427 0 4493 134 3 FreeSans 200 0 0 0 ENABLE_H
port 25 nsew signal input
flabel metal3 s 3927 0 3993 134 3 FreeSans 200 0 0 0 HLD_H_N
port 26 nsew signal input
flabel metal3 s 1754 0 1820 134 3 FreeSans 200 0 0 0 ENABLE_VDDA_H
port 27 nsew signal input
flabel metal3 s 1623 0 1689 134 3 FreeSans 200 0 0 0 ANALOG_EN
port 28 nsew signal input
flabel metal3 s 1422 0 1488 134 3 FreeSans 200 0 0 0 ENABLE_INP_H
port 29 nsew signal input
flabel metal3 s 4076 0 4142 134 3 FreeSans 200 0 0 0 IN
port 30 nsew signal output
flabel metal3 s 4876 0 4942 134 3 FreeSans 200 0 0 0 IN_H
port 31 nsew signal output
flabel metal3 s 8807 0 8873 134 3 FreeSans 200 0 0 0 VINREF
port 32 nsew signal input
flabel metal3 s 14825 0 14891 157 3 FreeSans 520 90 0 0 OUT
port 33 nsew signal input
flabel metal3 s 13047 0 13113 134 3 FreeSans 520 90 0 0 ANALOG_POL
port 34 nsew signal input
flabel metal3 s 10331 0 10397 156 3 FreeSans 520 90 0 0 ANALOG_SEL
port 35 nsew signal input
flabel metal3 s 25028 0 25094 134 3 FreeSans 520 90 0 0 SLOW
port 36 nsew signal input
flabel metal3 s 24889 0 24955 183 3 FreeSans 520 90 0 0 OE_N
port 37 nsew signal input
flabel metal3 s 25995 0 26061 166 3 FreeSans 520 270 0 0 TIE_HI_ESD
port 38 nsew signal output
flabel metal3 s 23058 0 23178 166 3 FreeSans 520 270 0 0 TIE_LO_ESD
port 39 nsew signal output
flabel metal3 s 321 0 440 166 3 FreeSans 520 90 0 0 PAD_A_ESD_0_H
port 40 nsew signal bidirectional
flabel metal3 s 66 0 186 166 3 FreeSans 520 90 0 0 PAD_A_ESD_1_H
port 41 nsew signal bidirectional
flabel metal3 s 577 0 697 166 3 FreeSans 520 90 0 0 PAD_A_NOESD_H
port 42 nsew signal bidirectional
flabel metal3 s 1153 0 1273 129 3 FreeSans 520 0 0 0 ENABLE_VSWITCH_H
port 43 nsew signal input
flabel metal3 s 19169 0 19243 74 3 FreeSans 520 90 0 0 ENABLE_VDDIO
port 44 nsew signal input
flabel comment s 27364 3338 27364 3338 0 FreeSans 200 0 0 0 DM_H_N<0>
flabel comment s 27364 3422 27364 3422 0 FreeSans 200 0 0 0 DM_H_N<1>
flabel comment s 27364 3500 27364 3500 0 FreeSans 200 0 0 0 DM_H_N<2>
flabel comment s 3811 3339 3811 3339 0 FreeSans 200 0 0 0 SLEW_CTL_H<0>
flabel comment s 3811 3416 3811 3416 0 FreeSans 200 0 0 0 SLEW_CTL_H<1>
flabel comment s 3811 3494 3811 3494 0 FreeSans 200 0 0 0 SLEW_CTL_H_N<0>
flabel comment s 3811 3581 3811 3581 0 FreeSans 200 0 0 0 SLEW_CTL_H_N<1>
flabel comment s 19013 3335 19013 3335 0 FreeSans 200 0 0 0 IB_MODE_SEL_H<0>
flabel comment s 19013 3417 19013 3417 0 FreeSans 200 0 0 0 IB_MODE_SEL_H<1>
flabel comment s 20264 3488 20264 3488 0 FreeSans 200 0 0 0 VTRIP_SEL_H
flabel comment s 21050 3577 21050 3577 0 FreeSans 200 0 0 0 INP_DIS_H_N
flabel comment s 27364 3580 27364 3580 0 FreeSans 200 0 0 0 DM_H<0>
flabel comment s 27364 3661 27364 3661 0 FreeSans 200 0 0 0 DM_H<1>
flabel comment s 27364 3736 27364 3736 0 FreeSans 200 0 0 0 DM_H<2>
flabel comment s 27364 4014 27364 4014 0 FreeSans 200 0 0 0 OD_I_H
flabel comment s 27364 4094 27364 4094 0 FreeSans 200 0 0 0 HLD_I_H_N
flabel comment s 27364 3817 27364 3817 0 FreeSans 200 0 0 0 HLD_I_OVR_H
flabel comment s 645 3227 645 3227 0 FreeSans 200 0 0 0 SLEW_CTL_H_N<1>
flabel comment s 645 3140 645 3140 0 FreeSans 200 0 0 0 SLEW_CTL_H_N<0>
flabel comment s 645 3062 645 3062 0 FreeSans 200 0 0 0 SLEW_CTL_H<1>
flabel comment s 645 2985 645 2985 0 FreeSans 200 0 0 0 SLEW_CTL_H<0>
flabel comment s 1943 2853 1943 2853 0 FreeSans 440 0 0 0 ANTENNA FIX
flabel comment s 1448 33476 1448 33476 0 FreeSans 400 90 0 0 SLEW_CTL_H_N<0>
flabel comment s 1323 33470 1323 33470 0 FreeSans 400 90 0 0 SLEW_CTL_H_N<1>
flabel comment s 2075 33462 2075 33462 0 FreeSans 400 90 0 0 SLEW_CTL_H<0>
flabel comment s 1559 33523 1559 33523 0 FreeSans 400 90 0 0 SLEW_CTL_H<1>
flabel comment s 1559 32055 1559 32055 0 FreeSans 400 90 0 0 SLEW_CTL_H<1>
flabel comment s 2075 11425 2075 11425 0 FreeSans 400 90 0 0 SLEW_CTL_H<0>
flabel comment s 1559 11486 1559 11486 0 FreeSans 400 90 0 0 SLEW_CTL_H<1>
flabel comment s 732 10300 732 10300 0 FreeSans 400 90 0 0 SLEW_CTL_H_N<0>
flabel comment s 607 10361 607 10361 0 FreeSans 400 90 0 0 SLEW_CTL_H_N<1>
flabel comment s 1303 3565 1303 3565 0 FreeSans 400 90 0 0 SLEW_CTL_H<0>
flabel comment s 1178 3626 1178 3626 0 FreeSans 400 90 0 0 SLEW_CTL_H<1>
flabel comment s 607 3626 607 3626 0 FreeSans 400 90 0 0 SLEW_CTL_H_N<1>
flabel comment s 24735 1646 24735 1646 0 FreeSans 440 0 0 0 ANTENNA FIX
flabel comment s 21351 1652 21351 1652 0 FreeSans 440 0 0 0 ANTENNA FIX
flabel comment s 12875 1651 12875 1651 0 FreeSans 440 0 0 0 ANTENNA FIX
flabel comment s 10549 1652 10549 1652 0 FreeSans 440 0 0 0 ANTENNA FIX
flabel comment s 8914 1649 8914 1649 0 FreeSans 440 0 0 0 ANTENNA FIX
flabel comment s 5318 2847 5318 2847 0 FreeSans 440 0 0 0 ANTENNA FIX
flabel comment s 1924 5044 1924 5044 0 FreeSans 440 0 0 0 ANTENNA FIX
flabel comment s 1783 3565 1783 3565 0 FreeSans 400 90 0 0 SLEW_CTL_H_N<0>
flabel comment s 19458 38439 19458 38439 0 FreeSans 200 0 0 0 M1_FLOAT
rlabel metal4 s 27746 10625 28000 11221 1 AMUXBUS_A
port 12 nsew signal bidirectional
rlabel metal4 s 27746 9673 28000 10269 1 AMUXBUS_B
port 13 nsew signal bidirectional
rlabel metal4 s 27746 2693 28000 2707 1 VCCD
port 10 nsew power bidirectional
rlabel metal4 s 27746 1777 28000 1786 1 VCCD
port 10 nsew power bidirectional
rlabel metal4 s 27651 1786 28000 2693 1 VCCD
port 10 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 1 VCCD
port 10 nsew power bidirectional
rlabel metal5 s 27746 1797 28000 2687 1 VCCD
port 10 nsew power bidirectional
rlabel metal4 s 27746 407 28000 1497 1 VCCHIB
port 9 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 1 VCCHIB
port 9 nsew power bidirectional
rlabel metal5 s 27746 427 28000 1477 1 VCCHIB
port 9 nsew power bidirectional
rlabel metal4 s 27807 2987 28000 3677 1 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 1 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 27807 3007 28000 3657 1 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 27746 3957 28000 4887 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 27746 14007 28000 19000 1 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 1 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 1 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 27746 3977 28000 4867 1 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 27746 14007 28000 18997 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 27746 12817 28000 13707 1 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 1 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal5 s 27746 12837 28000 13687 1 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal4 s 0 9547 254 9613 1 VSSA
port 5 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 1 VSSA
port 5 nsew ground bidirectional
rlabel metal4 s 0 11281 254 11347 1 VSSA
port 5 nsew ground bidirectional
rlabel metal4 s 27746 7347 28000 8037 1 VSSA
port 5 nsew ground bidirectional
rlabel metal4 s 27746 9547 28000 9613 1 VSSA
port 5 nsew ground bidirectional
rlabel metal4 s 27746 10329 28000 10565 1 VSSA
port 5 nsew ground bidirectional
rlabel metal4 s 27746 11281 28000 11347 1 VSSA
port 5 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 1 VSSA
port 5 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 1 VSSA
port 5 nsew ground bidirectional
rlabel metal5 s 27746 7368 28000 8017 1 VSSA
port 5 nsew ground bidirectional
rlabel metal5 s 27746 9547 28000 11347 1 VSSA
port 5 nsew ground bidirectional
rlabel metal4 s 27746 8317 28000 9247 1 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 1 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 27746 8337 28000 9227 1 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 1 VSSIO
port 3 nsew ground bidirectional
rlabel metal4 s 27746 35157 28000 40000 1 VSSIO
port 3 nsew ground bidirectional
rlabel metal4 s 27746 5167 28000 6097 1 VSSIO
port 3 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 1 VSSIO
port 3 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 1 VSSIO
port 3 nsew ground bidirectional
rlabel metal5 s 27746 35157 28000 40000 1 VSSIO
port 3 nsew ground bidirectional
rlabel metal5 s 27746 5187 28000 6077 1 VSSIO
port 3 nsew ground bidirectional
rlabel metal4 s 27746 11647 28000 12537 1 VSSIO_Q
port 1 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 1 VSSIO_Q
port 1 nsew ground bidirectional
rlabel metal5 s 27746 11667 28000 12517 1 VSSIO_Q
port 1 nsew ground bidirectional
rlabel metal4 s 27746 6377 28000 7067 1 VSWITCH
port 2 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 1 VSWITCH
port 2 nsew power bidirectional
rlabel metal5 s 27746 6397 28000 7047 1 VSWITCH
port 2 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 28000 40000
string GDS_END 43499818
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42873614
string LEFclass PAD
string LEFsymmetry X Y R90
<< end >>
