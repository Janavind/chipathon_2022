magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< dnwell >>
tri -700 6714 -614 6800 se
rect -614 6714 764 6800
tri 764 6714 850 6800 sw
rect -700 -714 850 6714
tri -700 -800 -614 -714 ne
rect -614 -800 764 -714
tri 764 -800 850 -714 nw
<< nwell >>
rect -10 0 160 6000
<< pwell >>
rect -1166 7074 1316 7208
rect -1166 6026 -1032 7074
rect 1182 6026 1316 7074
rect -1166 -26 -574 6026
rect 724 -26 1316 6026
rect -1166 -1074 -1032 -26
rect 1182 -1074 1316 -26
rect -1166 -1208 1316 -1074
<< obsactive >>
rect -1500 -1600 1700 7600
<< locali >>
rect -1140 7158 1290 7182
rect -1140 7124 -986 7158
rect -952 7124 -914 7158
rect -880 7124 -842 7158
rect -808 7124 -770 7158
rect -736 7124 -698 7158
rect -664 7124 -626 7158
rect -592 7124 -554 7158
rect -520 7124 -482 7158
rect -448 7124 -410 7158
rect -376 7124 -338 7158
rect -304 7124 -266 7158
rect -232 7124 -194 7158
rect -160 7124 -122 7158
rect -88 7124 -50 7158
rect -16 7124 22 7158
rect 56 7124 94 7158
rect 128 7124 166 7158
rect 200 7124 238 7158
rect 272 7124 310 7158
rect 344 7124 382 7158
rect 416 7124 454 7158
rect 488 7124 526 7158
rect 560 7124 598 7158
rect 632 7124 670 7158
rect 704 7124 742 7158
rect 776 7124 814 7158
rect 848 7124 886 7158
rect 920 7124 958 7158
rect 992 7124 1030 7158
rect 1064 7124 1102 7158
rect 1136 7124 1290 7158
rect -1140 7100 1290 7124
rect -1140 7085 -1058 7100
rect -1140 7051 -1116 7085
rect -1082 7051 -1058 7085
rect -1140 7013 -1058 7051
rect -1140 6979 -1116 7013
rect -1082 6979 -1058 7013
rect -1140 6941 -1058 6979
rect -1140 6907 -1116 6941
rect -1082 6907 -1058 6941
rect -1140 6869 -1058 6907
rect -1140 6835 -1116 6869
rect -1082 6835 -1058 6869
rect -1140 6797 -1058 6835
rect -1140 6763 -1116 6797
rect -1082 6763 -1058 6797
rect -1140 6725 -1058 6763
rect -1140 6691 -1116 6725
rect -1082 6691 -1058 6725
rect -1140 6653 -1058 6691
rect -1140 6619 -1116 6653
rect -1082 6619 -1058 6653
rect -1140 6581 -1058 6619
rect -1140 6547 -1116 6581
rect -1082 6547 -1058 6581
rect -1140 -547 -1058 6547
rect 1208 7085 1290 7100
rect 1208 7051 1232 7085
rect 1266 7051 1290 7085
rect 1208 7013 1290 7051
rect 1208 6979 1232 7013
rect 1266 6979 1290 7013
rect 1208 6941 1290 6979
rect 1208 6907 1232 6941
rect 1266 6907 1290 6941
rect 1208 6869 1290 6907
rect 1208 6835 1232 6869
rect 1266 6835 1290 6869
rect 1208 6797 1290 6835
rect 1208 6763 1232 6797
rect 1266 6763 1290 6797
rect 1208 6725 1290 6763
rect 1208 6691 1232 6725
rect 1266 6691 1290 6725
rect 1208 6653 1290 6691
rect 1208 6619 1232 6653
rect 1266 6619 1290 6653
rect 1208 6581 1290 6619
rect 1208 6547 1232 6581
rect 1266 6547 1290 6581
rect -962 5969 -896 5991
rect -962 5935 -946 5969
rect -912 5935 -896 5969
rect 1046 5969 1112 5991
rect -962 5897 -896 5935
rect -962 5863 -946 5897
rect -912 5863 -896 5897
rect -962 5825 -896 5863
rect -962 5791 -946 5825
rect -912 5791 -896 5825
rect -962 5753 -896 5791
rect -962 5719 -946 5753
rect -912 5719 -896 5753
rect -962 5681 -896 5719
rect -962 5647 -946 5681
rect -912 5647 -896 5681
rect -962 5609 -896 5647
rect -962 5575 -946 5609
rect -912 5575 -896 5609
rect -962 5537 -896 5575
rect -962 5503 -946 5537
rect -912 5503 -896 5537
rect -962 5465 -896 5503
rect -962 5431 -946 5465
rect -912 5431 -896 5465
rect -962 5393 -896 5431
rect -962 5359 -946 5393
rect -912 5359 -896 5393
rect -962 5321 -896 5359
rect -962 5287 -946 5321
rect -912 5287 -896 5321
rect -962 5249 -896 5287
rect -962 5215 -946 5249
rect -912 5215 -896 5249
rect -962 5177 -896 5215
rect -962 5143 -946 5177
rect -912 5143 -896 5177
rect -962 5105 -896 5143
rect -962 5071 -946 5105
rect -912 5071 -896 5105
rect -962 5033 -896 5071
rect -962 4999 -946 5033
rect -912 4999 -896 5033
rect -962 4961 -896 4999
rect -962 4927 -946 4961
rect -912 4927 -896 4961
rect -962 4889 -896 4927
rect -962 4855 -946 4889
rect -912 4855 -896 4889
rect -962 4817 -896 4855
rect -962 4783 -946 4817
rect -912 4783 -896 4817
rect -962 4745 -896 4783
rect -962 4711 -946 4745
rect -912 4711 -896 4745
rect -962 4673 -896 4711
rect -962 4639 -946 4673
rect -912 4639 -896 4673
rect -962 4601 -896 4639
rect -962 4567 -946 4601
rect -912 4567 -896 4601
rect -962 4529 -896 4567
rect -962 4495 -946 4529
rect -912 4495 -896 4529
rect -962 4457 -896 4495
rect -962 4423 -946 4457
rect -912 4423 -896 4457
rect -962 4385 -896 4423
rect -962 4351 -946 4385
rect -912 4351 -896 4385
rect -962 4313 -896 4351
rect -962 4279 -946 4313
rect -912 4279 -896 4313
rect -962 4241 -896 4279
rect -962 4207 -946 4241
rect -912 4207 -896 4241
rect -962 4169 -896 4207
rect -962 4135 -946 4169
rect -912 4135 -896 4169
rect -962 4097 -896 4135
rect -962 4063 -946 4097
rect -912 4063 -896 4097
rect -962 4025 -896 4063
rect -962 3991 -946 4025
rect -912 3991 -896 4025
rect -962 3953 -896 3991
rect -962 3919 -946 3953
rect -912 3919 -896 3953
rect -962 3881 -896 3919
rect -962 3847 -946 3881
rect -912 3847 -896 3881
rect -962 3809 -896 3847
rect -962 3775 -946 3809
rect -912 3775 -896 3809
rect -962 3737 -896 3775
rect -962 3703 -946 3737
rect -912 3703 -896 3737
rect -962 3665 -896 3703
rect -962 3631 -946 3665
rect -912 3631 -896 3665
rect -962 3593 -896 3631
rect -962 3559 -946 3593
rect -912 3559 -896 3593
rect -962 3521 -896 3559
rect -962 3487 -946 3521
rect -912 3487 -896 3521
rect -962 3449 -896 3487
rect -962 3415 -946 3449
rect -912 3415 -896 3449
rect -962 3377 -896 3415
rect -962 3343 -946 3377
rect -912 3343 -896 3377
rect -962 3305 -896 3343
rect -962 3271 -946 3305
rect -912 3271 -896 3305
rect -962 3233 -896 3271
rect -962 3199 -946 3233
rect -912 3199 -896 3233
rect -962 3161 -896 3199
rect -962 3127 -946 3161
rect -912 3127 -896 3161
rect -962 3089 -896 3127
rect -962 3055 -946 3089
rect -912 3055 -896 3089
rect -962 3017 -896 3055
rect -962 2983 -946 3017
rect -912 2983 -896 3017
rect -962 2945 -896 2983
rect -962 2911 -946 2945
rect -912 2911 -896 2945
rect -962 2873 -896 2911
rect -962 2839 -946 2873
rect -912 2839 -896 2873
rect -962 2801 -896 2839
rect -962 2767 -946 2801
rect -912 2767 -896 2801
rect -962 2729 -896 2767
rect -962 2695 -946 2729
rect -912 2695 -896 2729
rect -962 2657 -896 2695
rect -962 2623 -946 2657
rect -912 2623 -896 2657
rect -962 2585 -896 2623
rect -962 2551 -946 2585
rect -912 2551 -896 2585
rect -962 2513 -896 2551
rect -962 2479 -946 2513
rect -912 2479 -896 2513
rect -962 2441 -896 2479
rect -962 2407 -946 2441
rect -912 2407 -896 2441
rect -962 2369 -896 2407
rect -962 2335 -946 2369
rect -912 2335 -896 2369
rect -962 2297 -896 2335
rect -962 2263 -946 2297
rect -912 2263 -896 2297
rect -962 2225 -896 2263
rect -962 2191 -946 2225
rect -912 2191 -896 2225
rect -962 2153 -896 2191
rect -962 2119 -946 2153
rect -912 2119 -896 2153
rect -962 2081 -896 2119
rect -962 2047 -946 2081
rect -912 2047 -896 2081
rect -962 2009 -896 2047
rect -962 1975 -946 2009
rect -912 1975 -896 2009
rect -962 1937 -896 1975
rect -962 1903 -946 1937
rect -912 1903 -896 1937
rect -962 1865 -896 1903
rect -962 1831 -946 1865
rect -912 1831 -896 1865
rect -962 1793 -896 1831
rect -962 1759 -946 1793
rect -912 1759 -896 1793
rect -962 1721 -896 1759
rect -962 1687 -946 1721
rect -912 1687 -896 1721
rect -962 1649 -896 1687
rect -962 1615 -946 1649
rect -912 1615 -896 1649
rect -962 1577 -896 1615
rect -962 1543 -946 1577
rect -912 1543 -896 1577
rect -962 1505 -896 1543
rect -962 1471 -946 1505
rect -912 1471 -896 1505
rect -962 1433 -896 1471
rect -962 1399 -946 1433
rect -912 1399 -896 1433
rect -962 1361 -896 1399
rect -962 1327 -946 1361
rect -912 1327 -896 1361
rect -962 1289 -896 1327
rect -962 1255 -946 1289
rect -912 1255 -896 1289
rect -962 1217 -896 1255
rect -962 1183 -946 1217
rect -912 1183 -896 1217
rect -962 1145 -896 1183
rect -962 1111 -946 1145
rect -912 1111 -896 1145
rect -962 1073 -896 1111
rect -962 1039 -946 1073
rect -912 1039 -896 1073
rect -962 1001 -896 1039
rect -962 967 -946 1001
rect -912 967 -896 1001
rect -962 929 -896 967
rect -962 895 -946 929
rect -912 895 -896 929
rect -962 857 -896 895
rect -962 823 -946 857
rect -912 823 -896 857
rect -962 785 -896 823
rect -962 751 -946 785
rect -912 751 -896 785
rect -962 713 -896 751
rect -962 679 -946 713
rect -912 679 -896 713
rect -962 641 -896 679
rect -962 607 -946 641
rect -912 607 -896 641
rect -962 569 -896 607
rect -962 535 -946 569
rect -912 535 -896 569
rect -962 497 -896 535
rect -962 463 -946 497
rect -912 463 -896 497
rect -962 425 -896 463
rect -962 391 -946 425
rect -912 391 -896 425
rect -962 353 -896 391
rect -962 319 -946 353
rect -912 319 -896 353
rect -962 281 -896 319
rect -962 247 -946 281
rect -912 247 -896 281
rect -962 209 -896 247
rect -962 175 -946 209
rect -912 175 -896 209
rect -962 137 -896 175
rect -962 103 -946 137
rect -912 103 -896 137
rect -962 65 -896 103
rect -962 31 -946 65
rect -912 31 -896 65
rect 8 5933 142 5957
rect 8 67 22 5933
rect 128 67 142 5933
rect 8 43 142 67
rect 1046 5935 1062 5969
rect 1096 5935 1112 5969
rect 1046 5897 1112 5935
rect 1046 5863 1062 5897
rect 1096 5863 1112 5897
rect 1046 5825 1112 5863
rect 1046 5791 1062 5825
rect 1096 5791 1112 5825
rect 1046 5753 1112 5791
rect 1046 5719 1062 5753
rect 1096 5719 1112 5753
rect 1046 5681 1112 5719
rect 1046 5647 1062 5681
rect 1096 5647 1112 5681
rect 1046 5609 1112 5647
rect 1046 5575 1062 5609
rect 1096 5575 1112 5609
rect 1046 5537 1112 5575
rect 1046 5503 1062 5537
rect 1096 5503 1112 5537
rect 1046 5465 1112 5503
rect 1046 5431 1062 5465
rect 1096 5431 1112 5465
rect 1046 5393 1112 5431
rect 1046 5359 1062 5393
rect 1096 5359 1112 5393
rect 1046 5321 1112 5359
rect 1046 5287 1062 5321
rect 1096 5287 1112 5321
rect 1046 5249 1112 5287
rect 1046 5215 1062 5249
rect 1096 5215 1112 5249
rect 1046 5177 1112 5215
rect 1046 5143 1062 5177
rect 1096 5143 1112 5177
rect 1046 5105 1112 5143
rect 1046 5071 1062 5105
rect 1096 5071 1112 5105
rect 1046 5033 1112 5071
rect 1046 4999 1062 5033
rect 1096 4999 1112 5033
rect 1046 4961 1112 4999
rect 1046 4927 1062 4961
rect 1096 4927 1112 4961
rect 1046 4889 1112 4927
rect 1046 4855 1062 4889
rect 1096 4855 1112 4889
rect 1046 4817 1112 4855
rect 1046 4783 1062 4817
rect 1096 4783 1112 4817
rect 1046 4745 1112 4783
rect 1046 4711 1062 4745
rect 1096 4711 1112 4745
rect 1046 4673 1112 4711
rect 1046 4639 1062 4673
rect 1096 4639 1112 4673
rect 1046 4601 1112 4639
rect 1046 4567 1062 4601
rect 1096 4567 1112 4601
rect 1046 4529 1112 4567
rect 1046 4495 1062 4529
rect 1096 4495 1112 4529
rect 1046 4457 1112 4495
rect 1046 4423 1062 4457
rect 1096 4423 1112 4457
rect 1046 4385 1112 4423
rect 1046 4351 1062 4385
rect 1096 4351 1112 4385
rect 1046 4313 1112 4351
rect 1046 4279 1062 4313
rect 1096 4279 1112 4313
rect 1046 4241 1112 4279
rect 1046 4207 1062 4241
rect 1096 4207 1112 4241
rect 1046 4169 1112 4207
rect 1046 4135 1062 4169
rect 1096 4135 1112 4169
rect 1046 4097 1112 4135
rect 1046 4063 1062 4097
rect 1096 4063 1112 4097
rect 1046 4025 1112 4063
rect 1046 3991 1062 4025
rect 1096 3991 1112 4025
rect 1046 3953 1112 3991
rect 1046 3919 1062 3953
rect 1096 3919 1112 3953
rect 1046 3881 1112 3919
rect 1046 3847 1062 3881
rect 1096 3847 1112 3881
rect 1046 3809 1112 3847
rect 1046 3775 1062 3809
rect 1096 3775 1112 3809
rect 1046 3737 1112 3775
rect 1046 3703 1062 3737
rect 1096 3703 1112 3737
rect 1046 3665 1112 3703
rect 1046 3631 1062 3665
rect 1096 3631 1112 3665
rect 1046 3593 1112 3631
rect 1046 3559 1062 3593
rect 1096 3559 1112 3593
rect 1046 3521 1112 3559
rect 1046 3487 1062 3521
rect 1096 3487 1112 3521
rect 1046 3449 1112 3487
rect 1046 3415 1062 3449
rect 1096 3415 1112 3449
rect 1046 3377 1112 3415
rect 1046 3343 1062 3377
rect 1096 3343 1112 3377
rect 1046 3305 1112 3343
rect 1046 3271 1062 3305
rect 1096 3271 1112 3305
rect 1046 3233 1112 3271
rect 1046 3199 1062 3233
rect 1096 3199 1112 3233
rect 1046 3161 1112 3199
rect 1046 3127 1062 3161
rect 1096 3127 1112 3161
rect 1046 3089 1112 3127
rect 1046 3055 1062 3089
rect 1096 3055 1112 3089
rect 1046 3017 1112 3055
rect 1046 2983 1062 3017
rect 1096 2983 1112 3017
rect 1046 2945 1112 2983
rect 1046 2911 1062 2945
rect 1096 2911 1112 2945
rect 1046 2873 1112 2911
rect 1046 2839 1062 2873
rect 1096 2839 1112 2873
rect 1046 2801 1112 2839
rect 1046 2767 1062 2801
rect 1096 2767 1112 2801
rect 1046 2729 1112 2767
rect 1046 2695 1062 2729
rect 1096 2695 1112 2729
rect 1046 2657 1112 2695
rect 1046 2623 1062 2657
rect 1096 2623 1112 2657
rect 1046 2585 1112 2623
rect 1046 2551 1062 2585
rect 1096 2551 1112 2585
rect 1046 2513 1112 2551
rect 1046 2479 1062 2513
rect 1096 2479 1112 2513
rect 1046 2441 1112 2479
rect 1046 2407 1062 2441
rect 1096 2407 1112 2441
rect 1046 2369 1112 2407
rect 1046 2335 1062 2369
rect 1096 2335 1112 2369
rect 1046 2297 1112 2335
rect 1046 2263 1062 2297
rect 1096 2263 1112 2297
rect 1046 2225 1112 2263
rect 1046 2191 1062 2225
rect 1096 2191 1112 2225
rect 1046 2153 1112 2191
rect 1046 2119 1062 2153
rect 1096 2119 1112 2153
rect 1046 2081 1112 2119
rect 1046 2047 1062 2081
rect 1096 2047 1112 2081
rect 1046 2009 1112 2047
rect 1046 1975 1062 2009
rect 1096 1975 1112 2009
rect 1046 1937 1112 1975
rect 1046 1903 1062 1937
rect 1096 1903 1112 1937
rect 1046 1865 1112 1903
rect 1046 1831 1062 1865
rect 1096 1831 1112 1865
rect 1046 1793 1112 1831
rect 1046 1759 1062 1793
rect 1096 1759 1112 1793
rect 1046 1721 1112 1759
rect 1046 1687 1062 1721
rect 1096 1687 1112 1721
rect 1046 1649 1112 1687
rect 1046 1615 1062 1649
rect 1096 1615 1112 1649
rect 1046 1577 1112 1615
rect 1046 1543 1062 1577
rect 1096 1543 1112 1577
rect 1046 1505 1112 1543
rect 1046 1471 1062 1505
rect 1096 1471 1112 1505
rect 1046 1433 1112 1471
rect 1046 1399 1062 1433
rect 1096 1399 1112 1433
rect 1046 1361 1112 1399
rect 1046 1327 1062 1361
rect 1096 1327 1112 1361
rect 1046 1289 1112 1327
rect 1046 1255 1062 1289
rect 1096 1255 1112 1289
rect 1046 1217 1112 1255
rect 1046 1183 1062 1217
rect 1096 1183 1112 1217
rect 1046 1145 1112 1183
rect 1046 1111 1062 1145
rect 1096 1111 1112 1145
rect 1046 1073 1112 1111
rect 1046 1039 1062 1073
rect 1096 1039 1112 1073
rect 1046 1001 1112 1039
rect 1046 967 1062 1001
rect 1096 967 1112 1001
rect 1046 929 1112 967
rect 1046 895 1062 929
rect 1096 895 1112 929
rect 1046 857 1112 895
rect 1046 823 1062 857
rect 1096 823 1112 857
rect 1046 785 1112 823
rect 1046 751 1062 785
rect 1096 751 1112 785
rect 1046 713 1112 751
rect 1046 679 1062 713
rect 1096 679 1112 713
rect 1046 641 1112 679
rect 1046 607 1062 641
rect 1096 607 1112 641
rect 1046 569 1112 607
rect 1046 535 1062 569
rect 1096 535 1112 569
rect 1046 497 1112 535
rect 1046 463 1062 497
rect 1096 463 1112 497
rect 1046 425 1112 463
rect 1046 391 1062 425
rect 1096 391 1112 425
rect 1046 353 1112 391
rect 1046 319 1062 353
rect 1096 319 1112 353
rect 1046 281 1112 319
rect 1046 247 1062 281
rect 1096 247 1112 281
rect 1046 209 1112 247
rect 1046 175 1062 209
rect 1096 175 1112 209
rect 1046 137 1112 175
rect 1046 103 1062 137
rect 1096 103 1112 137
rect 1046 65 1112 103
rect -962 9 -896 31
rect 1046 31 1062 65
rect 1096 31 1112 65
rect 1046 9 1112 31
rect -1140 -581 -1116 -547
rect -1082 -581 -1058 -547
rect -1140 -619 -1058 -581
rect -1140 -653 -1116 -619
rect -1082 -653 -1058 -619
rect 1208 -547 1290 6547
rect 1208 -581 1232 -547
rect 1266 -581 1290 -547
rect 1208 -619 1290 -581
rect -1140 -691 -1058 -653
rect -1140 -725 -1116 -691
rect -1082 -725 -1058 -691
rect -1140 -763 -1058 -725
rect -1140 -797 -1116 -763
rect -1082 -797 -1058 -763
rect -1140 -835 -1058 -797
rect -1140 -869 -1116 -835
rect -1082 -869 -1058 -835
rect -296 -659 460 -643
rect -296 -693 -280 -659
rect -246 -693 -206 -659
rect -172 -693 -132 -659
rect -98 -693 -58 -659
rect -24 -693 16 -659
rect 50 -693 90 -659
rect 124 -693 164 -659
rect 198 -693 238 -659
rect 272 -693 312 -659
rect 346 -693 386 -659
rect 420 -693 460 -659
rect -296 -733 460 -693
rect -296 -767 -280 -733
rect -246 -767 -206 -733
rect -172 -767 -132 -733
rect -98 -767 -58 -733
rect -24 -767 16 -733
rect 50 -767 90 -733
rect 124 -767 164 -733
rect 198 -767 238 -733
rect 272 -767 312 -733
rect 346 -767 386 -733
rect 420 -767 460 -733
rect -296 -857 460 -767
rect 1208 -653 1232 -619
rect 1266 -653 1290 -619
rect 1208 -691 1290 -653
rect 1208 -725 1232 -691
rect 1266 -725 1290 -691
rect 1208 -763 1290 -725
rect 1208 -797 1232 -763
rect 1266 -797 1290 -763
rect 1208 -835 1290 -797
rect -1140 -907 -1058 -869
rect -1140 -941 -1116 -907
rect -1082 -941 -1058 -907
rect -1140 -979 -1058 -941
rect -1140 -1013 -1116 -979
rect -1082 -1013 -1058 -979
rect -1140 -1051 -1058 -1013
rect -1140 -1085 -1116 -1051
rect -1082 -1085 -1058 -1051
rect -1140 -1100 -1058 -1085
rect 1208 -869 1232 -835
rect 1266 -869 1290 -835
rect 1208 -907 1290 -869
rect 1208 -941 1232 -907
rect 1266 -941 1290 -907
rect 1208 -979 1290 -941
rect 1208 -1013 1232 -979
rect 1266 -1013 1290 -979
rect 1208 -1051 1290 -1013
rect 1208 -1085 1232 -1051
rect 1266 -1085 1290 -1051
rect 1208 -1100 1290 -1085
rect -1140 -1124 1290 -1100
rect -1140 -1158 -986 -1124
rect -952 -1158 -914 -1124
rect -880 -1158 -842 -1124
rect -808 -1158 -770 -1124
rect -736 -1158 -698 -1124
rect -664 -1158 -626 -1124
rect -592 -1158 -554 -1124
rect -520 -1158 -482 -1124
rect -448 -1158 -410 -1124
rect -376 -1158 -338 -1124
rect -304 -1158 -266 -1124
rect -232 -1158 -194 -1124
rect -160 -1158 -122 -1124
rect -88 -1158 -50 -1124
rect -16 -1158 22 -1124
rect 56 -1158 94 -1124
rect 128 -1158 166 -1124
rect 200 -1158 238 -1124
rect 272 -1158 310 -1124
rect 344 -1158 382 -1124
rect 416 -1158 454 -1124
rect 488 -1158 526 -1124
rect 560 -1158 598 -1124
rect 632 -1158 670 -1124
rect 704 -1158 742 -1124
rect 776 -1158 814 -1124
rect 848 -1158 886 -1124
rect 920 -1158 958 -1124
rect 992 -1158 1030 -1124
rect 1064 -1158 1102 -1124
rect 1136 -1158 1290 -1124
rect -1140 -1182 1290 -1158
<< viali >>
rect -986 7124 -952 7158
rect -914 7124 -880 7158
rect -842 7124 -808 7158
rect -770 7124 -736 7158
rect -698 7124 -664 7158
rect -626 7124 -592 7158
rect -554 7124 -520 7158
rect -482 7124 -448 7158
rect -410 7124 -376 7158
rect -338 7124 -304 7158
rect -266 7124 -232 7158
rect -194 7124 -160 7158
rect -122 7124 -88 7158
rect -50 7124 -16 7158
rect 22 7124 56 7158
rect 94 7124 128 7158
rect 166 7124 200 7158
rect 238 7124 272 7158
rect 310 7124 344 7158
rect 382 7124 416 7158
rect 454 7124 488 7158
rect 526 7124 560 7158
rect 598 7124 632 7158
rect 670 7124 704 7158
rect 742 7124 776 7158
rect 814 7124 848 7158
rect 886 7124 920 7158
rect 958 7124 992 7158
rect 1030 7124 1064 7158
rect 1102 7124 1136 7158
rect -1116 7051 -1082 7085
rect -1116 6979 -1082 7013
rect -1116 6907 -1082 6941
rect -1116 6835 -1082 6869
rect -1116 6763 -1082 6797
rect -1116 6691 -1082 6725
rect -1116 6619 -1082 6653
rect -1116 6547 -1082 6581
rect 1232 7051 1266 7085
rect 1232 6979 1266 7013
rect 1232 6907 1266 6941
rect 1232 6835 1266 6869
rect 1232 6763 1266 6797
rect 1232 6691 1266 6725
rect 1232 6619 1266 6653
rect 1232 6547 1266 6581
rect -946 5935 -912 5969
rect -946 5863 -912 5897
rect -946 5791 -912 5825
rect -946 5719 -912 5753
rect -946 5647 -912 5681
rect -946 5575 -912 5609
rect -946 5503 -912 5537
rect -946 5431 -912 5465
rect -946 5359 -912 5393
rect -946 5287 -912 5321
rect -946 5215 -912 5249
rect -946 5143 -912 5177
rect -946 5071 -912 5105
rect -946 4999 -912 5033
rect -946 4927 -912 4961
rect -946 4855 -912 4889
rect -946 4783 -912 4817
rect -946 4711 -912 4745
rect -946 4639 -912 4673
rect -946 4567 -912 4601
rect -946 4495 -912 4529
rect -946 4423 -912 4457
rect -946 4351 -912 4385
rect -946 4279 -912 4313
rect -946 4207 -912 4241
rect -946 4135 -912 4169
rect -946 4063 -912 4097
rect -946 3991 -912 4025
rect -946 3919 -912 3953
rect -946 3847 -912 3881
rect -946 3775 -912 3809
rect -946 3703 -912 3737
rect -946 3631 -912 3665
rect -946 3559 -912 3593
rect -946 3487 -912 3521
rect -946 3415 -912 3449
rect -946 3343 -912 3377
rect -946 3271 -912 3305
rect -946 3199 -912 3233
rect -946 3127 -912 3161
rect -946 3055 -912 3089
rect -946 2983 -912 3017
rect -946 2911 -912 2945
rect -946 2839 -912 2873
rect -946 2767 -912 2801
rect -946 2695 -912 2729
rect -946 2623 -912 2657
rect -946 2551 -912 2585
rect -946 2479 -912 2513
rect -946 2407 -912 2441
rect -946 2335 -912 2369
rect -946 2263 -912 2297
rect -946 2191 -912 2225
rect -946 2119 -912 2153
rect -946 2047 -912 2081
rect -946 1975 -912 2009
rect -946 1903 -912 1937
rect -946 1831 -912 1865
rect -946 1759 -912 1793
rect -946 1687 -912 1721
rect -946 1615 -912 1649
rect -946 1543 -912 1577
rect -946 1471 -912 1505
rect -946 1399 -912 1433
rect -946 1327 -912 1361
rect -946 1255 -912 1289
rect -946 1183 -912 1217
rect -946 1111 -912 1145
rect -946 1039 -912 1073
rect -946 967 -912 1001
rect -946 895 -912 929
rect -946 823 -912 857
rect -946 751 -912 785
rect -946 679 -912 713
rect -946 607 -912 641
rect -946 535 -912 569
rect -946 463 -912 497
rect -946 391 -912 425
rect -946 319 -912 353
rect -946 247 -912 281
rect -946 175 -912 209
rect -946 103 -912 137
rect -946 31 -912 65
rect 22 67 128 5933
rect 1062 5935 1096 5969
rect 1062 5863 1096 5897
rect 1062 5791 1096 5825
rect 1062 5719 1096 5753
rect 1062 5647 1096 5681
rect 1062 5575 1096 5609
rect 1062 5503 1096 5537
rect 1062 5431 1096 5465
rect 1062 5359 1096 5393
rect 1062 5287 1096 5321
rect 1062 5215 1096 5249
rect 1062 5143 1096 5177
rect 1062 5071 1096 5105
rect 1062 4999 1096 5033
rect 1062 4927 1096 4961
rect 1062 4855 1096 4889
rect 1062 4783 1096 4817
rect 1062 4711 1096 4745
rect 1062 4639 1096 4673
rect 1062 4567 1096 4601
rect 1062 4495 1096 4529
rect 1062 4423 1096 4457
rect 1062 4351 1096 4385
rect 1062 4279 1096 4313
rect 1062 4207 1096 4241
rect 1062 4135 1096 4169
rect 1062 4063 1096 4097
rect 1062 3991 1096 4025
rect 1062 3919 1096 3953
rect 1062 3847 1096 3881
rect 1062 3775 1096 3809
rect 1062 3703 1096 3737
rect 1062 3631 1096 3665
rect 1062 3559 1096 3593
rect 1062 3487 1096 3521
rect 1062 3415 1096 3449
rect 1062 3343 1096 3377
rect 1062 3271 1096 3305
rect 1062 3199 1096 3233
rect 1062 3127 1096 3161
rect 1062 3055 1096 3089
rect 1062 2983 1096 3017
rect 1062 2911 1096 2945
rect 1062 2839 1096 2873
rect 1062 2767 1096 2801
rect 1062 2695 1096 2729
rect 1062 2623 1096 2657
rect 1062 2551 1096 2585
rect 1062 2479 1096 2513
rect 1062 2407 1096 2441
rect 1062 2335 1096 2369
rect 1062 2263 1096 2297
rect 1062 2191 1096 2225
rect 1062 2119 1096 2153
rect 1062 2047 1096 2081
rect 1062 1975 1096 2009
rect 1062 1903 1096 1937
rect 1062 1831 1096 1865
rect 1062 1759 1096 1793
rect 1062 1687 1096 1721
rect 1062 1615 1096 1649
rect 1062 1543 1096 1577
rect 1062 1471 1096 1505
rect 1062 1399 1096 1433
rect 1062 1327 1096 1361
rect 1062 1255 1096 1289
rect 1062 1183 1096 1217
rect 1062 1111 1096 1145
rect 1062 1039 1096 1073
rect 1062 967 1096 1001
rect 1062 895 1096 929
rect 1062 823 1096 857
rect 1062 751 1096 785
rect 1062 679 1096 713
rect 1062 607 1096 641
rect 1062 535 1096 569
rect 1062 463 1096 497
rect 1062 391 1096 425
rect 1062 319 1096 353
rect 1062 247 1096 281
rect 1062 175 1096 209
rect 1062 103 1096 137
rect 1062 31 1096 65
rect -1116 -581 -1082 -547
rect -1116 -653 -1082 -619
rect 1232 -581 1266 -547
rect -1116 -725 -1082 -691
rect -1116 -797 -1082 -763
rect -1116 -869 -1082 -835
rect -280 -693 -246 -659
rect -206 -693 -172 -659
rect -132 -693 -98 -659
rect -58 -693 -24 -659
rect 16 -693 50 -659
rect 90 -693 124 -659
rect 164 -693 198 -659
rect 238 -693 272 -659
rect 312 -693 346 -659
rect 386 -693 420 -659
rect -280 -767 -246 -733
rect -206 -767 -172 -733
rect -132 -767 -98 -733
rect -58 -767 -24 -733
rect 16 -767 50 -733
rect 90 -767 124 -733
rect 164 -767 198 -733
rect 238 -767 272 -733
rect 312 -767 346 -733
rect 386 -767 420 -733
rect 1232 -653 1266 -619
rect 1232 -725 1266 -691
rect 1232 -797 1266 -763
rect -1116 -941 -1082 -907
rect -1116 -1013 -1082 -979
rect -1116 -1085 -1082 -1051
rect 1232 -869 1266 -835
rect 1232 -941 1266 -907
rect 1232 -1013 1266 -979
rect 1232 -1085 1266 -1051
rect -986 -1158 -952 -1124
rect -914 -1158 -880 -1124
rect -842 -1158 -808 -1124
rect -770 -1158 -736 -1124
rect -698 -1158 -664 -1124
rect -626 -1158 -592 -1124
rect -554 -1158 -520 -1124
rect -482 -1158 -448 -1124
rect -410 -1158 -376 -1124
rect -338 -1158 -304 -1124
rect -266 -1158 -232 -1124
rect -194 -1158 -160 -1124
rect -122 -1158 -88 -1124
rect -50 -1158 -16 -1124
rect 22 -1158 56 -1124
rect 94 -1158 128 -1124
rect 166 -1158 200 -1124
rect 238 -1158 272 -1124
rect 310 -1158 344 -1124
rect 382 -1158 416 -1124
rect 454 -1158 488 -1124
rect 526 -1158 560 -1124
rect 598 -1158 632 -1124
rect 670 -1158 704 -1124
rect 742 -1158 776 -1124
rect 814 -1158 848 -1124
rect 886 -1158 920 -1124
rect 958 -1158 992 -1124
rect 1030 -1158 1064 -1124
rect 1102 -1158 1136 -1124
<< metal1 >>
rect -1140 7158 1290 7182
rect -1140 7124 -986 7158
rect -952 7124 -914 7158
rect -880 7124 -842 7158
rect -808 7124 -770 7158
rect -736 7124 -698 7158
rect -664 7124 -626 7158
rect -592 7124 -554 7158
rect -520 7124 -482 7158
rect -448 7124 -410 7158
rect -376 7124 -338 7158
rect -304 7124 -266 7158
rect -232 7124 -194 7158
rect -160 7124 -122 7158
rect -88 7124 -50 7158
rect -16 7124 22 7158
rect 56 7124 94 7158
rect 128 7124 166 7158
rect 200 7124 238 7158
rect 272 7124 310 7158
rect 344 7124 382 7158
rect 416 7124 454 7158
rect 488 7124 526 7158
rect 560 7124 598 7158
rect 632 7124 670 7158
rect 704 7124 742 7158
rect 776 7124 814 7158
rect 848 7124 886 7158
rect 920 7124 958 7158
rect 992 7124 1030 7158
rect 1064 7124 1102 7158
rect 1136 7124 1290 7158
rect -1140 7100 1290 7124
rect -1140 7085 -492 7100
tri -492 7085 -477 7100 nw
tri 627 7085 642 7100 ne
rect 642 7085 1290 7100
rect -1140 7051 -1116 7085
rect -1082 7051 -526 7085
tri -526 7051 -492 7085 nw
tri 642 7051 676 7085 ne
rect 676 7051 1232 7085
rect 1266 7051 1290 7085
rect -1140 7013 -564 7051
tri -564 7013 -526 7051 nw
tri 676 7013 714 7051 ne
rect 714 7013 1290 7051
rect -1140 6979 -1116 7013
rect -1082 6979 -598 7013
tri -598 6979 -564 7013 nw
tri 714 6979 748 7013 ne
rect 748 6979 1232 7013
rect 1266 6979 1290 7013
rect -1140 6941 -636 6979
tri -636 6941 -598 6979 nw
tri 748 6941 786 6979 ne
rect 786 6941 1290 6979
rect -1140 6907 -1116 6941
rect -1082 6907 -670 6941
tri -670 6907 -636 6941 nw
tri 786 6907 820 6941 ne
rect 820 6907 1232 6941
rect 1266 6907 1290 6941
rect -1140 6869 -708 6907
tri -708 6869 -670 6907 nw
tri 820 6869 858 6907 ne
rect 858 6869 1290 6907
rect -1140 6835 -1116 6869
rect -1082 6835 -742 6869
tri -742 6835 -708 6869 nw
tri 858 6835 892 6869 ne
rect 892 6835 1232 6869
rect 1266 6835 1290 6869
rect -1140 6797 -780 6835
tri -780 6797 -742 6835 nw
tri 892 6797 930 6835 ne
rect 930 6797 1290 6835
rect -1140 6763 -1116 6797
rect -1082 6763 -814 6797
tri -814 6763 -780 6797 nw
tri 930 6763 964 6797 ne
rect 964 6763 1232 6797
rect 1266 6763 1290 6797
rect -1140 6725 -852 6763
tri -852 6725 -814 6763 nw
tri 964 6725 1002 6763 ne
rect 1002 6725 1290 6763
rect -1140 6691 -1116 6725
rect -1082 6691 -886 6725
tri -886 6691 -852 6725 nw
tri 1002 6691 1036 6725 ne
rect 1036 6691 1232 6725
rect 1266 6691 1290 6725
rect -1140 6653 -924 6691
tri -924 6653 -886 6691 nw
tri 1036 6653 1074 6691 ne
rect 1074 6653 1290 6691
rect -1140 6619 -1116 6653
rect -1082 6619 -958 6653
tri -958 6619 -924 6653 nw
tri 1074 6619 1108 6653 ne
rect 1108 6619 1232 6653
rect 1266 6619 1290 6653
rect -1140 6581 -996 6619
tri -996 6581 -958 6619 nw
tri 1108 6581 1146 6619 ne
rect 1146 6581 1290 6619
rect -1140 6547 -1116 6581
rect -1082 6547 -1030 6581
tri -1030 6547 -996 6581 nw
tri 1146 6547 1180 6581 ne
rect 1180 6547 1232 6581
rect 1266 6547 1290 6581
rect -1140 6519 -1058 6547
tri -1058 6519 -1030 6547 nw
tri 1180 6519 1208 6547 ne
rect 1208 6519 1290 6547
rect -958 5969 -900 5981
rect -958 5935 -946 5969
rect -912 5935 -900 5969
rect 1050 5969 1108 5981
rect -958 5897 -900 5935
rect -958 5863 -946 5897
rect -912 5863 -900 5897
rect -958 5825 -900 5863
rect -958 5791 -946 5825
rect -912 5791 -900 5825
rect -958 5753 -900 5791
rect -958 5719 -946 5753
rect -912 5719 -900 5753
rect -958 5681 -900 5719
rect -958 5647 -946 5681
rect -912 5647 -900 5681
rect -958 5609 -900 5647
rect -958 5575 -946 5609
rect -912 5575 -900 5609
rect -958 5537 -900 5575
rect -958 5503 -946 5537
rect -912 5503 -900 5537
rect -958 5465 -900 5503
rect -958 5431 -946 5465
rect -912 5431 -900 5465
rect -958 5393 -900 5431
rect -958 5359 -946 5393
rect -912 5359 -900 5393
rect -958 5321 -900 5359
rect -958 5287 -946 5321
rect -912 5287 -900 5321
rect -958 5249 -900 5287
rect -958 5215 -946 5249
rect -912 5215 -900 5249
rect -958 5177 -900 5215
rect -958 5143 -946 5177
rect -912 5143 -900 5177
rect -958 5105 -900 5143
rect -958 5071 -946 5105
rect -912 5071 -900 5105
rect -958 5033 -900 5071
rect -958 4999 -946 5033
rect -912 4999 -900 5033
rect -958 4961 -900 4999
rect -958 4927 -946 4961
rect -912 4927 -900 4961
rect -958 4889 -900 4927
rect -958 4855 -946 4889
rect -912 4855 -900 4889
rect -958 4817 -900 4855
rect -958 4783 -946 4817
rect -912 4783 -900 4817
rect -958 4745 -900 4783
rect -958 4711 -946 4745
rect -912 4711 -900 4745
rect -958 4673 -900 4711
rect -958 4639 -946 4673
rect -912 4639 -900 4673
rect -958 4601 -900 4639
rect -958 4567 -946 4601
rect -912 4567 -900 4601
rect -958 4529 -900 4567
rect -958 4495 -946 4529
rect -912 4495 -900 4529
rect -958 4457 -900 4495
rect -958 4423 -946 4457
rect -912 4423 -900 4457
rect -958 4385 -900 4423
rect -958 4351 -946 4385
rect -912 4351 -900 4385
rect -958 4313 -900 4351
rect -958 4279 -946 4313
rect -912 4279 -900 4313
rect -958 4241 -900 4279
rect -958 4207 -946 4241
rect -912 4207 -900 4241
rect -958 4169 -900 4207
rect -958 4135 -946 4169
rect -912 4135 -900 4169
rect -958 4097 -900 4135
rect -958 4063 -946 4097
rect -912 4063 -900 4097
rect -958 4025 -900 4063
rect -958 3991 -946 4025
rect -912 3991 -900 4025
rect -958 3953 -900 3991
rect -958 3919 -946 3953
rect -912 3919 -900 3953
rect -958 3881 -900 3919
rect -958 3847 -946 3881
rect -912 3847 -900 3881
rect -958 3809 -900 3847
rect -958 3775 -946 3809
rect -912 3775 -900 3809
rect -958 3737 -900 3775
rect -958 3703 -946 3737
rect -912 3703 -900 3737
rect -958 3665 -900 3703
rect -958 3631 -946 3665
rect -912 3631 -900 3665
rect -958 3593 -900 3631
rect -958 3559 -946 3593
rect -912 3559 -900 3593
rect -958 3521 -900 3559
rect -958 3487 -946 3521
rect -912 3487 -900 3521
rect -958 3449 -900 3487
rect -958 3415 -946 3449
rect -912 3415 -900 3449
rect -958 3377 -900 3415
rect -958 3343 -946 3377
rect -912 3343 -900 3377
rect -958 3305 -900 3343
rect -958 3271 -946 3305
rect -912 3271 -900 3305
rect -958 3233 -900 3271
rect -958 3199 -946 3233
rect -912 3199 -900 3233
rect -958 3161 -900 3199
rect -958 3127 -946 3161
rect -912 3127 -900 3161
rect -958 3089 -900 3127
rect -958 3055 -946 3089
rect -912 3055 -900 3089
rect -958 3017 -900 3055
rect -958 2983 -946 3017
rect -912 2983 -900 3017
rect -958 2945 -900 2983
rect -958 2911 -946 2945
rect -912 2911 -900 2945
rect -958 2873 -900 2911
rect -958 2839 -946 2873
rect -912 2839 -900 2873
rect -958 2801 -900 2839
rect -958 2767 -946 2801
rect -912 2767 -900 2801
rect -958 2729 -900 2767
rect -958 2695 -946 2729
rect -912 2695 -900 2729
rect -958 2657 -900 2695
rect -958 2623 -946 2657
rect -912 2623 -900 2657
rect -958 2585 -900 2623
rect -958 2551 -946 2585
rect -912 2551 -900 2585
rect -958 2513 -900 2551
rect -958 2479 -946 2513
rect -912 2479 -900 2513
rect -958 2441 -900 2479
rect -958 2407 -946 2441
rect -912 2407 -900 2441
rect -958 2369 -900 2407
rect -958 2335 -946 2369
rect -912 2335 -900 2369
rect -958 2297 -900 2335
rect -958 2263 -946 2297
rect -912 2263 -900 2297
rect -958 2225 -900 2263
rect -958 2191 -946 2225
rect -912 2191 -900 2225
rect -958 2153 -900 2191
rect -958 2119 -946 2153
rect -912 2119 -900 2153
rect -958 2081 -900 2119
rect -958 2047 -946 2081
rect -912 2047 -900 2081
rect -958 2009 -900 2047
rect -958 1975 -946 2009
rect -912 1975 -900 2009
rect -958 1937 -900 1975
rect -958 1903 -946 1937
rect -912 1903 -900 1937
rect -958 1865 -900 1903
rect -958 1831 -946 1865
rect -912 1831 -900 1865
rect -958 1793 -900 1831
rect -958 1759 -946 1793
rect -912 1759 -900 1793
rect -958 1721 -900 1759
rect -958 1687 -946 1721
rect -912 1687 -900 1721
rect -958 1649 -900 1687
rect -958 1615 -946 1649
rect -912 1615 -900 1649
rect -958 1577 -900 1615
rect -958 1543 -946 1577
rect -912 1543 -900 1577
rect -958 1505 -900 1543
rect -958 1471 -946 1505
rect -912 1471 -900 1505
rect -958 1433 -900 1471
rect -958 1399 -946 1433
rect -912 1399 -900 1433
rect -958 1361 -900 1399
rect -958 1327 -946 1361
rect -912 1327 -900 1361
rect -958 1289 -900 1327
rect -958 1255 -946 1289
rect -912 1255 -900 1289
rect -958 1217 -900 1255
rect -958 1183 -946 1217
rect -912 1183 -900 1217
rect -958 1145 -900 1183
rect -958 1111 -946 1145
rect -912 1111 -900 1145
rect -958 1073 -900 1111
rect -958 1039 -946 1073
rect -912 1039 -900 1073
rect -958 1001 -900 1039
rect -958 967 -946 1001
rect -912 967 -900 1001
rect -958 929 -900 967
rect -958 895 -946 929
rect -912 895 -900 929
rect -958 857 -900 895
rect -958 823 -946 857
rect -912 823 -900 857
rect -958 785 -900 823
rect -958 751 -946 785
rect -912 751 -900 785
rect -958 713 -900 751
rect -958 679 -946 713
rect -912 679 -900 713
rect -958 641 -900 679
rect -958 607 -946 641
rect -912 607 -900 641
rect -958 569 -900 607
rect -958 535 -946 569
rect -912 535 -900 569
rect -958 497 -900 535
rect -958 463 -946 497
rect -912 463 -900 497
rect -958 425 -900 463
rect -958 391 -946 425
rect -912 391 -900 425
rect -958 353 -900 391
rect -958 319 -946 353
rect -912 319 -900 353
rect -958 281 -900 319
rect -958 247 -946 281
rect -912 247 -900 281
rect -958 209 -900 247
rect -958 175 -946 209
rect -912 175 -900 209
rect -958 137 -900 175
rect -958 103 -946 137
rect -912 103 -900 137
rect -958 65 -900 103
rect -958 31 -946 65
rect -912 31 -900 65
rect 10 5939 140 5945
rect 10 63 17 5939
rect 133 63 140 5939
rect 10 55 140 63
rect 1050 5935 1062 5969
rect 1096 5935 1108 5969
rect 1050 5897 1108 5935
rect 1050 5863 1062 5897
rect 1096 5863 1108 5897
rect 1050 5825 1108 5863
rect 1050 5791 1062 5825
rect 1096 5791 1108 5825
rect 1050 5753 1108 5791
rect 1050 5719 1062 5753
rect 1096 5719 1108 5753
rect 1050 5681 1108 5719
rect 1050 5647 1062 5681
rect 1096 5647 1108 5681
rect 1050 5609 1108 5647
rect 1050 5575 1062 5609
rect 1096 5575 1108 5609
rect 1050 5537 1108 5575
rect 1050 5503 1062 5537
rect 1096 5503 1108 5537
rect 1050 5465 1108 5503
rect 1050 5431 1062 5465
rect 1096 5431 1108 5465
rect 1050 5393 1108 5431
rect 1050 5359 1062 5393
rect 1096 5359 1108 5393
rect 1050 5321 1108 5359
rect 1050 5287 1062 5321
rect 1096 5287 1108 5321
rect 1050 5249 1108 5287
rect 1050 5215 1062 5249
rect 1096 5215 1108 5249
rect 1050 5177 1108 5215
rect 1050 5143 1062 5177
rect 1096 5143 1108 5177
rect 1050 5105 1108 5143
rect 1050 5071 1062 5105
rect 1096 5071 1108 5105
rect 1050 5033 1108 5071
rect 1050 4999 1062 5033
rect 1096 4999 1108 5033
rect 1050 4961 1108 4999
rect 1050 4927 1062 4961
rect 1096 4927 1108 4961
rect 1050 4889 1108 4927
rect 1050 4855 1062 4889
rect 1096 4855 1108 4889
rect 1050 4817 1108 4855
rect 1050 4783 1062 4817
rect 1096 4783 1108 4817
rect 1050 4745 1108 4783
rect 1050 4711 1062 4745
rect 1096 4711 1108 4745
rect 1050 4673 1108 4711
rect 1050 4639 1062 4673
rect 1096 4639 1108 4673
rect 1050 4601 1108 4639
rect 1050 4567 1062 4601
rect 1096 4567 1108 4601
rect 1050 4529 1108 4567
rect 1050 4495 1062 4529
rect 1096 4495 1108 4529
rect 1050 4457 1108 4495
rect 1050 4423 1062 4457
rect 1096 4423 1108 4457
rect 1050 4385 1108 4423
rect 1050 4351 1062 4385
rect 1096 4351 1108 4385
rect 1050 4313 1108 4351
rect 1050 4279 1062 4313
rect 1096 4279 1108 4313
rect 1050 4241 1108 4279
rect 1050 4207 1062 4241
rect 1096 4207 1108 4241
rect 1050 4169 1108 4207
rect 1050 4135 1062 4169
rect 1096 4135 1108 4169
rect 1050 4097 1108 4135
rect 1050 4063 1062 4097
rect 1096 4063 1108 4097
rect 1050 4025 1108 4063
rect 1050 3991 1062 4025
rect 1096 3991 1108 4025
rect 1050 3953 1108 3991
rect 1050 3919 1062 3953
rect 1096 3919 1108 3953
rect 1050 3881 1108 3919
rect 1050 3847 1062 3881
rect 1096 3847 1108 3881
rect 1050 3809 1108 3847
rect 1050 3775 1062 3809
rect 1096 3775 1108 3809
rect 1050 3737 1108 3775
rect 1050 3703 1062 3737
rect 1096 3703 1108 3737
rect 1050 3665 1108 3703
rect 1050 3631 1062 3665
rect 1096 3631 1108 3665
rect 1050 3593 1108 3631
rect 1050 3559 1062 3593
rect 1096 3559 1108 3593
rect 1050 3521 1108 3559
rect 1050 3487 1062 3521
rect 1096 3487 1108 3521
rect 1050 3449 1108 3487
rect 1050 3415 1062 3449
rect 1096 3415 1108 3449
rect 1050 3377 1108 3415
rect 1050 3343 1062 3377
rect 1096 3343 1108 3377
rect 1050 3305 1108 3343
rect 1050 3271 1062 3305
rect 1096 3271 1108 3305
rect 1050 3233 1108 3271
rect 1050 3199 1062 3233
rect 1096 3199 1108 3233
rect 1050 3161 1108 3199
rect 1050 3127 1062 3161
rect 1096 3127 1108 3161
rect 1050 3089 1108 3127
rect 1050 3055 1062 3089
rect 1096 3055 1108 3089
rect 1050 3017 1108 3055
rect 1050 2983 1062 3017
rect 1096 2983 1108 3017
rect 1050 2945 1108 2983
rect 1050 2911 1062 2945
rect 1096 2911 1108 2945
rect 1050 2873 1108 2911
rect 1050 2839 1062 2873
rect 1096 2839 1108 2873
rect 1050 2801 1108 2839
rect 1050 2767 1062 2801
rect 1096 2767 1108 2801
rect 1050 2729 1108 2767
rect 1050 2695 1062 2729
rect 1096 2695 1108 2729
rect 1050 2657 1108 2695
rect 1050 2623 1062 2657
rect 1096 2623 1108 2657
rect 1050 2585 1108 2623
rect 1050 2551 1062 2585
rect 1096 2551 1108 2585
rect 1050 2513 1108 2551
rect 1050 2479 1062 2513
rect 1096 2479 1108 2513
rect 1050 2441 1108 2479
rect 1050 2407 1062 2441
rect 1096 2407 1108 2441
rect 1050 2369 1108 2407
rect 1050 2335 1062 2369
rect 1096 2335 1108 2369
rect 1050 2297 1108 2335
rect 1050 2263 1062 2297
rect 1096 2263 1108 2297
rect 1050 2225 1108 2263
rect 1050 2191 1062 2225
rect 1096 2191 1108 2225
rect 1050 2153 1108 2191
rect 1050 2119 1062 2153
rect 1096 2119 1108 2153
rect 1050 2081 1108 2119
rect 1050 2047 1062 2081
rect 1096 2047 1108 2081
rect 1050 2009 1108 2047
rect 1050 1975 1062 2009
rect 1096 1975 1108 2009
rect 1050 1937 1108 1975
rect 1050 1903 1062 1937
rect 1096 1903 1108 1937
rect 1050 1865 1108 1903
rect 1050 1831 1062 1865
rect 1096 1831 1108 1865
rect 1050 1793 1108 1831
rect 1050 1759 1062 1793
rect 1096 1759 1108 1793
rect 1050 1721 1108 1759
rect 1050 1687 1062 1721
rect 1096 1687 1108 1721
rect 1050 1649 1108 1687
rect 1050 1615 1062 1649
rect 1096 1615 1108 1649
rect 1050 1577 1108 1615
rect 1050 1543 1062 1577
rect 1096 1543 1108 1577
rect 1050 1505 1108 1543
rect 1050 1471 1062 1505
rect 1096 1471 1108 1505
rect 1050 1433 1108 1471
rect 1050 1399 1062 1433
rect 1096 1399 1108 1433
rect 1050 1361 1108 1399
rect 1050 1327 1062 1361
rect 1096 1327 1108 1361
rect 1050 1289 1108 1327
rect 1050 1255 1062 1289
rect 1096 1255 1108 1289
rect 1050 1217 1108 1255
rect 1050 1183 1062 1217
rect 1096 1183 1108 1217
rect 1050 1145 1108 1183
rect 1050 1111 1062 1145
rect 1096 1111 1108 1145
rect 1050 1073 1108 1111
rect 1050 1039 1062 1073
rect 1096 1039 1108 1073
rect 1050 1001 1108 1039
rect 1050 967 1062 1001
rect 1096 967 1108 1001
rect 1050 929 1108 967
rect 1050 895 1062 929
rect 1096 895 1108 929
rect 1050 857 1108 895
rect 1050 823 1062 857
rect 1096 823 1108 857
rect 1050 785 1108 823
rect 1050 751 1062 785
rect 1096 751 1108 785
rect 1050 713 1108 751
rect 1050 679 1062 713
rect 1096 679 1108 713
rect 1050 641 1108 679
rect 1050 607 1062 641
rect 1096 607 1108 641
rect 1050 569 1108 607
rect 1050 535 1062 569
rect 1096 535 1108 569
rect 1050 497 1108 535
rect 1050 463 1062 497
rect 1096 463 1108 497
rect 1050 425 1108 463
rect 1050 391 1062 425
rect 1096 391 1108 425
rect 1050 353 1108 391
rect 1050 319 1062 353
rect 1096 319 1108 353
rect 1050 281 1108 319
rect 1050 247 1062 281
rect 1096 247 1108 281
rect 1050 209 1108 247
rect 1050 175 1062 209
rect 1096 175 1108 209
rect 1050 137 1108 175
rect 1050 103 1062 137
rect 1096 103 1108 137
rect 1050 65 1108 103
rect -958 19 -900 31
rect 1050 31 1062 65
rect 1096 31 1108 65
rect 1050 19 1108 31
rect -1140 -547 -1058 -519
tri -1058 -547 -1030 -519 sw
tri 1180 -547 1208 -519 se
rect 1208 -547 1290 -519
rect -1140 -581 -1116 -547
rect -1082 -581 -1030 -547
tri -1030 -581 -996 -547 sw
tri 1146 -581 1180 -547 se
rect 1180 -581 1232 -547
rect 1266 -581 1290 -547
rect -1140 -619 -996 -581
tri -996 -619 -958 -581 sw
tri 1108 -619 1146 -581 se
rect 1146 -619 1290 -581
rect -1140 -653 -1116 -619
rect -1082 -643 -958 -619
tri -958 -643 -934 -619 sw
tri 1084 -643 1108 -619 se
rect 1108 -643 1232 -619
rect -1082 -653 -934 -643
tri -934 -653 -924 -643 sw
rect -296 -650 460 -643
rect -1140 -659 -924 -653
tri -924 -659 -918 -653 sw
rect -1140 -691 -918 -659
rect -1140 -725 -1116 -691
rect -1082 -693 -918 -691
tri -918 -693 -884 -659 sw
rect -1082 -725 -884 -693
tri -884 -725 -852 -693 sw
rect -296 -702 -289 -650
rect -237 -702 -215 -650
rect -163 -702 -141 -650
rect -89 -702 -67 -650
rect -15 -702 7 -650
rect 59 -702 81 -650
rect 133 -702 155 -650
rect 207 -702 229 -650
rect 281 -702 303 -650
rect 355 -702 377 -650
rect 429 -702 460 -650
tri 1074 -653 1084 -643 se
rect 1084 -653 1232 -643
rect 1266 -653 1290 -619
tri 1036 -691 1074 -653 se
rect 1074 -691 1290 -653
rect -296 -724 460 -702
rect -1140 -733 -852 -725
tri -852 -733 -844 -725 sw
rect -1140 -763 -844 -733
rect -1140 -797 -1116 -763
rect -1082 -767 -844 -763
tri -844 -767 -810 -733 sw
rect -1082 -785 -810 -767
tri -810 -785 -792 -767 sw
rect -296 -776 -289 -724
rect -237 -776 -215 -724
rect -163 -776 -141 -724
rect -89 -776 -67 -724
rect -15 -776 7 -724
rect 59 -776 81 -724
rect 133 -776 155 -724
rect 207 -776 229 -724
rect 281 -776 303 -724
rect 355 -776 377 -724
rect 429 -776 460 -724
tri 1002 -725 1036 -691 se
rect 1036 -725 1232 -691
rect 1266 -725 1290 -691
tri 964 -763 1002 -725 se
rect 1002 -763 1290 -725
rect -296 -785 460 -776
tri 942 -785 964 -763 se
rect 964 -785 1232 -763
rect -1082 -797 -792 -785
tri -792 -797 -780 -785 sw
tri 930 -797 942 -785 se
rect 942 -797 1232 -785
rect 1266 -797 1290 -763
rect -1140 -835 -780 -797
tri -780 -835 -742 -797 sw
tri 892 -835 930 -797 se
rect 930 -835 1290 -797
rect -1140 -869 -1116 -835
rect -1082 -869 -742 -835
tri -742 -869 -708 -835 sw
tri 858 -869 892 -835 se
rect 892 -869 1232 -835
rect 1266 -869 1290 -835
rect -1140 -907 -708 -869
tri -708 -907 -670 -869 sw
tri 820 -907 858 -869 se
rect 858 -907 1290 -869
rect -1140 -941 -1116 -907
rect -1082 -941 -670 -907
tri -670 -941 -636 -907 sw
tri 786 -941 820 -907 se
rect 820 -941 1232 -907
rect 1266 -941 1290 -907
rect -1140 -979 -636 -941
tri -636 -979 -598 -941 sw
tri 748 -979 786 -941 se
rect 786 -979 1290 -941
rect -1140 -1013 -1116 -979
rect -1082 -1013 -598 -979
tri -598 -1013 -564 -979 sw
tri 714 -1013 748 -979 se
rect 748 -1013 1232 -979
rect 1266 -1013 1290 -979
rect -1140 -1051 -564 -1013
tri -564 -1051 -526 -1013 sw
tri 676 -1051 714 -1013 se
rect 714 -1051 1290 -1013
rect -1140 -1085 -1116 -1051
rect -1082 -1085 -526 -1051
tri -526 -1085 -492 -1051 sw
tri 642 -1085 676 -1051 se
rect 676 -1085 1232 -1051
rect 1266 -1085 1290 -1051
rect -1140 -1097 -492 -1085
tri -492 -1097 -480 -1085 sw
tri 630 -1097 642 -1085 se
rect 642 -1097 1290 -1085
rect -1140 -1100 -480 -1097
tri -480 -1100 -477 -1097 sw
tri 627 -1100 630 -1097 se
rect 630 -1100 1290 -1097
rect -1140 -1124 1290 -1100
rect -1140 -1158 -986 -1124
rect -952 -1158 -914 -1124
rect -880 -1158 -842 -1124
rect -808 -1158 -770 -1124
rect -736 -1158 -698 -1124
rect -664 -1158 -626 -1124
rect -592 -1158 -554 -1124
rect -520 -1158 -482 -1124
rect -448 -1158 -410 -1124
rect -376 -1158 -338 -1124
rect -304 -1158 -266 -1124
rect -232 -1158 -194 -1124
rect -160 -1158 -122 -1124
rect -88 -1158 -50 -1124
rect -16 -1158 22 -1124
rect 56 -1158 94 -1124
rect 128 -1158 166 -1124
rect 200 -1158 238 -1124
rect 272 -1158 310 -1124
rect 344 -1158 382 -1124
rect 416 -1158 454 -1124
rect 488 -1158 526 -1124
rect 560 -1158 598 -1124
rect 632 -1158 670 -1124
rect 704 -1158 742 -1124
rect 776 -1158 814 -1124
rect 848 -1158 886 -1124
rect 920 -1158 958 -1124
rect 992 -1158 1030 -1124
rect 1064 -1158 1102 -1124
rect 1136 -1158 1290 -1124
rect -1140 -1182 1290 -1158
<< via1 >>
rect 17 5933 133 5939
rect 17 67 22 5933
rect 22 67 128 5933
rect 128 67 133 5933
rect 17 63 133 67
rect -289 -659 -237 -650
rect -289 -693 -280 -659
rect -280 -693 -246 -659
rect -246 -693 -237 -659
rect -289 -702 -237 -693
rect -215 -659 -163 -650
rect -215 -693 -206 -659
rect -206 -693 -172 -659
rect -172 -693 -163 -659
rect -215 -702 -163 -693
rect -141 -659 -89 -650
rect -141 -693 -132 -659
rect -132 -693 -98 -659
rect -98 -693 -89 -659
rect -141 -702 -89 -693
rect -67 -659 -15 -650
rect -67 -693 -58 -659
rect -58 -693 -24 -659
rect -24 -693 -15 -659
rect -67 -702 -15 -693
rect 7 -659 59 -650
rect 7 -693 16 -659
rect 16 -693 50 -659
rect 50 -693 59 -659
rect 7 -702 59 -693
rect 81 -659 133 -650
rect 81 -693 90 -659
rect 90 -693 124 -659
rect 124 -693 133 -659
rect 81 -702 133 -693
rect 155 -659 207 -650
rect 155 -693 164 -659
rect 164 -693 198 -659
rect 198 -693 207 -659
rect 155 -702 207 -693
rect 229 -659 281 -650
rect 229 -693 238 -659
rect 238 -693 272 -659
rect 272 -693 281 -659
rect 229 -702 281 -693
rect 303 -659 355 -650
rect 303 -693 312 -659
rect 312 -693 346 -659
rect 346 -693 355 -659
rect 303 -702 355 -693
rect 377 -659 429 -650
rect 377 -693 386 -659
rect 386 -693 420 -659
rect 420 -693 429 -659
rect 377 -702 429 -693
rect -289 -733 -237 -724
rect -289 -767 -280 -733
rect -280 -767 -246 -733
rect -246 -767 -237 -733
rect -289 -776 -237 -767
rect -215 -733 -163 -724
rect -215 -767 -206 -733
rect -206 -767 -172 -733
rect -172 -767 -163 -733
rect -215 -776 -163 -767
rect -141 -733 -89 -724
rect -141 -767 -132 -733
rect -132 -767 -98 -733
rect -98 -767 -89 -733
rect -141 -776 -89 -767
rect -67 -733 -15 -724
rect -67 -767 -58 -733
rect -58 -767 -24 -733
rect -24 -767 -15 -733
rect -67 -776 -15 -767
rect 7 -733 59 -724
rect 7 -767 16 -733
rect 16 -767 50 -733
rect 50 -767 59 -733
rect 7 -776 59 -767
rect 81 -733 133 -724
rect 81 -767 90 -733
rect 90 -767 124 -733
rect 124 -767 133 -733
rect 81 -776 133 -767
rect 155 -733 207 -724
rect 155 -767 164 -733
rect 164 -767 198 -733
rect 198 -767 207 -733
rect 155 -776 207 -767
rect 229 -733 281 -724
rect 229 -767 238 -733
rect 238 -767 272 -733
rect 272 -767 281 -733
rect 229 -776 281 -767
rect 303 -733 355 -724
rect 303 -767 312 -733
rect 312 -767 346 -733
rect 346 -767 355 -733
rect 303 -776 355 -767
rect 377 -733 429 -724
rect 377 -767 386 -733
rect 386 -767 420 -733
rect 420 -767 429 -733
rect 377 -776 429 -767
<< metal2 >>
rect 11 5939 139 5945
rect 11 63 17 5939
rect 133 63 139 5939
rect 11 57 139 63
rect -296 -650 460 -643
rect -296 -702 -289 -650
rect -237 -702 -215 -650
rect -163 -702 -141 -650
rect -89 -702 -67 -650
rect -15 -702 7 -650
rect 59 -702 81 -650
rect 133 -702 155 -650
rect 207 -702 229 -650
rect 281 -702 303 -650
rect 355 -702 377 -650
rect 429 -702 460 -650
rect -296 -724 460 -702
rect -296 -776 -289 -724
rect -237 -776 -215 -724
rect -163 -776 -141 -724
rect -89 -776 -67 -724
rect -15 -776 7 -724
rect 59 -776 81 -724
rect 133 -776 155 -724
rect 207 -776 229 -724
rect 281 -776 303 -724
rect 355 -776 377 -724
rect 429 -776 460 -724
rect -296 -857 460 -776
<< labels >>
flabel comment s 1085 159 1085 159 0 FreeSans 2000 0 0 0 S
flabel comment s -925 159 -925 159 0 FreeSans 2000 0 0 0 S
flabel comment s 67 159 67 159 0 FreeSans 2000 0 0 0 D
<< properties >>
string GDS_END 8334402
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8229130
<< end >>
