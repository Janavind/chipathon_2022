magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< locali >>
rect 1935 9564 1969 9580
rect 1935 9514 1969 9530
<< viali >>
rect 1935 9530 1969 9564
<< metal1 >>
rect 1923 9564 1981 9570
rect 1923 9530 1935 9564
rect 1969 9561 1981 9564
rect 40669 9561 40675 9573
rect 1969 9533 40675 9561
rect 1969 9530 1981 9533
rect 1923 9524 1981 9530
rect 40669 9521 40675 9533
rect 40727 9521 40733 9573
rect 1629 8649 1689 8705
rect 6621 8649 6681 8705
rect 11613 8649 11673 8705
rect 16605 8649 16665 8705
rect 21597 8649 21657 8705
rect 26589 8649 26649 8705
rect 31581 8649 31641 8705
rect 36573 8649 36633 8705
rect 40669 8615 40675 8624
rect 1473 8581 40675 8615
rect 40669 8572 40675 8581
rect 40727 8615 40733 8624
rect 40727 8581 40785 8615
rect 40727 8572 40733 8581
rect 1501 6632 1529 6698
rect 1501 6604 1601 6632
rect 1478 6192 1524 6446
rect 1573 5316 1601 6604
rect 1703 6552 1731 6698
rect 6493 6632 6521 6698
rect 6493 6604 6593 6632
rect 1646 6524 1731 6552
rect 1646 5304 1674 6524
rect 6470 6192 6516 6446
rect 6565 5316 6593 6604
rect 6695 6552 6723 6698
rect 11485 6632 11513 6698
rect 11485 6604 11585 6632
rect 6638 6524 6723 6552
rect 6638 5304 6666 6524
rect 11462 6192 11508 6446
rect 11557 5316 11585 6604
rect 11687 6552 11715 6698
rect 16477 6632 16505 6698
rect 16477 6604 16577 6632
rect 11630 6524 11715 6552
rect 11630 5304 11658 6524
rect 16454 6192 16500 6446
rect 16549 5316 16577 6604
rect 16679 6552 16707 6698
rect 21469 6632 21497 6698
rect 21469 6604 21569 6632
rect 16622 6524 16707 6552
rect 16622 5304 16650 6524
rect 21446 6192 21492 6446
rect 21541 5316 21569 6604
rect 21671 6552 21699 6698
rect 26461 6632 26489 6698
rect 26461 6604 26561 6632
rect 21614 6524 21699 6552
rect 21614 5304 21642 6524
rect 26438 6192 26484 6446
rect 26533 5316 26561 6604
rect 26663 6552 26691 6698
rect 31453 6632 31481 6698
rect 31453 6604 31553 6632
rect 26606 6524 26691 6552
rect 26606 5304 26634 6524
rect 31430 6192 31476 6446
rect 31525 5316 31553 6604
rect 31655 6552 31683 6698
rect 36445 6632 36473 6698
rect 36445 6604 36545 6632
rect 31598 6524 31683 6552
rect 31598 5304 31626 6524
rect 36422 6192 36468 6446
rect 36517 5316 36545 6604
rect 36647 6552 36675 6698
rect 36590 6524 36675 6552
rect 36590 5304 36618 6524
rect 1573 4124 1601 4190
rect 1454 4096 1601 4124
rect 1454 3690 1482 4096
rect 1646 4044 1674 4190
rect 6565 4124 6593 4190
rect 6446 4096 6593 4124
rect 1646 4016 1946 4044
rect 1918 3814 1946 4016
rect 6446 3690 6474 4096
rect 6638 4044 6666 4190
rect 11557 4124 11585 4190
rect 11438 4096 11585 4124
rect 6638 4016 6938 4044
rect 6910 3814 6938 4016
rect 11438 3690 11466 4096
rect 11630 4044 11658 4190
rect 16549 4124 16577 4190
rect 16430 4096 16577 4124
rect 11630 4016 11930 4044
rect 11902 3814 11930 4016
rect 16430 3690 16458 4096
rect 16622 4044 16650 4190
rect 21541 4124 21569 4190
rect 21422 4096 21569 4124
rect 16622 4016 16922 4044
rect 16894 3814 16922 4016
rect 21422 3690 21450 4096
rect 21614 4044 21642 4190
rect 26533 4124 26561 4190
rect 26414 4096 26561 4124
rect 21614 4016 21914 4044
rect 21886 3814 21914 4016
rect 26414 3690 26442 4096
rect 26606 4044 26634 4190
rect 31525 4124 31553 4190
rect 31406 4096 31553 4124
rect 26606 4016 26906 4044
rect 26878 3814 26906 4016
rect 31406 3690 31434 4096
rect 31598 4044 31626 4190
rect 36517 4124 36545 4190
rect 36398 4096 36545 4124
rect 31598 4016 31898 4044
rect 31870 3814 31898 4016
rect 36398 3690 36426 4096
rect 36590 4044 36618 4190
rect 36590 4016 36890 4044
rect 36862 3814 36890 4016
rect 1454 1192 1482 1258
rect 1440 1164 1482 1192
rect 816 252 844 1006
rect 1280 252 1308 1006
rect 1440 252 1468 1164
rect 1918 1112 1946 1258
rect 1904 1084 1946 1112
rect 2050 1112 2078 1258
rect 2514 1192 2542 1258
rect 2702 1192 2730 1258
rect 2514 1164 2556 1192
rect 2050 1084 2092 1112
rect 1904 252 1932 1084
rect 2064 252 2092 1084
rect 2528 252 2556 1164
rect 2688 1164 2730 1192
rect 2688 252 2716 1164
rect 3166 1112 3194 1258
rect 3152 1084 3194 1112
rect 3298 1112 3326 1258
rect 3762 1192 3790 1258
rect 3950 1192 3978 1258
rect 3762 1164 3804 1192
rect 3298 1084 3340 1112
rect 3152 252 3180 1084
rect 3312 252 3340 1084
rect 3776 252 3804 1164
rect 3936 1164 3978 1192
rect 3936 252 3964 1164
rect 4414 1112 4442 1258
rect 4400 1084 4442 1112
rect 4546 1112 4574 1258
rect 5010 1192 5038 1258
rect 5198 1192 5226 1258
rect 5010 1164 5052 1192
rect 4546 1084 4588 1112
rect 4400 252 4428 1084
rect 4560 252 4588 1084
rect 5024 252 5052 1164
rect 5184 1164 5226 1192
rect 5184 252 5212 1164
rect 5662 1112 5690 1258
rect 5648 1084 5690 1112
rect 5794 1112 5822 1258
rect 6258 1192 6286 1258
rect 6446 1192 6474 1258
rect 6258 1164 6300 1192
rect 5794 1084 5836 1112
rect 5648 252 5676 1084
rect 5808 252 5836 1084
rect 6272 252 6300 1164
rect 6432 1164 6474 1192
rect 6432 252 6460 1164
rect 6910 1112 6938 1258
rect 6896 1084 6938 1112
rect 7042 1112 7070 1258
rect 7506 1192 7534 1258
rect 7694 1192 7722 1258
rect 7506 1164 7548 1192
rect 7042 1084 7084 1112
rect 6896 252 6924 1084
rect 7056 252 7084 1084
rect 7520 252 7548 1164
rect 7680 1164 7722 1192
rect 7680 252 7708 1164
rect 8158 1112 8186 1258
rect 8144 1084 8186 1112
rect 8290 1112 8318 1258
rect 8754 1192 8782 1258
rect 8942 1192 8970 1258
rect 8754 1164 8796 1192
rect 8290 1084 8332 1112
rect 8144 252 8172 1084
rect 8304 252 8332 1084
rect 8768 252 8796 1164
rect 8928 1164 8970 1192
rect 8928 252 8956 1164
rect 9406 1112 9434 1258
rect 9392 1084 9434 1112
rect 9538 1112 9566 1258
rect 10002 1192 10030 1258
rect 10190 1192 10218 1258
rect 10002 1164 10044 1192
rect 9538 1084 9580 1112
rect 9392 252 9420 1084
rect 9552 252 9580 1084
rect 10016 252 10044 1164
rect 10176 1164 10218 1192
rect 10176 252 10204 1164
rect 10654 1112 10682 1258
rect 10640 1084 10682 1112
rect 10786 1112 10814 1258
rect 11250 1192 11278 1258
rect 11438 1192 11466 1258
rect 11250 1164 11292 1192
rect 10786 1084 10828 1112
rect 10640 252 10668 1084
rect 10800 252 10828 1084
rect 11264 252 11292 1164
rect 11424 1164 11466 1192
rect 11424 252 11452 1164
rect 11902 1112 11930 1258
rect 11888 1084 11930 1112
rect 12034 1112 12062 1258
rect 12498 1192 12526 1258
rect 12686 1192 12714 1258
rect 12498 1164 12540 1192
rect 12034 1084 12076 1112
rect 11888 252 11916 1084
rect 12048 252 12076 1084
rect 12512 252 12540 1164
rect 12672 1164 12714 1192
rect 12672 252 12700 1164
rect 13150 1112 13178 1258
rect 13136 1084 13178 1112
rect 13282 1112 13310 1258
rect 13746 1192 13774 1258
rect 13934 1192 13962 1258
rect 13746 1164 13788 1192
rect 13282 1084 13324 1112
rect 13136 252 13164 1084
rect 13296 252 13324 1084
rect 13760 252 13788 1164
rect 13920 1164 13962 1192
rect 13920 252 13948 1164
rect 14398 1112 14426 1258
rect 14384 1084 14426 1112
rect 14530 1112 14558 1258
rect 14994 1192 15022 1258
rect 15182 1192 15210 1258
rect 14994 1164 15036 1192
rect 14530 1084 14572 1112
rect 14384 252 14412 1084
rect 14544 252 14572 1084
rect 15008 252 15036 1164
rect 15168 1164 15210 1192
rect 15168 252 15196 1164
rect 15646 1112 15674 1258
rect 15632 1084 15674 1112
rect 15778 1112 15806 1258
rect 16242 1192 16270 1258
rect 16430 1192 16458 1258
rect 16242 1164 16284 1192
rect 15778 1084 15820 1112
rect 15632 252 15660 1084
rect 15792 252 15820 1084
rect 16256 252 16284 1164
rect 16416 1164 16458 1192
rect 16416 252 16444 1164
rect 16894 1112 16922 1258
rect 16880 1084 16922 1112
rect 17026 1112 17054 1258
rect 17490 1192 17518 1258
rect 17678 1192 17706 1258
rect 17490 1164 17532 1192
rect 17026 1084 17068 1112
rect 16880 252 16908 1084
rect 17040 252 17068 1084
rect 17504 252 17532 1164
rect 17664 1164 17706 1192
rect 17664 252 17692 1164
rect 18142 1112 18170 1258
rect 18128 1084 18170 1112
rect 18274 1112 18302 1258
rect 18738 1192 18766 1258
rect 18926 1192 18954 1258
rect 18738 1164 18780 1192
rect 18274 1084 18316 1112
rect 18128 252 18156 1084
rect 18288 252 18316 1084
rect 18752 252 18780 1164
rect 18912 1164 18954 1192
rect 18912 252 18940 1164
rect 19390 1112 19418 1258
rect 19376 1084 19418 1112
rect 19522 1112 19550 1258
rect 19986 1192 20014 1258
rect 20174 1192 20202 1258
rect 19986 1164 20028 1192
rect 19522 1084 19564 1112
rect 19376 252 19404 1084
rect 19536 252 19564 1084
rect 20000 252 20028 1164
rect 20160 1164 20202 1192
rect 20160 252 20188 1164
rect 20638 1112 20666 1258
rect 20624 1084 20666 1112
rect 20770 1112 20798 1258
rect 21234 1192 21262 1258
rect 21422 1192 21450 1258
rect 21234 1164 21276 1192
rect 20770 1084 20812 1112
rect 20624 252 20652 1084
rect 20784 252 20812 1084
rect 21248 252 21276 1164
rect 21408 1164 21450 1192
rect 21408 252 21436 1164
rect 21886 1112 21914 1258
rect 21872 1084 21914 1112
rect 22018 1112 22046 1258
rect 22482 1192 22510 1258
rect 22670 1192 22698 1258
rect 22482 1164 22524 1192
rect 22018 1084 22060 1112
rect 21872 252 21900 1084
rect 22032 252 22060 1084
rect 22496 252 22524 1164
rect 22656 1164 22698 1192
rect 22656 252 22684 1164
rect 23134 1112 23162 1258
rect 23120 1084 23162 1112
rect 23266 1112 23294 1258
rect 23730 1192 23758 1258
rect 23918 1192 23946 1258
rect 23730 1164 23772 1192
rect 23266 1084 23308 1112
rect 23120 252 23148 1084
rect 23280 252 23308 1084
rect 23744 252 23772 1164
rect 23904 1164 23946 1192
rect 23904 252 23932 1164
rect 24382 1112 24410 1258
rect 24368 1084 24410 1112
rect 24514 1112 24542 1258
rect 24978 1192 25006 1258
rect 25166 1192 25194 1258
rect 24978 1164 25020 1192
rect 24514 1084 24556 1112
rect 24368 252 24396 1084
rect 24528 252 24556 1084
rect 24992 252 25020 1164
rect 25152 1164 25194 1192
rect 25152 252 25180 1164
rect 25630 1112 25658 1258
rect 25616 1084 25658 1112
rect 25762 1112 25790 1258
rect 26226 1192 26254 1258
rect 26414 1192 26442 1258
rect 26226 1164 26268 1192
rect 25762 1084 25804 1112
rect 25616 252 25644 1084
rect 25776 252 25804 1084
rect 26240 252 26268 1164
rect 26400 1164 26442 1192
rect 26400 252 26428 1164
rect 26878 1112 26906 1258
rect 26864 1084 26906 1112
rect 27010 1112 27038 1258
rect 27474 1192 27502 1258
rect 27662 1192 27690 1258
rect 27474 1164 27516 1192
rect 27010 1084 27052 1112
rect 26864 252 26892 1084
rect 27024 252 27052 1084
rect 27488 252 27516 1164
rect 27648 1164 27690 1192
rect 27648 252 27676 1164
rect 28126 1112 28154 1258
rect 28112 1084 28154 1112
rect 28258 1112 28286 1258
rect 28722 1192 28750 1258
rect 28910 1192 28938 1258
rect 28722 1164 28764 1192
rect 28258 1084 28300 1112
rect 28112 252 28140 1084
rect 28272 252 28300 1084
rect 28736 252 28764 1164
rect 28896 1164 28938 1192
rect 28896 252 28924 1164
rect 29374 1112 29402 1258
rect 29360 1084 29402 1112
rect 29506 1112 29534 1258
rect 29970 1192 29998 1258
rect 30158 1192 30186 1258
rect 29970 1164 30012 1192
rect 29506 1084 29548 1112
rect 29360 252 29388 1084
rect 29520 252 29548 1084
rect 29984 252 30012 1164
rect 30144 1164 30186 1192
rect 30144 252 30172 1164
rect 30622 1112 30650 1258
rect 30608 1084 30650 1112
rect 30754 1112 30782 1258
rect 31218 1192 31246 1258
rect 31406 1192 31434 1258
rect 31218 1164 31260 1192
rect 30754 1084 30796 1112
rect 30608 252 30636 1084
rect 30768 252 30796 1084
rect 31232 252 31260 1164
rect 31392 1164 31434 1192
rect 31392 252 31420 1164
rect 31870 1112 31898 1258
rect 31856 1084 31898 1112
rect 32002 1112 32030 1258
rect 32466 1192 32494 1258
rect 32654 1192 32682 1258
rect 32466 1164 32508 1192
rect 32002 1084 32044 1112
rect 31856 252 31884 1084
rect 32016 252 32044 1084
rect 32480 252 32508 1164
rect 32640 1164 32682 1192
rect 32640 252 32668 1164
rect 33118 1112 33146 1258
rect 33104 1084 33146 1112
rect 33250 1112 33278 1258
rect 33714 1192 33742 1258
rect 33902 1192 33930 1258
rect 33714 1164 33756 1192
rect 33250 1084 33292 1112
rect 33104 252 33132 1084
rect 33264 252 33292 1084
rect 33728 252 33756 1164
rect 33888 1164 33930 1192
rect 33888 252 33916 1164
rect 34366 1112 34394 1258
rect 34352 1084 34394 1112
rect 34498 1112 34526 1258
rect 34962 1192 34990 1258
rect 35150 1192 35178 1258
rect 34962 1164 35004 1192
rect 34498 1084 34540 1112
rect 34352 252 34380 1084
rect 34512 252 34540 1084
rect 34976 252 35004 1164
rect 35136 1164 35178 1192
rect 35136 252 35164 1164
rect 35614 1112 35642 1258
rect 35600 1084 35642 1112
rect 35746 1112 35774 1258
rect 36210 1192 36238 1258
rect 36398 1192 36426 1258
rect 36210 1164 36252 1192
rect 35746 1084 35788 1112
rect 35600 252 35628 1084
rect 35760 252 35788 1084
rect 36224 252 36252 1164
rect 36384 1164 36426 1192
rect 36384 252 36412 1164
rect 36862 1112 36890 1258
rect 36848 1084 36890 1112
rect 36994 1112 37022 1258
rect 37458 1192 37486 1258
rect 37646 1192 37674 1258
rect 37458 1164 37500 1192
rect 36994 1084 37036 1112
rect 36848 252 36876 1084
rect 37008 252 37036 1084
rect 37472 252 37500 1164
rect 37632 1164 37674 1192
rect 37632 252 37660 1164
rect 38110 1112 38138 1258
rect 38096 1084 38138 1112
rect 38242 1112 38270 1258
rect 38706 1192 38734 1258
rect 38894 1192 38922 1258
rect 38706 1164 38748 1192
rect 38242 1084 38284 1112
rect 38096 252 38124 1084
rect 38256 252 38284 1084
rect 38720 252 38748 1164
rect 38880 1164 38922 1192
rect 38880 252 38908 1164
rect 39358 1112 39386 1258
rect 39344 1084 39386 1112
rect 39490 1112 39518 1258
rect 39954 1192 39982 1258
rect 40142 1192 40170 1258
rect 39954 1164 39996 1192
rect 39490 1084 39532 1112
rect 39344 252 39372 1084
rect 39504 252 39532 1084
rect 39968 252 39996 1164
rect 40128 1164 40170 1192
rect 40128 252 40156 1164
rect 40606 1112 40634 1258
rect 40592 1084 40634 1112
rect 40738 1112 40766 1258
rect 41202 1192 41230 1258
rect 41202 1164 41244 1192
rect 40738 1084 40780 1112
rect 40592 252 40620 1084
rect 40752 252 40780 1084
rect 41216 252 41244 1164
<< via1 >>
rect 40675 9521 40727 9573
rect 40675 8572 40727 8624
<< metal2 >>
rect 1360 9797 1388 9825
rect 40675 9573 40727 9579
rect 40675 9515 40727 9521
rect 40687 8630 40715 9515
rect 40675 8624 40727 8630
rect 40675 8566 40727 8572
<< metal3 >>
rect -49 10032 49 10130
rect 41261 10032 41359 10130
rect 0 9533 41310 9593
rect -49 8912 49 9010
rect 41261 8912 41359 9010
rect 1601 8469 1699 8567
rect 6593 8469 6691 8567
rect 11585 8469 11683 8567
rect 16577 8469 16675 8567
rect 21569 8469 21667 8567
rect 26561 8469 26659 8567
rect 31553 8469 31651 8567
rect 36545 8469 36643 8567
rect 1587 8053 1685 8151
rect 6579 8053 6677 8151
rect 11571 8053 11669 8151
rect 16563 8053 16661 8151
rect 21555 8053 21653 8151
rect 26547 8053 26645 8151
rect 31539 8053 31637 8151
rect 36531 8053 36629 8151
rect 1702 7851 1800 7949
rect 6694 7851 6792 7949
rect 11686 7851 11784 7949
rect 16678 7851 16776 7949
rect 21670 7851 21768 7949
rect 26662 7851 26760 7949
rect 31654 7851 31752 7949
rect 36646 7851 36744 7949
rect 1581 7519 1679 7617
rect 6573 7519 6671 7617
rect 11565 7519 11663 7617
rect 16557 7519 16655 7617
rect 21549 7519 21647 7617
rect 26541 7519 26639 7617
rect 31533 7519 31631 7617
rect 36525 7519 36623 7617
rect 1592 7082 1690 7180
rect 6584 7082 6682 7180
rect 11576 7082 11674 7180
rect 16568 7082 16666 7180
rect 21560 7082 21658 7180
rect 26552 7082 26650 7180
rect 31544 7082 31642 7180
rect 36536 7082 36634 7180
rect 1706 6289 1804 6387
rect 6698 6289 6796 6387
rect 11690 6289 11788 6387
rect 16682 6289 16780 6387
rect 21674 6289 21772 6387
rect 26666 6289 26764 6387
rect 31658 6289 31756 6387
rect 36650 6289 36748 6387
rect 1706 5967 1804 6065
rect 6698 5967 6796 6065
rect 11690 5967 11788 6065
rect 16682 5967 16780 6065
rect 21674 5967 21772 6065
rect 26666 5967 26764 6065
rect 31658 5967 31756 6065
rect 36650 5967 36748 6065
rect 1694 5129 1792 5227
rect 6686 5129 6784 5227
rect 11678 5129 11776 5227
rect 16670 5129 16768 5227
rect 21662 5129 21760 5227
rect 26654 5129 26752 5227
rect 31646 5129 31744 5227
rect 36638 5129 36736 5227
rect 1776 4355 1874 4453
rect 6768 4355 6866 4453
rect 11760 4355 11858 4453
rect 16752 4355 16850 4453
rect 21744 4355 21842 4453
rect 26736 4355 26834 4453
rect 31728 4355 31826 4453
rect 36720 4355 36818 4453
rect 0 4222 36818 4282
rect 0 3506 41310 3566
rect 0 3382 41310 3442
rect 0 3258 41310 3318
rect 0 3134 41310 3194
rect 0 3010 41310 3070
rect 0 2886 41310 2946
rect 0 2762 41310 2822
rect 0 2638 41310 2698
rect 1949 1862 2047 1960
rect 3197 1862 3295 1960
rect 4445 1862 4543 1960
rect 5693 1862 5791 1960
rect 6941 1862 7039 1960
rect 8189 1862 8287 1960
rect 9437 1862 9535 1960
rect 10685 1862 10783 1960
rect 11933 1862 12031 1960
rect 13181 1862 13279 1960
rect 14429 1862 14527 1960
rect 15677 1862 15775 1960
rect 16925 1862 17023 1960
rect 18173 1862 18271 1960
rect 19421 1862 19519 1960
rect 20669 1862 20767 1960
rect 21917 1862 22015 1960
rect 23165 1862 23263 1960
rect 24413 1862 24511 1960
rect 25661 1862 25759 1960
rect 26909 1862 27007 1960
rect 28157 1862 28255 1960
rect 29405 1862 29503 1960
rect 30653 1862 30751 1960
rect 31901 1862 31999 1960
rect 33149 1862 33247 1960
rect 34397 1862 34495 1960
rect 35645 1862 35743 1960
rect 36893 1862 36991 1960
rect 38141 1862 38239 1960
rect 39389 1862 39487 1960
rect 40637 1862 40735 1960
rect 0 951 41310 1011
rect 1132 313 1230 411
rect 1518 313 1616 411
rect 2380 313 2478 411
rect 2766 313 2864 411
rect 3628 313 3726 411
rect 4014 313 4112 411
rect 4876 313 4974 411
rect 5262 313 5360 411
rect 6124 313 6222 411
rect 6510 313 6608 411
rect 7372 313 7470 411
rect 7758 313 7856 411
rect 8620 313 8718 411
rect 9006 313 9104 411
rect 9868 313 9966 411
rect 10254 313 10352 411
rect 11116 313 11214 411
rect 11502 313 11600 411
rect 12364 313 12462 411
rect 12750 313 12848 411
rect 13612 313 13710 411
rect 13998 313 14096 411
rect 14860 313 14958 411
rect 15246 313 15344 411
rect 16108 313 16206 411
rect 16494 313 16592 411
rect 17356 313 17454 411
rect 17742 313 17840 411
rect 18604 313 18702 411
rect 18990 313 19088 411
rect 19852 313 19950 411
rect 20238 313 20336 411
rect 21100 313 21198 411
rect 21486 313 21584 411
rect 22348 313 22446 411
rect 22734 313 22832 411
rect 23596 313 23694 411
rect 23982 313 24080 411
rect 24844 313 24942 411
rect 25230 313 25328 411
rect 26092 313 26190 411
rect 26478 313 26576 411
rect 27340 313 27438 411
rect 27726 313 27824 411
rect 28588 313 28686 411
rect 28974 313 29072 411
rect 29836 313 29934 411
rect 30222 313 30320 411
rect 31084 313 31182 411
rect 31470 313 31568 411
rect 32332 313 32430 411
rect 32718 313 32816 411
rect 33580 313 33678 411
rect 33966 313 34064 411
rect 34828 313 34926 411
rect 35214 313 35312 411
rect 36076 313 36174 411
rect 36462 313 36560 411
rect 37324 313 37422 411
rect 37710 313 37808 411
rect 38572 313 38670 411
rect 38958 313 39056 411
rect 39820 313 39918 411
rect 40206 313 40304 411
rect 41068 313 41166 411
use sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_array  sky130_sram_1kbyte_1rw1r_8x1024_8_column_mux_array_0
timestamp 1666464484
transform 1 0 0 0 -1 3938
box 0 87 41310 2680
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_0
timestamp 1666464484
transform 1 0 1923 0 1 9514
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_0
timestamp 1666464484
transform 1 0 40669 0 1 9515
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_1
timestamp 1666464484
transform 1 0 40669 0 1 8566
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_precharge_array  sky130_sram_1kbyte_1rw1r_8x1024_8_precharge_array_0
timestamp 1666464484
transform 1 0 0 0 -1 1006
box 0 -12 41310 768
use sky130_sram_1kbyte_1rw1r_8x1024_8_sense_amp_array  sky130_sram_1kbyte_1rw1r_8x1024_8_sense_amp_array_0
timestamp 1666464484
transform 1 0 0 0 -1 6446
box 0 0 37255 2256
use sky130_sram_1kbyte_1rw1r_8x1024_8_write_driver_array  sky130_sram_1kbyte_1rw1r_8x1024_8_write_driver_array_0
timestamp 1666464484
transform 1 0 0 0 -1 8709
box 998 4 40785 2011
use sky130_sram_1kbyte_1rw1r_8x1024_8_write_mask_and_array  sky130_sram_1kbyte_1rw1r_8x1024_8_write_mask_and_array_0
timestamp 1666464484
transform 1 0 0 0 -1 10081
box -49 -49 41359 1177
<< labels >>
rlabel metal3 s 21674 5967 21772 6065 4 vdd
port 1 nsew
rlabel metal3 s 36638 5129 36736 5227 4 vdd
port 1 nsew
rlabel metal3 s 31533 7519 31631 7617 4 vdd
port 1 nsew
rlabel metal3 s 26666 5967 26764 6065 4 vdd
port 1 nsew
rlabel metal3 s 26541 7519 26639 7617 4 vdd
port 1 nsew
rlabel metal3 s 21662 5129 21760 5227 4 vdd
port 1 nsew
rlabel metal3 s 41261 8912 41359 9010 4 vdd
port 1 nsew
rlabel metal3 s 31646 5129 31744 5227 4 vdd
port 1 nsew
rlabel metal3 s 36525 7519 36623 7617 4 vdd
port 1 nsew
rlabel metal3 s 31658 5967 31756 6065 4 vdd
port 1 nsew
rlabel metal3 s 26561 8469 26659 8567 4 vdd
port 1 nsew
rlabel metal3 s 21549 7519 21647 7617 4 vdd
port 1 nsew
rlabel metal3 s 36545 8469 36643 8567 4 vdd
port 1 nsew
rlabel metal3 s 21569 8469 21667 8567 4 vdd
port 1 nsew
rlabel metal3 s 31553 8469 31651 8567 4 vdd
port 1 nsew
rlabel metal3 s 26654 5129 26752 5227 4 vdd
port 1 nsew
rlabel metal3 s 36650 5967 36748 6065 4 vdd
port 1 nsew
rlabel metal3 s 23165 1862 23263 1960 4 gnd
port 2 nsew
rlabel metal3 s 26736 4355 26834 4453 4 gnd
port 2 nsew
rlabel metal3 s 31728 4355 31826 4453 4 gnd
port 2 nsew
rlabel metal3 s 36646 7851 36744 7949 4 gnd
port 2 nsew
rlabel metal3 s 40637 1862 40735 1960 4 gnd
port 2 nsew
rlabel metal3 s 20669 1862 20767 1960 4 gnd
port 2 nsew
rlabel metal3 s 36650 6289 36748 6387 4 gnd
port 2 nsew
rlabel metal3 s 26547 8053 26645 8151 4 gnd
port 2 nsew
rlabel metal3 s 39389 1862 39487 1960 4 gnd
port 2 nsew
rlabel metal3 s 31901 1862 31999 1960 4 gnd
port 2 nsew
rlabel metal3 s 21674 6289 21772 6387 4 gnd
port 2 nsew
rlabel metal3 s 36893 1862 36991 1960 4 gnd
port 2 nsew
rlabel metal3 s 21917 1862 22015 1960 4 gnd
port 2 nsew
rlabel metal3 s 38141 1862 38239 1960 4 gnd
port 2 nsew
rlabel metal3 s 35645 1862 35743 1960 4 gnd
port 2 nsew
rlabel metal3 s 33149 1862 33247 1960 4 gnd
port 2 nsew
rlabel metal3 s 21560 7082 21658 7180 4 gnd
port 2 nsew
rlabel metal3 s 26552 7082 26650 7180 4 gnd
port 2 nsew
rlabel metal3 s 34397 1862 34495 1960 4 gnd
port 2 nsew
rlabel metal3 s 30653 1862 30751 1960 4 gnd
port 2 nsew
rlabel metal3 s 36531 8053 36629 8151 4 gnd
port 2 nsew
rlabel metal3 s 31539 8053 31637 8151 4 gnd
port 2 nsew
rlabel metal3 s 29405 1862 29503 1960 4 gnd
port 2 nsew
rlabel metal3 s 21744 4355 21842 4453 4 gnd
port 2 nsew
rlabel metal3 s 21670 7851 21768 7949 4 gnd
port 2 nsew
rlabel metal3 s 31544 7082 31642 7180 4 gnd
port 2 nsew
rlabel metal3 s 28157 1862 28255 1960 4 gnd
port 2 nsew
rlabel metal3 s 31654 7851 31752 7949 4 gnd
port 2 nsew
rlabel metal3 s 36536 7082 36634 7180 4 gnd
port 2 nsew
rlabel metal3 s 25661 1862 25759 1960 4 gnd
port 2 nsew
rlabel metal3 s 41261 10032 41359 10130 4 gnd
port 2 nsew
rlabel metal3 s 26666 6289 26764 6387 4 gnd
port 2 nsew
rlabel metal3 s 26909 1862 27007 1960 4 gnd
port 2 nsew
rlabel metal3 s 36720 4355 36818 4453 4 gnd
port 2 nsew
rlabel metal3 s 31658 6289 31756 6387 4 gnd
port 2 nsew
rlabel metal3 s 26662 7851 26760 7949 4 gnd
port 2 nsew
rlabel metal3 s 24413 1862 24511 1960 4 gnd
port 2 nsew
rlabel metal3 s 21555 8053 21653 8151 4 gnd
port 2 nsew
rlabel metal3 s 0 2638 41310 2698 4 sel_7
port 3 nsew
rlabel metal3 s 0 4222 36818 4282 4 s_en
port 4 nsew
rlabel metal3 s 0 9533 41310 9593 4 w_en
port 5 nsew
rlabel metal3 s 1706 5967 1804 6065 4 vdd
port 1 nsew
rlabel metal3 s 1694 5129 1792 5227 4 vdd
port 1 nsew
rlabel metal3 s 14429 1862 14527 1960 4 gnd
port 2 nsew
rlabel metal3 s 16563 8053 16661 8151 4 gnd
port 2 nsew
rlabel metal3 s 11565 7519 11663 7617 4 vdd
port 1 nsew
rlabel metal3 s 16682 5967 16780 6065 4 vdd
port 1 nsew
rlabel metal3 s 0 951 41310 1011 4 p_en_bar
port 6 nsew
rlabel metal3 s 11585 8469 11683 8567 4 vdd
port 1 nsew
rlabel metal3 s 16925 1862 17023 1960 4 gnd
port 2 nsew
rlabel metal3 s 18173 1862 18271 1960 4 gnd
port 2 nsew
rlabel metal3 s 0 3506 41310 3566 4 sel_0
port 7 nsew
rlabel metal3 s 19421 1862 19519 1960 4 gnd
port 2 nsew
rlabel metal3 s 6941 1862 7039 1960 4 gnd
port 2 nsew
rlabel metal3 s 0 3382 41310 3442 4 sel_1
port 8 nsew
rlabel metal3 s 6573 7519 6671 7617 4 vdd
port 1 nsew
rlabel metal3 s 16568 7082 16666 7180 4 gnd
port 2 nsew
rlabel metal3 s 0 3258 41310 3318 4 sel_2
port 9 nsew
rlabel metal3 s 11571 8053 11669 8151 4 gnd
port 2 nsew
rlabel metal3 s 6698 6289 6796 6387 4 gnd
port 2 nsew
rlabel metal3 s 11933 1862 12031 1960 4 gnd
port 2 nsew
rlabel metal3 s 16577 8469 16675 8567 4 vdd
port 1 nsew
rlabel metal3 s 6579 8053 6677 8151 4 gnd
port 2 nsew
rlabel metal3 s 1581 7519 1679 7617 4 vdd
port 1 nsew
rlabel metal3 s 1776 4355 1874 4453 4 gnd
port 2 nsew
rlabel metal3 s 6593 8469 6691 8567 4 vdd
port 1 nsew
rlabel metal3 s 16682 6289 16780 6387 4 gnd
port 2 nsew
rlabel metal3 s 11690 6289 11788 6387 4 gnd
port 2 nsew
rlabel metal3 s 16557 7519 16655 7617 4 vdd
port 1 nsew
rlabel metal3 s 0 3134 41310 3194 4 sel_3
port 10 nsew
rlabel metal3 s 11678 5129 11776 5227 4 vdd
port 1 nsew
rlabel metal3 s 6768 4355 6866 4453 4 gnd
port 2 nsew
rlabel metal3 s 1706 6289 1804 6387 4 gnd
port 2 nsew
rlabel metal3 s 6686 5129 6784 5227 4 vdd
port 1 nsew
rlabel metal3 s -49 8912 49 9010 4 vdd
port 1 nsew
rlabel metal3 s 6698 5967 6796 6065 4 vdd
port 1 nsew
rlabel metal3 s 6584 7082 6682 7180 4 gnd
port 2 nsew
rlabel metal3 s -49 10032 49 10130 4 gnd
port 2 nsew
rlabel metal3 s 1601 8469 1699 8567 4 vdd
port 1 nsew
rlabel metal3 s 11760 4355 11858 4453 4 gnd
port 2 nsew
rlabel metal3 s 16670 5129 16768 5227 4 vdd
port 1 nsew
rlabel metal3 s 1949 1862 2047 1960 4 gnd
port 2 nsew
rlabel metal3 s 9437 1862 9535 1960 4 gnd
port 2 nsew
rlabel metal3 s 11686 7851 11784 7949 4 gnd
port 2 nsew
rlabel metal3 s 1587 8053 1685 8151 4 gnd
port 2 nsew
rlabel metal3 s 1592 7082 1690 7180 4 gnd
port 2 nsew
rlabel metal3 s 6694 7851 6792 7949 4 gnd
port 2 nsew
rlabel metal3 s 4445 1862 4543 1960 4 gnd
port 2 nsew
rlabel metal3 s 5693 1862 5791 1960 4 gnd
port 2 nsew
rlabel metal3 s 0 3010 41310 3070 4 sel_4
port 11 nsew
rlabel metal3 s 15677 1862 15775 1960 4 gnd
port 2 nsew
rlabel metal3 s 11576 7082 11674 7180 4 gnd
port 2 nsew
rlabel metal3 s 8189 1862 8287 1960 4 gnd
port 2 nsew
rlabel metal3 s 16678 7851 16776 7949 4 gnd
port 2 nsew
rlabel metal3 s 1702 7851 1800 7949 4 gnd
port 2 nsew
rlabel metal3 s 0 2886 41310 2946 4 sel_5
port 12 nsew
rlabel metal3 s 13181 1862 13279 1960 4 gnd
port 2 nsew
rlabel metal3 s 0 2762 41310 2822 4 sel_6
port 13 nsew
rlabel metal3 s 16752 4355 16850 4453 4 gnd
port 2 nsew
rlabel metal3 s 3197 1862 3295 1960 4 gnd
port 2 nsew
rlabel metal3 s 11690 5967 11788 6065 4 vdd
port 1 nsew
rlabel metal3 s 10685 1862 10783 1960 4 gnd
port 2 nsew
rlabel metal3 s 3628 313 3726 411 4 vdd
port 1 nsew
rlabel metal3 s 12750 313 12848 411 4 vdd
port 1 nsew
rlabel metal3 s 5262 313 5360 411 4 vdd
port 1 nsew
rlabel metal3 s 15246 313 15344 411 4 vdd
port 1 nsew
rlabel metal3 s 6510 313 6608 411 4 vdd
port 1 nsew
rlabel metal3 s 11116 313 11214 411 4 vdd
port 1 nsew
rlabel metal3 s 13998 313 14096 411 4 vdd
port 1 nsew
rlabel metal3 s 9868 313 9966 411 4 vdd
port 1 nsew
rlabel metal3 s 11502 313 11600 411 4 vdd
port 1 nsew
rlabel metal3 s 16108 313 16206 411 4 vdd
port 1 nsew
rlabel metal3 s 2380 313 2478 411 4 vdd
port 1 nsew
rlabel metal3 s 2766 313 2864 411 4 vdd
port 1 nsew
rlabel metal3 s 1132 313 1230 411 4 vdd
port 1 nsew
rlabel metal3 s 12364 313 12462 411 4 vdd
port 1 nsew
rlabel metal3 s 8620 313 8718 411 4 vdd
port 1 nsew
rlabel metal3 s 20238 313 20336 411 4 vdd
port 1 nsew
rlabel metal3 s 1518 313 1616 411 4 vdd
port 1 nsew
rlabel metal3 s 16494 313 16592 411 4 vdd
port 1 nsew
rlabel metal3 s 18990 313 19088 411 4 vdd
port 1 nsew
rlabel metal3 s 19852 313 19950 411 4 vdd
port 1 nsew
rlabel metal3 s 13612 313 13710 411 4 vdd
port 1 nsew
rlabel metal3 s 17356 313 17454 411 4 vdd
port 1 nsew
rlabel metal3 s 7758 313 7856 411 4 vdd
port 1 nsew
rlabel metal3 s 17742 313 17840 411 4 vdd
port 1 nsew
rlabel metal3 s 4014 313 4112 411 4 vdd
port 1 nsew
rlabel metal3 s 6124 313 6222 411 4 vdd
port 1 nsew
rlabel metal3 s 18604 313 18702 411 4 vdd
port 1 nsew
rlabel metal3 s 14860 313 14958 411 4 vdd
port 1 nsew
rlabel metal3 s 10254 313 10352 411 4 vdd
port 1 nsew
rlabel metal3 s 4876 313 4974 411 4 vdd
port 1 nsew
rlabel metal3 s 9006 313 9104 411 4 vdd
port 1 nsew
rlabel metal3 s 7372 313 7470 411 4 vdd
port 1 nsew
rlabel metal3 s 33580 313 33678 411 4 vdd
port 1 nsew
rlabel metal3 s 34828 313 34926 411 4 vdd
port 1 nsew
rlabel metal3 s 23982 313 24080 411 4 vdd
port 1 nsew
rlabel metal3 s 30222 313 30320 411 4 vdd
port 1 nsew
rlabel metal3 s 22734 313 22832 411 4 vdd
port 1 nsew
rlabel metal3 s 32332 313 32430 411 4 vdd
port 1 nsew
rlabel metal3 s 27726 313 27824 411 4 vdd
port 1 nsew
rlabel metal3 s 40206 313 40304 411 4 vdd
port 1 nsew
rlabel metal3 s 23596 313 23694 411 4 vdd
port 1 nsew
rlabel metal3 s 39820 313 39918 411 4 vdd
port 1 nsew
rlabel metal3 s 41068 313 41166 411 4 vdd
port 1 nsew
rlabel metal3 s 29836 313 29934 411 4 vdd
port 1 nsew
rlabel metal3 s 21486 313 21584 411 4 vdd
port 1 nsew
rlabel metal3 s 31084 313 31182 411 4 vdd
port 1 nsew
rlabel metal3 s 28974 313 29072 411 4 vdd
port 1 nsew
rlabel metal3 s 27340 313 27438 411 4 vdd
port 1 nsew
rlabel metal3 s 28588 313 28686 411 4 vdd
port 1 nsew
rlabel metal3 s 36076 313 36174 411 4 vdd
port 1 nsew
rlabel metal3 s 38572 313 38670 411 4 vdd
port 1 nsew
rlabel metal3 s 37324 313 37422 411 4 vdd
port 1 nsew
rlabel metal3 s 26092 313 26190 411 4 vdd
port 1 nsew
rlabel metal3 s 31470 313 31568 411 4 vdd
port 1 nsew
rlabel metal3 s 38958 313 39056 411 4 vdd
port 1 nsew
rlabel metal3 s 35214 313 35312 411 4 vdd
port 1 nsew
rlabel metal3 s 33966 313 34064 411 4 vdd
port 1 nsew
rlabel metal3 s 22348 313 22446 411 4 vdd
port 1 nsew
rlabel metal3 s 26478 313 26576 411 4 vdd
port 1 nsew
rlabel metal3 s 21100 313 21198 411 4 vdd
port 1 nsew
rlabel metal3 s 25230 313 25328 411 4 vdd
port 1 nsew
rlabel metal3 s 32718 313 32816 411 4 vdd
port 1 nsew
rlabel metal3 s 36462 313 36560 411 4 vdd
port 1 nsew
rlabel metal3 s 37710 313 37808 411 4 vdd
port 1 nsew
rlabel metal3 s 24844 313 24942 411 4 vdd
port 1 nsew
rlabel metal2 s 1360 9797 1388 9825 4 bank_wmask_0
port 14 nsew
rlabel metal1 s 1473 8581 40785 8615 4 wdriver_sel_0
port 15 nsew
rlabel metal1 s 21597 8649 21657 8705 4 din_4
port 16 nsew
rlabel metal1 s 26589 8649 26649 8705 4 din_5
port 17 nsew
rlabel metal1 s 31581 8649 31641 8705 4 din_6
port 18 nsew
rlabel metal1 s 36573 8649 36633 8705 4 din_7
port 19 nsew
rlabel metal1 s 21446 6192 21492 6446 4 dout_4
port 20 nsew
rlabel metal1 s 26438 6192 26484 6446 4 dout_5
port 21 nsew
rlabel metal1 s 31430 6192 31476 6446 4 dout_6
port 22 nsew
rlabel metal1 s 36422 6192 36468 6446 4 dout_7
port 23 nsew
rlabel metal1 s 1478 6192 1524 6446 4 dout_0
port 24 nsew
rlabel metal1 s 6470 6192 6516 6446 4 dout_1
port 25 nsew
rlabel metal1 s 11462 6192 11508 6446 4 dout_2
port 26 nsew
rlabel metal1 s 16454 6192 16500 6446 4 dout_3
port 27 nsew
rlabel metal1 s 1629 8649 1689 8705 4 din_0
port 28 nsew
rlabel metal1 s 6621 8649 6681 8705 4 din_1
port 29 nsew
rlabel metal1 s 11613 8649 11673 8705 4 din_2
port 30 nsew
rlabel metal1 s 16605 8649 16665 8705 4 din_3
port 31 nsew
rlabel metal1 s 1280 252 1308 1006 4 rbl_bl
port 32 nsew
rlabel metal1 s 816 252 844 1006 4 rbl_br
port 33 nsew
rlabel metal1 s 1440 252 1468 1006 4 bl_0
port 34 nsew
rlabel metal1 s 1904 252 1932 1006 4 br_0
port 35 nsew
rlabel metal1 s 2528 252 2556 1006 4 bl_1
port 36 nsew
rlabel metal1 s 2064 252 2092 1006 4 br_1
port 37 nsew
rlabel metal1 s 2688 252 2716 1006 4 bl_2
port 38 nsew
rlabel metal1 s 3152 252 3180 1006 4 br_2
port 39 nsew
rlabel metal1 s 3776 252 3804 1006 4 bl_3
port 40 nsew
rlabel metal1 s 3312 252 3340 1006 4 br_3
port 41 nsew
rlabel metal1 s 3936 252 3964 1006 4 bl_4
port 42 nsew
rlabel metal1 s 4400 252 4428 1006 4 br_4
port 43 nsew
rlabel metal1 s 5024 252 5052 1006 4 bl_5
port 44 nsew
rlabel metal1 s 4560 252 4588 1006 4 br_5
port 45 nsew
rlabel metal1 s 5184 252 5212 1006 4 bl_6
port 46 nsew
rlabel metal1 s 5648 252 5676 1006 4 br_6
port 47 nsew
rlabel metal1 s 6272 252 6300 1006 4 bl_7
port 48 nsew
rlabel metal1 s 5808 252 5836 1006 4 br_7
port 49 nsew
rlabel metal1 s 6432 252 6460 1006 4 bl_8
port 50 nsew
rlabel metal1 s 6896 252 6924 1006 4 br_8
port 51 nsew
rlabel metal1 s 7520 252 7548 1006 4 bl_9
port 52 nsew
rlabel metal1 s 7056 252 7084 1006 4 br_9
port 53 nsew
rlabel metal1 s 7680 252 7708 1006 4 bl_10
port 54 nsew
rlabel metal1 s 8144 252 8172 1006 4 br_10
port 55 nsew
rlabel metal1 s 8768 252 8796 1006 4 bl_11
port 56 nsew
rlabel metal1 s 8304 252 8332 1006 4 br_11
port 57 nsew
rlabel metal1 s 8928 252 8956 1006 4 bl_12
port 58 nsew
rlabel metal1 s 9392 252 9420 1006 4 br_12
port 59 nsew
rlabel metal1 s 10016 252 10044 1006 4 bl_13
port 60 nsew
rlabel metal1 s 9552 252 9580 1006 4 br_13
port 61 nsew
rlabel metal1 s 10176 252 10204 1006 4 bl_14
port 62 nsew
rlabel metal1 s 10640 252 10668 1006 4 br_14
port 63 nsew
rlabel metal1 s 11264 252 11292 1006 4 bl_15
port 64 nsew
rlabel metal1 s 10800 252 10828 1006 4 br_15
port 65 nsew
rlabel metal1 s 11424 252 11452 1006 4 bl_16
port 66 nsew
rlabel metal1 s 11888 252 11916 1006 4 br_16
port 67 nsew
rlabel metal1 s 12512 252 12540 1006 4 bl_17
port 68 nsew
rlabel metal1 s 12048 252 12076 1006 4 br_17
port 69 nsew
rlabel metal1 s 12672 252 12700 1006 4 bl_18
port 70 nsew
rlabel metal1 s 13136 252 13164 1006 4 br_18
port 71 nsew
rlabel metal1 s 13760 252 13788 1006 4 bl_19
port 72 nsew
rlabel metal1 s 13296 252 13324 1006 4 br_19
port 73 nsew
rlabel metal1 s 13920 252 13948 1006 4 bl_20
port 74 nsew
rlabel metal1 s 14384 252 14412 1006 4 br_20
port 75 nsew
rlabel metal1 s 15008 252 15036 1006 4 bl_21
port 76 nsew
rlabel metal1 s 14544 252 14572 1006 4 br_21
port 77 nsew
rlabel metal1 s 15168 252 15196 1006 4 bl_22
port 78 nsew
rlabel metal1 s 15632 252 15660 1006 4 br_22
port 79 nsew
rlabel metal1 s 16256 252 16284 1006 4 bl_23
port 80 nsew
rlabel metal1 s 15792 252 15820 1006 4 br_23
port 81 nsew
rlabel metal1 s 16416 252 16444 1006 4 bl_24
port 82 nsew
rlabel metal1 s 16880 252 16908 1006 4 br_24
port 83 nsew
rlabel metal1 s 17504 252 17532 1006 4 bl_25
port 84 nsew
rlabel metal1 s 17040 252 17068 1006 4 br_25
port 85 nsew
rlabel metal1 s 17664 252 17692 1006 4 bl_26
port 86 nsew
rlabel metal1 s 18128 252 18156 1006 4 br_26
port 87 nsew
rlabel metal1 s 18752 252 18780 1006 4 bl_27
port 88 nsew
rlabel metal1 s 18288 252 18316 1006 4 br_27
port 89 nsew
rlabel metal1 s 18912 252 18940 1006 4 bl_28
port 90 nsew
rlabel metal1 s 19376 252 19404 1006 4 br_28
port 91 nsew
rlabel metal1 s 20000 252 20028 1006 4 bl_29
port 92 nsew
rlabel metal1 s 19536 252 19564 1006 4 br_29
port 93 nsew
rlabel metal1 s 20160 252 20188 1006 4 bl_30
port 94 nsew
rlabel metal1 s 20624 252 20652 1006 4 br_30
port 95 nsew
rlabel metal1 s 20784 252 20812 1006 4 br_31
port 96 nsew
rlabel metal1 s 21248 252 21276 1006 4 bl_31
port 97 nsew
rlabel metal1 s 21408 252 21436 1006 4 bl_32
port 98 nsew
rlabel metal1 s 21872 252 21900 1006 4 br_32
port 99 nsew
rlabel metal1 s 22496 252 22524 1006 4 bl_33
port 100 nsew
rlabel metal1 s 22032 252 22060 1006 4 br_33
port 101 nsew
rlabel metal1 s 22656 252 22684 1006 4 bl_34
port 102 nsew
rlabel metal1 s 23120 252 23148 1006 4 br_34
port 103 nsew
rlabel metal1 s 23744 252 23772 1006 4 bl_35
port 104 nsew
rlabel metal1 s 23280 252 23308 1006 4 br_35
port 105 nsew
rlabel metal1 s 23904 252 23932 1006 4 bl_36
port 106 nsew
rlabel metal1 s 24368 252 24396 1006 4 br_36
port 107 nsew
rlabel metal1 s 24992 252 25020 1006 4 bl_37
port 108 nsew
rlabel metal1 s 24528 252 24556 1006 4 br_37
port 109 nsew
rlabel metal1 s 25152 252 25180 1006 4 bl_38
port 110 nsew
rlabel metal1 s 25616 252 25644 1006 4 br_38
port 111 nsew
rlabel metal1 s 26240 252 26268 1006 4 bl_39
port 112 nsew
rlabel metal1 s 25776 252 25804 1006 4 br_39
port 113 nsew
rlabel metal1 s 26400 252 26428 1006 4 bl_40
port 114 nsew
rlabel metal1 s 26864 252 26892 1006 4 br_40
port 115 nsew
rlabel metal1 s 27488 252 27516 1006 4 bl_41
port 116 nsew
rlabel metal1 s 27024 252 27052 1006 4 br_41
port 117 nsew
rlabel metal1 s 27648 252 27676 1006 4 bl_42
port 118 nsew
rlabel metal1 s 28112 252 28140 1006 4 br_42
port 119 nsew
rlabel metal1 s 28736 252 28764 1006 4 bl_43
port 120 nsew
rlabel metal1 s 28272 252 28300 1006 4 br_43
port 121 nsew
rlabel metal1 s 28896 252 28924 1006 4 bl_44
port 122 nsew
rlabel metal1 s 29360 252 29388 1006 4 br_44
port 123 nsew
rlabel metal1 s 29984 252 30012 1006 4 bl_45
port 124 nsew
rlabel metal1 s 29520 252 29548 1006 4 br_45
port 125 nsew
rlabel metal1 s 30144 252 30172 1006 4 bl_46
port 126 nsew
rlabel metal1 s 30608 252 30636 1006 4 br_46
port 127 nsew
rlabel metal1 s 31232 252 31260 1006 4 bl_47
port 128 nsew
rlabel metal1 s 30768 252 30796 1006 4 br_47
port 129 nsew
rlabel metal1 s 31392 252 31420 1006 4 bl_48
port 130 nsew
rlabel metal1 s 31856 252 31884 1006 4 br_48
port 131 nsew
rlabel metal1 s 32480 252 32508 1006 4 bl_49
port 132 nsew
rlabel metal1 s 32016 252 32044 1006 4 br_49
port 133 nsew
rlabel metal1 s 32640 252 32668 1006 4 bl_50
port 134 nsew
rlabel metal1 s 33104 252 33132 1006 4 br_50
port 135 nsew
rlabel metal1 s 33728 252 33756 1006 4 bl_51
port 136 nsew
rlabel metal1 s 33264 252 33292 1006 4 br_51
port 137 nsew
rlabel metal1 s 33888 252 33916 1006 4 bl_52
port 138 nsew
rlabel metal1 s 34352 252 34380 1006 4 br_52
port 139 nsew
rlabel metal1 s 34976 252 35004 1006 4 bl_53
port 140 nsew
rlabel metal1 s 34512 252 34540 1006 4 br_53
port 141 nsew
rlabel metal1 s 35136 252 35164 1006 4 bl_54
port 142 nsew
rlabel metal1 s 35600 252 35628 1006 4 br_54
port 143 nsew
rlabel metal1 s 36224 252 36252 1006 4 bl_55
port 144 nsew
rlabel metal1 s 35760 252 35788 1006 4 br_55
port 145 nsew
rlabel metal1 s 36384 252 36412 1006 4 bl_56
port 146 nsew
rlabel metal1 s 36848 252 36876 1006 4 br_56
port 147 nsew
rlabel metal1 s 37472 252 37500 1006 4 bl_57
port 148 nsew
rlabel metal1 s 37008 252 37036 1006 4 br_57
port 149 nsew
rlabel metal1 s 37632 252 37660 1006 4 bl_58
port 150 nsew
rlabel metal1 s 38096 252 38124 1006 4 br_58
port 151 nsew
rlabel metal1 s 38720 252 38748 1006 4 bl_59
port 152 nsew
rlabel metal1 s 38256 252 38284 1006 4 br_59
port 153 nsew
rlabel metal1 s 38880 252 38908 1006 4 bl_60
port 154 nsew
rlabel metal1 s 39344 252 39372 1006 4 br_60
port 155 nsew
rlabel metal1 s 39968 252 39996 1006 4 bl_61
port 156 nsew
rlabel metal1 s 39504 252 39532 1006 4 br_61
port 157 nsew
rlabel metal1 s 40128 252 40156 1006 4 bl_62
port 158 nsew
rlabel metal1 s 40592 252 40620 1006 4 br_62
port 159 nsew
rlabel metal1 s 41216 252 41244 1006 4 bl_63
port 160 nsew
rlabel metal1 s 40752 252 40780 1006 4 br_63
port 161 nsew
rlabel locali s 1952 9547 1952 9547 4 wdriver_sel_0
port 15 nsew
<< properties >>
string FIXED_BBOX 0 0 41310 10081
string GDS_END 6720960
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 6610694
<< end >>
