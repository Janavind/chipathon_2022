magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 21 964 157
rect 29 -17 63 21
<< locali >>
rect 284 347 336 492
rect 456 347 508 492
rect 628 347 680 492
rect 800 347 852 492
rect 284 299 946 347
rect 17 143 80 265
rect 752 181 946 299
rect 284 147 946 181
rect 284 56 336 147
rect 456 56 508 147
rect 628 56 680 147
rect 800 56 852 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 19 459 78 493
rect 19 425 35 459
rect 69 425 78 459
rect 19 305 78 425
rect 114 265 164 492
rect 198 459 250 493
rect 198 425 207 459
rect 241 425 250 459
rect 198 305 250 425
rect 370 459 422 493
rect 370 425 378 459
rect 412 425 422 459
rect 370 381 422 425
rect 542 459 594 493
rect 542 425 548 459
rect 582 425 594 459
rect 542 381 594 425
rect 714 459 766 493
rect 714 425 724 459
rect 758 425 766 459
rect 714 381 766 425
rect 886 459 945 493
rect 886 425 896 459
rect 930 425 945 459
rect 886 381 945 425
rect 114 215 718 265
rect 29 17 78 109
rect 114 53 164 215
rect 198 17 250 122
rect 370 17 422 113
rect 542 17 594 113
rect 714 17 766 113
rect 886 17 946 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 35 425 69 459
rect 207 425 241 459
rect 378 425 412 459
rect 548 425 582 459
rect 724 425 758 459
rect 896 425 930 459
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 14 459 998 468
rect 14 428 35 459
rect 23 425 35 428
rect 69 428 207 459
rect 69 425 81 428
rect 23 416 81 425
rect 195 425 207 428
rect 241 428 378 459
rect 241 425 253 428
rect 195 416 253 425
rect 366 425 378 428
rect 412 428 548 459
rect 412 425 424 428
rect 366 416 424 425
rect 536 425 548 428
rect 582 428 724 459
rect 582 425 594 428
rect 536 416 594 425
rect 712 425 724 428
rect 758 428 896 459
rect 758 425 770 428
rect 712 416 770 425
rect 884 425 896 428
rect 930 428 998 459
rect 930 425 942 428
rect 884 416 942 425
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 17 143 80 265 6 A
port 1 nsew signal input
rlabel metal1 s 884 416 942 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 712 416 770 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 536 416 594 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 366 416 424 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 195 416 253 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 23 416 81 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 14 428 998 468 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 -48 1012 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 964 157 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1050 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 800 56 852 147 6 X
port 7 nsew signal output
rlabel locali s 628 56 680 147 6 X
port 7 nsew signal output
rlabel locali s 456 56 508 147 6 X
port 7 nsew signal output
rlabel locali s 284 56 336 147 6 X
port 7 nsew signal output
rlabel locali s 284 147 946 181 6 X
port 7 nsew signal output
rlabel locali s 752 181 946 299 6 X
port 7 nsew signal output
rlabel locali s 284 299 946 347 6 X
port 7 nsew signal output
rlabel locali s 800 347 852 492 6 X
port 7 nsew signal output
rlabel locali s 628 347 680 492 6 X
port 7 nsew signal output
rlabel locali s 456 347 508 492 6 X
port 7 nsew signal output
rlabel locali s 284 347 336 492 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1012 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2261880
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2253036
<< end >>
