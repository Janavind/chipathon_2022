magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect 1018 673 3074 722
rect 1018 391 3186 673
rect 1018 390 3074 391
rect 1018 -130 2908 390
rect 1073 -316 2908 -130
rect 2102 -422 2908 -316
<< pwell >>
rect 1322 -683 2656 -647
rect 1213 -1263 2656 -683
rect 1322 -1299 2656 -1263
<< mvnmos >>
rect 1401 -1273 1521 -673
rect 1577 -1273 1697 -673
rect 1753 -1273 1873 -673
rect 1929 -1273 2049 -673
rect 2105 -1273 2225 -673
rect 2281 -1273 2401 -673
rect 2457 -1273 2577 -673
<< mvpmos >>
rect 1761 456 1861 540
rect 1917 456 2017 540
rect 2197 456 2297 540
rect 2353 456 2453 540
rect 2699 456 2799 656
rect 2855 456 2955 656
rect 1192 172 1592 256
rect 1648 172 2048 256
rect 2104 172 2504 256
rect 1192 -250 1992 -166
rect 2221 -356 2321 -56
rect 2377 -356 2477 -56
rect 2533 -356 2633 -56
rect 2689 -356 2789 -56
<< mvndiff >>
rect 1348 -751 1401 -673
rect 1348 -785 1356 -751
rect 1390 -785 1401 -751
rect 1348 -819 1401 -785
rect 1348 -853 1356 -819
rect 1390 -853 1401 -819
rect 1348 -887 1401 -853
rect 1348 -921 1356 -887
rect 1390 -921 1401 -887
rect 1348 -955 1401 -921
rect 1348 -989 1356 -955
rect 1390 -989 1401 -955
rect 1348 -1023 1401 -989
rect 1348 -1057 1356 -1023
rect 1390 -1057 1401 -1023
rect 1348 -1091 1401 -1057
rect 1348 -1125 1356 -1091
rect 1390 -1125 1401 -1091
rect 1348 -1159 1401 -1125
rect 1348 -1193 1356 -1159
rect 1390 -1193 1401 -1159
rect 1348 -1227 1401 -1193
rect 1348 -1261 1356 -1227
rect 1390 -1261 1401 -1227
rect 1348 -1273 1401 -1261
rect 1521 -751 1577 -673
rect 1521 -785 1532 -751
rect 1566 -785 1577 -751
rect 1521 -819 1577 -785
rect 1521 -853 1532 -819
rect 1566 -853 1577 -819
rect 1521 -887 1577 -853
rect 1521 -921 1532 -887
rect 1566 -921 1577 -887
rect 1521 -955 1577 -921
rect 1521 -989 1532 -955
rect 1566 -989 1577 -955
rect 1521 -1023 1577 -989
rect 1521 -1057 1532 -1023
rect 1566 -1057 1577 -1023
rect 1521 -1091 1577 -1057
rect 1521 -1125 1532 -1091
rect 1566 -1125 1577 -1091
rect 1521 -1159 1577 -1125
rect 1521 -1193 1532 -1159
rect 1566 -1193 1577 -1159
rect 1521 -1227 1577 -1193
rect 1521 -1261 1532 -1227
rect 1566 -1261 1577 -1227
rect 1521 -1273 1577 -1261
rect 1697 -751 1753 -673
rect 1697 -785 1708 -751
rect 1742 -785 1753 -751
rect 1697 -819 1753 -785
rect 1697 -853 1708 -819
rect 1742 -853 1753 -819
rect 1697 -887 1753 -853
rect 1697 -921 1708 -887
rect 1742 -921 1753 -887
rect 1697 -955 1753 -921
rect 1697 -989 1708 -955
rect 1742 -989 1753 -955
rect 1697 -1023 1753 -989
rect 1697 -1057 1708 -1023
rect 1742 -1057 1753 -1023
rect 1697 -1091 1753 -1057
rect 1697 -1125 1708 -1091
rect 1742 -1125 1753 -1091
rect 1697 -1159 1753 -1125
rect 1697 -1193 1708 -1159
rect 1742 -1193 1753 -1159
rect 1697 -1227 1753 -1193
rect 1697 -1261 1708 -1227
rect 1742 -1261 1753 -1227
rect 1697 -1273 1753 -1261
rect 1873 -751 1929 -673
rect 1873 -785 1884 -751
rect 1918 -785 1929 -751
rect 1873 -819 1929 -785
rect 1873 -853 1884 -819
rect 1918 -853 1929 -819
rect 1873 -887 1929 -853
rect 1873 -921 1884 -887
rect 1918 -921 1929 -887
rect 1873 -955 1929 -921
rect 1873 -989 1884 -955
rect 1918 -989 1929 -955
rect 1873 -1023 1929 -989
rect 1873 -1057 1884 -1023
rect 1918 -1057 1929 -1023
rect 1873 -1091 1929 -1057
rect 1873 -1125 1884 -1091
rect 1918 -1125 1929 -1091
rect 1873 -1159 1929 -1125
rect 1873 -1193 1884 -1159
rect 1918 -1193 1929 -1159
rect 1873 -1227 1929 -1193
rect 1873 -1261 1884 -1227
rect 1918 -1261 1929 -1227
rect 1873 -1273 1929 -1261
rect 2049 -751 2105 -673
rect 2049 -785 2060 -751
rect 2094 -785 2105 -751
rect 2049 -819 2105 -785
rect 2049 -853 2060 -819
rect 2094 -853 2105 -819
rect 2049 -887 2105 -853
rect 2049 -921 2060 -887
rect 2094 -921 2105 -887
rect 2049 -955 2105 -921
rect 2049 -989 2060 -955
rect 2094 -989 2105 -955
rect 2049 -1023 2105 -989
rect 2049 -1057 2060 -1023
rect 2094 -1057 2105 -1023
rect 2049 -1091 2105 -1057
rect 2049 -1125 2060 -1091
rect 2094 -1125 2105 -1091
rect 2049 -1159 2105 -1125
rect 2049 -1193 2060 -1159
rect 2094 -1193 2105 -1159
rect 2049 -1227 2105 -1193
rect 2049 -1261 2060 -1227
rect 2094 -1261 2105 -1227
rect 2049 -1273 2105 -1261
rect 2225 -751 2281 -673
rect 2225 -785 2236 -751
rect 2270 -785 2281 -751
rect 2225 -819 2281 -785
rect 2225 -853 2236 -819
rect 2270 -853 2281 -819
rect 2225 -887 2281 -853
rect 2225 -921 2236 -887
rect 2270 -921 2281 -887
rect 2225 -955 2281 -921
rect 2225 -989 2236 -955
rect 2270 -989 2281 -955
rect 2225 -1023 2281 -989
rect 2225 -1057 2236 -1023
rect 2270 -1057 2281 -1023
rect 2225 -1091 2281 -1057
rect 2225 -1125 2236 -1091
rect 2270 -1125 2281 -1091
rect 2225 -1159 2281 -1125
rect 2225 -1193 2236 -1159
rect 2270 -1193 2281 -1159
rect 2225 -1227 2281 -1193
rect 2225 -1261 2236 -1227
rect 2270 -1261 2281 -1227
rect 2225 -1273 2281 -1261
rect 2401 -751 2457 -673
rect 2401 -785 2412 -751
rect 2446 -785 2457 -751
rect 2401 -819 2457 -785
rect 2401 -853 2412 -819
rect 2446 -853 2457 -819
rect 2401 -887 2457 -853
rect 2401 -921 2412 -887
rect 2446 -921 2457 -887
rect 2401 -955 2457 -921
rect 2401 -989 2412 -955
rect 2446 -989 2457 -955
rect 2401 -1023 2457 -989
rect 2401 -1057 2412 -1023
rect 2446 -1057 2457 -1023
rect 2401 -1091 2457 -1057
rect 2401 -1125 2412 -1091
rect 2446 -1125 2457 -1091
rect 2401 -1159 2457 -1125
rect 2401 -1193 2412 -1159
rect 2446 -1193 2457 -1159
rect 2401 -1227 2457 -1193
rect 2401 -1261 2412 -1227
rect 2446 -1261 2457 -1227
rect 2401 -1273 2457 -1261
rect 2577 -751 2630 -673
rect 2577 -785 2588 -751
rect 2622 -785 2630 -751
rect 2577 -819 2630 -785
rect 2577 -853 2588 -819
rect 2622 -853 2630 -819
rect 2577 -887 2630 -853
rect 2577 -921 2588 -887
rect 2622 -921 2630 -887
rect 2577 -955 2630 -921
rect 2577 -989 2588 -955
rect 2622 -989 2630 -955
rect 2577 -1023 2630 -989
rect 2577 -1057 2588 -1023
rect 2622 -1057 2630 -1023
rect 2577 -1091 2630 -1057
rect 2577 -1125 2588 -1091
rect 2622 -1125 2630 -1091
rect 2577 -1159 2630 -1125
rect 2577 -1193 2588 -1159
rect 2622 -1193 2630 -1159
rect 2577 -1227 2630 -1193
rect 2577 -1261 2588 -1227
rect 2622 -1261 2630 -1227
rect 2577 -1273 2630 -1261
<< mvpdiff >>
rect 2646 638 2699 656
rect 2646 604 2654 638
rect 2688 604 2699 638
rect 2646 570 2699 604
rect 1708 502 1761 540
rect 1708 468 1716 502
rect 1750 468 1761 502
rect 1708 456 1761 468
rect 1861 502 1917 540
rect 1861 468 1872 502
rect 1906 468 1917 502
rect 1861 456 1917 468
rect 2017 502 2070 540
rect 2017 468 2028 502
rect 2062 468 2070 502
rect 2017 456 2070 468
rect 2144 502 2197 540
rect 2144 468 2152 502
rect 2186 468 2197 502
rect 2144 456 2197 468
rect 2297 502 2353 540
rect 2297 468 2308 502
rect 2342 468 2353 502
rect 2297 456 2353 468
rect 2453 502 2506 540
rect 2453 468 2464 502
rect 2498 468 2506 502
rect 2453 456 2506 468
rect 2646 536 2654 570
rect 2688 536 2699 570
rect 2646 502 2699 536
rect 2646 468 2654 502
rect 2688 468 2699 502
rect 2646 456 2699 468
rect 2799 638 2855 656
rect 2799 604 2810 638
rect 2844 604 2855 638
rect 2799 570 2855 604
rect 2799 536 2810 570
rect 2844 536 2855 570
rect 2799 502 2855 536
rect 2799 468 2810 502
rect 2844 468 2855 502
rect 2799 456 2855 468
rect 2955 638 3008 656
rect 2955 604 2966 638
rect 3000 604 3008 638
rect 2955 570 3008 604
rect 2955 536 2966 570
rect 3000 536 3008 570
rect 2955 502 3008 536
rect 2955 468 2966 502
rect 3000 468 3008 502
rect 2955 456 3008 468
rect 1139 218 1192 256
rect 1139 184 1147 218
rect 1181 184 1192 218
rect 1139 172 1192 184
rect 1592 218 1648 256
rect 1592 184 1603 218
rect 1637 184 1648 218
rect 1592 172 1648 184
rect 2048 218 2104 256
rect 2048 184 2059 218
rect 2093 184 2104 218
rect 2048 172 2104 184
rect 2504 218 2557 256
rect 2504 184 2515 218
rect 2549 184 2557 218
rect 2504 172 2557 184
rect 2168 -106 2221 -56
rect 2168 -140 2176 -106
rect 2210 -140 2221 -106
rect 1139 -204 1192 -166
rect 1139 -238 1147 -204
rect 1181 -238 1192 -204
rect 1139 -250 1192 -238
rect 1992 -204 2045 -166
rect 1992 -238 2003 -204
rect 2037 -238 2045 -204
rect 1992 -250 2045 -238
rect 2168 -174 2221 -140
rect 2168 -208 2176 -174
rect 2210 -208 2221 -174
rect 2168 -242 2221 -208
rect 2168 -276 2176 -242
rect 2210 -276 2221 -242
rect 2168 -310 2221 -276
rect 2168 -344 2176 -310
rect 2210 -344 2221 -310
rect 2168 -356 2221 -344
rect 2321 -106 2377 -56
rect 2321 -140 2332 -106
rect 2366 -140 2377 -106
rect 2321 -174 2377 -140
rect 2321 -208 2332 -174
rect 2366 -208 2377 -174
rect 2321 -242 2377 -208
rect 2321 -276 2332 -242
rect 2366 -276 2377 -242
rect 2321 -310 2377 -276
rect 2321 -344 2332 -310
rect 2366 -344 2377 -310
rect 2321 -356 2377 -344
rect 2477 -106 2533 -56
rect 2477 -140 2488 -106
rect 2522 -140 2533 -106
rect 2477 -174 2533 -140
rect 2477 -208 2488 -174
rect 2522 -208 2533 -174
rect 2477 -242 2533 -208
rect 2477 -276 2488 -242
rect 2522 -276 2533 -242
rect 2477 -310 2533 -276
rect 2477 -344 2488 -310
rect 2522 -344 2533 -310
rect 2477 -356 2533 -344
rect 2633 -106 2689 -56
rect 2633 -140 2644 -106
rect 2678 -140 2689 -106
rect 2633 -174 2689 -140
rect 2633 -208 2644 -174
rect 2678 -208 2689 -174
rect 2633 -242 2689 -208
rect 2633 -276 2644 -242
rect 2678 -276 2689 -242
rect 2633 -310 2689 -276
rect 2633 -344 2644 -310
rect 2678 -344 2689 -310
rect 2633 -356 2689 -344
rect 2789 -106 2842 -56
rect 2789 -140 2800 -106
rect 2834 -140 2842 -106
rect 2789 -174 2842 -140
rect 2789 -208 2800 -174
rect 2834 -208 2842 -174
rect 2789 -242 2842 -208
rect 2789 -276 2800 -242
rect 2834 -276 2842 -242
rect 2789 -310 2842 -276
rect 2789 -344 2800 -310
rect 2834 -344 2842 -310
rect 2789 -356 2842 -344
<< mvndiffc >>
rect 1356 -785 1390 -751
rect 1356 -853 1390 -819
rect 1356 -921 1390 -887
rect 1356 -989 1390 -955
rect 1356 -1057 1390 -1023
rect 1356 -1125 1390 -1091
rect 1356 -1193 1390 -1159
rect 1356 -1261 1390 -1227
rect 1532 -785 1566 -751
rect 1532 -853 1566 -819
rect 1532 -921 1566 -887
rect 1532 -989 1566 -955
rect 1532 -1057 1566 -1023
rect 1532 -1125 1566 -1091
rect 1532 -1193 1566 -1159
rect 1532 -1261 1566 -1227
rect 1708 -785 1742 -751
rect 1708 -853 1742 -819
rect 1708 -921 1742 -887
rect 1708 -989 1742 -955
rect 1708 -1057 1742 -1023
rect 1708 -1125 1742 -1091
rect 1708 -1193 1742 -1159
rect 1708 -1261 1742 -1227
rect 1884 -785 1918 -751
rect 1884 -853 1918 -819
rect 1884 -921 1918 -887
rect 1884 -989 1918 -955
rect 1884 -1057 1918 -1023
rect 1884 -1125 1918 -1091
rect 1884 -1193 1918 -1159
rect 1884 -1261 1918 -1227
rect 2060 -785 2094 -751
rect 2060 -853 2094 -819
rect 2060 -921 2094 -887
rect 2060 -989 2094 -955
rect 2060 -1057 2094 -1023
rect 2060 -1125 2094 -1091
rect 2060 -1193 2094 -1159
rect 2060 -1261 2094 -1227
rect 2236 -785 2270 -751
rect 2236 -853 2270 -819
rect 2236 -921 2270 -887
rect 2236 -989 2270 -955
rect 2236 -1057 2270 -1023
rect 2236 -1125 2270 -1091
rect 2236 -1193 2270 -1159
rect 2236 -1261 2270 -1227
rect 2412 -785 2446 -751
rect 2412 -853 2446 -819
rect 2412 -921 2446 -887
rect 2412 -989 2446 -955
rect 2412 -1057 2446 -1023
rect 2412 -1125 2446 -1091
rect 2412 -1193 2446 -1159
rect 2412 -1261 2446 -1227
rect 2588 -785 2622 -751
rect 2588 -853 2622 -819
rect 2588 -921 2622 -887
rect 2588 -989 2622 -955
rect 2588 -1057 2622 -1023
rect 2588 -1125 2622 -1091
rect 2588 -1193 2622 -1159
rect 2588 -1261 2622 -1227
<< mvpdiffc >>
rect 2654 604 2688 638
rect 1716 468 1750 502
rect 1872 468 1906 502
rect 2028 468 2062 502
rect 2152 468 2186 502
rect 2308 468 2342 502
rect 2464 468 2498 502
rect 2654 536 2688 570
rect 2654 468 2688 502
rect 2810 604 2844 638
rect 2810 536 2844 570
rect 2810 468 2844 502
rect 2966 604 3000 638
rect 2966 536 3000 570
rect 2966 468 3000 502
rect 1147 184 1181 218
rect 1603 184 1637 218
rect 2059 184 2093 218
rect 2515 184 2549 218
rect 2176 -140 2210 -106
rect 1147 -238 1181 -204
rect 2003 -238 2037 -204
rect 2176 -208 2210 -174
rect 2176 -276 2210 -242
rect 2176 -344 2210 -310
rect 2332 -140 2366 -106
rect 2332 -208 2366 -174
rect 2332 -276 2366 -242
rect 2332 -344 2366 -310
rect 2488 -140 2522 -106
rect 2488 -208 2522 -174
rect 2488 -276 2522 -242
rect 2488 -344 2522 -310
rect 2644 -140 2678 -106
rect 2644 -208 2678 -174
rect 2644 -276 2678 -242
rect 2644 -344 2678 -310
rect 2800 -140 2834 -106
rect 2800 -208 2834 -174
rect 2800 -276 2834 -242
rect 2800 -344 2834 -310
<< psubdiff >>
rect 1239 -733 1273 -709
rect 1239 -807 1273 -767
rect 1239 -881 1273 -841
rect 1239 -955 1273 -915
rect 1239 -1029 1273 -989
rect 1239 -1104 1273 -1063
rect 1239 -1179 1273 -1138
rect 1239 -1237 1273 -1213
<< mvnsubdiff >>
rect 3086 583 3120 607
rect 3086 515 3120 549
rect 3086 457 3120 481
<< psubdiffcont >>
rect 1239 -767 1273 -733
rect 1239 -841 1273 -807
rect 1239 -915 1273 -881
rect 1239 -989 1273 -955
rect 1239 -1063 1273 -1029
rect 1239 -1138 1273 -1104
rect 1239 -1213 1273 -1179
<< mvnsubdiffcont >>
rect 3086 549 3120 583
rect 3086 481 3120 515
<< poly >>
rect 2699 656 2799 688
rect 2855 656 2955 688
rect 1761 540 1861 572
rect 1917 540 2017 572
rect 2197 540 2297 572
rect 2353 540 2453 572
rect 1761 424 1861 456
rect 1917 424 2017 456
rect 2197 424 2297 456
rect 2353 424 2453 456
rect 2699 424 2799 456
rect 2855 424 2955 456
rect 1605 408 2017 424
rect 1605 374 1621 408
rect 1655 374 1690 408
rect 1724 374 1759 408
rect 1793 374 1828 408
rect 1862 374 1897 408
rect 1931 374 1967 408
rect 2001 374 2017 408
rect 1605 358 2017 374
rect 2164 408 2298 424
rect 2164 374 2180 408
rect 2214 374 2248 408
rect 2282 374 2298 408
rect 2164 358 2298 374
rect 2353 408 2487 424
rect 2353 374 2369 408
rect 2403 374 2437 408
rect 2471 374 2487 408
rect 2353 358 2487 374
rect 2699 408 2955 424
rect 2699 374 2715 408
rect 2749 374 2810 408
rect 2844 374 2905 408
rect 2939 374 2955 408
rect 2699 358 2955 374
rect 1192 256 1592 288
rect 1648 256 2048 288
rect 2104 256 2504 288
rect 1192 124 1592 172
rect 1192 90 1208 124
rect 1242 90 1291 124
rect 1325 90 1374 124
rect 1408 90 1458 124
rect 1492 90 1542 124
rect 1576 90 1592 124
rect 1192 18 1592 90
rect 1648 140 2048 172
rect 2104 140 2504 172
rect 1648 124 2504 140
rect 1648 90 1664 124
rect 1698 90 1734 124
rect 1768 90 1804 124
rect 1838 90 1874 124
rect 1908 90 1944 124
rect 1978 90 2014 124
rect 2048 90 2084 124
rect 2118 90 2153 124
rect 2187 90 2222 124
rect 2256 90 2291 124
rect 2325 90 2360 124
rect 2394 90 2429 124
rect 2463 90 2504 124
rect 1648 74 2504 90
rect 1192 -16 1372 18
rect 1406 -16 1450 18
rect 1484 -16 1529 18
rect 1563 -16 1592 18
rect 1192 -68 1592 -16
rect 2221 -56 2321 -24
rect 2377 -56 2477 -24
rect 2533 -56 2633 -24
rect 2689 -56 2789 -24
rect 1192 -84 1992 -68
rect 1192 -118 1208 -84
rect 1242 -118 1282 -84
rect 1316 -118 1356 -84
rect 1390 -118 1430 -84
rect 1464 -118 1504 -84
rect 1538 -118 1577 -84
rect 1611 -118 1650 -84
rect 1684 -118 1723 -84
rect 1757 -118 1796 -84
rect 1830 -118 1869 -84
rect 1903 -118 1942 -84
rect 1976 -118 1992 -84
rect 1192 -166 1992 -118
rect 1192 -298 1992 -250
rect 1192 -332 1252 -298
rect 1286 -332 1321 -298
rect 1355 -332 1390 -298
rect 1424 -332 1459 -298
rect 1493 -332 1528 -298
rect 1562 -332 1597 -298
rect 1631 -332 1666 -298
rect 1700 -332 1735 -298
rect 1769 -332 1804 -298
rect 1838 -332 1873 -298
rect 1907 -332 1942 -298
rect 1976 -332 1992 -298
rect 1192 -348 1992 -332
rect 2221 -413 2321 -356
rect 2221 -447 2254 -413
rect 2288 -447 2321 -413
rect 2221 -481 2321 -447
rect 2221 -515 2254 -481
rect 2288 -515 2321 -481
rect 2221 -531 2321 -515
rect 2377 -413 2477 -356
rect 2377 -447 2413 -413
rect 2447 -447 2477 -413
rect 2377 -481 2477 -447
rect 2533 -388 2633 -356
rect 2689 -388 2789 -356
rect 2533 -404 2789 -388
rect 2533 -438 2549 -404
rect 2583 -438 2644 -404
rect 2678 -438 2739 -404
rect 2773 -438 2789 -404
rect 2533 -454 2789 -438
rect 2377 -515 2413 -481
rect 2447 -515 2477 -481
rect 2377 -531 2477 -515
rect 1401 -591 1697 -575
rect 1401 -625 1417 -591
rect 1451 -625 1493 -591
rect 1527 -625 1570 -591
rect 1604 -625 1647 -591
rect 1681 -625 1697 -591
rect 1401 -641 1697 -625
rect 1401 -673 1521 -641
rect 1577 -673 1697 -641
rect 1753 -591 2577 -575
rect 1753 -625 1769 -591
rect 1803 -625 1837 -591
rect 1871 -625 1906 -591
rect 1940 -625 1975 -591
rect 2009 -625 2044 -591
rect 2078 -625 2113 -591
rect 2147 -625 2182 -591
rect 2216 -625 2251 -591
rect 2285 -625 2320 -591
rect 2354 -625 2389 -591
rect 2423 -625 2458 -591
rect 2492 -625 2527 -591
rect 2561 -625 2577 -591
rect 1753 -641 2577 -625
rect 1753 -673 1873 -641
rect 1929 -673 2049 -641
rect 2105 -673 2225 -641
rect 2281 -673 2401 -641
rect 2457 -673 2577 -641
rect 1401 -1305 1521 -1273
rect 1577 -1305 1697 -1273
rect 1753 -1305 1873 -1273
rect 1929 -1305 2049 -1273
rect 2105 -1305 2225 -1273
rect 2281 -1305 2401 -1273
rect 2457 -1305 2577 -1273
<< polycont >>
rect 1621 374 1655 408
rect 1690 374 1724 408
rect 1759 374 1793 408
rect 1828 374 1862 408
rect 1897 374 1931 408
rect 1967 374 2001 408
rect 2180 374 2214 408
rect 2248 374 2282 408
rect 2369 374 2403 408
rect 2437 374 2471 408
rect 2715 374 2749 408
rect 2810 374 2844 408
rect 2905 374 2939 408
rect 1208 90 1242 124
rect 1291 90 1325 124
rect 1374 90 1408 124
rect 1458 90 1492 124
rect 1542 90 1576 124
rect 1664 90 1698 124
rect 1734 90 1768 124
rect 1804 90 1838 124
rect 1874 90 1908 124
rect 1944 90 1978 124
rect 2014 90 2048 124
rect 2084 90 2118 124
rect 2153 90 2187 124
rect 2222 90 2256 124
rect 2291 90 2325 124
rect 2360 90 2394 124
rect 2429 90 2463 124
rect 1372 -16 1406 18
rect 1450 -16 1484 18
rect 1529 -16 1563 18
rect 1208 -118 1242 -84
rect 1282 -118 1316 -84
rect 1356 -118 1390 -84
rect 1430 -118 1464 -84
rect 1504 -118 1538 -84
rect 1577 -118 1611 -84
rect 1650 -118 1684 -84
rect 1723 -118 1757 -84
rect 1796 -118 1830 -84
rect 1869 -118 1903 -84
rect 1942 -118 1976 -84
rect 1252 -332 1286 -298
rect 1321 -332 1355 -298
rect 1390 -332 1424 -298
rect 1459 -332 1493 -298
rect 1528 -332 1562 -298
rect 1597 -332 1631 -298
rect 1666 -332 1700 -298
rect 1735 -332 1769 -298
rect 1804 -332 1838 -298
rect 1873 -332 1907 -298
rect 1942 -332 1976 -298
rect 2254 -447 2288 -413
rect 2254 -515 2288 -481
rect 2413 -447 2447 -413
rect 2549 -438 2583 -404
rect 2644 -438 2678 -404
rect 2739 -438 2773 -404
rect 2413 -515 2447 -481
rect 1417 -625 1451 -591
rect 1493 -625 1527 -591
rect 1570 -625 1604 -591
rect 1647 -625 1681 -591
rect 1769 -625 1803 -591
rect 1837 -625 1871 -591
rect 1906 -625 1940 -591
rect 1975 -625 2009 -591
rect 2044 -625 2078 -591
rect 2113 -625 2147 -591
rect 2182 -625 2216 -591
rect 2251 -625 2285 -591
rect 2320 -625 2354 -591
rect 2389 -625 2423 -591
rect 2458 -625 2492 -591
rect 2527 -625 2561 -591
<< locali >>
rect 2654 638 2688 654
rect 1871 579 1909 613
rect 2151 579 2189 613
rect 2459 579 2497 613
rect 2652 604 2654 613
rect 2810 638 2844 654
rect 2688 604 2690 613
rect 2652 579 2690 604
rect 2966 638 3000 654
rect 1714 502 1752 523
rect 1714 489 1716 502
rect 1750 489 1752 502
rect 1872 502 1906 579
rect 1716 452 1750 468
rect 2026 502 2064 523
rect 2026 489 2028 502
rect 1872 452 1906 468
rect 2062 489 2064 502
rect 2152 502 2186 579
rect 2028 452 2062 468
rect 2308 502 2346 523
rect 2152 452 2186 468
rect 2342 489 2346 502
rect 2464 502 2498 579
rect 2308 452 2342 468
rect 2464 452 2498 468
rect 2654 570 2688 579
rect 2654 502 2688 536
rect 2810 570 2844 604
rect 2964 604 2966 613
rect 3000 604 3002 613
rect 2964 579 3002 604
rect 3086 583 3120 607
rect 2810 523 2844 536
rect 2966 570 3000 579
rect 2808 502 2846 523
rect 2808 489 2810 502
rect 2654 452 2688 468
rect 2844 489 2846 502
rect 2966 502 3000 536
rect 2810 452 2844 468
rect 2966 452 3000 468
rect 3086 523 3120 549
rect 3086 515 3094 523
rect 3128 489 3166 523
rect 3086 457 3120 481
rect 1605 374 1621 408
rect 1655 374 1690 408
rect 1724 374 1759 408
rect 1793 374 1828 408
rect 1862 374 1897 408
rect 1931 374 1967 408
rect 2001 374 2017 408
rect 2164 403 2180 408
rect 2214 374 2248 408
rect 2282 403 2298 408
rect 2295 374 2298 403
rect 2353 374 2369 408
rect 2403 407 2437 408
rect 2471 407 2487 408
rect 2403 374 2434 407
rect 2471 374 2506 407
rect 1151 266 1189 300
rect 1117 218 1223 266
rect 1117 184 1147 218
rect 1181 184 1223 218
rect 1117 168 1223 184
rect 1603 218 1637 234
rect 1603 168 1637 184
rect 1711 124 1909 374
rect 2186 369 2261 374
rect 2468 373 2506 374
rect 2699 374 2715 408
rect 2749 403 2810 408
rect 2844 403 2905 408
rect 2755 374 2810 403
rect 2755 369 2811 374
rect 2845 369 2900 403
rect 2939 374 2955 408
rect 2025 264 2063 298
rect 2643 264 2681 298
rect 2059 218 2093 264
rect 2059 168 2093 184
rect 2515 218 2579 234
rect 2549 184 2579 218
rect 1192 90 1208 124
rect 1242 90 1291 124
rect 1325 90 1374 124
rect 1408 90 1458 124
rect 1492 90 1542 124
rect 1576 90 1592 124
rect 1648 90 1656 124
rect 1698 90 1734 124
rect 1768 90 1804 124
rect 1846 90 1874 124
rect 1924 90 1944 124
rect 2002 90 2014 124
rect 2080 90 2084 124
rect 2118 90 2124 124
rect 2187 90 2203 124
rect 2256 90 2282 124
rect 2325 90 2360 124
rect 2395 90 2429 124
rect 2474 90 2479 124
rect 1325 18 1592 90
rect 2515 56 2579 184
rect 1325 -16 1372 18
rect 1406 -16 1450 18
rect 1484 -16 1529 18
rect 1563 -16 1592 18
rect 1325 -38 1592 -16
rect 2029 -1 2579 56
rect 1325 -72 1338 -38
rect 1372 -72 1419 -38
rect 1453 -72 1500 -38
rect 1534 -72 1581 -38
rect 1615 -72 1697 -57
rect 1325 -84 1697 -72
rect 1192 -118 1208 -84
rect 1242 -118 1282 -84
rect 1316 -118 1356 -84
rect 1390 -118 1430 -84
rect 1464 -118 1504 -84
rect 1538 -118 1577 -84
rect 1611 -118 1650 -84
rect 1684 -118 1723 -84
rect 1757 -118 1796 -84
rect 1830 -118 1869 -84
rect 1903 -118 1942 -84
rect 1976 -118 1992 -84
rect 1325 -120 1697 -118
rect 1325 -154 1338 -120
rect 1372 -154 1419 -120
rect 1453 -154 1500 -120
rect 1534 -154 1581 -120
rect 1615 -154 1697 -120
rect 1147 -204 1181 -188
rect 1147 -288 1181 -250
rect 1325 -298 1697 -154
rect 2029 -188 2095 -1
rect 2003 -204 2095 -188
rect 2037 -238 2095 -204
rect 2003 -254 2095 -238
rect 2144 -106 2250 -90
rect 2144 -135 2176 -106
rect 2210 -135 2250 -106
rect 2210 -140 2216 -135
rect 2178 -169 2216 -140
rect 2144 -174 2250 -169
rect 2144 -208 2176 -174
rect 2210 -208 2250 -174
rect 2144 -242 2250 -208
rect 2144 -276 2176 -242
rect 2210 -276 2250 -242
rect 1236 -332 1252 -298
rect 1286 -332 1321 -298
rect 1355 -332 1390 -298
rect 1424 -332 1459 -298
rect 1493 -332 1528 -298
rect 1562 -332 1597 -298
rect 1631 -332 1666 -298
rect 1700 -332 1735 -298
rect 1769 -332 1804 -298
rect 1838 -332 1873 -298
rect 1907 -332 1942 -298
rect 1976 -332 1992 -298
rect 2144 -310 2250 -276
rect 1401 -591 1697 -332
rect 2144 -344 2176 -310
rect 2210 -344 2250 -310
rect 2144 -360 2250 -344
rect 2332 -106 2366 -90
rect 2332 -174 2366 -140
rect 2332 -217 2366 -208
rect 2332 -289 2366 -276
rect 2332 -360 2366 -344
rect 2488 -106 2522 -90
rect 2488 -174 2522 -140
rect 2488 -242 2522 -208
rect 2488 -310 2522 -276
rect 2488 -360 2522 -344
rect 2644 -106 2704 264
rect 2678 -140 2704 -106
rect 2644 -174 2704 -140
rect 2678 -208 2704 -174
rect 2644 -242 2704 -208
rect 2678 -276 2704 -242
rect 2644 -310 2704 -276
rect 2678 -344 2704 -310
rect 2644 -361 2704 -344
rect 2739 -106 2845 -90
rect 2739 -135 2800 -106
rect 2834 -135 2845 -106
rect 2773 -140 2800 -135
rect 2773 -169 2811 -140
rect 2739 -174 2845 -169
rect 2739 -208 2800 -174
rect 2834 -208 2845 -174
rect 2739 -242 2845 -208
rect 2739 -276 2800 -242
rect 2834 -276 2845 -242
rect 2739 -310 2845 -276
rect 2739 -344 2800 -310
rect 2834 -344 2845 -310
rect 2739 -360 2845 -344
rect 2254 -413 2288 -397
rect 2383 -413 2489 -397
rect 2383 -443 2413 -413
rect 2447 -443 2489 -413
rect 2254 -479 2267 -447
rect 2254 -481 2301 -479
rect 2288 -515 2301 -481
rect 2254 -517 2301 -515
rect 2254 -531 2267 -517
rect 2447 -447 2455 -443
rect 2417 -477 2455 -447
rect 2383 -481 2489 -477
rect 2383 -515 2413 -481
rect 2447 -515 2489 -481
rect 2383 -531 2489 -515
rect 2533 -438 2549 -404
rect 2583 -438 2644 -404
rect 2678 -438 2739 -404
rect 2773 -438 2789 -404
rect 2533 -439 2789 -438
rect 2533 -473 2587 -439
rect 2621 -473 2660 -439
rect 2694 -473 2733 -439
rect 2767 -473 2789 -439
rect 2533 -591 2789 -473
rect 1401 -625 1417 -591
rect 1451 -625 1493 -591
rect 1527 -625 1570 -591
rect 1604 -625 1647 -591
rect 1681 -625 1697 -591
rect 1753 -625 1769 -591
rect 1803 -625 1837 -591
rect 1871 -625 1906 -591
rect 1940 -625 1975 -591
rect 2009 -625 2044 -591
rect 2078 -625 2113 -591
rect 2147 -625 2182 -591
rect 2216 -625 2251 -591
rect 2285 -625 2320 -591
rect 2354 -625 2389 -591
rect 2423 -625 2458 -591
rect 2492 -625 2527 -591
rect 2561 -625 2789 -591
rect 1239 -733 1356 -709
rect 1273 -735 1356 -733
rect 1273 -741 1390 -735
rect 1273 -767 1356 -741
rect 1239 -785 1356 -767
rect 1239 -807 1390 -785
rect 1273 -813 1390 -807
rect 1273 -841 1356 -813
rect 1239 -853 1356 -841
rect 1239 -881 1390 -853
rect 1273 -885 1390 -881
rect 1273 -915 1356 -885
rect 1239 -921 1356 -915
rect 1239 -955 1390 -921
rect 1273 -989 1356 -955
rect 1239 -1023 1390 -989
rect 1239 -1029 1356 -1023
rect 1273 -1057 1356 -1029
rect 1273 -1063 1390 -1057
rect 1239 -1091 1390 -1063
rect 1239 -1104 1356 -1091
rect 1273 -1125 1356 -1104
rect 1273 -1138 1390 -1125
rect 1239 -1159 1390 -1138
rect 1239 -1179 1356 -1159
rect 1273 -1193 1356 -1179
rect 1273 -1213 1390 -1193
rect 1239 -1227 1390 -1213
rect 1239 -1237 1356 -1227
rect 1356 -1277 1390 -1261
rect 1488 -751 1600 -735
rect 1488 -785 1532 -751
rect 1566 -785 1600 -751
rect 1488 -819 1600 -785
rect 1488 -853 1532 -819
rect 1566 -853 1600 -819
rect 1488 -887 1600 -853
rect 1488 -921 1532 -887
rect 1566 -921 1600 -887
rect 1488 -955 1600 -921
rect 1488 -965 1532 -955
rect 1488 -999 1494 -965
rect 1528 -989 1532 -965
rect 1566 -965 1600 -955
rect 1528 -999 1566 -989
rect 1488 -1023 1600 -999
rect 1488 -1057 1532 -1023
rect 1566 -1057 1600 -1023
rect 1488 -1091 1600 -1057
rect 1488 -1125 1532 -1091
rect 1566 -1125 1600 -1091
rect 1488 -1159 1600 -1125
rect 1488 -1193 1532 -1159
rect 1566 -1193 1600 -1159
rect 1488 -1227 1600 -1193
rect 1488 -1261 1532 -1227
rect 1566 -1261 1600 -1227
rect 1488 -1277 1600 -1261
rect 1708 -741 1742 -735
rect 1708 -813 1742 -785
rect 1708 -885 1742 -853
rect 1708 -955 1742 -921
rect 1708 -1023 1742 -989
rect 1708 -1091 1742 -1057
rect 1708 -1159 1742 -1125
rect 1708 -1227 1742 -1193
rect 1708 -1277 1742 -1261
rect 1835 -751 1947 -735
rect 1835 -785 1884 -751
rect 1918 -785 1947 -751
rect 1835 -819 1947 -785
rect 1835 -853 1884 -819
rect 1918 -853 1947 -819
rect 1835 -887 1947 -853
rect 1835 -921 1884 -887
rect 1918 -921 1947 -887
rect 1835 -955 1947 -921
rect 1835 -965 1884 -955
rect 1918 -965 1947 -955
rect 1869 -989 1884 -965
rect 1869 -999 1913 -989
rect 1835 -1023 1947 -999
rect 1835 -1057 1884 -1023
rect 1918 -1057 1947 -1023
rect 1835 -1091 1947 -1057
rect 1835 -1125 1884 -1091
rect 1918 -1125 1947 -1091
rect 1835 -1159 1947 -1125
rect 1835 -1193 1884 -1159
rect 1918 -1193 1947 -1159
rect 1835 -1227 1947 -1193
rect 1835 -1261 1884 -1227
rect 1918 -1261 1947 -1227
rect 1835 -1277 1947 -1261
rect 2060 -741 2094 -735
rect 2060 -813 2094 -785
rect 2060 -885 2094 -853
rect 2060 -955 2094 -921
rect 2236 -751 2270 -735
rect 2236 -819 2270 -785
rect 2236 -887 2270 -853
rect 2236 -955 2270 -921
rect 2060 -1023 2094 -989
rect 2232 -989 2236 -965
rect 2412 -741 2446 -735
rect 2412 -813 2446 -785
rect 2412 -885 2446 -853
rect 2412 -955 2446 -921
rect 2232 -999 2270 -989
rect 2588 -751 2622 -735
rect 2588 -819 2622 -785
rect 2588 -887 2622 -853
rect 2588 -955 2622 -921
rect 2060 -1091 2094 -1057
rect 2060 -1159 2094 -1125
rect 2060 -1227 2094 -1193
rect 2060 -1277 2094 -1261
rect 2236 -1023 2270 -999
rect 2236 -1091 2270 -1057
rect 2236 -1159 2270 -1125
rect 2236 -1227 2270 -1193
rect 2236 -1277 2270 -1261
rect 2412 -1023 2446 -989
rect 2530 -999 2568 -965
rect 2602 -999 2622 -989
rect 2412 -1091 2446 -1057
rect 2412 -1159 2446 -1125
rect 2412 -1227 2446 -1193
rect 2412 -1277 2446 -1261
rect 2588 -1023 2622 -999
rect 2588 -1091 2622 -1057
rect 2588 -1159 2622 -1125
rect 2588 -1227 2622 -1193
rect 2588 -1277 2622 -1261
<< viali >>
rect 1837 579 1871 613
rect 1909 579 1943 613
rect 2117 579 2151 613
rect 2189 579 2223 613
rect 2425 579 2459 613
rect 2497 579 2531 613
rect 2618 579 2652 613
rect 2690 579 2724 613
rect 1680 489 1714 523
rect 1752 489 1786 523
rect 1992 489 2026 523
rect 2064 489 2098 523
rect 2274 489 2308 523
rect 2346 489 2380 523
rect 2930 579 2964 613
rect 3002 579 3036 613
rect 2774 489 2808 523
rect 2846 489 2880 523
rect 3094 515 3128 523
rect 3094 489 3120 515
rect 3120 489 3128 515
rect 3166 489 3200 523
rect 2152 374 2180 403
rect 2180 374 2186 403
rect 2261 374 2282 403
rect 2282 374 2295 403
rect 2434 374 2437 407
rect 2437 374 2468 407
rect 1117 266 1151 300
rect 1189 266 1223 300
rect 2152 369 2186 374
rect 2261 369 2295 374
rect 2434 373 2468 374
rect 2506 373 2540 407
rect 2721 374 2749 403
rect 2749 374 2755 403
rect 2811 374 2844 403
rect 2844 374 2845 403
rect 2721 369 2755 374
rect 2811 369 2845 374
rect 2900 374 2905 403
rect 2905 374 2934 403
rect 2900 369 2934 374
rect 1991 264 2025 298
rect 2063 264 2097 298
rect 2609 264 2643 298
rect 2681 264 2715 298
rect 1656 90 1664 124
rect 1664 90 1690 124
rect 1734 90 1768 124
rect 1812 90 1838 124
rect 1838 90 1846 124
rect 1890 90 1908 124
rect 1908 90 1924 124
rect 1968 90 1978 124
rect 1978 90 2002 124
rect 2046 90 2048 124
rect 2048 90 2080 124
rect 2124 90 2153 124
rect 2153 90 2158 124
rect 2203 90 2222 124
rect 2222 90 2237 124
rect 2282 90 2291 124
rect 2291 90 2316 124
rect 2361 90 2394 124
rect 2394 90 2395 124
rect 2440 90 2463 124
rect 2463 90 2474 124
rect 1338 -72 1372 -38
rect 1419 -72 1453 -38
rect 1500 -72 1534 -38
rect 1581 -72 1615 -38
rect 1338 -154 1372 -120
rect 1419 -154 1453 -120
rect 1500 -154 1534 -120
rect 1581 -154 1615 -120
rect 1147 -238 1181 -216
rect 1147 -250 1181 -238
rect 1147 -322 1181 -288
rect 2144 -140 2176 -135
rect 2176 -140 2178 -135
rect 2144 -169 2178 -140
rect 2216 -169 2250 -135
rect 2332 -242 2366 -217
rect 2332 -251 2366 -242
rect 2332 -310 2366 -289
rect 2332 -323 2366 -310
rect 2739 -169 2773 -135
rect 2811 -140 2834 -135
rect 2834 -140 2845 -135
rect 2811 -169 2845 -140
rect 2267 -447 2288 -445
rect 2288 -447 2301 -445
rect 2267 -479 2301 -447
rect 2267 -551 2301 -517
rect 2383 -447 2413 -443
rect 2413 -447 2417 -443
rect 2383 -477 2417 -447
rect 2455 -477 2489 -443
rect 2587 -473 2621 -439
rect 2660 -473 2694 -439
rect 2733 -473 2767 -439
rect 1356 -751 1390 -741
rect 1356 -775 1390 -751
rect 1356 -819 1390 -813
rect 1356 -847 1390 -819
rect 1356 -887 1390 -885
rect 1356 -919 1390 -887
rect 1494 -999 1528 -965
rect 1566 -999 1600 -965
rect 1708 -751 1742 -741
rect 1708 -775 1742 -751
rect 1708 -819 1742 -813
rect 1708 -847 1742 -819
rect 1708 -887 1742 -885
rect 1708 -919 1742 -887
rect 1835 -999 1869 -965
rect 1913 -989 1918 -965
rect 1918 -989 1947 -965
rect 1913 -999 1947 -989
rect 2060 -751 2094 -741
rect 2060 -775 2094 -751
rect 2060 -819 2094 -813
rect 2060 -847 2094 -819
rect 2060 -887 2094 -885
rect 2060 -919 2094 -887
rect 2198 -999 2232 -965
rect 2412 -751 2446 -741
rect 2412 -775 2446 -751
rect 2412 -819 2446 -813
rect 2412 -847 2446 -819
rect 2412 -887 2446 -885
rect 2412 -919 2446 -887
rect 2270 -999 2304 -965
rect 2496 -999 2530 -965
rect 2568 -989 2588 -965
rect 2588 -989 2602 -965
rect 2568 -999 2602 -989
<< metal1 >>
rect 1167 623 1173 675
rect 1225 623 1237 675
rect 1289 647 2037 675
rect 1289 623 1295 647
tri 1295 623 1319 647 nw
tri 1999 623 2023 647 ne
rect 2023 623 2037 647
tri 2037 623 2089 675 sw
tri 2023 619 2027 623 ne
rect 2027 619 2089 623
tri 2089 619 2093 623 sw
rect 1819 567 1825 619
rect 1877 567 1889 619
rect 1941 613 1955 619
tri 2027 613 2033 619 ne
rect 2033 613 3048 619
rect 1943 579 1955 613
tri 2033 609 2037 613 ne
rect 2037 609 2117 613
tri 2037 579 2067 609 ne
rect 2067 579 2117 609
rect 2151 579 2189 613
rect 2223 579 2425 613
rect 2459 579 2497 613
rect 2531 579 2618 613
rect 2652 579 2690 613
rect 2724 579 2930 613
rect 2964 579 3002 613
rect 3036 579 3048 613
rect 1941 567 1955 579
tri 2067 573 2073 579 ne
rect 2073 573 3048 579
rect 1668 523 2392 529
rect 1668 489 1680 523
rect 1714 489 1752 523
rect 1786 489 1992 523
rect 2026 489 2064 523
rect 2098 489 2274 523
rect 2308 489 2346 523
rect 2380 489 2392 523
rect 1668 483 2392 489
rect 2762 523 3212 529
rect 2762 489 2774 523
rect 2808 489 2846 523
rect 2880 489 3094 523
rect 3128 489 3166 523
rect 3200 489 3212 523
rect 2762 483 3212 489
rect 2140 403 2262 415
rect 2140 369 2152 403
rect 2186 369 2261 403
rect 2140 363 2262 369
rect 2314 363 2326 415
rect 2378 363 2384 415
tri 3470 413 3472 415 se
rect 2415 361 2421 413
rect 2473 361 2485 413
rect 2537 407 2552 413
tri 3466 409 3470 413 se
rect 3470 409 3472 413
rect 2540 373 2552 407
rect 2537 363 2552 373
rect 2709 403 3472 409
rect 2709 369 2721 403
rect 2755 369 2811 403
rect 2845 369 2900 403
rect 2934 369 3472 403
rect 2709 363 3472 369
rect 2537 361 2543 363
tri 2543 361 2545 363 nw
tri 1161 306 1167 312 se
rect 1167 306 1173 312
rect 1105 300 1173 306
rect 1105 266 1117 300
rect 1151 266 1173 300
rect 1105 260 1173 266
rect 1225 260 1237 312
rect 1289 260 1295 312
rect 1819 258 1825 310
rect 1877 258 1889 310
rect 1941 304 1947 310
tri 1947 304 1953 310 sw
rect 1941 298 2727 304
rect 1941 264 1991 298
rect 2025 264 2063 298
rect 2097 264 2609 298
rect 2643 264 2681 298
rect 2715 264 2727 298
rect 1941 258 2727 264
rect 1644 124 2581 130
rect 1644 90 1656 124
rect 1690 90 1734 124
rect 1768 90 1812 124
rect 1846 90 1890 124
rect 1924 90 1968 124
rect 2002 90 2046 124
rect 2080 90 2124 124
rect 2158 90 2203 124
rect 2237 90 2282 124
rect 2316 90 2361 124
rect 2395 90 2440 124
rect 2474 90 2581 124
rect 1644 84 2581 90
tri 2569 78 2575 84 ne
rect 2575 78 2581 84
rect 2633 78 2646 130
rect 2698 78 2704 130
rect 1326 -38 1627 -32
rect 1326 -72 1338 -38
rect 1372 -72 1419 -38
rect 1453 -72 1500 -38
rect 1534 -72 1581 -38
rect 1615 -72 1627 -38
rect 1326 -120 1627 -72
rect 1326 -154 1338 -120
rect 1372 -154 1419 -120
rect 1453 -154 1500 -120
rect 1534 -154 1581 -120
rect 1615 -154 1627 -120
rect 1326 -160 1627 -154
rect 2132 -135 2857 -129
rect 2132 -169 2144 -135
rect 2178 -169 2216 -135
rect 2250 -169 2739 -135
rect 2773 -169 2811 -135
rect 2845 -169 2857 -135
rect 2132 -175 2857 -169
rect 1141 -205 2326 -204
rect 1141 -216 2372 -205
rect 1141 -250 1147 -216
rect 1181 -217 2372 -216
rect 1181 -250 2332 -217
rect 1141 -251 2332 -250
rect 2366 -251 2372 -217
rect 1141 -288 2372 -251
rect 1141 -322 1147 -288
rect 1181 -289 2372 -288
rect 1181 -322 2332 -289
rect 1141 -323 2332 -322
rect 2366 -323 2372 -289
rect 1141 -334 2372 -323
rect 2326 -335 2372 -334
rect 2256 -439 2308 -433
rect 2371 -485 2381 -433
rect 2433 -485 2445 -433
rect 2497 -485 2503 -433
rect 2575 -485 2581 -433
rect 2633 -485 2651 -433
rect 2703 -485 2721 -433
rect 2773 -485 2779 -433
rect 2256 -503 2308 -491
rect 2256 -561 2308 -555
rect 2261 -563 2307 -561
rect 1350 -741 2452 -729
rect 1350 -775 1356 -741
rect 1390 -775 1708 -741
rect 1742 -775 2060 -741
rect 2094 -775 2412 -741
rect 2446 -775 2452 -741
rect 1350 -813 2452 -775
rect 1350 -847 1356 -813
rect 1390 -847 1708 -813
rect 1742 -847 2060 -813
rect 2094 -847 2412 -813
rect 2446 -847 2452 -813
rect 1350 -885 2452 -847
rect 1350 -919 1356 -885
rect 1390 -919 1708 -885
rect 1742 -919 2060 -885
rect 2094 -919 2412 -885
rect 2446 -919 2452 -885
rect 1350 -931 2452 -919
rect 1470 -965 2615 -959
rect 1470 -999 1494 -965
rect 1528 -999 1566 -965
rect 1600 -999 1835 -965
rect 1869 -999 1913 -965
rect 1947 -999 1957 -965
rect 1470 -1005 1957 -999
tri 1905 -1057 1957 -1005 ne
rect 2009 -999 2198 -965
rect 2232 -999 2270 -965
rect 2304 -999 2496 -965
rect 2530 -999 2568 -965
rect 2602 -999 2615 -965
rect 2009 -1005 2615 -999
rect 1957 -1036 2009 -1017
tri 2009 -1057 2061 -1005 nw
rect 1957 -1094 2009 -1088
<< via1 >>
rect 1173 623 1225 675
rect 1237 623 1289 675
rect 1825 613 1877 619
rect 1825 579 1837 613
rect 1837 579 1871 613
rect 1871 579 1877 613
rect 1825 567 1877 579
rect 1889 613 1941 619
rect 1889 579 1909 613
rect 1909 579 1941 613
rect 1889 567 1941 579
rect 2262 403 2314 415
rect 2262 369 2295 403
rect 2295 369 2314 403
rect 2262 363 2314 369
rect 2326 363 2378 415
rect 2421 407 2473 413
rect 2421 373 2434 407
rect 2434 373 2468 407
rect 2468 373 2473 407
rect 2421 361 2473 373
rect 2485 407 2537 413
rect 2485 373 2506 407
rect 2506 373 2537 407
rect 2485 361 2537 373
rect 1173 300 1225 312
rect 1173 266 1189 300
rect 1189 266 1223 300
rect 1223 266 1225 300
rect 1173 260 1225 266
rect 1237 260 1289 312
rect 1825 258 1877 310
rect 1889 258 1941 310
rect 2581 78 2633 130
rect 2646 78 2698 130
rect 2256 -445 2308 -439
rect 2256 -479 2267 -445
rect 2267 -479 2301 -445
rect 2301 -479 2308 -445
rect 2256 -491 2308 -479
rect 2381 -443 2433 -433
rect 2381 -477 2383 -443
rect 2383 -477 2417 -443
rect 2417 -477 2433 -443
rect 2381 -485 2433 -477
rect 2445 -443 2497 -433
rect 2445 -477 2455 -443
rect 2455 -477 2489 -443
rect 2489 -477 2497 -443
rect 2445 -485 2497 -477
rect 2581 -439 2633 -433
rect 2581 -473 2587 -439
rect 2587 -473 2621 -439
rect 2621 -473 2633 -439
rect 2581 -485 2633 -473
rect 2651 -439 2703 -433
rect 2651 -473 2660 -439
rect 2660 -473 2694 -439
rect 2694 -473 2703 -439
rect 2651 -485 2703 -473
rect 2721 -439 2773 -433
rect 2721 -473 2733 -439
rect 2733 -473 2767 -439
rect 2767 -473 2773 -439
rect 2721 -485 2773 -473
rect 2256 -517 2308 -503
rect 2256 -551 2267 -517
rect 2267 -551 2301 -517
rect 2301 -551 2308 -517
rect 2256 -555 2308 -551
rect 1957 -1017 2009 -965
rect 1957 -1088 2009 -1036
<< metal2 >>
rect 1167 623 1173 675
rect 1225 623 1237 675
rect 1289 623 1295 675
tri 1211 619 1215 623 ne
rect 1215 619 1295 623
tri 1215 585 1249 619 ne
tri 1234 363 1249 378 se
rect 1249 363 1295 619
tri 1232 361 1234 363 se
rect 1234 361 1295 363
tri 1183 312 1232 361 se
rect 1232 312 1295 361
rect 1167 260 1173 312
rect 1225 260 1237 312
rect 1289 260 1295 312
rect 1819 567 1825 619
rect 1877 567 1889 619
rect 1941 567 1947 619
rect 1819 310 1947 567
rect 1819 258 1825 310
rect 1877 258 1889 310
rect 1941 258 1947 310
rect 1819 -596 1868 258
tri 1868 179 1947 258 nw
rect 2256 363 2262 415
rect 2314 363 2326 415
rect 2378 363 2384 415
rect 2256 361 2343 363
tri 2343 361 2345 363 nw
rect 2415 361 2421 413
rect 2473 361 2485 413
rect 2537 361 2543 413
rect 2256 -439 2308 361
tri 2308 326 2343 361 nw
rect 2256 -503 2308 -491
tri 2375 -433 2415 -393 se
rect 2415 -433 2467 361
tri 2467 305 2523 361 nw
rect 2575 78 2581 130
rect 2633 78 2646 130
rect 2698 78 2704 130
rect 2575 -397 2628 78
tri 2628 40 2666 78 nw
tri 2628 -397 2649 -376 sw
tri 2467 -433 2503 -397 sw
rect 2375 -485 2381 -433
rect 2433 -485 2445 -433
rect 2497 -485 2503 -433
rect 2575 -433 2649 -397
tri 2649 -433 2685 -397 sw
rect 2575 -485 2581 -433
rect 2633 -485 2651 -433
rect 2703 -485 2721 -433
rect 2773 -485 2779 -433
tri 2375 -525 2415 -485 ne
rect 2458 -525 2463 -485
tri 2463 -525 2503 -485 nw
tri 2458 -530 2463 -525 nw
rect 2256 -561 2308 -555
tri 1819 -638 1861 -596 ne
rect 1861 -638 1868 -596
tri 1868 -638 1935 -571 sw
tri 1861 -645 1868 -638 ne
rect 1868 -645 1935 -638
tri 1868 -712 1935 -645 ne
tri 1935 -712 2009 -638 sw
tri 1935 -734 1957 -712 ne
rect 1957 -965 2009 -712
rect 1957 -1036 2009 -1017
rect 1957 -1094 2009 -1088
use sky130_fd_pr__nfet_01v8__example_55959141808637  sky130_fd_pr__nfet_01v8__example_55959141808637_0
timestamp 1666199351
transform 1 0 1401 0 1 -1273
box -1 0 297 1
use sky130_fd_pr__nfet_01v8__example_55959141808638  sky130_fd_pr__nfet_01v8__example_55959141808638_0
timestamp 1666199351
transform 1 0 1753 0 1 -1273
box -1 0 825 1
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_0
timestamp 1666199351
transform 1 0 2377 0 1 -356
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_1
timestamp 1666199351
transform 1 0 2533 0 1 -356
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_2
timestamp 1666199351
transform -1 0 2789 0 1 -356
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_3
timestamp 1666199351
transform -1 0 2321 0 1 -356
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808630  sky130_fd_pr__pfet_01v8__example_55959141808630_0
timestamp 1666199351
transform 1 0 1192 0 1 -250
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808632  sky130_fd_pr__pfet_01v8__example_55959141808632_0
timestamp 1666199351
transform -1 0 2017 0 1 456
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808634  sky130_fd_pr__pfet_01v8__example_55959141808634_0
timestamp 1666199351
transform 1 0 2197 0 1 456
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808634  sky130_fd_pr__pfet_01v8__example_55959141808634_1
timestamp 1666199351
transform -1 0 2453 0 1 456
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808635  sky130_fd_pr__pfet_01v8__example_55959141808635_0
timestamp 1666199351
transform 1 0 2699 0 1 456
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808636  sky130_fd_pr__pfet_01v8__example_55959141808636_0
timestamp 1666199351
transform 1 0 1192 0 1 172
box -1 0 401 1
use sky130_fd_pr__pfet_01v8__example_55959141808636  sky130_fd_pr__pfet_01v8__example_55959141808636_1
timestamp 1666199351
transform -1 0 2504 0 1 172
box -1 0 401 1
use sky130_fd_pr__pfet_01v8__example_55959141808636  sky130_fd_pr__pfet_01v8__example_55959141808636_2
timestamp 1666199351
transform 1 0 1648 0 1 172
box -1 0 401 1
<< labels >>
flabel metal1 s 2216 373 2244 401 3 FreeSans 280 0 0 0 EN_FAST_N[0]
port 1 nsew
flabel metal1 s 2413 -472 2441 -444 3 FreeSans 280 0 0 0 EN_FAST_N[1]
port 2 nsew
flabel metal1 s 2735 372 2763 400 3 FreeSans 280 0 0 0 I2C_MODE_H
port 3 nsew
flabel metal1 s 1378 -131 1406 -103 3 FreeSans 280 0 0 0 PDEN_H_N
port 4 nsew
flabel metal1 s 2605 -467 2633 -439 3 FreeSans 280 0 0 0 DRVLO_H_N
port 5 nsew
flabel metal1 s 1811 -1003 1839 -975 3 FreeSans 280 0 0 0 PD_H
port 6 nsew
flabel metal1 s 1834 -252 1862 -224 3 FreeSans 280 0 0 0 VCC_IO
port 7 nsew
flabel metal1 s 2075 -855 2103 -827 3 FreeSans 280 0 0 0 VGND_IO
port 8 nsew
flabel metal1 s 2863 495 2891 523 3 FreeSans 280 0 0 0 VCC_IO
port 7 nsew
flabel comment s 2887 519 2887 519 0 FreeSans 440 0 0 0 INT1
flabel comment s 2211 604 2211 604 0 FreeSans 440 0 0 0 INT2
<< properties >>
string GDS_END 48976646
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48948528
<< end >>
