magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< pwell >>
rect 10 76 514 730
<< nmos >>
rect 204 102 234 704
rect 290 102 320 704
<< ndiff >>
rect 148 692 204 704
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 234 692 290 704
rect 234 658 245 692
rect 279 658 290 692
rect 234 624 290 658
rect 234 590 245 624
rect 279 590 290 624
rect 234 556 290 590
rect 234 522 245 556
rect 279 522 290 556
rect 234 488 290 522
rect 234 454 245 488
rect 279 454 290 488
rect 234 420 290 454
rect 234 386 245 420
rect 279 386 290 420
rect 234 352 290 386
rect 234 318 245 352
rect 279 318 290 352
rect 234 284 290 318
rect 234 250 245 284
rect 279 250 290 284
rect 234 216 290 250
rect 234 182 245 216
rect 279 182 290 216
rect 234 148 290 182
rect 234 114 245 148
rect 279 114 290 148
rect 234 102 290 114
rect 320 692 376 704
rect 320 658 331 692
rect 365 658 376 692
rect 320 624 376 658
rect 320 590 331 624
rect 365 590 376 624
rect 320 556 376 590
rect 320 522 331 556
rect 365 522 376 556
rect 320 488 376 522
rect 320 454 331 488
rect 365 454 376 488
rect 320 420 376 454
rect 320 386 331 420
rect 365 386 376 420
rect 320 352 376 386
rect 320 318 331 352
rect 365 318 376 352
rect 320 284 376 318
rect 320 250 331 284
rect 365 250 376 284
rect 320 216 376 250
rect 320 182 331 216
rect 365 182 376 216
rect 320 148 376 182
rect 320 114 331 148
rect 365 114 376 148
rect 320 102 376 114
<< ndiffc >>
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 245 658 279 692
rect 245 590 279 624
rect 245 522 279 556
rect 245 454 279 488
rect 245 386 279 420
rect 245 318 279 352
rect 245 250 279 284
rect 245 182 279 216
rect 245 114 279 148
rect 331 658 365 692
rect 331 590 365 624
rect 331 522 365 556
rect 331 454 365 488
rect 331 386 365 420
rect 331 318 365 352
rect 331 250 365 284
rect 331 182 365 216
rect 331 114 365 148
<< psubdiff >>
rect 36 658 94 704
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 430 658 488 704
rect 430 624 442 658
rect 476 624 488 658
rect 430 590 488 624
rect 430 556 442 590
rect 476 556 488 590
rect 430 522 488 556
rect 430 488 442 522
rect 476 488 488 522
rect 430 454 488 488
rect 430 420 442 454
rect 476 420 488 454
rect 430 386 488 420
rect 430 352 442 386
rect 476 352 488 386
rect 430 318 488 352
rect 430 284 442 318
rect 476 284 488 318
rect 430 250 488 284
rect 430 216 442 250
rect 476 216 488 250
rect 430 182 488 216
rect 430 148 442 182
rect 476 148 488 182
rect 430 102 488 148
<< psubdiffcont >>
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 442 624 476 658
rect 442 556 476 590
rect 442 488 476 522
rect 442 420 476 454
rect 442 352 476 386
rect 442 284 476 318
rect 442 216 476 250
rect 442 148 476 182
<< poly >>
rect 161 776 363 796
rect 161 742 177 776
rect 211 742 245 776
rect 279 742 313 776
rect 347 742 363 776
rect 161 726 363 742
rect 204 704 234 726
rect 290 704 320 726
rect 204 80 234 102
rect 290 80 320 102
rect 161 64 363 80
rect 161 30 177 64
rect 211 30 245 64
rect 279 30 313 64
rect 347 30 363 64
rect 161 10 363 30
<< polycont >>
rect 177 742 211 776
rect 245 742 279 776
rect 313 742 347 776
rect 177 30 211 64
rect 245 30 279 64
rect 313 30 347 64
<< locali >>
rect 161 742 173 776
rect 211 742 245 776
rect 279 742 313 776
rect 351 742 363 776
rect 159 692 193 708
rect 48 672 82 674
rect 48 600 82 624
rect 48 528 82 556
rect 48 456 82 488
rect 48 386 82 420
rect 48 318 82 350
rect 48 250 82 278
rect 48 182 82 206
rect 48 132 82 134
rect 159 624 193 638
rect 159 556 193 566
rect 159 488 193 494
rect 159 420 193 422
rect 159 384 193 386
rect 159 312 193 318
rect 159 240 193 250
rect 159 168 193 182
rect 159 98 193 114
rect 245 692 279 708
rect 245 624 279 638
rect 245 556 279 566
rect 245 488 279 494
rect 245 420 279 422
rect 245 384 279 386
rect 245 312 279 318
rect 245 240 279 250
rect 245 168 279 182
rect 245 98 279 114
rect 331 692 365 708
rect 331 624 365 638
rect 331 556 365 566
rect 331 488 365 494
rect 331 420 365 422
rect 331 384 365 386
rect 331 312 365 318
rect 331 240 365 250
rect 331 168 365 182
rect 442 672 476 674
rect 442 600 476 624
rect 442 528 476 556
rect 442 456 476 488
rect 442 386 476 420
rect 442 318 476 350
rect 442 250 476 278
rect 442 182 476 206
rect 442 132 476 134
rect 331 98 365 114
rect 161 30 173 64
rect 211 30 245 64
rect 279 30 313 64
rect 351 30 363 64
<< viali >>
rect 173 742 177 776
rect 177 742 207 776
rect 245 742 279 776
rect 317 742 347 776
rect 347 742 351 776
rect 48 658 82 672
rect 48 638 82 658
rect 48 590 82 600
rect 48 566 82 590
rect 48 522 82 528
rect 48 494 82 522
rect 48 454 82 456
rect 48 422 82 454
rect 48 352 82 384
rect 48 350 82 352
rect 48 284 82 312
rect 48 278 82 284
rect 48 216 82 240
rect 48 206 82 216
rect 48 148 82 168
rect 48 134 82 148
rect 159 658 193 672
rect 159 638 193 658
rect 159 590 193 600
rect 159 566 193 590
rect 159 522 193 528
rect 159 494 193 522
rect 159 454 193 456
rect 159 422 193 454
rect 159 352 193 384
rect 159 350 193 352
rect 159 284 193 312
rect 159 278 193 284
rect 159 216 193 240
rect 159 206 193 216
rect 159 148 193 168
rect 159 134 193 148
rect 245 658 279 672
rect 245 638 279 658
rect 245 590 279 600
rect 245 566 279 590
rect 245 522 279 528
rect 245 494 279 522
rect 245 454 279 456
rect 245 422 279 454
rect 245 352 279 384
rect 245 350 279 352
rect 245 284 279 312
rect 245 278 279 284
rect 245 216 279 240
rect 245 206 279 216
rect 245 148 279 168
rect 245 134 279 148
rect 331 658 365 672
rect 331 638 365 658
rect 331 590 365 600
rect 331 566 365 590
rect 331 522 365 528
rect 331 494 365 522
rect 331 454 365 456
rect 331 422 365 454
rect 331 352 365 384
rect 331 350 365 352
rect 331 284 365 312
rect 331 278 365 284
rect 331 216 365 240
rect 331 206 365 216
rect 331 148 365 168
rect 331 134 365 148
rect 442 658 476 672
rect 442 638 476 658
rect 442 590 476 600
rect 442 566 476 590
rect 442 522 476 528
rect 442 494 476 522
rect 442 454 476 456
rect 442 422 476 454
rect 442 352 476 384
rect 442 350 476 352
rect 442 284 476 312
rect 442 278 476 284
rect 442 216 476 240
rect 442 206 476 216
rect 442 148 476 168
rect 442 134 476 148
rect 173 30 177 64
rect 177 30 207 64
rect 245 30 279 64
rect 317 30 347 64
rect 347 30 351 64
<< metal1 >>
rect 161 776 363 796
rect 161 742 173 776
rect 207 742 245 776
rect 279 742 317 776
rect 351 742 363 776
rect 161 730 363 742
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 150 672 202 684
rect 150 638 159 672
rect 193 638 202 672
rect 150 600 202 638
rect 150 566 159 600
rect 193 566 202 600
rect 150 528 202 566
rect 150 494 159 528
rect 193 494 202 528
rect 150 456 202 494
rect 150 422 159 456
rect 193 422 202 456
rect 150 384 202 422
rect 150 372 159 384
rect 193 372 202 384
rect 150 312 202 320
rect 150 308 159 312
rect 193 308 202 312
rect 150 244 202 256
rect 150 180 202 192
rect 150 122 202 128
rect 236 678 288 684
rect 236 614 288 626
rect 236 550 288 562
rect 236 494 245 498
rect 279 494 288 498
rect 236 486 288 494
rect 236 422 245 434
rect 279 422 288 434
rect 236 384 288 422
rect 236 350 245 384
rect 279 350 288 384
rect 236 312 288 350
rect 236 278 245 312
rect 279 278 288 312
rect 236 240 288 278
rect 236 206 245 240
rect 279 206 288 240
rect 236 168 288 206
rect 236 134 245 168
rect 279 134 288 168
rect 236 122 288 134
rect 322 672 374 684
rect 322 638 331 672
rect 365 638 374 672
rect 322 600 374 638
rect 322 566 331 600
rect 365 566 374 600
rect 322 528 374 566
rect 322 494 331 528
rect 365 494 374 528
rect 322 456 374 494
rect 322 422 331 456
rect 365 422 374 456
rect 322 384 374 422
rect 322 372 331 384
rect 365 372 374 384
rect 322 312 374 320
rect 322 308 331 312
rect 365 308 374 312
rect 322 244 374 256
rect 322 180 374 192
rect 322 122 374 128
rect 430 672 488 684
rect 430 638 442 672
rect 476 638 488 672
rect 430 600 488 638
rect 430 566 442 600
rect 476 566 488 600
rect 430 528 488 566
rect 430 494 442 528
rect 476 494 488 528
rect 430 456 488 494
rect 430 422 442 456
rect 476 422 488 456
rect 430 384 488 422
rect 430 350 442 384
rect 476 350 488 384
rect 430 312 488 350
rect 430 278 442 312
rect 476 278 488 312
rect 430 240 488 278
rect 430 206 442 240
rect 476 206 488 240
rect 430 168 488 206
rect 430 134 442 168
rect 476 134 488 168
rect 430 122 488 134
rect 161 64 363 76
rect 161 30 173 64
rect 207 30 245 64
rect 279 30 317 64
rect 351 30 363 64
rect 161 10 363 30
<< via1 >>
rect 150 350 159 372
rect 159 350 193 372
rect 193 350 202 372
rect 150 320 202 350
rect 150 278 159 308
rect 159 278 193 308
rect 193 278 202 308
rect 150 256 202 278
rect 150 240 202 244
rect 150 206 159 240
rect 159 206 193 240
rect 193 206 202 240
rect 150 192 202 206
rect 150 168 202 180
rect 150 134 159 168
rect 159 134 193 168
rect 193 134 202 168
rect 150 128 202 134
rect 236 672 288 678
rect 236 638 245 672
rect 245 638 279 672
rect 279 638 288 672
rect 236 626 288 638
rect 236 600 288 614
rect 236 566 245 600
rect 245 566 279 600
rect 279 566 288 600
rect 236 562 288 566
rect 236 528 288 550
rect 236 498 245 528
rect 245 498 279 528
rect 279 498 288 528
rect 236 456 288 486
rect 236 434 245 456
rect 245 434 279 456
rect 279 434 288 456
rect 322 350 331 372
rect 331 350 365 372
rect 365 350 374 372
rect 322 320 374 350
rect 322 278 331 308
rect 331 278 365 308
rect 365 278 374 308
rect 322 256 374 278
rect 322 240 374 244
rect 322 206 331 240
rect 331 206 365 240
rect 365 206 374 240
rect 322 192 374 206
rect 322 168 374 180
rect 322 134 331 168
rect 331 134 365 168
rect 365 134 374 168
rect 322 128 374 134
<< metal2 >>
rect 10 678 514 684
rect 10 626 236 678
rect 288 626 514 678
rect 10 614 514 626
rect 10 562 236 614
rect 288 562 514 614
rect 10 550 514 562
rect 10 498 236 550
rect 288 498 514 550
rect 10 486 514 498
rect 10 434 236 486
rect 288 434 514 486
rect 10 428 514 434
rect 10 372 514 378
rect 10 320 150 372
rect 202 320 322 372
rect 374 320 514 372
rect 10 308 514 320
rect 10 256 150 308
rect 202 256 322 308
rect 374 256 514 308
rect 10 244 514 256
rect 10 192 150 244
rect 202 192 322 244
rect 374 192 514 244
rect 10 180 514 192
rect 10 128 150 180
rect 202 128 322 180
rect 374 128 514 180
rect 10 122 514 128
<< labels >>
flabel metal2 s 10 428 30 684 7 FreeSans 300 180 0 0 DRAIN
port 1 nsew
flabel metal2 s 10 122 30 378 7 FreeSans 300 180 0 0 SOURCE
port 2 nsew
flabel metal1 s 430 122 488 138 3 FreeSans 300 90 0 0 SUBSTRATE
port 3 nsew
flabel metal1 s 161 10 363 76 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 36 122 94 138 3 FreeSans 300 90 0 0 SUBSTRATE
port 3 nsew
flabel metal1 s 161 730 363 796 0 FreeSans 300 0 0 0 GATE
port 4 nsew
<< properties >>
string GDS_END 1617378
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 1606514
<< end >>
