magic
tech sky130A
timestamp 1666199351
<< properties >>
string GDS_END 3190980
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3190464
<< end >>
