magic
tech sky130B
magscale 1 2
timestamp 1669704864
<< viali >>
rect 4721 47209 4755 47243
rect 5365 47209 5399 47243
rect 6009 47209 6043 47243
rect 7113 47209 7147 47243
rect 7757 47209 7791 47243
rect 8401 47209 8435 47243
rect 9137 47209 9171 47243
rect 10241 47209 10275 47243
rect 11161 47209 11195 47243
rect 12449 47209 12483 47243
rect 13553 47209 13587 47243
rect 15025 47209 15059 47243
rect 16313 47209 16347 47243
rect 20085 47209 20119 47243
rect 22109 47209 22143 47243
rect 29745 47209 29779 47243
rect 39129 47209 39163 47243
rect 42625 47209 42659 47243
rect 43913 47209 43947 47243
rect 44557 47209 44591 47243
rect 45201 47209 45235 47243
rect 45845 47209 45879 47243
rect 46489 47209 46523 47243
rect 15669 47141 15703 47175
rect 16957 47141 16991 47175
rect 17601 47141 17635 47175
rect 18889 47141 18923 47175
rect 19533 47141 19567 47175
rect 22569 47141 22603 47175
rect 36185 47141 36219 47175
rect 41981 47141 42015 47175
rect 18245 47073 18279 47107
rect 24685 47073 24719 47107
rect 26065 47073 26099 47107
rect 28733 47073 28767 47107
rect 32321 47073 32355 47107
rect 33793 47073 33827 47107
rect 35541 47073 35575 47107
rect 37565 47073 37599 47107
rect 19441 47005 19475 47039
rect 19963 47005 19997 47039
rect 21189 47005 21223 47039
rect 21281 47005 21315 47039
rect 22293 47005 22327 47039
rect 22385 47005 22419 47039
rect 22661 47005 22695 47039
rect 23673 47005 23707 47039
rect 23857 47005 23891 47039
rect 24869 47005 24903 47039
rect 25881 47005 25915 47039
rect 26157 47005 26191 47039
rect 27261 47005 27295 47039
rect 27353 47005 27387 47039
rect 27813 47005 27847 47039
rect 28825 47005 28859 47039
rect 29101 47005 29135 47039
rect 30757 47005 30791 47039
rect 31493 47005 31527 47039
rect 32873 47005 32907 47039
rect 33609 47005 33643 47039
rect 33885 47005 33919 47039
rect 34897 47005 34931 47039
rect 36829 47005 36863 47039
rect 37473 47005 37507 47039
rect 37841 47005 37875 47039
rect 38025 47005 38059 47039
rect 38485 47005 38519 47039
rect 40049 47005 40083 47039
rect 40693 47005 40727 47039
rect 41521 47005 41555 47039
rect 43269 47005 43303 47039
rect 21005 46937 21039 46971
rect 23121 46937 23155 46971
rect 24041 46937 24075 46971
rect 25145 46937 25179 46971
rect 30573 46937 30607 46971
rect 31033 46937 31067 46971
rect 32505 46937 32539 46971
rect 33425 46937 33459 46971
rect 19901 46869 19935 46903
rect 25053 46869 25087 46903
rect 25697 46869 25731 46903
rect 30941 46869 30975 46903
rect 32597 46869 32631 46903
rect 32689 46869 32723 46903
rect 41337 46869 41371 46903
rect 17325 46665 17359 46699
rect 21189 46665 21223 46699
rect 24961 46665 24995 46699
rect 25145 46665 25179 46699
rect 25237 46665 25271 46699
rect 25973 46665 26007 46699
rect 26157 46665 26191 46699
rect 29653 46665 29687 46699
rect 34713 46665 34747 46699
rect 35633 46665 35667 46699
rect 23857 46597 23891 46631
rect 24317 46597 24351 46631
rect 25421 46597 25455 46631
rect 28273 46597 28307 46631
rect 28457 46597 28491 46631
rect 33057 46597 33091 46631
rect 6929 46529 6963 46563
rect 14657 46529 14691 46563
rect 17141 46529 17175 46563
rect 17877 46529 17911 46563
rect 17969 46529 18003 46563
rect 18429 46529 18463 46563
rect 19901 46529 19935 46563
rect 20085 46529 20119 46563
rect 20729 46529 20763 46563
rect 21191 46529 21225 46563
rect 22477 46529 22511 46563
rect 22661 46529 22695 46563
rect 23121 46529 23155 46563
rect 23304 46529 23338 46563
rect 23397 46529 23431 46563
rect 23673 46529 23707 46563
rect 25053 46529 25087 46563
rect 26155 46529 26189 46563
rect 26617 46529 26651 46563
rect 27445 46529 27479 46563
rect 27537 46529 27571 46563
rect 27721 46529 27755 46563
rect 27813 46529 27847 46563
rect 28641 46529 28675 46563
rect 29285 46529 29319 46563
rect 29469 46529 29503 46563
rect 29745 46529 29779 46563
rect 30205 46529 30239 46563
rect 30481 46529 30515 46563
rect 30757 46529 30791 46563
rect 31677 46529 31711 46563
rect 32505 46529 32539 46563
rect 32965 46529 32999 46563
rect 33517 46529 33551 46563
rect 33793 46529 33827 46563
rect 34529 46529 34563 46563
rect 34641 46529 34675 46563
rect 34897 46529 34931 46563
rect 35631 46529 35665 46563
rect 37841 46529 37875 46563
rect 38117 46529 38151 46563
rect 39221 46529 39255 46563
rect 40969 46529 41003 46563
rect 41797 46529 41831 46563
rect 43269 46529 43303 46563
rect 43913 46529 43947 46563
rect 44557 46529 44591 46563
rect 16313 46461 16347 46495
rect 19257 46461 19291 46495
rect 19717 46461 19751 46495
rect 23489 46461 23523 46495
rect 31033 46461 31067 46495
rect 33149 46461 33183 46495
rect 34345 46461 34379 46495
rect 36093 46461 36127 46495
rect 38761 46461 38795 46495
rect 38945 46461 38979 46495
rect 40325 46461 40359 46495
rect 18613 46393 18647 46427
rect 20821 46393 20855 46427
rect 22385 46393 22419 46427
rect 30297 46393 30331 46427
rect 37937 46393 37971 46427
rect 38025 46393 38059 46427
rect 39129 46393 39163 46427
rect 42625 46393 42659 46427
rect 21373 46325 21407 46359
rect 26525 46325 26559 46359
rect 27261 46325 27295 46359
rect 31493 46325 31527 46359
rect 32321 46325 32355 46359
rect 35449 46325 35483 46359
rect 36001 46325 36035 46359
rect 36553 46325 36587 46359
rect 37657 46325 37691 46359
rect 39681 46325 39715 46359
rect 41705 46325 41739 46359
rect 17417 46121 17451 46155
rect 23305 46121 23339 46155
rect 25789 46121 25823 46155
rect 27629 46121 27663 46155
rect 30757 46121 30791 46155
rect 35173 46121 35207 46155
rect 37381 46121 37415 46155
rect 38485 46121 38519 46155
rect 41337 46121 41371 46155
rect 41981 46121 42015 46155
rect 42625 46121 42659 46155
rect 43361 46121 43395 46155
rect 20085 46053 20119 46087
rect 25145 46053 25179 46087
rect 27997 46053 28031 46087
rect 31953 46053 31987 46087
rect 37749 46053 37783 46087
rect 40693 46053 40727 46087
rect 23489 45985 23523 46019
rect 23673 45985 23707 46019
rect 23765 45985 23799 46019
rect 26525 45985 26559 46019
rect 28641 45985 28675 46019
rect 29193 45985 29227 46019
rect 31493 45985 31527 46019
rect 32045 45985 32079 46019
rect 35357 45985 35391 46019
rect 35541 45985 35575 46019
rect 36277 45985 36311 46019
rect 40049 45985 40083 46019
rect 17877 45917 17911 45951
rect 18613 45917 18647 45951
rect 18889 45917 18923 45951
rect 19448 45917 19482 45951
rect 19579 45917 19613 45951
rect 19903 45917 19937 45951
rect 20821 45917 20855 45951
rect 21097 45917 21131 45951
rect 21741 45917 21775 45951
rect 21925 45917 21959 45951
rect 22385 45917 22419 45951
rect 23581 45917 23615 45951
rect 23949 45917 23983 45951
rect 24961 45917 24995 45951
rect 25237 45917 25271 45951
rect 26709 45917 26743 45951
rect 26801 45917 26835 45951
rect 27813 45917 27847 45951
rect 28089 45917 28123 45951
rect 28825 45917 28859 45951
rect 30021 45917 30055 45951
rect 30205 45917 30239 45951
rect 30297 45917 30331 45951
rect 31677 45917 31711 45951
rect 32505 45917 32539 45951
rect 33793 45917 33827 45951
rect 33885 45917 33919 45951
rect 35633 45917 35667 45951
rect 36461 45917 36495 45951
rect 36553 45917 36587 45951
rect 36737 45917 36771 45951
rect 36829 45917 36863 45951
rect 37565 45917 37599 45951
rect 37841 45917 37875 45951
rect 38393 45917 38427 45951
rect 38853 45917 38887 45951
rect 39497 45917 39531 45951
rect 18521 45849 18555 45883
rect 20729 45849 20763 45883
rect 22569 45849 22603 45883
rect 22753 45849 22787 45883
rect 26341 45849 26375 45883
rect 16773 45781 16807 45815
rect 18061 45781 18095 45815
rect 19901 45781 19935 45815
rect 21833 45781 21867 45815
rect 24777 45781 24811 45815
rect 29101 45781 29135 45815
rect 29837 45781 29871 45815
rect 33241 45781 33275 45815
rect 18153 45577 18187 45611
rect 24593 45577 24627 45611
rect 25421 45577 25455 45611
rect 33977 45577 34011 45611
rect 35081 45577 35115 45611
rect 42717 45577 42751 45611
rect 17693 45509 17727 45543
rect 18889 45509 18923 45543
rect 21281 45509 21315 45543
rect 23765 45509 23799 45543
rect 24725 45509 24759 45543
rect 30573 45509 30607 45543
rect 32781 45509 32815 45543
rect 35173 45509 35207 45543
rect 18337 45441 18371 45475
rect 18981 45441 19015 45475
rect 19625 45441 19659 45475
rect 20177 45441 20211 45475
rect 20453 45441 20487 45475
rect 21097 45441 21131 45475
rect 21465 45441 21499 45475
rect 22569 45441 22603 45475
rect 22753 45441 22787 45475
rect 23489 45441 23523 45475
rect 23627 45441 23661 45475
rect 24501 45441 24535 45475
rect 24869 45441 24903 45475
rect 25605 45441 25639 45475
rect 26065 45441 26099 45475
rect 27261 45441 27295 45475
rect 27813 45441 27847 45475
rect 27997 45441 28031 45475
rect 28273 45441 28307 45475
rect 29159 45441 29193 45475
rect 29561 45441 29595 45475
rect 30113 45441 30147 45475
rect 30297 45441 30331 45475
rect 30389 45441 30423 45475
rect 31585 45441 31619 45475
rect 32597 45441 32631 45475
rect 32873 45441 32907 45475
rect 33609 45441 33643 45475
rect 34069 45441 34103 45475
rect 34713 45441 34747 45475
rect 34897 45441 34931 45475
rect 36185 45441 36219 45475
rect 36645 45441 36679 45475
rect 37841 45441 37875 45475
rect 38300 45441 38334 45475
rect 39129 45441 39163 45475
rect 39773 45441 39807 45475
rect 40417 45441 40451 45475
rect 20085 45373 20119 45407
rect 22201 45373 22235 45407
rect 22385 45373 22419 45407
rect 23857 45373 23891 45407
rect 29469 45373 29503 45407
rect 31309 45373 31343 45407
rect 33868 45373 33902 45407
rect 34161 45373 34195 45407
rect 35725 45373 35759 45407
rect 37933 45373 37967 45407
rect 24317 45305 24351 45339
rect 30205 45305 30239 45339
rect 36737 45305 36771 45339
rect 38945 45305 38979 45339
rect 40233 45305 40267 45339
rect 40877 45305 40911 45339
rect 19533 45237 19567 45271
rect 26249 45237 26283 45271
rect 26525 45237 26559 45271
rect 27905 45237 27939 45271
rect 29009 45237 29043 45271
rect 31217 45237 31251 45271
rect 32413 45237 32447 45271
rect 33425 45237 33459 45271
rect 35909 45237 35943 45271
rect 38393 45237 38427 45271
rect 39589 45237 39623 45271
rect 41521 45237 41555 45271
rect 19809 45033 19843 45067
rect 23489 45033 23523 45067
rect 31861 45033 31895 45067
rect 38209 45033 38243 45067
rect 39221 45033 39255 45067
rect 40049 45033 40083 45067
rect 40601 45033 40635 45067
rect 41705 45033 41739 45067
rect 42349 45033 42383 45067
rect 20453 44965 20487 44999
rect 33517 44965 33551 44999
rect 25973 44897 26007 44931
rect 26985 44897 27019 44931
rect 27905 44897 27939 44931
rect 29745 44897 29779 44931
rect 30573 44897 30607 44931
rect 38761 44897 38795 44931
rect 18705 44829 18739 44863
rect 19993 44829 20027 44863
rect 20637 44829 20671 44863
rect 21189 44829 21223 44863
rect 21465 44829 21499 44863
rect 22385 44829 22419 44863
rect 22845 44829 22879 44863
rect 23673 44829 23707 44863
rect 23765 44829 23799 44863
rect 23949 44829 23983 44863
rect 24041 44829 24075 44863
rect 24593 44829 24627 44863
rect 25743 44829 25777 44863
rect 26065 44829 26099 44863
rect 26525 44829 26559 44863
rect 26801 44829 26835 44863
rect 27537 44829 27571 44863
rect 27813 44829 27847 44863
rect 28181 44829 28215 44863
rect 28641 44829 28675 44863
rect 28917 44829 28951 44863
rect 30389 44829 30423 44863
rect 32045 44829 32079 44863
rect 32137 44829 32171 44863
rect 32321 44829 32355 44863
rect 32413 44829 32447 44863
rect 33425 44829 33459 44863
rect 33793 44829 33827 44863
rect 33977 44829 34011 44863
rect 35725 44829 35759 44863
rect 35909 44829 35943 44863
rect 37013 44829 37047 44863
rect 37197 44829 37231 44863
rect 37473 44829 37507 44863
rect 38302 44829 38336 44863
rect 38669 44829 38703 44863
rect 41153 44829 41187 44863
rect 21097 44761 21131 44795
rect 22661 44761 22695 44795
rect 24685 44761 24719 44795
rect 25329 44761 25363 44795
rect 25513 44761 25547 44795
rect 26617 44761 26651 44795
rect 28733 44761 28767 44795
rect 29101 44761 29135 44795
rect 32873 44761 32907 44795
rect 37657 44761 37691 44795
rect 18797 44693 18831 44727
rect 25881 44693 25915 44727
rect 34897 44693 34931 44727
rect 19901 44489 19935 44523
rect 20729 44489 20763 44523
rect 21373 44489 21407 44523
rect 25513 44489 25547 44523
rect 27261 44489 27295 44523
rect 30297 44489 30331 44523
rect 36553 44489 36587 44523
rect 38669 44489 38703 44523
rect 40141 44489 40175 44523
rect 41337 44489 41371 44523
rect 22937 44421 22971 44455
rect 24869 44421 24903 44455
rect 27169 44421 27203 44455
rect 33701 44421 33735 44455
rect 34345 44421 34379 44455
rect 40693 44421 40727 44455
rect 18981 44353 19015 44387
rect 19809 44353 19843 44387
rect 20821 44353 20855 44387
rect 21281 44353 21315 44387
rect 22477 44353 22511 44387
rect 23121 44353 23155 44387
rect 23305 44353 23339 44387
rect 24133 44353 24167 44387
rect 25513 44353 25547 44387
rect 26341 44353 26375 44387
rect 27445 44353 27479 44387
rect 29469 44353 29503 44387
rect 29653 44353 29687 44387
rect 31125 44353 31159 44387
rect 34161 44353 34195 44387
rect 34529 44353 34563 44387
rect 35725 44353 35759 44387
rect 37473 44353 37507 44387
rect 37657 44353 37691 44387
rect 38117 44353 38151 44387
rect 38853 44353 38887 44387
rect 39037 44353 39071 44387
rect 39129 44353 39163 44387
rect 39589 44353 39623 44387
rect 23765 44285 23799 44319
rect 24317 44285 24351 44319
rect 25329 44285 25363 44319
rect 25881 44285 25915 44319
rect 27629 44285 27663 44319
rect 28641 44285 28675 44319
rect 30941 44285 30975 44319
rect 32873 44285 32907 44319
rect 35817 44285 35851 44319
rect 19165 44217 19199 44251
rect 23857 44217 23891 44251
rect 22385 44149 22419 44183
rect 37565 44149 37599 44183
rect 21189 43945 21223 43979
rect 26157 43945 26191 43979
rect 29009 43945 29043 43979
rect 29745 43945 29779 43979
rect 30941 43945 30975 43979
rect 31769 43945 31803 43979
rect 34253 43945 34287 43979
rect 35541 43945 35575 43979
rect 36553 43945 36587 43979
rect 36829 43945 36863 43979
rect 39037 43945 39071 43979
rect 40141 43945 40175 43979
rect 20637 43877 20671 43911
rect 21833 43877 21867 43911
rect 33149 43877 33183 43911
rect 38577 43877 38611 43911
rect 22661 43809 22695 43843
rect 24869 43809 24903 43843
rect 26801 43809 26835 43843
rect 34989 43809 35023 43843
rect 21649 43741 21683 43775
rect 22937 43741 22971 43775
rect 23397 43741 23431 43775
rect 27169 43741 27203 43775
rect 27629 43741 27663 43775
rect 28365 43741 28399 43775
rect 29193 43741 29227 43775
rect 31033 43741 31067 43775
rect 31677 43741 31711 43775
rect 31861 43741 31895 43775
rect 32505 43741 32539 43775
rect 32689 43741 32723 43775
rect 33517 43741 33551 43775
rect 33977 43741 34011 43775
rect 34161 43741 34195 43775
rect 35725 43741 35759 43775
rect 35909 43741 35943 43775
rect 37013 43741 37047 43775
rect 37565 43741 37599 43775
rect 37749 43741 37783 43775
rect 38025 43741 38059 43775
rect 25697 43673 25731 43707
rect 28457 43673 28491 43707
rect 32321 43673 32355 43707
rect 33333 43673 33367 43707
rect 36001 43673 36035 43707
rect 37933 43673 37967 43707
rect 22477 43401 22511 43435
rect 23581 43401 23615 43435
rect 27629 43401 27663 43435
rect 33241 43401 33275 43435
rect 35173 43401 35207 43435
rect 35725 43401 35759 43435
rect 36829 43401 36863 43435
rect 37565 43401 37599 43435
rect 38117 43401 38151 43435
rect 39129 43401 39163 43435
rect 24961 43333 24995 43367
rect 25145 43333 25179 43367
rect 25789 43333 25823 43367
rect 26157 43333 26191 43367
rect 29285 43333 29319 43367
rect 32321 43333 32355 43367
rect 32689 43333 32723 43367
rect 36185 43333 36219 43367
rect 38669 43333 38703 43367
rect 23673 43265 23707 43299
rect 24133 43265 24167 43299
rect 24317 43265 24351 43299
rect 24501 43265 24535 43299
rect 25329 43265 25363 43299
rect 25973 43265 26007 43299
rect 27169 43265 27203 43299
rect 31217 43265 31251 43299
rect 31769 43265 31803 43299
rect 32505 43265 32539 43299
rect 33149 43265 33183 43299
rect 33793 43265 33827 43299
rect 34437 43265 34471 43299
rect 36921 43265 36955 43299
rect 23029 43197 23063 43231
rect 28641 43197 28675 43231
rect 29193 43197 29227 43231
rect 29745 43129 29779 43163
rect 27445 43061 27479 43095
rect 30389 43061 30423 43095
rect 24685 42857 24719 42891
rect 25789 42857 25823 42891
rect 26249 42857 26283 42891
rect 29745 42857 29779 42891
rect 32873 42857 32907 42891
rect 33425 42857 33459 42891
rect 33977 42857 34011 42891
rect 35449 42857 35483 42891
rect 25145 42789 25179 42823
rect 34989 42789 35023 42823
rect 36001 42789 36035 42823
rect 24041 42721 24075 42755
rect 27261 42721 27295 42755
rect 27721 42721 27755 42755
rect 28457 42721 28491 42755
rect 30389 42721 30423 42755
rect 36645 42721 36679 42755
rect 31953 42653 31987 42687
rect 30941 42585 30975 42619
rect 22937 42517 22971 42551
rect 29009 42517 29043 42551
rect 31493 42517 31527 42551
rect 25237 42313 25271 42347
rect 26341 42313 26375 42347
rect 27261 42313 27295 42347
rect 27721 42313 27755 42347
rect 29929 42313 29963 42347
rect 32321 42313 32355 42347
rect 34253 42313 34287 42347
rect 36001 42313 36035 42347
rect 25789 42245 25823 42279
rect 28273 42245 28307 42279
rect 30757 42245 30791 42279
rect 35541 42245 35575 42279
rect 29285 41973 29319 42007
rect 25329 41769 25363 41803
rect 29745 41769 29779 41803
rect 22937 6749 22971 6783
rect 24593 6749 24627 6783
rect 21925 6613 21959 6647
rect 22385 6613 22419 6647
rect 24685 6613 24719 6647
rect 24777 6341 24811 6375
rect 26065 6341 26099 6375
rect 22201 6273 22235 6307
rect 22661 6273 22695 6307
rect 28181 6273 28215 6307
rect 24133 6205 24167 6239
rect 24685 6205 24719 6239
rect 25973 6205 26007 6239
rect 25237 6137 25271 6171
rect 26525 6137 26559 6171
rect 20821 6069 20855 6103
rect 21281 6069 21315 6103
rect 22017 6069 22051 6103
rect 22753 6069 22787 6103
rect 23489 6069 23523 6103
rect 27353 6069 27387 6103
rect 28089 6069 28123 6103
rect 25973 5865 26007 5899
rect 26709 5865 26743 5899
rect 21925 5797 21959 5831
rect 23857 5797 23891 5831
rect 27997 5797 28031 5831
rect 21373 5729 21407 5763
rect 22753 5729 22787 5763
rect 23305 5729 23339 5763
rect 24685 5729 24719 5763
rect 24961 5729 24995 5763
rect 27445 5729 27479 5763
rect 20637 5661 20671 5695
rect 26617 5661 26651 5695
rect 20729 5593 20763 5627
rect 21465 5593 21499 5627
rect 23397 5593 23431 5627
rect 24777 5593 24811 5627
rect 27537 5593 27571 5627
rect 20177 5525 20211 5559
rect 21373 5321 21407 5355
rect 24501 5321 24535 5355
rect 23029 5253 23063 5287
rect 23121 5253 23155 5287
rect 25881 5253 25915 5287
rect 27813 5253 27847 5287
rect 19993 5185 20027 5219
rect 20821 5185 20855 5219
rect 21281 5185 21315 5219
rect 22477 5185 22511 5219
rect 24409 5185 24443 5219
rect 25237 5117 25271 5151
rect 25789 5117 25823 5151
rect 27629 5117 27663 5151
rect 27905 5117 27939 5151
rect 28457 5117 28491 5151
rect 20637 5049 20671 5083
rect 22293 5049 22327 5083
rect 23581 5049 23615 5083
rect 26341 5049 26375 5083
rect 19441 4981 19475 5015
rect 20085 4981 20119 5015
rect 29101 4981 29135 5015
rect 22109 4777 22143 4811
rect 25789 4777 25823 4811
rect 27537 4777 27571 4811
rect 25053 4709 25087 4743
rect 18889 4641 18923 4675
rect 20913 4641 20947 4675
rect 22845 4641 22879 4675
rect 23305 4641 23339 4675
rect 28825 4641 28859 4675
rect 29101 4641 29135 4675
rect 18061 4573 18095 4607
rect 19717 4573 19751 4607
rect 20177 4573 20211 4607
rect 22293 4573 22327 4607
rect 25237 4573 25271 4607
rect 25697 4573 25731 4607
rect 26985 4573 27019 4607
rect 27629 4573 27663 4607
rect 29745 4573 29779 4607
rect 30573 4573 30607 4607
rect 21005 4505 21039 4539
rect 21557 4505 21591 4539
rect 22937 4505 22971 4539
rect 29009 4505 29043 4539
rect 30481 4505 30515 4539
rect 19625 4437 19659 4471
rect 20269 4437 20303 4471
rect 26801 4437 26835 4471
rect 29929 4437 29963 4471
rect 20545 4165 20579 4199
rect 22201 4165 22235 4199
rect 24317 4165 24351 4199
rect 25513 4165 25547 4199
rect 27353 4165 27387 4199
rect 29101 4165 29135 4199
rect 29837 4165 29871 4199
rect 29929 4097 29963 4131
rect 18613 4029 18647 4063
rect 20453 4029 20487 4063
rect 21097 4029 21131 4063
rect 22109 4029 22143 4063
rect 22385 4029 22419 4063
rect 24225 4029 24259 4063
rect 25421 4029 25455 4063
rect 26065 4029 26099 4063
rect 27261 4029 27295 4063
rect 27537 4029 27571 4063
rect 28917 4029 28951 4063
rect 29193 4029 29227 4063
rect 30389 4029 30423 4063
rect 19257 3961 19291 3995
rect 23673 3961 23707 3995
rect 24777 3961 24811 3995
rect 15025 3893 15059 3927
rect 16129 3893 16163 3927
rect 17233 3893 17267 3927
rect 17969 3893 18003 3927
rect 19901 3893 19935 3927
rect 23397 3689 23431 3723
rect 23949 3689 23983 3723
rect 25881 3689 25915 3723
rect 16313 3621 16347 3655
rect 33609 3621 33643 3655
rect 37473 3621 37507 3655
rect 15025 3553 15059 3587
rect 17601 3553 17635 3587
rect 20361 3553 20395 3587
rect 24961 3553 24995 3587
rect 27077 3553 27111 3587
rect 28273 3553 28307 3587
rect 31033 3553 31067 3587
rect 35541 3553 35575 3587
rect 4261 3485 4295 3519
rect 5181 3485 5215 3519
rect 6009 3485 6043 3519
rect 6837 3485 6871 3519
rect 7665 3485 7699 3519
rect 8493 3485 8527 3519
rect 9321 3485 9355 3519
rect 10149 3485 10183 3519
rect 10977 3485 11011 3519
rect 11713 3485 11747 3519
rect 12357 3485 12391 3519
rect 13001 3485 13035 3519
rect 13645 3485 13679 3519
rect 15669 3485 15703 3519
rect 16957 3485 16991 3519
rect 18245 3485 18279 3519
rect 18705 3485 18739 3519
rect 19625 3485 19659 3519
rect 20453 3485 20487 3519
rect 20913 3485 20947 3519
rect 23857 3485 23891 3519
rect 25973 3485 26007 3519
rect 29929 3485 29963 3519
rect 30389 3485 30423 3519
rect 31677 3485 31711 3519
rect 32321 3485 32355 3519
rect 32965 3485 32999 3519
rect 34897 3485 34931 3519
rect 36185 3485 36219 3519
rect 36829 3485 36863 3519
rect 38117 3485 38151 3519
rect 38761 3485 38795 3519
rect 40049 3485 40083 3519
rect 40693 3485 40727 3519
rect 41337 3485 41371 3519
rect 41981 3485 42015 3519
rect 42901 3485 42935 3519
rect 43361 3485 43395 3519
rect 45201 3485 45235 3519
rect 45845 3485 45879 3519
rect 46489 3485 46523 3519
rect 47133 3485 47167 3519
rect 47777 3485 47811 3519
rect 21649 3417 21683 3451
rect 21741 3417 21775 3451
rect 22293 3417 22327 3451
rect 24685 3417 24719 3451
rect 24777 3417 24811 3451
rect 27261 3417 27295 3451
rect 27353 3417 27387 3451
rect 28457 3417 28491 3451
rect 28549 3417 28583 3451
rect 18797 3349 18831 3383
rect 19717 3349 19751 3383
rect 21005 3349 21039 3383
rect 29837 3349 29871 3383
rect 18153 3145 18187 3179
rect 19441 3145 19475 3179
rect 20821 3077 20855 3111
rect 22753 3077 22787 3111
rect 24133 3077 24167 3111
rect 25329 3077 25363 3111
rect 27721 3077 27755 3111
rect 28917 3077 28951 3111
rect 29009 3077 29043 3111
rect 30113 3077 30147 3111
rect 31493 3077 31527 3111
rect 18245 3009 18279 3043
rect 19533 3009 19567 3043
rect 20177 3009 20211 3043
rect 26617 3009 26651 3043
rect 30757 3009 30791 3043
rect 31401 3009 31435 3043
rect 34253 3009 34287 3043
rect 4721 2941 4755 2975
rect 7297 2941 7331 2975
rect 9229 2941 9263 2975
rect 14381 2941 14415 2975
rect 15669 2941 15703 2975
rect 20729 2941 20763 2975
rect 21373 2941 21407 2975
rect 22661 2941 22695 2975
rect 22937 2941 22971 2975
rect 24041 2941 24075 2975
rect 24409 2941 24443 2975
rect 25237 2941 25271 2975
rect 25513 2941 25547 2975
rect 27169 2941 27203 2975
rect 27813 2941 27847 2975
rect 28549 2941 28583 2975
rect 29561 2941 29595 2975
rect 30205 2941 30239 2975
rect 33609 2941 33643 2975
rect 35541 2941 35575 2975
rect 38117 2941 38151 2975
rect 39405 2941 39439 2975
rect 41337 2941 41371 2975
rect 43269 2941 43303 2975
rect 45201 2941 45235 2975
rect 4077 2873 4111 2907
rect 5365 2873 5399 2907
rect 10517 2873 10551 2907
rect 12449 2873 12483 2907
rect 13737 2873 13771 2907
rect 15025 2873 15059 2907
rect 18889 2873 18923 2907
rect 32965 2873 32999 2907
rect 34897 2873 34931 2907
rect 36185 2873 36219 2907
rect 2789 2805 2823 2839
rect 3433 2805 3467 2839
rect 6009 2805 6043 2839
rect 7941 2805 7975 2839
rect 8585 2805 8619 2839
rect 9873 2805 9907 2839
rect 11161 2805 11195 2839
rect 13093 2805 13127 2839
rect 16313 2805 16347 2839
rect 17601 2805 17635 2839
rect 32321 2805 32355 2839
rect 37473 2805 37507 2839
rect 38761 2805 38795 2839
rect 40049 2805 40083 2839
rect 40693 2805 40727 2839
rect 42625 2805 42659 2839
rect 43913 2805 43947 2839
rect 44557 2805 44591 2839
rect 45845 2805 45879 2839
rect 46489 2805 46523 2839
rect 47777 2805 47811 2839
rect 15669 2601 15703 2635
rect 20821 2601 20855 2635
rect 22201 2601 22235 2635
rect 27261 2601 27295 2635
rect 27813 2601 27847 2635
rect 28549 2601 28583 2635
rect 30481 2601 30515 2635
rect 31033 2601 31067 2635
rect 5365 2533 5399 2567
rect 7941 2533 7975 2567
rect 9873 2533 9907 2567
rect 12449 2533 12483 2567
rect 18245 2533 18279 2567
rect 20085 2533 20119 2567
rect 21465 2533 21499 2567
rect 26525 2533 26559 2567
rect 29745 2533 29779 2567
rect 32321 2533 32355 2567
rect 34897 2533 34931 2567
rect 37473 2533 37507 2567
rect 40049 2533 40083 2567
rect 43913 2533 43947 2567
rect 46489 2533 46523 2567
rect 2789 2465 2823 2499
rect 7297 2465 7331 2499
rect 8585 2465 8619 2499
rect 11161 2465 11195 2499
rect 13093 2465 13127 2499
rect 15025 2465 15059 2499
rect 18889 2465 18923 2499
rect 22753 2465 22787 2499
rect 23029 2465 23063 2499
rect 23949 2465 23983 2499
rect 25329 2465 25363 2499
rect 25789 2465 25823 2499
rect 33609 2465 33643 2499
rect 36185 2465 36219 2499
rect 38761 2465 38795 2499
rect 40693 2465 40727 2499
rect 42625 2465 42659 2499
rect 45201 2465 45235 2499
rect 2145 2397 2179 2431
rect 3433 2397 3467 2431
rect 4721 2397 4755 2431
rect 6009 2397 6043 2431
rect 10517 2397 10551 2431
rect 13737 2397 13771 2431
rect 16313 2397 16347 2431
rect 17601 2397 17635 2431
rect 19993 2397 20027 2431
rect 24041 2397 24075 2431
rect 24593 2397 24627 2431
rect 26617 2397 26651 2431
rect 27169 2397 27203 2431
rect 28457 2397 28491 2431
rect 30573 2397 30607 2431
rect 32965 2397 32999 2431
rect 35541 2397 35575 2431
rect 38117 2397 38151 2431
rect 41337 2397 41371 2431
rect 43269 2397 43303 2431
rect 45845 2397 45879 2431
rect 47777 2397 47811 2431
rect 22845 2329 22879 2363
rect 25421 2329 25455 2363
rect 24685 2261 24719 2295
<< metal1 >>
rect 19426 47744 19432 47796
rect 19484 47784 19490 47796
rect 23934 47784 23940 47796
rect 19484 47756 23940 47784
rect 19484 47744 19490 47756
rect 23934 47744 23940 47756
rect 23992 47744 23998 47796
rect 16942 47676 16948 47728
rect 17000 47716 17006 47728
rect 23750 47716 23756 47728
rect 17000 47688 23756 47716
rect 17000 47676 17006 47688
rect 23750 47676 23756 47688
rect 23808 47676 23814 47728
rect 18874 47608 18880 47660
rect 18932 47648 18938 47660
rect 24578 47648 24584 47660
rect 18932 47620 24584 47648
rect 18932 47608 18938 47620
rect 24578 47608 24584 47620
rect 24636 47608 24642 47660
rect 5074 47540 5080 47592
rect 5132 47580 5138 47592
rect 22094 47580 22100 47592
rect 5132 47552 22100 47580
rect 5132 47540 5138 47552
rect 22094 47540 22100 47552
rect 22152 47540 22158 47592
rect 28994 47540 29000 47592
rect 29052 47580 29058 47592
rect 34698 47580 34704 47592
rect 29052 47552 34704 47580
rect 29052 47540 29058 47552
rect 34698 47540 34704 47552
rect 34756 47540 34762 47592
rect 36446 47540 36452 47592
rect 36504 47580 36510 47592
rect 41230 47580 41236 47592
rect 36504 47552 41236 47580
rect 36504 47540 36510 47552
rect 41230 47540 41236 47552
rect 41288 47540 41294 47592
rect 17586 47472 17592 47524
rect 17644 47512 17650 47524
rect 21266 47512 21272 47524
rect 17644 47484 21272 47512
rect 17644 47472 17650 47484
rect 21266 47472 21272 47484
rect 21324 47472 21330 47524
rect 23750 47472 23756 47524
rect 23808 47512 23814 47524
rect 24762 47512 24768 47524
rect 23808 47484 24768 47512
rect 23808 47472 23814 47484
rect 24762 47472 24768 47484
rect 24820 47512 24826 47524
rect 27522 47512 27528 47524
rect 24820 47484 27528 47512
rect 24820 47472 24826 47484
rect 27522 47472 27528 47484
rect 27580 47472 27586 47524
rect 33594 47472 33600 47524
rect 33652 47512 33658 47524
rect 36354 47512 36360 47524
rect 33652 47484 36360 47512
rect 33652 47472 33658 47484
rect 36354 47472 36360 47484
rect 36412 47512 36418 47524
rect 36412 47484 38654 47512
rect 36412 47472 36418 47484
rect 11698 47404 11704 47456
rect 11756 47444 11762 47456
rect 20070 47444 20076 47456
rect 11756 47416 20076 47444
rect 11756 47404 11762 47416
rect 20070 47404 20076 47416
rect 20128 47404 20134 47456
rect 22186 47404 22192 47456
rect 22244 47444 22250 47456
rect 29638 47444 29644 47456
rect 22244 47416 29644 47444
rect 22244 47404 22250 47416
rect 29638 47404 29644 47416
rect 29696 47404 29702 47456
rect 31570 47404 31576 47456
rect 31628 47444 31634 47456
rect 36538 47444 36544 47456
rect 31628 47416 36544 47444
rect 31628 47404 31634 47416
rect 36538 47404 36544 47416
rect 36596 47404 36602 47456
rect 38626 47444 38654 47484
rect 41966 47444 41972 47456
rect 38626 47416 41972 47444
rect 41966 47404 41972 47416
rect 42024 47404 42030 47456
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 4706 47240 4712 47252
rect 4667 47212 4712 47240
rect 4706 47200 4712 47212
rect 4764 47200 4770 47252
rect 5353 47243 5411 47249
rect 5353 47209 5365 47243
rect 5399 47240 5411 47243
rect 5810 47240 5816 47252
rect 5399 47212 5816 47240
rect 5399 47209 5411 47212
rect 5353 47203 5411 47209
rect 5810 47200 5816 47212
rect 5868 47200 5874 47252
rect 5994 47240 6000 47252
rect 5955 47212 6000 47240
rect 5994 47200 6000 47212
rect 6052 47200 6058 47252
rect 7098 47240 7104 47252
rect 7059 47212 7104 47240
rect 7098 47200 7104 47212
rect 7156 47200 7162 47252
rect 7742 47240 7748 47252
rect 7703 47212 7748 47240
rect 7742 47200 7748 47212
rect 7800 47200 7806 47252
rect 8386 47240 8392 47252
rect 8347 47212 8392 47240
rect 8386 47200 8392 47212
rect 8444 47200 8450 47252
rect 9122 47240 9128 47252
rect 9083 47212 9128 47240
rect 9122 47200 9128 47212
rect 9180 47200 9186 47252
rect 10226 47240 10232 47252
rect 10187 47212 10232 47240
rect 10226 47200 10232 47212
rect 10284 47200 10290 47252
rect 11146 47240 11152 47252
rect 11107 47212 11152 47240
rect 11146 47200 11152 47212
rect 11204 47200 11210 47252
rect 12434 47200 12440 47252
rect 12492 47240 12498 47252
rect 13538 47240 13544 47252
rect 12492 47212 12537 47240
rect 13499 47212 13544 47240
rect 12492 47200 12498 47212
rect 13538 47200 13544 47212
rect 13596 47200 13602 47252
rect 15013 47243 15071 47249
rect 15013 47209 15025 47243
rect 15059 47240 15071 47243
rect 15746 47240 15752 47252
rect 15059 47212 15752 47240
rect 15059 47209 15071 47212
rect 15013 47203 15071 47209
rect 15746 47200 15752 47212
rect 15804 47200 15810 47252
rect 16301 47243 16359 47249
rect 16301 47209 16313 47243
rect 16347 47240 16359 47243
rect 19058 47240 19064 47252
rect 16347 47212 19064 47240
rect 16347 47209 16359 47212
rect 16301 47203 16359 47209
rect 19058 47200 19064 47212
rect 19116 47200 19122 47252
rect 20070 47240 20076 47252
rect 20031 47212 20076 47240
rect 20070 47200 20076 47212
rect 20128 47200 20134 47252
rect 22094 47200 22100 47252
rect 22152 47240 22158 47252
rect 22152 47212 22197 47240
rect 22152 47200 22158 47212
rect 26786 47200 26792 47252
rect 26844 47240 26850 47252
rect 29733 47243 29791 47249
rect 29733 47240 29745 47243
rect 26844 47212 29745 47240
rect 26844 47200 26850 47212
rect 29733 47209 29745 47212
rect 29779 47209 29791 47243
rect 29733 47203 29791 47209
rect 32674 47200 32680 47252
rect 32732 47240 32738 47252
rect 39117 47243 39175 47249
rect 39117 47240 39129 47243
rect 32732 47212 39129 47240
rect 32732 47200 32738 47212
rect 39117 47209 39129 47212
rect 39163 47209 39175 47243
rect 39117 47203 39175 47209
rect 39298 47200 39304 47252
rect 39356 47240 39362 47252
rect 42613 47243 42671 47249
rect 42613 47240 42625 47243
rect 39356 47212 42625 47240
rect 39356 47200 39362 47212
rect 42613 47209 42625 47212
rect 42659 47209 42671 47243
rect 42613 47203 42671 47209
rect 43346 47200 43352 47252
rect 43404 47240 43410 47252
rect 43901 47243 43959 47249
rect 43901 47240 43913 47243
rect 43404 47212 43913 47240
rect 43404 47200 43410 47212
rect 43901 47209 43913 47212
rect 43947 47209 43959 47243
rect 43901 47203 43959 47209
rect 44082 47200 44088 47252
rect 44140 47240 44146 47252
rect 44545 47243 44603 47249
rect 44545 47240 44557 47243
rect 44140 47212 44557 47240
rect 44140 47200 44146 47212
rect 44545 47209 44557 47212
rect 44591 47209 44603 47243
rect 44545 47203 44603 47209
rect 44818 47200 44824 47252
rect 44876 47240 44882 47252
rect 45189 47243 45247 47249
rect 45189 47240 45201 47243
rect 44876 47212 45201 47240
rect 44876 47200 44882 47212
rect 45189 47209 45201 47212
rect 45235 47209 45247 47243
rect 45830 47240 45836 47252
rect 45791 47212 45836 47240
rect 45189 47203 45247 47209
rect 45830 47200 45836 47212
rect 45888 47200 45894 47252
rect 45922 47200 45928 47252
rect 45980 47240 45986 47252
rect 46477 47243 46535 47249
rect 46477 47240 46489 47243
rect 45980 47212 46489 47240
rect 45980 47200 45986 47212
rect 46477 47209 46489 47212
rect 46523 47209 46535 47243
rect 46477 47203 46535 47209
rect 15657 47175 15715 47181
rect 15657 47141 15669 47175
rect 15703 47172 15715 47175
rect 16850 47172 16856 47184
rect 15703 47144 16856 47172
rect 15703 47141 15715 47144
rect 15657 47135 15715 47141
rect 16850 47132 16856 47144
rect 16908 47132 16914 47184
rect 16942 47132 16948 47184
rect 17000 47172 17006 47184
rect 17586 47172 17592 47184
rect 17000 47144 17045 47172
rect 17547 47144 17592 47172
rect 17000 47132 17006 47144
rect 17586 47132 17592 47144
rect 17644 47132 17650 47184
rect 18874 47172 18880 47184
rect 18835 47144 18880 47172
rect 18874 47132 18880 47144
rect 18932 47132 18938 47184
rect 19334 47132 19340 47184
rect 19392 47172 19398 47184
rect 19521 47175 19579 47181
rect 19521 47172 19533 47175
rect 19392 47144 19533 47172
rect 19392 47132 19398 47144
rect 19521 47141 19533 47144
rect 19567 47172 19579 47175
rect 19978 47172 19984 47184
rect 19567 47144 19984 47172
rect 19567 47141 19579 47144
rect 19521 47135 19579 47141
rect 19978 47132 19984 47144
rect 20036 47132 20042 47184
rect 22370 47172 22376 47184
rect 20180 47144 22376 47172
rect 18233 47107 18291 47113
rect 18233 47073 18245 47107
rect 18279 47104 18291 47107
rect 20180 47104 20208 47144
rect 22370 47132 22376 47144
rect 22428 47132 22434 47184
rect 22557 47175 22615 47181
rect 22557 47141 22569 47175
rect 22603 47172 22615 47175
rect 28258 47172 28264 47184
rect 22603 47144 28264 47172
rect 22603 47141 22615 47144
rect 22557 47135 22615 47141
rect 28258 47132 28264 47144
rect 28316 47132 28322 47184
rect 30466 47132 30472 47184
rect 30524 47172 30530 47184
rect 36173 47175 36231 47181
rect 36173 47172 36185 47175
rect 30524 47144 36185 47172
rect 30524 47132 30530 47144
rect 36173 47141 36185 47144
rect 36219 47141 36231 47175
rect 36173 47135 36231 47141
rect 36814 47132 36820 47184
rect 36872 47172 36878 47184
rect 41874 47172 41880 47184
rect 36872 47144 41880 47172
rect 36872 47132 36878 47144
rect 41874 47132 41880 47144
rect 41932 47132 41938 47184
rect 41966 47132 41972 47184
rect 42024 47172 42030 47184
rect 42024 47144 42069 47172
rect 42024 47132 42030 47144
rect 18279 47076 20208 47104
rect 21008 47076 21312 47104
rect 18279 47073 18291 47076
rect 18233 47067 18291 47073
rect 19058 47036 19064 47048
rect 17880 47008 19064 47036
rect 16114 46860 16120 46912
rect 16172 46900 16178 46912
rect 17880 46900 17908 47008
rect 19058 46996 19064 47008
rect 19116 47036 19122 47048
rect 19429 47039 19487 47045
rect 19429 47036 19441 47039
rect 19116 47008 19441 47036
rect 19116 46996 19122 47008
rect 19429 47005 19441 47008
rect 19475 47005 19487 47039
rect 19429 46999 19487 47005
rect 19951 47039 20009 47045
rect 19951 47005 19963 47039
rect 19997 47036 20009 47039
rect 21008 47036 21036 47076
rect 21284 47048 21312 47076
rect 21358 47064 21364 47116
rect 21416 47104 21422 47116
rect 21416 47076 22692 47104
rect 21416 47064 21422 47076
rect 19997 47008 21036 47036
rect 21177 47039 21235 47045
rect 19997 47005 20009 47008
rect 19951 46999 20009 47005
rect 21177 47005 21189 47039
rect 21223 47005 21235 47039
rect 21177 46999 21235 47005
rect 17954 46928 17960 46980
rect 18012 46968 18018 46980
rect 20993 46971 21051 46977
rect 20993 46968 21005 46971
rect 18012 46940 21005 46968
rect 18012 46928 18018 46940
rect 20993 46937 21005 46940
rect 21039 46937 21051 46971
rect 21192 46968 21220 46999
rect 21266 46996 21272 47048
rect 21324 47036 21330 47048
rect 21324 47008 21417 47036
rect 21324 46996 21330 47008
rect 22186 46996 22192 47048
rect 22244 47036 22250 47048
rect 22281 47039 22339 47045
rect 22281 47036 22293 47039
rect 22244 47008 22293 47036
rect 22244 46996 22250 47008
rect 22281 47005 22293 47008
rect 22327 47005 22339 47039
rect 22281 46999 22339 47005
rect 22370 46996 22376 47048
rect 22428 47036 22434 47048
rect 22664 47045 22692 47076
rect 23382 47064 23388 47116
rect 23440 47104 23446 47116
rect 24673 47107 24731 47113
rect 24673 47104 24685 47107
rect 23440 47076 24685 47104
rect 23440 47064 23446 47076
rect 24673 47073 24685 47076
rect 24719 47073 24731 47107
rect 24673 47067 24731 47073
rect 25774 47064 25780 47116
rect 25832 47104 25838 47116
rect 26053 47107 26111 47113
rect 26053 47104 26065 47107
rect 25832 47076 26065 47104
rect 25832 47064 25838 47076
rect 26053 47073 26065 47076
rect 26099 47073 26111 47107
rect 28718 47104 28724 47116
rect 26053 47067 26111 47073
rect 27356 47076 27936 47104
rect 28679 47076 28724 47104
rect 27356 47048 27384 47076
rect 22649 47039 22707 47045
rect 22428 47008 22473 47036
rect 22428 46996 22434 47008
rect 22649 47005 22661 47039
rect 22695 47005 22707 47039
rect 22649 46999 22707 47005
rect 23566 46996 23572 47048
rect 23624 47036 23630 47048
rect 23661 47039 23719 47045
rect 23661 47036 23673 47039
rect 23624 47008 23673 47036
rect 23624 46996 23630 47008
rect 23661 47005 23673 47008
rect 23707 47005 23719 47039
rect 23661 46999 23719 47005
rect 23750 46996 23756 47048
rect 23808 47036 23814 47048
rect 23845 47039 23903 47045
rect 23845 47036 23857 47039
rect 23808 47008 23857 47036
rect 23808 46996 23814 47008
rect 23845 47005 23857 47008
rect 23891 47005 23903 47039
rect 24857 47039 24915 47045
rect 23845 46999 23903 47005
rect 23952 47008 24808 47036
rect 21818 46968 21824 46980
rect 21192 46940 21824 46968
rect 20993 46931 21051 46937
rect 21818 46928 21824 46940
rect 21876 46968 21882 46980
rect 22922 46968 22928 46980
rect 21876 46940 22928 46968
rect 21876 46928 21882 46940
rect 22922 46928 22928 46940
rect 22980 46928 22986 46980
rect 23109 46971 23167 46977
rect 23109 46937 23121 46971
rect 23155 46968 23167 46971
rect 23952 46968 23980 47008
rect 23155 46940 23980 46968
rect 24029 46971 24087 46977
rect 23155 46937 23167 46940
rect 23109 46931 23167 46937
rect 24029 46937 24041 46971
rect 24075 46968 24087 46971
rect 24578 46968 24584 46980
rect 24075 46940 24584 46968
rect 24075 46937 24087 46940
rect 24029 46931 24087 46937
rect 24578 46928 24584 46940
rect 24636 46928 24642 46980
rect 24780 46968 24808 47008
rect 24857 47005 24869 47039
rect 24903 47036 24915 47039
rect 25866 47036 25872 47048
rect 24903 47008 25728 47036
rect 25827 47008 25872 47036
rect 24903 47005 24915 47008
rect 24857 46999 24915 47005
rect 25130 46968 25136 46980
rect 24780 46940 24992 46968
rect 25091 46940 25136 46968
rect 16172 46872 17908 46900
rect 16172 46860 16178 46872
rect 18506 46860 18512 46912
rect 18564 46900 18570 46912
rect 19794 46900 19800 46912
rect 18564 46872 19800 46900
rect 18564 46860 18570 46872
rect 19794 46860 19800 46872
rect 19852 46860 19858 46912
rect 19889 46903 19947 46909
rect 19889 46869 19901 46903
rect 19935 46900 19947 46903
rect 20070 46900 20076 46912
rect 19935 46872 20076 46900
rect 19935 46869 19947 46872
rect 19889 46863 19947 46869
rect 20070 46860 20076 46872
rect 20128 46860 20134 46912
rect 22738 46860 22744 46912
rect 22796 46900 22802 46912
rect 23658 46900 23664 46912
rect 22796 46872 23664 46900
rect 22796 46860 22802 46872
rect 23658 46860 23664 46872
rect 23716 46860 23722 46912
rect 24964 46900 24992 46940
rect 25130 46928 25136 46940
rect 25188 46928 25194 46980
rect 25700 46968 25728 47008
rect 25866 46996 25872 47008
rect 25924 46996 25930 47048
rect 26145 47039 26203 47045
rect 26145 47005 26157 47039
rect 26191 47036 26203 47039
rect 26510 47036 26516 47048
rect 26191 47008 26516 47036
rect 26191 47005 26203 47008
rect 26145 46999 26203 47005
rect 26510 46996 26516 47008
rect 26568 46996 26574 47048
rect 27249 47039 27307 47045
rect 27249 47036 27261 47039
rect 26620 47008 27261 47036
rect 26620 46980 26648 47008
rect 27249 47005 27261 47008
rect 27295 47005 27307 47039
rect 27249 46999 27307 47005
rect 27338 46996 27344 47048
rect 27396 47036 27402 47048
rect 27801 47039 27859 47045
rect 27396 47008 27489 47036
rect 27396 46996 27402 47008
rect 27801 47005 27813 47039
rect 27847 47005 27859 47039
rect 27801 46999 27859 47005
rect 26602 46968 26608 46980
rect 25700 46940 26608 46968
rect 26602 46928 26608 46940
rect 26660 46928 26666 46980
rect 27816 46968 27844 46999
rect 27172 46940 27844 46968
rect 27908 46968 27936 47076
rect 28718 47064 28724 47076
rect 28776 47064 28782 47116
rect 29270 47064 29276 47116
rect 29328 47104 29334 47116
rect 32309 47107 32367 47113
rect 32309 47104 32321 47107
rect 29328 47076 32321 47104
rect 29328 47064 29334 47076
rect 32309 47073 32321 47076
rect 32355 47073 32367 47107
rect 33781 47107 33839 47113
rect 32309 47067 32367 47073
rect 32692 47076 33548 47104
rect 28810 47036 28816 47048
rect 28771 47008 28816 47036
rect 28810 46996 28816 47008
rect 28868 46996 28874 47048
rect 29086 47036 29092 47048
rect 29047 47008 29092 47036
rect 29086 46996 29092 47008
rect 29144 46996 29150 47048
rect 30650 46996 30656 47048
rect 30708 47036 30714 47048
rect 30745 47039 30803 47045
rect 30745 47036 30757 47039
rect 30708 47008 30757 47036
rect 30708 46996 30714 47008
rect 30745 47005 30757 47008
rect 30791 47005 30803 47039
rect 31481 47039 31539 47045
rect 31481 47036 31493 47039
rect 30745 46999 30803 47005
rect 30852 47008 31493 47036
rect 29104 46968 29132 46996
rect 30558 46968 30564 46980
rect 27908 46940 29132 46968
rect 30519 46940 30564 46968
rect 25038 46900 25044 46912
rect 24951 46872 25044 46900
rect 25038 46860 25044 46872
rect 25096 46860 25102 46912
rect 25682 46900 25688 46912
rect 25643 46872 25688 46900
rect 25682 46860 25688 46872
rect 25740 46860 25746 46912
rect 26050 46860 26056 46912
rect 26108 46900 26114 46912
rect 27172 46900 27200 46940
rect 30558 46928 30564 46940
rect 30616 46928 30622 46980
rect 30852 46968 30880 47008
rect 31481 47005 31493 47008
rect 31527 47005 31539 47039
rect 31481 46999 31539 47005
rect 32030 46996 32036 47048
rect 32088 47036 32094 47048
rect 32692 47036 32720 47076
rect 32088 47008 32720 47036
rect 32088 46996 32094 47008
rect 31018 46968 31024 46980
rect 30760 46940 30880 46968
rect 30979 46940 31024 46968
rect 26108 46872 27200 46900
rect 26108 46860 26114 46872
rect 27246 46860 27252 46912
rect 27304 46900 27310 46912
rect 30760 46900 30788 46940
rect 31018 46928 31024 46940
rect 31076 46928 31082 46980
rect 32493 46971 32551 46977
rect 32493 46968 32505 46971
rect 31496 46940 32505 46968
rect 31496 46912 31524 46940
rect 32493 46937 32505 46940
rect 32539 46937 32551 46971
rect 32493 46931 32551 46937
rect 30926 46900 30932 46912
rect 27304 46872 30788 46900
rect 30887 46872 30932 46900
rect 27304 46860 27310 46872
rect 30926 46860 30932 46872
rect 30984 46860 30990 46912
rect 31478 46860 31484 46912
rect 31536 46860 31542 46912
rect 31754 46860 31760 46912
rect 31812 46900 31818 46912
rect 32692 46909 32720 47008
rect 32861 47039 32919 47045
rect 32861 47005 32873 47039
rect 32907 47036 32919 47039
rect 33318 47036 33324 47048
rect 32907 47008 33324 47036
rect 32907 47005 32919 47008
rect 32861 46999 32919 47005
rect 33318 46996 33324 47008
rect 33376 46996 33382 47048
rect 33226 46928 33232 46980
rect 33284 46968 33290 46980
rect 33413 46971 33471 46977
rect 33413 46968 33425 46971
rect 33284 46940 33425 46968
rect 33284 46928 33290 46940
rect 33413 46937 33425 46940
rect 33459 46937 33471 46971
rect 33520 46968 33548 47076
rect 33781 47073 33793 47107
rect 33827 47104 33839 47107
rect 34238 47104 34244 47116
rect 33827 47076 34244 47104
rect 33827 47073 33839 47076
rect 33781 47067 33839 47073
rect 34238 47064 34244 47076
rect 34296 47064 34302 47116
rect 34514 47064 34520 47116
rect 34572 47104 34578 47116
rect 35529 47107 35587 47113
rect 35529 47104 35541 47107
rect 34572 47076 35541 47104
rect 34572 47064 34578 47076
rect 35529 47073 35541 47076
rect 35575 47073 35587 47107
rect 37553 47107 37611 47113
rect 37553 47104 37565 47107
rect 35529 47067 35587 47073
rect 35634 47076 37565 47104
rect 33594 46996 33600 47048
rect 33652 47036 33658 47048
rect 33870 47036 33876 47048
rect 33652 47008 33697 47036
rect 33831 47008 33876 47036
rect 33652 46996 33658 47008
rect 33870 46996 33876 47008
rect 33928 46996 33934 47048
rect 34698 46996 34704 47048
rect 34756 47036 34762 47048
rect 34885 47039 34943 47045
rect 34885 47036 34897 47039
rect 34756 47008 34897 47036
rect 34756 46996 34762 47008
rect 34885 47005 34897 47008
rect 34931 47005 34943 47039
rect 34885 46999 34943 47005
rect 35634 46968 35662 47076
rect 37553 47073 37565 47076
rect 37599 47073 37611 47107
rect 37553 47067 37611 47073
rect 37734 47064 37740 47116
rect 37792 47104 37798 47116
rect 39482 47104 39488 47116
rect 37792 47076 39488 47104
rect 37792 47064 37798 47076
rect 35894 46996 35900 47048
rect 35952 47036 35958 47048
rect 36814 47036 36820 47048
rect 35952 47008 36820 47036
rect 35952 46996 35958 47008
rect 36814 46996 36820 47008
rect 36872 46996 36878 47048
rect 37461 47039 37519 47045
rect 37461 47005 37473 47039
rect 37507 47036 37519 47039
rect 37642 47036 37648 47048
rect 37507 47008 37648 47036
rect 37507 47005 37519 47008
rect 37461 46999 37519 47005
rect 37642 46996 37648 47008
rect 37700 46996 37706 47048
rect 37844 47045 37872 47076
rect 39482 47064 39488 47076
rect 39540 47064 39546 47116
rect 37829 47039 37887 47045
rect 37829 47005 37841 47039
rect 37875 47005 37887 47039
rect 38010 47036 38016 47048
rect 37971 47008 38016 47036
rect 37829 46999 37887 47005
rect 38010 46996 38016 47008
rect 38068 46996 38074 47048
rect 38473 47039 38531 47045
rect 38473 47005 38485 47039
rect 38519 47005 38531 47039
rect 38473 46999 38531 47005
rect 40037 47039 40095 47045
rect 40037 47005 40049 47039
rect 40083 47036 40095 47039
rect 40126 47036 40132 47048
rect 40083 47008 40132 47036
rect 40083 47005 40095 47008
rect 40037 46999 40095 47005
rect 38488 46968 38516 46999
rect 40126 46996 40132 47008
rect 40184 46996 40190 47048
rect 40678 47036 40684 47048
rect 40639 47008 40684 47036
rect 40678 46996 40684 47008
rect 40736 46996 40742 47048
rect 41509 47039 41567 47045
rect 41509 47036 41521 47039
rect 41156 47008 41521 47036
rect 33520 46940 35662 46968
rect 36740 46940 38516 46968
rect 33413 46931 33471 46937
rect 32585 46903 32643 46909
rect 32585 46900 32597 46903
rect 31812 46872 32597 46900
rect 31812 46860 31818 46872
rect 32585 46869 32597 46872
rect 32631 46869 32643 46903
rect 32585 46863 32643 46869
rect 32677 46903 32735 46909
rect 32677 46869 32689 46903
rect 32723 46869 32735 46903
rect 32677 46863 32735 46869
rect 32766 46860 32772 46912
rect 32824 46900 32830 46912
rect 36740 46900 36768 46940
rect 32824 46872 36768 46900
rect 32824 46860 32830 46872
rect 37734 46860 37740 46912
rect 37792 46900 37798 46912
rect 38378 46900 38384 46912
rect 37792 46872 38384 46900
rect 37792 46860 37798 46872
rect 38378 46860 38384 46872
rect 38436 46900 38442 46912
rect 39666 46900 39672 46912
rect 38436 46872 39672 46900
rect 38436 46860 38442 46872
rect 39666 46860 39672 46872
rect 39724 46860 39730 46912
rect 40218 46860 40224 46912
rect 40276 46900 40282 46912
rect 41156 46900 41184 47008
rect 41509 47005 41521 47008
rect 41555 47005 41567 47039
rect 43254 47036 43260 47048
rect 43215 47008 43260 47036
rect 41509 46999 41567 47005
rect 41230 46928 41236 46980
rect 41288 46968 41294 46980
rect 41524 46968 41552 46999
rect 43254 46996 43260 47008
rect 43312 46996 43318 47048
rect 44082 46968 44088 46980
rect 41288 46940 41368 46968
rect 41524 46940 44088 46968
rect 41288 46928 41294 46940
rect 41340 46909 41368 46940
rect 44082 46928 44088 46940
rect 44140 46928 44146 46980
rect 40276 46872 41184 46900
rect 41325 46903 41383 46909
rect 40276 46860 40282 46872
rect 41325 46869 41337 46903
rect 41371 46869 41383 46903
rect 41325 46863 41383 46869
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 17313 46699 17371 46705
rect 17313 46665 17325 46699
rect 17359 46696 17371 46699
rect 19334 46696 19340 46708
rect 17359 46668 19340 46696
rect 17359 46665 17371 46668
rect 17313 46659 17371 46665
rect 19334 46656 19340 46668
rect 19392 46656 19398 46708
rect 19426 46656 19432 46708
rect 19484 46656 19490 46708
rect 19886 46656 19892 46708
rect 19944 46696 19950 46708
rect 21177 46699 21235 46705
rect 19944 46668 20576 46696
rect 19944 46656 19950 46668
rect 18322 46588 18328 46640
rect 18380 46628 18386 46640
rect 19444 46628 19472 46656
rect 20438 46628 20444 46640
rect 18380 46600 19472 46628
rect 19720 46600 20444 46628
rect 18380 46588 18386 46600
rect 6914 46520 6920 46572
rect 6972 46560 6978 46572
rect 14642 46560 14648 46572
rect 6972 46532 7017 46560
rect 14603 46532 14648 46560
rect 6972 46520 6978 46532
rect 14642 46520 14648 46532
rect 14700 46520 14706 46572
rect 17129 46563 17187 46569
rect 17129 46529 17141 46563
rect 17175 46560 17187 46563
rect 17865 46563 17923 46569
rect 17865 46560 17877 46563
rect 17175 46532 17877 46560
rect 17175 46529 17187 46532
rect 17129 46523 17187 46529
rect 17865 46529 17877 46532
rect 17911 46529 17923 46563
rect 17865 46523 17923 46529
rect 17954 46520 17960 46572
rect 18012 46560 18018 46572
rect 18417 46563 18475 46569
rect 18012 46532 18057 46560
rect 18012 46520 18018 46532
rect 18417 46529 18429 46563
rect 18463 46560 18475 46563
rect 18966 46560 18972 46572
rect 18463 46532 18972 46560
rect 18463 46529 18475 46532
rect 18417 46523 18475 46529
rect 18966 46520 18972 46532
rect 19024 46520 19030 46572
rect 19720 46560 19748 46600
rect 20438 46588 20444 46600
rect 20496 46588 20502 46640
rect 20548 46572 20576 46668
rect 21177 46665 21189 46699
rect 21223 46665 21235 46699
rect 21177 46659 21235 46665
rect 21192 46628 21220 46659
rect 21266 46656 21272 46708
rect 21324 46696 21330 46708
rect 24949 46699 25007 46705
rect 24949 46696 24961 46699
rect 21324 46668 24961 46696
rect 21324 46656 21330 46668
rect 24949 46665 24961 46668
rect 24995 46665 25007 46699
rect 24949 46659 25007 46665
rect 25133 46699 25191 46705
rect 25133 46665 25145 46699
rect 25179 46665 25191 46699
rect 25133 46659 25191 46665
rect 21450 46628 21456 46640
rect 21192 46600 21456 46628
rect 21450 46588 21456 46600
rect 21508 46588 21514 46640
rect 23474 46628 23480 46640
rect 21560 46600 23480 46628
rect 19168 46532 19748 46560
rect 16301 46495 16359 46501
rect 16301 46461 16313 46495
rect 16347 46492 16359 46495
rect 18046 46492 18052 46504
rect 16347 46464 18052 46492
rect 16347 46461 16359 46464
rect 16301 46455 16359 46461
rect 18046 46452 18052 46464
rect 18104 46452 18110 46504
rect 19168 46492 19196 46532
rect 19886 46520 19892 46572
rect 19944 46560 19950 46572
rect 20073 46564 20131 46569
rect 20073 46563 20208 46564
rect 19944 46532 19989 46560
rect 19944 46520 19950 46532
rect 20073 46529 20085 46563
rect 20119 46560 20208 46563
rect 20254 46560 20260 46572
rect 20119 46536 20260 46560
rect 20119 46529 20131 46536
rect 20180 46532 20260 46536
rect 20073 46523 20131 46529
rect 20254 46520 20260 46532
rect 20312 46520 20318 46572
rect 20530 46520 20536 46572
rect 20588 46560 20594 46572
rect 20717 46563 20775 46569
rect 20717 46560 20729 46563
rect 20588 46532 20729 46560
rect 20588 46520 20594 46532
rect 20717 46529 20729 46532
rect 20763 46529 20775 46563
rect 20717 46523 20775 46529
rect 21174 46520 21180 46572
rect 21232 46560 21238 46572
rect 21232 46532 21277 46560
rect 21232 46520 21238 46532
rect 18524 46464 19196 46492
rect 19245 46495 19303 46501
rect 15010 46384 15016 46436
rect 15068 46424 15074 46436
rect 18524 46424 18552 46464
rect 19245 46461 19257 46495
rect 19291 46492 19303 46495
rect 19702 46492 19708 46504
rect 19291 46464 19610 46492
rect 19663 46464 19708 46492
rect 19291 46461 19303 46464
rect 19245 46455 19303 46461
rect 15068 46396 18552 46424
rect 18601 46427 18659 46433
rect 15068 46384 15074 46396
rect 18601 46393 18613 46427
rect 18647 46424 18659 46427
rect 19582 46424 19610 46464
rect 19702 46452 19708 46464
rect 19760 46452 19766 46504
rect 21560 46492 21588 46600
rect 23474 46588 23480 46600
rect 23532 46588 23538 46640
rect 23842 46628 23848 46640
rect 23803 46600 23848 46628
rect 23842 46588 23848 46600
rect 23900 46588 23906 46640
rect 24302 46628 24308 46640
rect 24263 46600 24308 46628
rect 24302 46588 24308 46600
rect 24360 46588 24366 46640
rect 24854 46628 24860 46640
rect 24767 46600 24860 46628
rect 22465 46563 22523 46569
rect 22465 46529 22477 46563
rect 22511 46560 22523 46563
rect 22649 46563 22707 46569
rect 22511 46532 22600 46560
rect 22511 46529 22523 46532
rect 22465 46523 22523 46529
rect 19906 46464 21588 46492
rect 22572 46492 22600 46532
rect 22649 46529 22661 46563
rect 22695 46560 22707 46563
rect 22738 46560 22744 46572
rect 22695 46532 22744 46560
rect 22695 46529 22707 46532
rect 22649 46523 22707 46529
rect 22738 46520 22744 46532
rect 22796 46520 22802 46572
rect 22922 46520 22928 46572
rect 22980 46560 22986 46572
rect 23109 46563 23167 46569
rect 23109 46560 23121 46563
rect 22980 46532 23121 46560
rect 22980 46520 22986 46532
rect 23109 46529 23121 46532
rect 23155 46529 23167 46563
rect 23290 46560 23296 46572
rect 23251 46532 23296 46560
rect 23109 46523 23167 46529
rect 23290 46520 23296 46532
rect 23348 46520 23354 46572
rect 23382 46520 23388 46572
rect 23440 46560 23446 46572
rect 23658 46560 23664 46572
rect 23440 46532 23485 46560
rect 23619 46532 23664 46560
rect 23440 46520 23446 46532
rect 23658 46520 23664 46532
rect 23716 46560 23722 46572
rect 24780 46560 24808 46600
rect 24854 46588 24860 46600
rect 24912 46628 24918 46640
rect 25148 46628 25176 46659
rect 25222 46656 25228 46708
rect 25280 46696 25286 46708
rect 25280 46668 25325 46696
rect 25280 46656 25286 46668
rect 25866 46656 25872 46708
rect 25924 46696 25930 46708
rect 25961 46699 26019 46705
rect 25961 46696 25973 46699
rect 25924 46668 25973 46696
rect 25924 46656 25930 46668
rect 25961 46665 25973 46668
rect 26007 46665 26019 46699
rect 25961 46659 26019 46665
rect 26145 46699 26203 46705
rect 26145 46665 26157 46699
rect 26191 46665 26203 46699
rect 26145 46659 26203 46665
rect 24912 46600 25176 46628
rect 25409 46631 25467 46637
rect 24912 46588 24918 46600
rect 25409 46597 25421 46631
rect 25455 46628 25467 46631
rect 25682 46628 25688 46640
rect 25455 46600 25688 46628
rect 25455 46597 25467 46600
rect 25409 46591 25467 46597
rect 25682 46588 25688 46600
rect 25740 46588 25746 46640
rect 26160 46628 26188 46659
rect 28626 46656 28632 46708
rect 28684 46696 28690 46708
rect 28684 46668 29592 46696
rect 28684 46656 28690 46668
rect 28258 46628 28264 46640
rect 25976 46600 26188 46628
rect 27448 46600 28028 46628
rect 28219 46600 28264 46628
rect 23716 46532 24808 46560
rect 25041 46563 25099 46569
rect 23716 46520 23722 46532
rect 25041 46529 25053 46563
rect 25087 46560 25099 46563
rect 25774 46560 25780 46572
rect 25087 46532 25780 46560
rect 25087 46529 25099 46532
rect 25041 46523 25099 46529
rect 23198 46492 23204 46504
rect 22572 46464 23204 46492
rect 19906 46424 19934 46464
rect 23198 46452 23204 46464
rect 23256 46492 23262 46504
rect 23477 46495 23535 46501
rect 23477 46492 23489 46495
rect 23256 46464 23489 46492
rect 23256 46452 23262 46464
rect 23477 46461 23489 46464
rect 23523 46461 23535 46495
rect 23477 46455 23535 46461
rect 24302 46452 24308 46504
rect 24360 46492 24366 46504
rect 25056 46492 25084 46523
rect 25774 46520 25780 46532
rect 25832 46560 25838 46572
rect 25976 46560 26004 46600
rect 25832 46532 26004 46560
rect 26143 46563 26201 46569
rect 25832 46520 25838 46532
rect 26143 46529 26155 46563
rect 26189 46529 26201 46563
rect 26602 46560 26608 46572
rect 26563 46532 26608 46560
rect 26143 46523 26201 46529
rect 24360 46464 25084 46492
rect 24360 46452 24366 46464
rect 25222 46452 25228 46504
rect 25280 46492 25286 46504
rect 26160 46492 26188 46523
rect 26602 46520 26608 46532
rect 26660 46520 26666 46572
rect 26878 46520 26884 46572
rect 26936 46560 26942 46572
rect 27448 46569 27476 46600
rect 27433 46563 27491 46569
rect 27433 46560 27445 46563
rect 26936 46532 27445 46560
rect 26936 46520 26942 46532
rect 27433 46529 27445 46532
rect 27479 46529 27491 46563
rect 27433 46523 27491 46529
rect 27522 46520 27528 46572
rect 27580 46560 27586 46572
rect 27709 46563 27767 46569
rect 27580 46532 27625 46560
rect 27580 46520 27586 46532
rect 27709 46529 27721 46563
rect 27755 46529 27767 46563
rect 27709 46523 27767 46529
rect 26510 46492 26516 46504
rect 25280 46464 26516 46492
rect 25280 46452 25286 46464
rect 26510 46452 26516 46464
rect 26568 46452 26574 46504
rect 26620 46492 26648 46520
rect 27724 46492 27752 46523
rect 27798 46520 27804 46572
rect 27856 46560 27862 46572
rect 27856 46532 27901 46560
rect 27856 46520 27862 46532
rect 26620 46464 27752 46492
rect 28000 46492 28028 46600
rect 28258 46588 28264 46600
rect 28316 46588 28322 46640
rect 28445 46631 28503 46637
rect 28445 46597 28457 46631
rect 28491 46628 28503 46631
rect 29564 46628 29592 46668
rect 29638 46656 29644 46708
rect 29696 46696 29702 46708
rect 29696 46668 29741 46696
rect 29696 46656 29702 46668
rect 30098 46656 30104 46708
rect 30156 46696 30162 46708
rect 34514 46696 34520 46708
rect 30156 46668 34520 46696
rect 30156 46656 30162 46668
rect 34514 46656 34520 46668
rect 34572 46656 34578 46708
rect 34701 46699 34759 46705
rect 34701 46665 34713 46699
rect 34747 46696 34759 46699
rect 34974 46696 34980 46708
rect 34747 46668 34980 46696
rect 34747 46665 34759 46668
rect 34701 46659 34759 46665
rect 34974 46656 34980 46668
rect 35032 46656 35038 46708
rect 35621 46699 35679 46705
rect 35621 46665 35633 46699
rect 35667 46665 35679 46699
rect 35621 46659 35679 46665
rect 30282 46628 30288 46640
rect 28491 46600 29500 46628
rect 29564 46600 30288 46628
rect 28491 46597 28503 46600
rect 28445 46591 28503 46597
rect 29472 46572 29500 46600
rect 30282 46588 30288 46600
rect 30340 46588 30346 46640
rect 30650 46628 30656 46640
rect 30484 46600 30656 46628
rect 28629 46563 28687 46569
rect 28629 46529 28641 46563
rect 28675 46560 28687 46563
rect 29270 46560 29276 46572
rect 28675 46532 29276 46560
rect 28675 46529 28687 46532
rect 28629 46523 28687 46529
rect 29270 46520 29276 46532
rect 29328 46520 29334 46572
rect 29454 46560 29460 46572
rect 29415 46532 29460 46560
rect 29454 46520 29460 46532
rect 29512 46520 29518 46572
rect 29733 46563 29791 46569
rect 29733 46529 29745 46563
rect 29779 46560 29791 46563
rect 29822 46560 29828 46572
rect 29779 46532 29828 46560
rect 29779 46529 29791 46532
rect 29733 46523 29791 46529
rect 29822 46520 29828 46532
rect 29880 46560 29886 46572
rect 30484 46569 30512 46600
rect 30650 46588 30656 46600
rect 30708 46628 30714 46640
rect 33045 46631 33103 46637
rect 33045 46628 33057 46631
rect 30708 46600 33057 46628
rect 30708 46588 30714 46600
rect 33045 46597 33057 46600
rect 33091 46597 33103 46631
rect 33045 46591 33103 46597
rect 33134 46588 33140 46640
rect 33192 46628 33198 46640
rect 35526 46628 35532 46640
rect 33192 46600 35532 46628
rect 33192 46588 33198 46600
rect 30193 46563 30251 46569
rect 30193 46560 30205 46563
rect 29880 46532 30205 46560
rect 29880 46520 29886 46532
rect 30193 46529 30205 46532
rect 30239 46529 30251 46563
rect 30193 46523 30251 46529
rect 30469 46563 30527 46569
rect 30469 46529 30481 46563
rect 30515 46529 30527 46563
rect 30469 46523 30527 46529
rect 30745 46563 30803 46569
rect 30745 46529 30757 46563
rect 30791 46560 30803 46563
rect 30926 46560 30932 46572
rect 30791 46532 30932 46560
rect 30791 46529 30803 46532
rect 30745 46523 30803 46529
rect 30926 46520 30932 46532
rect 30984 46560 30990 46572
rect 31662 46560 31668 46572
rect 30984 46532 31524 46560
rect 31623 46532 31668 46560
rect 30984 46520 30990 46532
rect 31018 46492 31024 46504
rect 28000 46464 30788 46492
rect 30979 46464 31024 46492
rect 20809 46427 20867 46433
rect 20809 46424 20821 46427
rect 18647 46396 19472 46424
rect 19582 46396 19934 46424
rect 19966 46396 20821 46424
rect 18647 46393 18659 46396
rect 18601 46387 18659 46393
rect 13906 46316 13912 46368
rect 13964 46356 13970 46368
rect 19288 46356 19294 46368
rect 13964 46328 19294 46356
rect 13964 46316 13970 46328
rect 19288 46316 19294 46328
rect 19346 46316 19352 46368
rect 19444 46356 19472 46396
rect 19966 46356 19994 46396
rect 20809 46393 20821 46396
rect 20855 46424 20867 46427
rect 22370 46424 22376 46436
rect 20855 46396 21496 46424
rect 22331 46396 22376 46424
rect 20855 46393 20867 46396
rect 20809 46387 20867 46393
rect 19444 46328 19994 46356
rect 20070 46316 20076 46368
rect 20128 46356 20134 46368
rect 21361 46359 21419 46365
rect 21361 46356 21373 46359
rect 20128 46328 21373 46356
rect 20128 46316 20134 46328
rect 21361 46325 21373 46328
rect 21407 46325 21419 46359
rect 21468 46356 21496 46396
rect 22370 46384 22376 46396
rect 22428 46384 22434 46436
rect 23934 46384 23940 46436
rect 23992 46424 23998 46436
rect 30285 46427 30343 46433
rect 30285 46424 30297 46427
rect 23992 46396 30297 46424
rect 23992 46384 23998 46396
rect 30285 46393 30297 46396
rect 30331 46393 30343 46427
rect 30285 46387 30343 46393
rect 22830 46356 22836 46368
rect 21468 46328 22836 46356
rect 21361 46319 21419 46325
rect 22830 46316 22836 46328
rect 22888 46316 22894 46368
rect 22922 46316 22928 46368
rect 22980 46356 22986 46368
rect 23750 46356 23756 46368
rect 22980 46328 23756 46356
rect 22980 46316 22986 46328
rect 23750 46316 23756 46328
rect 23808 46316 23814 46368
rect 26513 46359 26571 46365
rect 26513 46325 26525 46359
rect 26559 46356 26571 46359
rect 27062 46356 27068 46368
rect 26559 46328 27068 46356
rect 26559 46325 26571 46328
rect 26513 46319 26571 46325
rect 27062 46316 27068 46328
rect 27120 46316 27126 46368
rect 27246 46356 27252 46368
rect 27207 46328 27252 46356
rect 27246 46316 27252 46328
rect 27304 46316 27310 46368
rect 30760 46356 30788 46464
rect 31018 46452 31024 46464
rect 31076 46452 31082 46504
rect 31496 46492 31524 46532
rect 31662 46520 31668 46532
rect 31720 46520 31726 46572
rect 32490 46560 32496 46572
rect 31772 46532 32168 46560
rect 32451 46532 32496 46560
rect 31772 46492 31800 46532
rect 31496 46464 31800 46492
rect 32140 46492 32168 46532
rect 32490 46520 32496 46532
rect 32548 46520 32554 46572
rect 32953 46563 33011 46569
rect 32953 46529 32965 46563
rect 32999 46560 33011 46563
rect 33226 46560 33232 46572
rect 32999 46532 33232 46560
rect 32999 46529 33011 46532
rect 32953 46523 33011 46529
rect 33226 46520 33232 46532
rect 33284 46520 33290 46572
rect 33505 46563 33563 46569
rect 33505 46529 33517 46563
rect 33551 46529 33563 46563
rect 33505 46523 33563 46529
rect 33781 46563 33839 46569
rect 33781 46529 33793 46563
rect 33827 46560 33839 46563
rect 34238 46560 34244 46572
rect 33827 46532 34244 46560
rect 33827 46529 33839 46532
rect 33781 46523 33839 46529
rect 33137 46495 33195 46501
rect 33137 46492 33149 46495
rect 32140 46464 33149 46492
rect 33137 46461 33149 46464
rect 33183 46461 33195 46495
rect 33520 46492 33548 46523
rect 34238 46520 34244 46532
rect 34296 46520 34302 46572
rect 34532 46569 34560 46600
rect 35526 46588 35532 46600
rect 35584 46628 35590 46640
rect 35636 46628 35664 46659
rect 36722 46656 36728 46708
rect 36780 46696 36786 46708
rect 39942 46696 39948 46708
rect 36780 46668 39948 46696
rect 36780 46656 36786 46668
rect 39942 46656 39948 46668
rect 40000 46656 40006 46708
rect 40034 46656 40040 46708
rect 40092 46696 40098 46708
rect 43254 46696 43260 46708
rect 40092 46668 43260 46696
rect 40092 46656 40098 46668
rect 43254 46656 43260 46668
rect 43312 46656 43318 46708
rect 35584 46600 35664 46628
rect 35584 46588 35590 46600
rect 37090 46588 37096 46640
rect 37148 46628 37154 46640
rect 37148 46600 41000 46628
rect 37148 46588 37154 46600
rect 34517 46563 34575 46569
rect 34517 46529 34529 46563
rect 34563 46529 34575 46563
rect 34517 46523 34575 46529
rect 34606 46520 34612 46572
rect 34664 46569 34670 46572
rect 34664 46563 34687 46569
rect 34675 46529 34687 46563
rect 34664 46523 34687 46529
rect 34664 46520 34670 46523
rect 34790 46520 34796 46572
rect 34848 46560 34854 46572
rect 34885 46563 34943 46569
rect 34885 46560 34897 46563
rect 34848 46532 34897 46560
rect 34848 46520 34854 46532
rect 34885 46529 34897 46532
rect 34931 46529 34943 46563
rect 34885 46523 34943 46529
rect 34974 46520 34980 46572
rect 35032 46560 35038 46572
rect 35618 46560 35624 46572
rect 35032 46532 35624 46560
rect 35032 46520 35038 46532
rect 35618 46520 35624 46532
rect 35676 46520 35682 46572
rect 35986 46520 35992 46572
rect 36044 46560 36050 46572
rect 37182 46560 37188 46572
rect 36044 46532 37188 46560
rect 36044 46520 36050 46532
rect 37182 46520 37188 46532
rect 37240 46520 37246 46572
rect 37734 46520 37740 46572
rect 37792 46564 37798 46572
rect 37829 46564 37887 46569
rect 37792 46563 37887 46564
rect 37792 46536 37841 46563
rect 37792 46520 37798 46536
rect 37829 46529 37841 46536
rect 37875 46529 37887 46563
rect 37829 46523 37887 46529
rect 38010 46520 38016 46572
rect 38068 46564 38074 46572
rect 38105 46564 38163 46569
rect 38068 46563 38163 46564
rect 38068 46536 38117 46563
rect 38068 46520 38074 46536
rect 38105 46529 38117 46536
rect 38151 46529 38163 46563
rect 39022 46560 39028 46572
rect 38105 46523 38163 46529
rect 38212 46532 39028 46560
rect 33870 46492 33876 46504
rect 33520 46464 33876 46492
rect 33137 46455 33195 46461
rect 33152 46424 33180 46455
rect 33870 46452 33876 46464
rect 33928 46452 33934 46504
rect 34330 46492 34336 46504
rect 34291 46464 34336 46492
rect 34330 46452 34336 46464
rect 34388 46452 34394 46504
rect 36081 46495 36139 46501
rect 36081 46492 36093 46495
rect 34440 46464 36093 46492
rect 34440 46424 34468 46464
rect 36081 46461 36093 46464
rect 36127 46492 36139 46495
rect 36722 46492 36728 46504
rect 36127 46464 36728 46492
rect 36127 46461 36139 46464
rect 36081 46455 36139 46461
rect 36722 46452 36728 46464
rect 36780 46452 36786 46504
rect 37458 46452 37464 46504
rect 37516 46492 37522 46504
rect 37516 46464 37872 46492
rect 37516 46452 37522 46464
rect 33152 46396 34468 46424
rect 34882 46384 34888 46436
rect 34940 46424 34946 46436
rect 37844 46424 37872 46464
rect 37925 46427 37983 46433
rect 37925 46424 37937 46427
rect 34940 46396 37780 46424
rect 37844 46396 37937 46424
rect 34940 46384 34946 46396
rect 31481 46359 31539 46365
rect 31481 46356 31493 46359
rect 30760 46328 31493 46356
rect 31481 46325 31493 46328
rect 31527 46325 31539 46359
rect 31481 46319 31539 46325
rect 31662 46316 31668 46368
rect 31720 46356 31726 46368
rect 32309 46359 32367 46365
rect 32309 46356 32321 46359
rect 31720 46328 32321 46356
rect 31720 46316 31726 46328
rect 32309 46325 32321 46328
rect 32355 46325 32367 46359
rect 32309 46319 32367 46325
rect 35342 46316 35348 46368
rect 35400 46356 35406 46368
rect 35437 46359 35495 46365
rect 35437 46356 35449 46359
rect 35400 46328 35449 46356
rect 35400 46316 35406 46328
rect 35437 46325 35449 46328
rect 35483 46325 35495 46359
rect 35986 46356 35992 46368
rect 35947 46328 35992 46356
rect 35437 46319 35495 46325
rect 35986 46316 35992 46328
rect 36044 46316 36050 46368
rect 36538 46356 36544 46368
rect 36499 46328 36544 46356
rect 36538 46316 36544 46328
rect 36596 46316 36602 46368
rect 37642 46356 37648 46368
rect 37603 46328 37648 46356
rect 37642 46316 37648 46328
rect 37700 46316 37706 46368
rect 37752 46356 37780 46396
rect 37925 46393 37937 46396
rect 37971 46393 37983 46427
rect 37925 46387 37983 46393
rect 38013 46427 38071 46433
rect 38013 46393 38025 46427
rect 38059 46424 38071 46427
rect 38212 46424 38240 46532
rect 39022 46520 39028 46532
rect 39080 46560 39086 46572
rect 40972 46569 41000 46600
rect 39209 46563 39267 46569
rect 39209 46560 39221 46563
rect 39080 46532 39221 46560
rect 39080 46520 39086 46532
rect 39209 46529 39221 46532
rect 39255 46529 39267 46563
rect 39209 46523 39267 46529
rect 40957 46563 41015 46569
rect 40957 46529 40969 46563
rect 41003 46529 41015 46563
rect 40957 46523 41015 46529
rect 41785 46563 41843 46569
rect 41785 46529 41797 46563
rect 41831 46529 41843 46563
rect 41785 46523 41843 46529
rect 38470 46452 38476 46504
rect 38528 46492 38534 46504
rect 38749 46495 38807 46501
rect 38749 46492 38761 46495
rect 38528 46464 38761 46492
rect 38528 46452 38534 46464
rect 38749 46461 38761 46464
rect 38795 46461 38807 46495
rect 38749 46455 38807 46461
rect 38838 46452 38844 46504
rect 38896 46492 38902 46504
rect 38933 46495 38991 46501
rect 38933 46492 38945 46495
rect 38896 46464 38945 46492
rect 38896 46452 38902 46464
rect 38933 46461 38945 46464
rect 38979 46461 38991 46495
rect 40313 46495 40371 46501
rect 40313 46492 40325 46495
rect 38933 46455 38991 46461
rect 39040 46464 40325 46492
rect 38059 46396 38240 46424
rect 38059 46393 38071 46396
rect 38013 46387 38071 46393
rect 38286 46384 38292 46436
rect 38344 46424 38350 46436
rect 39040 46424 39068 46464
rect 40313 46461 40325 46464
rect 40359 46461 40371 46495
rect 41800 46492 41828 46523
rect 42610 46520 42616 46572
rect 42668 46560 42674 46572
rect 43257 46563 43315 46569
rect 43257 46560 43269 46563
rect 42668 46532 43269 46560
rect 42668 46520 42674 46532
rect 43257 46529 43269 46532
rect 43303 46529 43315 46563
rect 43898 46560 43904 46572
rect 43859 46532 43904 46560
rect 43257 46523 43315 46529
rect 43898 46520 43904 46532
rect 43956 46520 43962 46572
rect 44542 46560 44548 46572
rect 44503 46532 44548 46560
rect 44542 46520 44548 46532
rect 44600 46520 44606 46572
rect 42702 46492 42708 46504
rect 41800 46464 42708 46492
rect 40313 46455 40371 46461
rect 42702 46452 42708 46464
rect 42760 46492 42766 46504
rect 45186 46492 45192 46504
rect 42760 46464 45192 46492
rect 42760 46452 42766 46464
rect 45186 46452 45192 46464
rect 45244 46452 45250 46504
rect 38344 46396 39068 46424
rect 38344 46384 38350 46396
rect 39114 46384 39120 46436
rect 39172 46424 39178 46436
rect 40034 46424 40040 46436
rect 39172 46396 40040 46424
rect 39172 46384 39178 46396
rect 40034 46384 40040 46396
rect 40092 46384 40098 46436
rect 41138 46384 41144 46436
rect 41196 46424 41202 46436
rect 42613 46427 42671 46433
rect 42613 46424 42625 46427
rect 41196 46396 42625 46424
rect 41196 46384 41202 46396
rect 42613 46393 42625 46396
rect 42659 46393 42671 46427
rect 42613 46387 42671 46393
rect 39669 46359 39727 46365
rect 39669 46356 39681 46359
rect 37752 46328 39681 46356
rect 39669 46325 39681 46328
rect 39715 46325 39727 46359
rect 41690 46356 41696 46368
rect 41651 46328 41696 46356
rect 39669 46319 39727 46325
rect 41690 46316 41696 46328
rect 41748 46316 41754 46368
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 17405 46155 17463 46161
rect 17405 46121 17417 46155
rect 17451 46152 17463 46155
rect 18506 46152 18512 46164
rect 17451 46124 18512 46152
rect 17451 46121 17463 46124
rect 17405 46115 17463 46121
rect 18506 46112 18512 46124
rect 18564 46112 18570 46164
rect 19702 46112 19708 46164
rect 19760 46152 19766 46164
rect 19760 46124 20208 46152
rect 19760 46112 19766 46124
rect 12802 46044 12808 46096
rect 12860 46084 12866 46096
rect 19288 46084 19294 46096
rect 12860 46056 19294 46084
rect 12860 46044 12866 46056
rect 19288 46044 19294 46056
rect 19346 46044 19352 46096
rect 19886 46044 19892 46096
rect 19944 46044 19950 46096
rect 20070 46084 20076 46096
rect 20031 46056 20076 46084
rect 20070 46044 20076 46056
rect 20128 46044 20134 46096
rect 20180 46084 20208 46124
rect 20438 46112 20444 46164
rect 20496 46152 20502 46164
rect 23293 46155 23351 46161
rect 23293 46152 23305 46155
rect 20496 46124 23305 46152
rect 20496 46112 20502 46124
rect 23293 46121 23305 46124
rect 23339 46121 23351 46155
rect 23293 46115 23351 46121
rect 25777 46155 25835 46161
rect 25777 46121 25789 46155
rect 25823 46152 25835 46155
rect 26418 46152 26424 46164
rect 25823 46124 26424 46152
rect 25823 46121 25835 46124
rect 25777 46115 25835 46121
rect 26418 46112 26424 46124
rect 26476 46112 26482 46164
rect 27062 46112 27068 46164
rect 27120 46152 27126 46164
rect 27617 46155 27675 46161
rect 27120 46124 27568 46152
rect 27120 46112 27126 46124
rect 21634 46084 21640 46096
rect 20180 46056 21640 46084
rect 21634 46044 21640 46056
rect 21692 46044 21698 46096
rect 23382 46084 23388 46096
rect 22066 46056 23388 46084
rect 19904 46016 19932 46044
rect 20162 46016 20168 46028
rect 18616 45988 20168 46016
rect 17865 45951 17923 45957
rect 17865 45917 17877 45951
rect 17911 45948 17923 45951
rect 18414 45948 18420 45960
rect 17911 45920 18420 45948
rect 17911 45917 17923 45920
rect 17865 45911 17923 45917
rect 18414 45908 18420 45920
rect 18472 45908 18478 45960
rect 18616 45957 18644 45988
rect 20162 45976 20168 45988
rect 20220 46016 20226 46028
rect 22066 46016 22094 46056
rect 23382 46044 23388 46056
rect 23440 46044 23446 46096
rect 25130 46084 25136 46096
rect 25043 46056 25136 46084
rect 25130 46044 25136 46056
rect 25188 46084 25194 46096
rect 25188 46056 25544 46084
rect 25188 46044 25194 46056
rect 20220 45988 20852 46016
rect 20220 45976 20226 45988
rect 18601 45951 18659 45957
rect 18601 45917 18613 45951
rect 18647 45917 18659 45951
rect 18874 45948 18880 45960
rect 18835 45920 18880 45948
rect 18601 45911 18659 45917
rect 18874 45908 18880 45920
rect 18932 45908 18938 45960
rect 19610 45958 19616 45960
rect 19582 45957 19616 45958
rect 19436 45951 19494 45957
rect 19436 45926 19448 45951
rect 19482 45926 19494 45951
rect 18509 45883 18567 45889
rect 18509 45849 18521 45883
rect 18555 45880 18567 45883
rect 18690 45880 18696 45892
rect 18555 45852 18696 45880
rect 18555 45849 18567 45852
rect 18509 45843 18567 45849
rect 18690 45840 18696 45852
rect 18748 45840 18754 45892
rect 19426 45874 19432 45926
rect 19484 45911 19494 45926
rect 19567 45951 19616 45957
rect 19567 45917 19579 45951
rect 19613 45917 19616 45951
rect 19567 45911 19616 45917
rect 19484 45874 19490 45911
rect 19610 45908 19616 45911
rect 19668 45908 19674 45960
rect 19891 45951 19949 45957
rect 19891 45917 19903 45951
rect 19937 45917 19949 45951
rect 20438 45948 20444 45960
rect 19891 45911 19949 45917
rect 20180 45920 20444 45948
rect 19904 45880 19932 45911
rect 20180 45880 20208 45920
rect 20438 45908 20444 45920
rect 20496 45908 20502 45960
rect 20824 45957 20852 45988
rect 21744 45988 22094 46016
rect 20809 45951 20867 45957
rect 20809 45917 20821 45951
rect 20855 45917 20867 45951
rect 20809 45911 20867 45917
rect 21085 45951 21143 45957
rect 21085 45917 21097 45951
rect 21131 45948 21143 45951
rect 21174 45948 21180 45960
rect 21131 45920 21180 45948
rect 21131 45917 21143 45920
rect 21085 45911 21143 45917
rect 21174 45908 21180 45920
rect 21232 45908 21238 45960
rect 21744 45957 21772 45988
rect 22646 45976 22652 46028
rect 22704 46016 22710 46028
rect 23477 46019 23535 46025
rect 23477 46016 23489 46019
rect 22704 45988 23489 46016
rect 22704 45976 22710 45988
rect 23477 45985 23489 45988
rect 23523 45985 23535 46019
rect 23658 46016 23664 46028
rect 23619 45988 23664 46016
rect 23477 45979 23535 45985
rect 23658 45976 23664 45988
rect 23716 45976 23722 46028
rect 23753 46019 23811 46025
rect 23753 45985 23765 46019
rect 23799 46016 23811 46019
rect 23842 46016 23848 46028
rect 23799 45988 23848 46016
rect 23799 45985 23811 45988
rect 23753 45979 23811 45985
rect 23842 45976 23848 45988
rect 23900 45976 23906 46028
rect 25516 46016 25544 46056
rect 25590 46044 25596 46096
rect 25648 46084 25654 46096
rect 27540 46084 27568 46124
rect 27617 46121 27629 46155
rect 27663 46152 27675 46155
rect 27798 46152 27804 46164
rect 27663 46124 27804 46152
rect 27663 46121 27675 46124
rect 27617 46115 27675 46121
rect 27798 46112 27804 46124
rect 27856 46112 27862 46164
rect 27890 46112 27896 46164
rect 27948 46152 27954 46164
rect 30745 46155 30803 46161
rect 30745 46152 30757 46155
rect 27948 46124 30757 46152
rect 27948 46112 27954 46124
rect 30745 46121 30757 46124
rect 30791 46121 30803 46155
rect 30745 46115 30803 46121
rect 34790 46112 34796 46164
rect 34848 46152 34854 46164
rect 35161 46155 35219 46161
rect 35161 46152 35173 46155
rect 34848 46124 35173 46152
rect 34848 46112 34854 46124
rect 35161 46121 35173 46124
rect 35207 46121 35219 46155
rect 37366 46152 37372 46164
rect 37327 46124 37372 46152
rect 35161 46115 35219 46121
rect 37366 46112 37372 46124
rect 37424 46112 37430 46164
rect 38010 46112 38016 46164
rect 38068 46152 38074 46164
rect 38473 46155 38531 46161
rect 38473 46152 38485 46155
rect 38068 46124 38485 46152
rect 38068 46112 38074 46124
rect 38473 46121 38485 46124
rect 38519 46121 38531 46155
rect 38473 46115 38531 46121
rect 38930 46112 38936 46164
rect 38988 46152 38994 46164
rect 41325 46155 41383 46161
rect 41325 46152 41337 46155
rect 38988 46124 41337 46152
rect 38988 46112 38994 46124
rect 41325 46121 41337 46124
rect 41371 46121 41383 46155
rect 41325 46115 41383 46121
rect 41506 46112 41512 46164
rect 41564 46152 41570 46164
rect 41969 46155 42027 46161
rect 41969 46152 41981 46155
rect 41564 46124 41981 46152
rect 41564 46112 41570 46124
rect 41969 46121 41981 46124
rect 42015 46121 42027 46155
rect 41969 46115 42027 46121
rect 42242 46112 42248 46164
rect 42300 46152 42306 46164
rect 42613 46155 42671 46161
rect 42613 46152 42625 46155
rect 42300 46124 42625 46152
rect 42300 46112 42306 46124
rect 42613 46121 42625 46124
rect 42659 46121 42671 46155
rect 42613 46115 42671 46121
rect 43349 46155 43407 46161
rect 43349 46121 43361 46155
rect 43395 46152 43407 46155
rect 44082 46152 44088 46164
rect 43395 46124 44088 46152
rect 43395 46121 43407 46124
rect 43349 46115 43407 46121
rect 44082 46112 44088 46124
rect 44140 46112 44146 46164
rect 27985 46087 28043 46093
rect 27985 46084 27997 46087
rect 25648 46056 27476 46084
rect 27540 46056 27997 46084
rect 25648 46044 25654 46056
rect 26326 46016 26332 46028
rect 25516 45988 26332 46016
rect 26326 45976 26332 45988
rect 26384 45976 26390 46028
rect 26513 46019 26571 46025
rect 26513 45985 26525 46019
rect 26559 46016 26571 46019
rect 27246 46016 27252 46028
rect 26559 45988 27252 46016
rect 26559 45985 26571 45988
rect 26513 45979 26571 45985
rect 27246 45976 27252 45988
rect 27304 45976 27310 46028
rect 27448 45960 27476 46056
rect 27985 46053 27997 46056
rect 28031 46084 28043 46087
rect 28810 46084 28816 46096
rect 28031 46056 28816 46084
rect 28031 46053 28043 46056
rect 27985 46047 28043 46053
rect 28810 46044 28816 46056
rect 28868 46044 28874 46096
rect 29454 46044 29460 46096
rect 29512 46084 29518 46096
rect 31941 46087 31999 46093
rect 31941 46084 31953 46087
rect 29512 46056 31953 46084
rect 29512 46044 29518 46056
rect 31941 46053 31953 46056
rect 31987 46053 31999 46087
rect 31941 46047 31999 46053
rect 35986 46044 35992 46096
rect 36044 46084 36050 46096
rect 36044 46056 37688 46084
rect 36044 46044 36050 46056
rect 27522 45976 27528 46028
rect 27580 46016 27586 46028
rect 28629 46019 28687 46025
rect 27580 45988 28120 46016
rect 27580 45976 27586 45988
rect 21729 45951 21787 45957
rect 21729 45917 21741 45951
rect 21775 45917 21787 45951
rect 21910 45948 21916 45960
rect 21871 45920 21916 45948
rect 21729 45911 21787 45917
rect 21910 45908 21916 45920
rect 21968 45908 21974 45960
rect 22370 45948 22376 45960
rect 22331 45920 22376 45948
rect 22370 45908 22376 45920
rect 22428 45908 22434 45960
rect 22830 45908 22836 45960
rect 22888 45908 22894 45960
rect 23569 45951 23627 45957
rect 23569 45948 23581 45951
rect 22940 45920 23581 45948
rect 20714 45880 20720 45892
rect 19904 45852 20208 45880
rect 20675 45852 20720 45880
rect 20714 45840 20720 45852
rect 20772 45840 20778 45892
rect 22557 45883 22615 45889
rect 22557 45849 22569 45883
rect 22603 45880 22615 45883
rect 22646 45880 22652 45892
rect 22603 45852 22652 45880
rect 22603 45849 22615 45852
rect 22557 45843 22615 45849
rect 22646 45840 22652 45852
rect 22704 45840 22710 45892
rect 22741 45883 22799 45889
rect 22741 45849 22753 45883
rect 22787 45880 22799 45883
rect 22848 45880 22876 45908
rect 22787 45852 22876 45880
rect 22787 45849 22799 45852
rect 22741 45843 22799 45849
rect 16761 45815 16819 45821
rect 16761 45781 16773 45815
rect 16807 45812 16819 45815
rect 17862 45812 17868 45824
rect 16807 45784 17868 45812
rect 16807 45781 16819 45784
rect 16761 45775 16819 45781
rect 17862 45772 17868 45784
rect 17920 45772 17926 45824
rect 18049 45815 18107 45821
rect 18049 45781 18061 45815
rect 18095 45812 18107 45815
rect 19702 45812 19708 45824
rect 18095 45784 19708 45812
rect 18095 45781 18107 45784
rect 18049 45775 18107 45781
rect 19702 45772 19708 45784
rect 19760 45772 19766 45824
rect 19889 45815 19947 45821
rect 19889 45781 19901 45815
rect 19935 45812 19947 45815
rect 20346 45812 20352 45824
rect 19935 45784 20352 45812
rect 19935 45781 19947 45784
rect 19889 45775 19947 45781
rect 20346 45772 20352 45784
rect 20404 45772 20410 45824
rect 21821 45815 21879 45821
rect 21821 45781 21833 45815
rect 21867 45812 21879 45815
rect 22940 45812 22968 45920
rect 23569 45917 23581 45920
rect 23615 45917 23627 45951
rect 23934 45948 23940 45960
rect 23895 45920 23940 45948
rect 23569 45911 23627 45917
rect 23934 45908 23940 45920
rect 23992 45908 23998 45960
rect 24762 45908 24768 45960
rect 24820 45948 24826 45960
rect 24949 45951 25007 45957
rect 24949 45948 24961 45951
rect 24820 45920 24961 45948
rect 24820 45908 24826 45920
rect 24949 45917 24961 45920
rect 24995 45917 25007 45951
rect 24949 45911 25007 45917
rect 25038 45908 25044 45960
rect 25096 45948 25102 45960
rect 25225 45951 25283 45957
rect 25225 45948 25237 45951
rect 25096 45920 25237 45948
rect 25096 45908 25102 45920
rect 25225 45917 25237 45920
rect 25271 45948 25283 45951
rect 26694 45948 26700 45960
rect 25271 45920 26556 45948
rect 26655 45920 26700 45948
rect 25271 45917 25283 45920
rect 25225 45911 25283 45917
rect 23014 45840 23020 45892
rect 23072 45880 23078 45892
rect 26329 45883 26387 45889
rect 26329 45880 26341 45883
rect 23072 45852 26341 45880
rect 23072 45840 23078 45852
rect 26329 45849 26341 45852
rect 26375 45849 26387 45883
rect 26528 45880 26556 45920
rect 26694 45908 26700 45920
rect 26752 45908 26758 45960
rect 26786 45908 26792 45960
rect 26844 45948 26850 45960
rect 27430 45948 27436 45960
rect 26844 45920 26889 45948
rect 27343 45920 27436 45948
rect 26844 45908 26850 45920
rect 27430 45908 27436 45920
rect 27488 45948 27494 45960
rect 28092 45957 28120 45988
rect 28629 45985 28641 46019
rect 28675 46016 28687 46019
rect 28718 46016 28724 46028
rect 28675 45988 28724 46016
rect 28675 45985 28687 45988
rect 28629 45979 28687 45985
rect 28718 45976 28724 45988
rect 28776 46016 28782 46028
rect 29181 46019 29239 46025
rect 28776 45988 29132 46016
rect 28776 45976 28782 45988
rect 27801 45951 27859 45957
rect 27801 45948 27813 45951
rect 27488 45920 27813 45948
rect 27488 45908 27494 45920
rect 27801 45917 27813 45920
rect 27847 45917 27859 45951
rect 27801 45911 27859 45917
rect 28077 45951 28135 45957
rect 28077 45917 28089 45951
rect 28123 45917 28135 45951
rect 28813 45951 28871 45957
rect 28813 45948 28825 45951
rect 28077 45911 28135 45917
rect 28184 45920 28825 45948
rect 28184 45880 28212 45920
rect 28813 45917 28825 45920
rect 28859 45948 28871 45951
rect 28902 45948 28908 45960
rect 28859 45920 28908 45948
rect 28859 45917 28871 45920
rect 28813 45911 28871 45917
rect 28902 45908 28908 45920
rect 28960 45908 28966 45960
rect 29104 45948 29132 45988
rect 29181 45985 29193 46019
rect 29227 46016 29239 46019
rect 30558 46016 30564 46028
rect 29227 45988 30564 46016
rect 29227 45985 29239 45988
rect 29181 45979 29239 45985
rect 30558 45976 30564 45988
rect 30616 45976 30622 46028
rect 31478 46016 31484 46028
rect 31439 45988 31484 46016
rect 31478 45976 31484 45988
rect 31536 45976 31542 46028
rect 31754 46016 31760 46028
rect 31680 45988 31760 46016
rect 30009 45951 30067 45957
rect 30009 45948 30021 45951
rect 29104 45920 30021 45948
rect 30009 45917 30021 45920
rect 30055 45917 30067 45951
rect 30190 45948 30196 45960
rect 30151 45920 30196 45948
rect 30009 45911 30067 45917
rect 30190 45908 30196 45920
rect 30248 45908 30254 45960
rect 30282 45908 30288 45960
rect 30340 45948 30346 45960
rect 31680 45957 31708 45988
rect 31754 45976 31760 45988
rect 31812 45976 31818 46028
rect 32030 46016 32036 46028
rect 31991 45988 32036 46016
rect 32030 45976 32036 45988
rect 32088 45976 32094 46028
rect 35342 46016 35348 46028
rect 35303 45988 35348 46016
rect 35342 45976 35348 45988
rect 35400 45976 35406 46028
rect 35526 46016 35532 46028
rect 35487 45988 35532 46016
rect 35526 45976 35532 45988
rect 35584 45976 35590 46028
rect 36265 46019 36323 46025
rect 36265 45985 36277 46019
rect 36311 46016 36323 46019
rect 37660 46016 37688 46056
rect 37734 46044 37740 46096
rect 37792 46084 37798 46096
rect 37792 46056 37837 46084
rect 37792 46044 37798 46056
rect 38194 46044 38200 46096
rect 38252 46084 38258 46096
rect 40681 46087 40739 46093
rect 40681 46084 40693 46087
rect 38252 46056 40693 46084
rect 38252 46044 38258 46056
rect 40681 46053 40693 46056
rect 40727 46053 40739 46087
rect 40681 46047 40739 46053
rect 39114 46016 39120 46028
rect 36311 45988 37044 46016
rect 37660 45988 38424 46016
rect 36311 45985 36323 45988
rect 36265 45979 36323 45985
rect 31665 45951 31723 45957
rect 30340 45920 30385 45948
rect 30340 45908 30346 45920
rect 31665 45917 31677 45951
rect 31711 45917 31723 45951
rect 31665 45911 31723 45917
rect 32493 45951 32551 45957
rect 32493 45917 32505 45951
rect 32539 45917 32551 45951
rect 32493 45911 32551 45917
rect 33781 45951 33839 45957
rect 33781 45917 33793 45951
rect 33827 45917 33839 45951
rect 33781 45911 33839 45917
rect 26528 45852 28212 45880
rect 26329 45843 26387 45849
rect 28534 45840 28540 45892
rect 28592 45880 28598 45892
rect 28592 45852 30052 45880
rect 28592 45840 28598 45852
rect 21867 45784 22968 45812
rect 21867 45781 21879 45784
rect 21821 45775 21879 45781
rect 23290 45772 23296 45824
rect 23348 45812 23354 45824
rect 24765 45815 24823 45821
rect 24765 45812 24777 45815
rect 23348 45784 24777 45812
rect 23348 45772 23354 45784
rect 24765 45781 24777 45784
rect 24811 45781 24823 45815
rect 24765 45775 24823 45781
rect 24854 45772 24860 45824
rect 24912 45812 24918 45824
rect 26786 45812 26792 45824
rect 24912 45784 26792 45812
rect 24912 45772 24918 45784
rect 26786 45772 26792 45784
rect 26844 45772 26850 45824
rect 28994 45772 29000 45824
rect 29052 45812 29058 45824
rect 29089 45815 29147 45821
rect 29089 45812 29101 45815
rect 29052 45784 29101 45812
rect 29052 45772 29058 45784
rect 29089 45781 29101 45784
rect 29135 45781 29147 45815
rect 29089 45775 29147 45781
rect 29638 45772 29644 45824
rect 29696 45812 29702 45824
rect 29825 45815 29883 45821
rect 29825 45812 29837 45815
rect 29696 45784 29837 45812
rect 29696 45772 29702 45784
rect 29825 45781 29837 45784
rect 29871 45781 29883 45815
rect 30024 45812 30052 45852
rect 32508 45812 32536 45911
rect 33796 45880 33824 45911
rect 33870 45908 33876 45960
rect 33928 45948 33934 45960
rect 35618 45948 35624 45960
rect 33928 45920 33973 45948
rect 35531 45920 35624 45948
rect 33928 45908 33934 45920
rect 35618 45908 35624 45920
rect 35676 45948 35682 45960
rect 36170 45948 36176 45960
rect 35676 45920 36176 45948
rect 35676 45908 35682 45920
rect 36170 45908 36176 45920
rect 36228 45908 36234 45960
rect 36446 45948 36452 45960
rect 36407 45920 36452 45948
rect 36446 45908 36452 45920
rect 36504 45908 36510 45960
rect 36538 45908 36544 45960
rect 36596 45948 36602 45960
rect 36722 45948 36728 45960
rect 36596 45920 36641 45948
rect 36683 45920 36728 45948
rect 36596 45908 36602 45920
rect 36722 45908 36728 45920
rect 36780 45908 36786 45960
rect 36814 45908 36820 45960
rect 36872 45948 36878 45960
rect 37016 45948 37044 45988
rect 37553 45951 37611 45957
rect 37553 45948 37565 45951
rect 36872 45920 36917 45948
rect 37016 45920 37565 45948
rect 36872 45908 36878 45920
rect 37553 45917 37565 45920
rect 37599 45917 37611 45951
rect 37553 45911 37611 45917
rect 37829 45951 37887 45957
rect 37829 45917 37841 45951
rect 37875 45948 37887 45951
rect 38102 45948 38108 45960
rect 37875 45920 38108 45948
rect 37875 45917 37887 45920
rect 37829 45911 37887 45917
rect 38102 45908 38108 45920
rect 38160 45908 38166 45960
rect 38396 45957 38424 45988
rect 38764 45988 39120 46016
rect 38381 45951 38439 45957
rect 38381 45917 38393 45951
rect 38427 45948 38439 45951
rect 38764 45948 38792 45988
rect 39114 45976 39120 45988
rect 39172 45976 39178 46028
rect 39942 45976 39948 46028
rect 40000 46016 40006 46028
rect 40037 46019 40095 46025
rect 40037 46016 40049 46019
rect 40000 45988 40049 46016
rect 40000 45976 40006 45988
rect 40037 45985 40049 45988
rect 40083 45985 40095 46019
rect 40037 45979 40095 45985
rect 38427 45920 38792 45948
rect 38841 45951 38899 45957
rect 38427 45917 38439 45920
rect 38381 45911 38439 45917
rect 38841 45917 38853 45951
rect 38887 45917 38899 45951
rect 39482 45948 39488 45960
rect 39395 45920 39488 45948
rect 38841 45911 38899 45917
rect 37642 45880 37648 45892
rect 33796 45852 37648 45880
rect 37642 45840 37648 45852
rect 37700 45840 37706 45892
rect 38856 45880 38884 45911
rect 39482 45908 39488 45920
rect 39540 45948 39546 45960
rect 40770 45948 40776 45960
rect 39540 45920 40776 45948
rect 39540 45908 39546 45920
rect 40770 45908 40776 45920
rect 40828 45908 40834 45960
rect 40310 45880 40316 45892
rect 38856 45852 40316 45880
rect 40310 45840 40316 45852
rect 40368 45840 40374 45892
rect 30024 45784 32536 45812
rect 29825 45775 29883 45781
rect 32674 45772 32680 45824
rect 32732 45812 32738 45824
rect 33229 45815 33287 45821
rect 33229 45812 33241 45815
rect 32732 45784 33241 45812
rect 32732 45772 32738 45784
rect 33229 45781 33241 45784
rect 33275 45781 33287 45815
rect 33229 45775 33287 45781
rect 34146 45772 34152 45824
rect 34204 45812 34210 45824
rect 35802 45812 35808 45824
rect 34204 45784 35808 45812
rect 34204 45772 34210 45784
rect 35802 45772 35808 45784
rect 35860 45772 35866 45824
rect 36538 45772 36544 45824
rect 36596 45812 36602 45824
rect 36998 45812 37004 45824
rect 36596 45784 37004 45812
rect 36596 45772 36602 45784
rect 36998 45772 37004 45784
rect 37056 45812 37062 45824
rect 39022 45812 39028 45824
rect 37056 45784 39028 45812
rect 37056 45772 37062 45784
rect 39022 45772 39028 45784
rect 39080 45772 39086 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 17218 45568 17224 45620
rect 17276 45608 17282 45620
rect 18141 45611 18199 45617
rect 18141 45608 18153 45611
rect 17276 45580 18153 45608
rect 17276 45568 17282 45580
rect 18141 45577 18153 45580
rect 18187 45608 18199 45611
rect 19426 45608 19432 45620
rect 18187 45580 19432 45608
rect 18187 45577 18199 45580
rect 18141 45571 18199 45577
rect 19426 45568 19432 45580
rect 19484 45568 19490 45620
rect 23014 45608 23020 45620
rect 21008 45580 23020 45608
rect 17681 45543 17739 45549
rect 17681 45509 17693 45543
rect 17727 45540 17739 45543
rect 17862 45540 17868 45552
rect 17727 45512 17868 45540
rect 17727 45509 17739 45512
rect 17681 45503 17739 45509
rect 17862 45500 17868 45512
rect 17920 45500 17926 45552
rect 18414 45500 18420 45552
rect 18472 45540 18478 45552
rect 18877 45543 18935 45549
rect 18877 45540 18889 45543
rect 18472 45512 18889 45540
rect 18472 45500 18478 45512
rect 18877 45509 18889 45512
rect 18923 45509 18935 45543
rect 20714 45540 20720 45552
rect 18877 45503 18935 45509
rect 19628 45512 20720 45540
rect 18322 45472 18328 45484
rect 18283 45444 18328 45472
rect 18322 45432 18328 45444
rect 18380 45432 18386 45484
rect 19628 45481 19656 45512
rect 20714 45500 20720 45512
rect 20772 45500 20778 45552
rect 18969 45475 19027 45481
rect 18969 45441 18981 45475
rect 19015 45441 19027 45475
rect 18969 45435 19027 45441
rect 19613 45475 19671 45481
rect 19613 45441 19625 45475
rect 19659 45441 19671 45475
rect 20162 45472 20168 45484
rect 20123 45444 20168 45472
rect 19613 45435 19671 45441
rect 9674 45364 9680 45416
rect 9732 45404 9738 45416
rect 18984 45404 19012 45435
rect 20162 45432 20168 45444
rect 20220 45432 20226 45484
rect 20438 45432 20444 45484
rect 20496 45472 20502 45484
rect 21008 45472 21036 45580
rect 23014 45568 23020 45580
rect 23072 45568 23078 45620
rect 24581 45611 24639 45617
rect 24581 45577 24593 45611
rect 24627 45577 24639 45611
rect 24581 45571 24639 45577
rect 21269 45543 21327 45549
rect 21269 45509 21281 45543
rect 21315 45540 21327 45543
rect 23753 45543 23811 45549
rect 23753 45540 23765 45543
rect 21315 45512 23765 45540
rect 21315 45509 21327 45512
rect 21269 45503 21327 45509
rect 20496 45444 21036 45472
rect 21085 45475 21143 45481
rect 20496 45432 20502 45444
rect 21085 45441 21097 45475
rect 21131 45472 21143 45475
rect 21358 45472 21364 45484
rect 21131 45444 21364 45472
rect 21131 45441 21143 45444
rect 21085 45435 21143 45441
rect 21358 45432 21364 45444
rect 21416 45432 21422 45484
rect 22572 45481 22600 45512
rect 23753 45509 23765 45512
rect 23799 45509 23811 45543
rect 23753 45503 23811 45509
rect 23842 45500 23848 45552
rect 23900 45540 23906 45552
rect 24596 45540 24624 45571
rect 24854 45568 24860 45620
rect 24912 45608 24918 45620
rect 25409 45611 25467 45617
rect 25409 45608 25421 45611
rect 24912 45580 25421 45608
rect 24912 45568 24918 45580
rect 25409 45577 25421 45580
rect 25455 45577 25467 45611
rect 25409 45571 25467 45577
rect 26326 45568 26332 45620
rect 26384 45608 26390 45620
rect 26878 45608 26884 45620
rect 26384 45580 26884 45608
rect 26384 45568 26390 45580
rect 26878 45568 26884 45580
rect 26936 45568 26942 45620
rect 27982 45568 27988 45620
rect 28040 45608 28046 45620
rect 28040 45580 29132 45608
rect 28040 45568 28046 45580
rect 24713 45543 24771 45549
rect 24713 45540 24725 45543
rect 23900 45512 24624 45540
rect 23900 45500 23906 45512
rect 24688 45509 24725 45540
rect 24759 45540 24771 45543
rect 28994 45540 29000 45552
rect 24759 45512 29000 45540
rect 24759 45509 24771 45512
rect 24688 45503 24771 45509
rect 21453 45475 21511 45481
rect 21453 45441 21465 45475
rect 21499 45472 21511 45475
rect 22557 45475 22615 45481
rect 21499 45444 22416 45472
rect 21499 45441 21511 45444
rect 21453 45435 21511 45441
rect 20073 45407 20131 45413
rect 20073 45404 20085 45407
rect 9732 45376 12434 45404
rect 18984 45376 20085 45404
rect 9732 45364 9738 45376
rect 12406 45336 12434 45376
rect 20073 45373 20085 45376
rect 20119 45373 20131 45407
rect 22189 45407 22247 45413
rect 22189 45404 22201 45407
rect 20073 45367 20131 45373
rect 22066 45376 22201 45404
rect 22066 45336 22094 45376
rect 22189 45373 22201 45376
rect 22235 45404 22247 45407
rect 22278 45404 22284 45416
rect 22235 45376 22284 45404
rect 22235 45373 22247 45376
rect 22189 45367 22247 45373
rect 22278 45364 22284 45376
rect 22336 45364 22342 45416
rect 22388 45413 22416 45444
rect 22557 45441 22569 45475
rect 22603 45441 22615 45475
rect 22738 45472 22744 45484
rect 22699 45444 22744 45472
rect 22557 45435 22615 45441
rect 22738 45432 22744 45444
rect 22796 45432 22802 45484
rect 23477 45475 23535 45481
rect 23477 45441 23489 45475
rect 23523 45441 23535 45475
rect 23477 45435 23535 45441
rect 22373 45407 22431 45413
rect 22373 45373 22385 45407
rect 22419 45373 22431 45407
rect 22373 45367 22431 45373
rect 12406 45308 22094 45336
rect 22388 45336 22416 45367
rect 22462 45364 22468 45416
rect 22520 45404 22526 45416
rect 23492 45404 23520 45435
rect 23566 45432 23572 45484
rect 23624 45481 23630 45484
rect 23624 45475 23673 45481
rect 23624 45441 23627 45475
rect 23661 45472 23673 45475
rect 24489 45475 24547 45481
rect 24489 45472 24501 45475
rect 23661 45444 24501 45472
rect 23661 45441 23673 45444
rect 23624 45435 23673 45441
rect 24489 45441 24501 45444
rect 24535 45441 24547 45475
rect 24489 45435 24547 45441
rect 23624 45432 23630 45435
rect 23750 45404 23756 45416
rect 22520 45376 23756 45404
rect 22520 45364 22526 45376
rect 23750 45364 23756 45376
rect 23808 45364 23814 45416
rect 23845 45407 23903 45413
rect 23845 45373 23857 45407
rect 23891 45404 23903 45407
rect 24688 45404 24716 45503
rect 28994 45500 29000 45512
rect 29052 45500 29058 45552
rect 29104 45540 29132 45580
rect 29270 45568 29276 45620
rect 29328 45608 29334 45620
rect 29822 45608 29828 45620
rect 29328 45580 29828 45608
rect 29328 45568 29334 45580
rect 29822 45568 29828 45580
rect 29880 45568 29886 45620
rect 31662 45608 31668 45620
rect 30392 45580 31668 45608
rect 30392 45540 30420 45580
rect 31662 45568 31668 45580
rect 31720 45568 31726 45620
rect 33318 45568 33324 45620
rect 33376 45608 33382 45620
rect 33965 45611 34023 45617
rect 33965 45608 33977 45611
rect 33376 45580 33977 45608
rect 33376 45568 33382 45580
rect 33965 45577 33977 45580
rect 34011 45608 34023 45611
rect 34606 45608 34612 45620
rect 34011 45580 34612 45608
rect 34011 45577 34023 45580
rect 33965 45571 34023 45577
rect 34606 45568 34612 45580
rect 34664 45568 34670 45620
rect 35069 45611 35127 45617
rect 35069 45577 35081 45611
rect 35115 45608 35127 45611
rect 36446 45608 36452 45620
rect 35115 45580 36452 45608
rect 35115 45577 35127 45580
rect 35069 45571 35127 45577
rect 30558 45540 30564 45552
rect 29104 45512 30420 45540
rect 30519 45512 30564 45540
rect 30558 45500 30564 45512
rect 30616 45500 30622 45552
rect 32769 45543 32827 45549
rect 32769 45509 32781 45543
rect 32815 45540 32827 45543
rect 33134 45540 33140 45552
rect 32815 45512 33140 45540
rect 32815 45509 32827 45512
rect 32769 45503 32827 45509
rect 33134 45500 33140 45512
rect 33192 45500 33198 45552
rect 34514 45540 34520 45552
rect 33428 45512 34520 45540
rect 24854 45472 24860 45484
rect 24815 45444 24860 45472
rect 24854 45432 24860 45444
rect 24912 45432 24918 45484
rect 25593 45475 25651 45481
rect 25593 45441 25605 45475
rect 25639 45472 25651 45475
rect 26053 45475 26111 45481
rect 25639 45444 25820 45472
rect 25639 45441 25651 45444
rect 25593 45435 25651 45441
rect 23891 45376 24716 45404
rect 23891 45373 23903 45376
rect 23845 45367 23903 45373
rect 24305 45339 24363 45345
rect 24305 45336 24317 45339
rect 22388 45308 24317 45336
rect 24305 45305 24317 45308
rect 24351 45305 24363 45339
rect 25792 45336 25820 45444
rect 26053 45441 26065 45475
rect 26099 45441 26111 45475
rect 26053 45435 26111 45441
rect 27249 45475 27307 45481
rect 27249 45441 27261 45475
rect 27295 45472 27307 45475
rect 27338 45472 27344 45484
rect 27295 45444 27344 45472
rect 27295 45441 27307 45444
rect 27249 45435 27307 45441
rect 26068 45404 26096 45435
rect 27338 45432 27344 45444
rect 27396 45432 27402 45484
rect 27614 45432 27620 45484
rect 27672 45472 27678 45484
rect 27801 45475 27859 45481
rect 27801 45472 27813 45475
rect 27672 45444 27813 45472
rect 27672 45432 27678 45444
rect 27801 45441 27813 45444
rect 27847 45441 27859 45475
rect 27982 45472 27988 45484
rect 27943 45444 27988 45472
rect 27801 45435 27859 45441
rect 27982 45432 27988 45444
rect 28040 45432 28046 45484
rect 28261 45475 28319 45481
rect 28261 45441 28273 45475
rect 28307 45472 28319 45475
rect 28718 45472 28724 45484
rect 28307 45444 28724 45472
rect 28307 45441 28319 45444
rect 28261 45435 28319 45441
rect 28718 45432 28724 45444
rect 28776 45432 28782 45484
rect 29178 45481 29184 45484
rect 29147 45475 29184 45481
rect 29147 45441 29159 45475
rect 29147 45435 29184 45441
rect 29178 45432 29184 45435
rect 29236 45432 29242 45484
rect 29549 45475 29607 45481
rect 29549 45472 29561 45475
rect 29288 45444 29561 45472
rect 26510 45404 26516 45416
rect 26068 45376 26516 45404
rect 26510 45364 26516 45376
rect 26568 45404 26574 45416
rect 28000 45404 28028 45432
rect 26568 45376 28028 45404
rect 28736 45404 28764 45432
rect 29288 45404 29316 45444
rect 29549 45441 29561 45444
rect 29595 45472 29607 45475
rect 30101 45475 30159 45481
rect 30101 45472 30113 45475
rect 29595 45444 30113 45472
rect 29595 45441 29607 45444
rect 29549 45435 29607 45441
rect 30101 45441 30113 45444
rect 30147 45441 30159 45475
rect 30282 45472 30288 45484
rect 30243 45444 30288 45472
rect 30101 45435 30159 45441
rect 30282 45432 30288 45444
rect 30340 45432 30346 45484
rect 30377 45475 30435 45481
rect 30377 45441 30389 45475
rect 30423 45472 30435 45475
rect 30742 45472 30748 45484
rect 30423 45444 30748 45472
rect 30423 45441 30435 45444
rect 30377 45435 30435 45441
rect 30742 45432 30748 45444
rect 30800 45432 30806 45484
rect 31573 45475 31631 45481
rect 31573 45441 31585 45475
rect 31619 45472 31631 45475
rect 32306 45472 32312 45484
rect 31619 45444 32312 45472
rect 31619 45441 31631 45444
rect 31573 45435 31631 45441
rect 32306 45432 32312 45444
rect 32364 45432 32370 45484
rect 32585 45475 32643 45481
rect 32585 45441 32597 45475
rect 32631 45441 32643 45475
rect 32585 45435 32643 45441
rect 32861 45475 32919 45481
rect 32861 45441 32873 45475
rect 32907 45472 32919 45475
rect 33428 45472 33456 45512
rect 34514 45500 34520 45512
rect 34572 45500 34578 45552
rect 35084 45540 35112 45571
rect 36446 45568 36452 45580
rect 36504 45568 36510 45620
rect 37826 45568 37832 45620
rect 37884 45608 37890 45620
rect 39206 45608 39212 45620
rect 37884 45580 39212 45608
rect 37884 45568 37890 45580
rect 39206 45568 39212 45580
rect 39264 45568 39270 45620
rect 42702 45608 42708 45620
rect 42615 45580 42708 45608
rect 42702 45568 42708 45580
rect 42760 45568 42766 45620
rect 34808 45512 35112 45540
rect 35161 45543 35219 45549
rect 33594 45472 33600 45484
rect 32907 45444 33456 45472
rect 33555 45444 33600 45472
rect 32907 45441 32919 45444
rect 32861 45435 32919 45441
rect 28736 45376 29316 45404
rect 29457 45407 29515 45413
rect 26568 45364 26574 45376
rect 29457 45373 29469 45407
rect 29503 45404 29515 45407
rect 30300 45404 30328 45432
rect 29503 45376 30328 45404
rect 31297 45407 31355 45413
rect 29503 45373 29515 45376
rect 29457 45367 29515 45373
rect 31297 45373 31309 45407
rect 31343 45404 31355 45407
rect 31754 45404 31760 45416
rect 31343 45376 31760 45404
rect 31343 45373 31355 45376
rect 31297 45367 31355 45373
rect 31754 45364 31760 45376
rect 31812 45404 31818 45416
rect 32122 45404 32128 45416
rect 31812 45376 32128 45404
rect 31812 45364 31818 45376
rect 32122 45364 32128 45376
rect 32180 45364 32186 45416
rect 32600 45404 32628 45435
rect 33594 45432 33600 45444
rect 33652 45432 33658 45484
rect 34057 45475 34115 45481
rect 34057 45441 34069 45475
rect 34103 45472 34115 45475
rect 34701 45475 34759 45481
rect 34701 45472 34713 45475
rect 34103 45444 34713 45472
rect 34103 45441 34115 45444
rect 34057 45435 34115 45441
rect 34701 45441 34713 45444
rect 34747 45441 34759 45475
rect 34701 45435 34759 45441
rect 33226 45404 33232 45416
rect 32600 45376 33232 45404
rect 33226 45364 33232 45376
rect 33284 45364 33290 45416
rect 33856 45407 33914 45413
rect 33856 45373 33868 45407
rect 33902 45404 33914 45407
rect 33962 45404 33968 45416
rect 33902 45376 33968 45404
rect 33902 45373 33914 45376
rect 33856 45367 33914 45373
rect 33962 45364 33968 45376
rect 34020 45364 34026 45416
rect 34146 45404 34152 45416
rect 34107 45376 34152 45404
rect 34146 45364 34152 45376
rect 34204 45364 34210 45416
rect 34238 45364 34244 45416
rect 34296 45404 34302 45416
rect 34808 45404 34836 45512
rect 35161 45509 35173 45543
rect 35207 45540 35219 45543
rect 35434 45540 35440 45552
rect 35207 45512 35440 45540
rect 35207 45509 35219 45512
rect 35161 45503 35219 45509
rect 35434 45500 35440 45512
rect 35492 45500 35498 45552
rect 42720 45540 42748 45568
rect 38580 45512 39804 45540
rect 38580 45484 38608 45512
rect 34885 45475 34943 45481
rect 34885 45441 34897 45475
rect 34931 45441 34943 45475
rect 34885 45435 34943 45441
rect 34296 45376 34836 45404
rect 34900 45404 34928 45435
rect 36170 45432 36176 45484
rect 36228 45472 36234 45484
rect 36630 45472 36636 45484
rect 36228 45444 36321 45472
rect 36591 45444 36636 45472
rect 36228 45432 36234 45444
rect 36630 45432 36636 45444
rect 36688 45432 36694 45484
rect 37829 45475 37887 45481
rect 37829 45441 37841 45475
rect 37875 45472 37887 45475
rect 38010 45472 38016 45484
rect 37875 45444 38016 45472
rect 37875 45441 37887 45444
rect 37829 45435 37887 45441
rect 38010 45432 38016 45444
rect 38068 45432 38074 45484
rect 38286 45472 38292 45484
rect 38199 45444 38292 45472
rect 38286 45432 38292 45444
rect 38344 45472 38350 45484
rect 38562 45472 38568 45484
rect 38344 45444 38568 45472
rect 38344 45432 38350 45444
rect 38562 45432 38568 45444
rect 38620 45432 38626 45484
rect 38654 45432 38660 45484
rect 38712 45472 38718 45484
rect 39776 45481 39804 45512
rect 41386 45512 42748 45540
rect 39117 45475 39175 45481
rect 39117 45472 39129 45475
rect 38712 45444 39129 45472
rect 38712 45432 38718 45444
rect 39117 45441 39129 45444
rect 39163 45441 39175 45475
rect 39117 45435 39175 45441
rect 39761 45475 39819 45481
rect 39761 45441 39773 45475
rect 39807 45472 39819 45475
rect 40126 45472 40132 45484
rect 39807 45444 40132 45472
rect 39807 45441 39819 45444
rect 39761 45435 39819 45441
rect 40126 45432 40132 45444
rect 40184 45432 40190 45484
rect 40310 45432 40316 45484
rect 40368 45472 40374 45484
rect 40405 45475 40463 45481
rect 40405 45472 40417 45475
rect 40368 45444 40417 45472
rect 40368 45432 40374 45444
rect 40405 45441 40417 45444
rect 40451 45472 40463 45475
rect 41386 45472 41414 45512
rect 40451 45444 41414 45472
rect 40451 45441 40463 45444
rect 40405 45435 40463 45441
rect 35618 45404 35624 45416
rect 34900 45376 35624 45404
rect 34296 45364 34302 45376
rect 35618 45364 35624 45376
rect 35676 45364 35682 45416
rect 35713 45407 35771 45413
rect 35713 45373 35725 45407
rect 35759 45404 35771 45407
rect 35894 45404 35900 45416
rect 35759 45376 35900 45404
rect 35759 45373 35771 45376
rect 35713 45367 35771 45373
rect 35894 45364 35900 45376
rect 35952 45364 35958 45416
rect 36188 45404 36216 45432
rect 36188 45376 37228 45404
rect 37200 45348 37228 45376
rect 37458 45364 37464 45416
rect 37516 45404 37522 45416
rect 37918 45404 37924 45416
rect 37516 45376 37924 45404
rect 37516 45364 37522 45376
rect 37918 45364 37924 45376
rect 37976 45364 37982 45416
rect 38102 45364 38108 45416
rect 38160 45404 38166 45416
rect 38160 45376 40264 45404
rect 38160 45364 38166 45376
rect 25866 45336 25872 45348
rect 25779 45308 25872 45336
rect 24305 45299 24363 45305
rect 25866 45296 25872 45308
rect 25924 45336 25930 45348
rect 27338 45336 27344 45348
rect 25924 45308 27344 45336
rect 25924 45296 25930 45308
rect 27338 45296 27344 45308
rect 27396 45296 27402 45348
rect 27614 45296 27620 45348
rect 27672 45336 27678 45348
rect 29086 45336 29092 45348
rect 27672 45308 29092 45336
rect 27672 45296 27678 45308
rect 29086 45296 29092 45308
rect 29144 45336 29150 45348
rect 30190 45336 30196 45348
rect 29144 45308 30196 45336
rect 29144 45296 29150 45308
rect 30190 45296 30196 45308
rect 30248 45296 30254 45348
rect 36722 45336 36728 45348
rect 36683 45308 36728 45336
rect 36722 45296 36728 45308
rect 36780 45296 36786 45348
rect 37182 45296 37188 45348
rect 37240 45336 37246 45348
rect 40236 45345 40264 45376
rect 38933 45339 38991 45345
rect 38933 45336 38945 45339
rect 37240 45308 38945 45336
rect 37240 45296 37246 45308
rect 38933 45305 38945 45308
rect 38979 45305 38991 45339
rect 38933 45299 38991 45305
rect 40221 45339 40279 45345
rect 40221 45305 40233 45339
rect 40267 45305 40279 45339
rect 40221 45299 40279 45305
rect 40402 45296 40408 45348
rect 40460 45336 40466 45348
rect 40865 45339 40923 45345
rect 40865 45336 40877 45339
rect 40460 45308 40877 45336
rect 40460 45296 40466 45308
rect 40865 45305 40877 45308
rect 40911 45305 40923 45339
rect 40865 45299 40923 45305
rect 18966 45228 18972 45280
rect 19024 45268 19030 45280
rect 19521 45271 19579 45277
rect 19521 45268 19533 45271
rect 19024 45240 19533 45268
rect 19024 45228 19030 45240
rect 19521 45237 19533 45240
rect 19567 45237 19579 45271
rect 19521 45231 19579 45237
rect 25774 45228 25780 45280
rect 25832 45268 25838 45280
rect 26237 45271 26295 45277
rect 26237 45268 26249 45271
rect 25832 45240 26249 45268
rect 25832 45228 25838 45240
rect 26237 45237 26249 45240
rect 26283 45268 26295 45271
rect 26326 45268 26332 45280
rect 26283 45240 26332 45268
rect 26283 45237 26295 45240
rect 26237 45231 26295 45237
rect 26326 45228 26332 45240
rect 26384 45228 26390 45280
rect 26510 45268 26516 45280
rect 26471 45240 26516 45268
rect 26510 45228 26516 45240
rect 26568 45228 26574 45280
rect 27798 45228 27804 45280
rect 27856 45268 27862 45280
rect 27893 45271 27951 45277
rect 27893 45268 27905 45271
rect 27856 45240 27905 45268
rect 27856 45228 27862 45240
rect 27893 45237 27905 45240
rect 27939 45237 27951 45271
rect 27893 45231 27951 45237
rect 28626 45228 28632 45280
rect 28684 45268 28690 45280
rect 28997 45271 29055 45277
rect 28997 45268 29009 45271
rect 28684 45240 29009 45268
rect 28684 45228 28690 45240
rect 28997 45237 29009 45240
rect 29043 45237 29055 45271
rect 28997 45231 29055 45237
rect 29178 45228 29184 45280
rect 29236 45268 29242 45280
rect 29730 45268 29736 45280
rect 29236 45240 29736 45268
rect 29236 45228 29242 45240
rect 29730 45228 29736 45240
rect 29788 45228 29794 45280
rect 31018 45228 31024 45280
rect 31076 45268 31082 45280
rect 31205 45271 31263 45277
rect 31205 45268 31217 45271
rect 31076 45240 31217 45268
rect 31076 45228 31082 45240
rect 31205 45237 31217 45240
rect 31251 45237 31263 45271
rect 32398 45268 32404 45280
rect 32359 45240 32404 45268
rect 31205 45231 31263 45237
rect 32398 45228 32404 45240
rect 32456 45228 32462 45280
rect 32582 45228 32588 45280
rect 32640 45268 32646 45280
rect 33413 45271 33471 45277
rect 33413 45268 33425 45271
rect 32640 45240 33425 45268
rect 32640 45228 32646 45240
rect 33413 45237 33425 45240
rect 33459 45237 33471 45271
rect 33413 45231 33471 45237
rect 35526 45228 35532 45280
rect 35584 45268 35590 45280
rect 35897 45271 35955 45277
rect 35897 45268 35909 45271
rect 35584 45240 35909 45268
rect 35584 45228 35590 45240
rect 35897 45237 35909 45240
rect 35943 45237 35955 45271
rect 38378 45268 38384 45280
rect 38339 45240 38384 45268
rect 35897 45231 35955 45237
rect 38378 45228 38384 45240
rect 38436 45228 38442 45280
rect 39022 45228 39028 45280
rect 39080 45268 39086 45280
rect 39577 45271 39635 45277
rect 39577 45268 39589 45271
rect 39080 45240 39589 45268
rect 39080 45228 39086 45240
rect 39577 45237 39589 45240
rect 39623 45237 39635 45271
rect 39577 45231 39635 45237
rect 41138 45228 41144 45280
rect 41196 45268 41202 45280
rect 41509 45271 41567 45277
rect 41509 45268 41521 45271
rect 41196 45240 41521 45268
rect 41196 45228 41202 45240
rect 41509 45237 41521 45240
rect 41555 45237 41567 45271
rect 41509 45231 41567 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 19797 45067 19855 45073
rect 19797 45033 19809 45067
rect 19843 45064 19855 45067
rect 20530 45064 20536 45076
rect 19843 45036 20536 45064
rect 19843 45033 19855 45036
rect 19797 45027 19855 45033
rect 20530 45024 20536 45036
rect 20588 45024 20594 45076
rect 23477 45067 23535 45073
rect 23477 45033 23489 45067
rect 23523 45064 23535 45067
rect 23566 45064 23572 45076
rect 23523 45036 23572 45064
rect 23523 45033 23535 45036
rect 23477 45027 23535 45033
rect 23566 45024 23572 45036
rect 23624 45024 23630 45076
rect 25424 45036 29776 45064
rect 20162 44956 20168 45008
rect 20220 44996 20226 45008
rect 20441 44999 20499 45005
rect 20441 44996 20453 44999
rect 20220 44968 20453 44996
rect 20220 44956 20226 44968
rect 20441 44965 20453 44968
rect 20487 44965 20499 44999
rect 20441 44959 20499 44965
rect 20456 44928 20484 44959
rect 23658 44956 23664 45008
rect 23716 44996 23722 45008
rect 25424 44996 25452 45036
rect 23716 44968 25452 44996
rect 27540 44968 28948 44996
rect 23716 44956 23722 44968
rect 25038 44928 25044 44940
rect 20456 44900 21220 44928
rect 18690 44860 18696 44872
rect 18651 44832 18696 44860
rect 18690 44820 18696 44832
rect 18748 44820 18754 44872
rect 19978 44860 19984 44872
rect 19939 44832 19984 44860
rect 19978 44820 19984 44832
rect 20036 44820 20042 44872
rect 20625 44863 20683 44869
rect 20625 44829 20637 44863
rect 20671 44860 20683 44863
rect 20990 44860 20996 44872
rect 20671 44832 20996 44860
rect 20671 44829 20683 44832
rect 20625 44823 20683 44829
rect 20990 44820 20996 44832
rect 21048 44820 21054 44872
rect 21192 44869 21220 44900
rect 23676 44900 25044 44928
rect 21177 44863 21235 44869
rect 21177 44829 21189 44863
rect 21223 44829 21235 44863
rect 21450 44860 21456 44872
rect 21411 44832 21456 44860
rect 21177 44823 21235 44829
rect 21450 44820 21456 44832
rect 21508 44820 21514 44872
rect 22370 44860 22376 44872
rect 22331 44832 22376 44860
rect 22370 44820 22376 44832
rect 22428 44820 22434 44872
rect 23676 44869 23704 44900
rect 25038 44888 25044 44900
rect 25096 44888 25102 44940
rect 25961 44931 26019 44937
rect 25961 44897 25973 44931
rect 26007 44928 26019 44931
rect 26973 44931 27031 44937
rect 26973 44928 26985 44931
rect 26007 44900 26985 44928
rect 26007 44897 26019 44900
rect 25961 44891 26019 44897
rect 26973 44897 26985 44900
rect 27019 44897 27031 44931
rect 26973 44891 27031 44897
rect 22833 44863 22891 44869
rect 22833 44829 22845 44863
rect 22879 44829 22891 44863
rect 22833 44823 22891 44829
rect 23661 44863 23719 44869
rect 23661 44829 23673 44863
rect 23707 44829 23719 44863
rect 23661 44823 23719 44829
rect 20806 44752 20812 44804
rect 20864 44792 20870 44804
rect 21085 44795 21143 44801
rect 21085 44792 21097 44795
rect 20864 44764 21097 44792
rect 20864 44752 20870 44764
rect 21085 44761 21097 44764
rect 21131 44761 21143 44795
rect 21085 44755 21143 44761
rect 22462 44752 22468 44804
rect 22520 44792 22526 44804
rect 22649 44795 22707 44801
rect 22649 44792 22661 44795
rect 22520 44764 22661 44792
rect 22520 44752 22526 44764
rect 22649 44761 22661 44764
rect 22695 44761 22707 44795
rect 22848 44792 22876 44823
rect 23750 44820 23756 44872
rect 23808 44860 23814 44872
rect 23937 44863 23995 44869
rect 23808 44832 23853 44860
rect 23808 44820 23814 44832
rect 23937 44829 23949 44863
rect 23983 44829 23995 44863
rect 23937 44823 23995 44829
rect 23952 44792 23980 44823
rect 24026 44820 24032 44872
rect 24084 44860 24090 44872
rect 24578 44860 24584 44872
rect 24084 44832 24129 44860
rect 24539 44832 24584 44860
rect 24084 44820 24090 44832
rect 24578 44820 24584 44832
rect 24636 44820 24642 44872
rect 25590 44820 25596 44872
rect 25648 44860 25654 44872
rect 25731 44863 25789 44869
rect 25731 44860 25743 44863
rect 25648 44832 25743 44860
rect 25648 44820 25654 44832
rect 25731 44829 25743 44832
rect 25777 44829 25789 44863
rect 26050 44860 26056 44872
rect 26011 44832 26056 44860
rect 25731 44823 25789 44829
rect 26050 44820 26056 44832
rect 26108 44820 26114 44872
rect 26418 44820 26424 44872
rect 26476 44860 26482 44872
rect 26513 44863 26571 44869
rect 26513 44860 26525 44863
rect 26476 44832 26525 44860
rect 26476 44820 26482 44832
rect 26513 44829 26525 44832
rect 26559 44829 26571 44863
rect 26513 44823 26571 44829
rect 26789 44863 26847 44869
rect 26789 44829 26801 44863
rect 26835 44860 26847 44863
rect 27338 44860 27344 44872
rect 26835 44832 27344 44860
rect 26835 44829 26847 44832
rect 26789 44823 26847 44829
rect 27338 44820 27344 44832
rect 27396 44820 27402 44872
rect 27430 44820 27436 44872
rect 27488 44860 27494 44872
rect 27540 44869 27568 44968
rect 27893 44931 27951 44937
rect 27893 44897 27905 44931
rect 27939 44928 27951 44931
rect 28350 44928 28356 44940
rect 27939 44900 28356 44928
rect 27939 44897 27951 44900
rect 27893 44891 27951 44897
rect 28350 44888 28356 44900
rect 28408 44888 28414 44940
rect 27525 44863 27583 44869
rect 27525 44860 27537 44863
rect 27488 44832 27537 44860
rect 27488 44820 27494 44832
rect 27525 44829 27537 44832
rect 27571 44829 27583 44863
rect 27798 44860 27804 44872
rect 27759 44832 27804 44860
rect 27525 44823 27583 44829
rect 27798 44820 27804 44832
rect 27856 44820 27862 44872
rect 28169 44863 28227 44869
rect 28169 44829 28181 44863
rect 28215 44860 28227 44863
rect 28626 44860 28632 44872
rect 28215 44832 28632 44860
rect 28215 44829 28227 44832
rect 28169 44823 28227 44829
rect 28626 44820 28632 44832
rect 28684 44820 28690 44872
rect 28920 44869 28948 44968
rect 29748 44937 29776 45036
rect 31478 45024 31484 45076
rect 31536 45064 31542 45076
rect 31849 45067 31907 45073
rect 31849 45064 31861 45067
rect 31536 45036 31861 45064
rect 31536 45024 31542 45036
rect 31849 45033 31861 45036
rect 31895 45033 31907 45067
rect 31849 45027 31907 45033
rect 35618 45024 35624 45076
rect 35676 45064 35682 45076
rect 38102 45064 38108 45076
rect 35676 45036 38108 45064
rect 35676 45024 35682 45036
rect 33505 44999 33563 45005
rect 32048 44968 33272 44996
rect 29733 44931 29791 44937
rect 29733 44897 29745 44931
rect 29779 44897 29791 44931
rect 30558 44928 30564 44940
rect 30519 44900 30564 44928
rect 29733 44891 29791 44897
rect 30558 44888 30564 44900
rect 30616 44888 30622 44940
rect 28905 44863 28963 44869
rect 28905 44829 28917 44863
rect 28951 44829 28963 44863
rect 28905 44823 28963 44829
rect 28994 44820 29000 44872
rect 29052 44860 29058 44872
rect 30377 44863 30435 44869
rect 30377 44860 30389 44863
rect 29052 44832 30389 44860
rect 29052 44820 29058 44832
rect 30377 44829 30389 44832
rect 30423 44860 30435 44863
rect 31754 44860 31760 44872
rect 30423 44832 31760 44860
rect 30423 44829 30435 44832
rect 30377 44823 30435 44829
rect 31754 44820 31760 44832
rect 31812 44860 31818 44872
rect 31938 44860 31944 44872
rect 31812 44832 31944 44860
rect 31812 44820 31818 44832
rect 31938 44820 31944 44832
rect 31996 44820 32002 44872
rect 32048 44869 32076 44968
rect 33134 44928 33140 44940
rect 32140 44900 33140 44928
rect 32140 44869 32168 44900
rect 33134 44888 33140 44900
rect 33192 44888 33198 44940
rect 33244 44928 33272 44968
rect 33505 44965 33517 44999
rect 33551 44996 33563 44999
rect 33594 44996 33600 45008
rect 33551 44968 33600 44996
rect 33551 44965 33563 44968
rect 33505 44959 33563 44965
rect 33594 44956 33600 44968
rect 33652 44956 33658 45008
rect 33244 44900 34008 44928
rect 32033 44863 32091 44869
rect 32033 44829 32045 44863
rect 32079 44829 32091 44863
rect 32033 44823 32091 44829
rect 32125 44863 32183 44869
rect 32125 44829 32137 44863
rect 32171 44829 32183 44863
rect 32306 44860 32312 44872
rect 32267 44832 32312 44860
rect 32125 44823 32183 44829
rect 32306 44820 32312 44832
rect 32364 44820 32370 44872
rect 32401 44863 32459 44869
rect 32401 44829 32413 44863
rect 32447 44860 32459 44863
rect 33226 44860 33232 44872
rect 32447 44832 33232 44860
rect 32447 44829 32459 44832
rect 32401 44823 32459 44829
rect 33226 44820 33232 44832
rect 33284 44820 33290 44872
rect 33318 44820 33324 44872
rect 33376 44860 33382 44872
rect 33413 44863 33471 44869
rect 33413 44860 33425 44863
rect 33376 44832 33425 44860
rect 33376 44820 33382 44832
rect 33413 44829 33425 44832
rect 33459 44829 33471 44863
rect 33778 44860 33784 44872
rect 33739 44832 33784 44860
rect 33413 44823 33471 44829
rect 33778 44820 33784 44832
rect 33836 44820 33842 44872
rect 33980 44869 34008 44900
rect 33965 44863 34023 44869
rect 33965 44829 33977 44863
rect 34011 44860 34023 44863
rect 34514 44860 34520 44872
rect 34011 44832 34520 44860
rect 34011 44829 34023 44832
rect 33965 44823 34023 44829
rect 34514 44820 34520 44832
rect 34572 44820 34578 44872
rect 35728 44869 35756 45036
rect 38102 45024 38108 45036
rect 38160 45024 38166 45076
rect 38197 45067 38255 45073
rect 38197 45033 38209 45067
rect 38243 45064 38255 45067
rect 38378 45064 38384 45076
rect 38243 45036 38384 45064
rect 38243 45033 38255 45036
rect 38197 45027 38255 45033
rect 38378 45024 38384 45036
rect 38436 45024 38442 45076
rect 39206 45064 39212 45076
rect 39167 45036 39212 45064
rect 39206 45024 39212 45036
rect 39264 45024 39270 45076
rect 40034 45064 40040 45076
rect 39995 45036 40040 45064
rect 40034 45024 40040 45036
rect 40092 45024 40098 45076
rect 40126 45024 40132 45076
rect 40184 45064 40190 45076
rect 40589 45067 40647 45073
rect 40589 45064 40601 45067
rect 40184 45036 40601 45064
rect 40184 45024 40190 45036
rect 40589 45033 40601 45036
rect 40635 45033 40647 45067
rect 40589 45027 40647 45033
rect 40770 45024 40776 45076
rect 40828 45064 40834 45076
rect 41693 45067 41751 45073
rect 41693 45064 41705 45067
rect 40828 45036 41705 45064
rect 40828 45024 40834 45036
rect 41693 45033 41705 45036
rect 41739 45033 41751 45067
rect 41693 45027 41751 45033
rect 42337 45067 42395 45073
rect 42337 45033 42349 45067
rect 42383 45064 42395 45067
rect 42702 45064 42708 45076
rect 42383 45036 42708 45064
rect 42383 45033 42395 45036
rect 42337 45027 42395 45033
rect 42702 45024 42708 45036
rect 42760 45024 42766 45076
rect 35802 44956 35808 45008
rect 35860 44996 35866 45008
rect 37458 44996 37464 45008
rect 35860 44968 37464 44996
rect 35860 44956 35866 44968
rect 37458 44956 37464 44968
rect 37516 44996 37522 45008
rect 38838 44996 38844 45008
rect 37516 44968 38844 44996
rect 37516 44956 37522 44968
rect 38838 44956 38844 44968
rect 38896 44956 38902 45008
rect 38010 44928 38016 44940
rect 37476 44900 38016 44928
rect 35713 44863 35771 44869
rect 35713 44829 35725 44863
rect 35759 44829 35771 44863
rect 35713 44823 35771 44829
rect 35897 44863 35955 44869
rect 35897 44829 35909 44863
rect 35943 44829 35955 44863
rect 36998 44860 37004 44872
rect 36959 44832 37004 44860
rect 35897 44823 35955 44829
rect 24673 44795 24731 44801
rect 24673 44792 24685 44795
rect 22848 44764 24685 44792
rect 22649 44755 22707 44761
rect 24673 44761 24685 44764
rect 24719 44761 24731 44795
rect 25317 44795 25375 44801
rect 25317 44792 25329 44795
rect 24673 44755 24731 44761
rect 24780 44764 25329 44792
rect 18785 44727 18843 44733
rect 18785 44693 18797 44727
rect 18831 44724 18843 44727
rect 18966 44724 18972 44736
rect 18831 44696 18972 44724
rect 18831 44693 18843 44696
rect 18785 44687 18843 44693
rect 18966 44684 18972 44696
rect 19024 44684 19030 44736
rect 21174 44684 21180 44736
rect 21232 44724 21238 44736
rect 24780 44724 24808 44764
rect 25317 44761 25329 44764
rect 25363 44761 25375 44795
rect 25498 44792 25504 44804
rect 25459 44764 25504 44792
rect 25317 44755 25375 44761
rect 25498 44752 25504 44764
rect 25556 44752 25562 44804
rect 26605 44795 26663 44801
rect 26605 44761 26617 44795
rect 26651 44792 26663 44795
rect 26878 44792 26884 44804
rect 26651 44764 26884 44792
rect 26651 44761 26663 44764
rect 26605 44755 26663 44761
rect 26878 44752 26884 44764
rect 26936 44752 26942 44804
rect 27706 44792 27712 44804
rect 26988 44764 27712 44792
rect 21232 44696 24808 44724
rect 21232 44684 21238 44696
rect 24854 44684 24860 44736
rect 24912 44724 24918 44736
rect 25866 44724 25872 44736
rect 24912 44696 25872 44724
rect 24912 44684 24918 44696
rect 25866 44684 25872 44696
rect 25924 44684 25930 44736
rect 25958 44684 25964 44736
rect 26016 44724 26022 44736
rect 26988 44724 27016 44764
rect 27706 44752 27712 44764
rect 27764 44752 27770 44804
rect 27816 44792 27844 44820
rect 28721 44795 28779 44801
rect 28721 44792 28733 44795
rect 27816 44764 28733 44792
rect 28721 44761 28733 44764
rect 28767 44761 28779 44795
rect 28721 44755 28779 44761
rect 29089 44795 29147 44801
rect 29089 44761 29101 44795
rect 29135 44761 29147 44795
rect 29089 44755 29147 44761
rect 26016 44696 27016 44724
rect 26016 44684 26022 44696
rect 27246 44684 27252 44736
rect 27304 44724 27310 44736
rect 29104 44724 29132 44755
rect 29178 44752 29184 44804
rect 29236 44792 29242 44804
rect 32861 44795 32919 44801
rect 32861 44792 32873 44795
rect 29236 44764 32873 44792
rect 29236 44752 29242 44764
rect 32861 44761 32873 44764
rect 32907 44761 32919 44795
rect 32861 44755 32919 44761
rect 27304 44696 29132 44724
rect 27304 44684 27310 44696
rect 33042 44684 33048 44736
rect 33100 44724 33106 44736
rect 34885 44727 34943 44733
rect 34885 44724 34897 44727
rect 33100 44696 34897 44724
rect 33100 44684 33106 44696
rect 34885 44693 34897 44696
rect 34931 44693 34943 44727
rect 35912 44724 35940 44823
rect 36998 44820 37004 44832
rect 37056 44820 37062 44872
rect 37182 44860 37188 44872
rect 37143 44832 37188 44860
rect 37182 44820 37188 44832
rect 37240 44820 37246 44872
rect 37476 44869 37504 44900
rect 38010 44888 38016 44900
rect 38068 44928 38074 44940
rect 38562 44928 38568 44940
rect 38068 44900 38568 44928
rect 38068 44888 38074 44900
rect 38562 44888 38568 44900
rect 38620 44928 38626 44940
rect 38749 44931 38807 44937
rect 38749 44928 38761 44931
rect 38620 44900 38761 44928
rect 38620 44888 38626 44900
rect 38749 44897 38761 44900
rect 38795 44897 38807 44931
rect 38749 44891 38807 44897
rect 37461 44863 37519 44869
rect 37461 44829 37473 44863
rect 37507 44829 37519 44863
rect 37461 44823 37519 44829
rect 38286 44820 38292 44872
rect 38344 44860 38350 44872
rect 38657 44863 38715 44869
rect 38344 44832 38389 44860
rect 38344 44820 38350 44832
rect 38657 44829 38669 44863
rect 38703 44860 38715 44863
rect 41138 44860 41144 44872
rect 38703 44832 41144 44860
rect 38703 44829 38715 44832
rect 38657 44823 38715 44829
rect 37642 44792 37648 44804
rect 37603 44764 37648 44792
rect 37642 44752 37648 44764
rect 37700 44752 37706 44804
rect 37918 44752 37924 44804
rect 37976 44792 37982 44804
rect 38470 44792 38476 44804
rect 37976 44764 38476 44792
rect 37976 44752 37982 44764
rect 38470 44752 38476 44764
rect 38528 44792 38534 44804
rect 38672 44792 38700 44823
rect 41138 44820 41144 44832
rect 41196 44820 41202 44872
rect 38528 44764 38700 44792
rect 38528 44752 38534 44764
rect 38654 44724 38660 44736
rect 35912 44696 38660 44724
rect 34885 44687 34943 44693
rect 38654 44684 38660 44696
rect 38712 44684 38718 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 18322 44480 18328 44532
rect 18380 44520 18386 44532
rect 19889 44523 19947 44529
rect 19889 44520 19901 44523
rect 18380 44492 19901 44520
rect 18380 44480 18386 44492
rect 19889 44489 19901 44492
rect 19935 44489 19947 44523
rect 19889 44483 19947 44489
rect 19978 44480 19984 44532
rect 20036 44520 20042 44532
rect 20717 44523 20775 44529
rect 20717 44520 20729 44523
rect 20036 44492 20729 44520
rect 20036 44480 20042 44492
rect 20717 44489 20729 44492
rect 20763 44489 20775 44523
rect 20717 44483 20775 44489
rect 21361 44523 21419 44529
rect 21361 44489 21373 44523
rect 21407 44520 21419 44523
rect 22738 44520 22744 44532
rect 21407 44492 22744 44520
rect 21407 44489 21419 44492
rect 21361 44483 21419 44489
rect 22738 44480 22744 44492
rect 22796 44520 22802 44532
rect 25498 44520 25504 44532
rect 22796 44492 25360 44520
rect 25459 44492 25504 44520
rect 22796 44480 22802 44492
rect 22925 44455 22983 44461
rect 22925 44421 22937 44455
rect 22971 44452 22983 44455
rect 23750 44452 23756 44464
rect 22971 44424 23756 44452
rect 22971 44421 22983 44424
rect 22925 44415 22983 44421
rect 23750 44412 23756 44424
rect 23808 44452 23814 44464
rect 24854 44452 24860 44464
rect 23808 44424 24256 44452
rect 24815 44424 24860 44452
rect 23808 44412 23814 44424
rect 18966 44384 18972 44396
rect 18927 44356 18972 44384
rect 18966 44344 18972 44356
rect 19024 44344 19030 44396
rect 19797 44387 19855 44393
rect 19797 44353 19809 44387
rect 19843 44384 19855 44387
rect 20070 44384 20076 44396
rect 19843 44356 20076 44384
rect 19843 44353 19855 44356
rect 19797 44347 19855 44353
rect 20070 44344 20076 44356
rect 20128 44344 20134 44396
rect 20806 44384 20812 44396
rect 20767 44356 20812 44384
rect 20806 44344 20812 44356
rect 20864 44344 20870 44396
rect 20990 44344 20996 44396
rect 21048 44384 21054 44396
rect 21269 44387 21327 44393
rect 21269 44384 21281 44387
rect 21048 44356 21281 44384
rect 21048 44344 21054 44356
rect 21269 44353 21281 44356
rect 21315 44353 21327 44387
rect 22462 44384 22468 44396
rect 22423 44356 22468 44384
rect 21269 44347 21327 44353
rect 22462 44344 22468 44356
rect 22520 44344 22526 44396
rect 23106 44384 23112 44396
rect 23067 44356 23112 44384
rect 23106 44344 23112 44356
rect 23164 44344 23170 44396
rect 23293 44387 23351 44393
rect 23293 44353 23305 44387
rect 23339 44384 23351 44387
rect 23474 44384 23480 44396
rect 23339 44356 23480 44384
rect 23339 44353 23351 44356
rect 23293 44347 23351 44353
rect 23474 44344 23480 44356
rect 23532 44344 23538 44396
rect 24121 44387 24179 44393
rect 24121 44353 24133 44387
rect 24167 44382 24179 44387
rect 24228 44382 24256 44424
rect 24854 44412 24860 44424
rect 24912 44412 24918 44464
rect 25332 44452 25360 44492
rect 25498 44480 25504 44492
rect 25556 44480 25562 44532
rect 27246 44520 27252 44532
rect 27207 44492 27252 44520
rect 27246 44480 27252 44492
rect 27304 44480 27310 44532
rect 27338 44480 27344 44532
rect 27396 44520 27402 44532
rect 30285 44523 30343 44529
rect 27396 44492 29500 44520
rect 27396 44480 27402 44492
rect 25332 44424 26464 44452
rect 25498 44384 25504 44396
rect 24167 44354 24256 44382
rect 25459 44356 25504 44384
rect 24167 44353 24179 44354
rect 24121 44347 24179 44353
rect 25498 44344 25504 44356
rect 25556 44344 25562 44396
rect 25608 44356 26004 44384
rect 23566 44276 23572 44328
rect 23624 44316 23630 44328
rect 23753 44319 23811 44325
rect 23753 44316 23765 44319
rect 23624 44288 23765 44316
rect 23624 44276 23630 44288
rect 23753 44285 23765 44288
rect 23799 44316 23811 44319
rect 24026 44316 24032 44328
rect 23799 44288 24032 44316
rect 23799 44285 23811 44288
rect 23753 44279 23811 44285
rect 24026 44276 24032 44288
rect 24084 44276 24090 44328
rect 24305 44319 24363 44325
rect 24305 44285 24317 44319
rect 24351 44316 24363 44319
rect 25038 44316 25044 44328
rect 24351 44288 25044 44316
rect 24351 44285 24363 44288
rect 24305 44279 24363 44285
rect 25038 44276 25044 44288
rect 25096 44316 25102 44328
rect 25317 44319 25375 44325
rect 25317 44316 25329 44319
rect 25096 44288 25329 44316
rect 25096 44276 25102 44288
rect 25317 44285 25329 44288
rect 25363 44316 25375 44319
rect 25608 44316 25636 44356
rect 25866 44316 25872 44328
rect 25363 44288 25636 44316
rect 25827 44288 25872 44316
rect 25363 44285 25375 44288
rect 25317 44279 25375 44285
rect 25866 44276 25872 44288
rect 25924 44276 25930 44328
rect 25976 44316 26004 44356
rect 26234 44344 26240 44396
rect 26292 44384 26298 44396
rect 26329 44387 26387 44393
rect 26329 44384 26341 44387
rect 26292 44356 26341 44384
rect 26292 44344 26298 44356
rect 26329 44353 26341 44356
rect 26375 44353 26387 44387
rect 26436 44384 26464 44424
rect 26510 44412 26516 44464
rect 26568 44452 26574 44464
rect 27154 44452 27160 44464
rect 26568 44424 27160 44452
rect 26568 44412 26574 44424
rect 27154 44412 27160 44424
rect 27212 44412 27218 44464
rect 29270 44452 29276 44464
rect 27356 44424 29276 44452
rect 27356 44384 27384 44424
rect 29270 44412 29276 44424
rect 29328 44412 29334 44464
rect 26436 44356 27384 44384
rect 26329 44347 26387 44353
rect 27430 44344 27436 44396
rect 27488 44384 27494 44396
rect 29472 44393 29500 44492
rect 30285 44489 30297 44523
rect 30331 44520 30343 44523
rect 30926 44520 30932 44532
rect 30331 44492 30932 44520
rect 30331 44489 30343 44492
rect 30285 44483 30343 44489
rect 30926 44480 30932 44492
rect 30984 44480 30990 44532
rect 36541 44523 36599 44529
rect 36541 44489 36553 44523
rect 36587 44520 36599 44523
rect 37734 44520 37740 44532
rect 36587 44492 37740 44520
rect 36587 44489 36599 44492
rect 36541 44483 36599 44489
rect 37734 44480 37740 44492
rect 37792 44480 37798 44532
rect 38654 44520 38660 44532
rect 38615 44492 38660 44520
rect 38654 44480 38660 44492
rect 38712 44480 38718 44532
rect 40126 44520 40132 44532
rect 40087 44492 40132 44520
rect 40126 44480 40132 44492
rect 40184 44480 40190 44532
rect 41325 44523 41383 44529
rect 41325 44489 41337 44523
rect 41371 44520 41383 44523
rect 42702 44520 42708 44532
rect 41371 44492 42708 44520
rect 41371 44489 41383 44492
rect 41325 44483 41383 44489
rect 42702 44480 42708 44492
rect 42760 44480 42766 44532
rect 32582 44452 32588 44464
rect 31036 44424 32588 44452
rect 29457 44387 29515 44393
rect 27488 44356 27533 44384
rect 27488 44344 27494 44356
rect 29457 44353 29469 44387
rect 29503 44353 29515 44387
rect 29638 44384 29644 44396
rect 29599 44356 29644 44384
rect 29457 44347 29515 44353
rect 27617 44319 27675 44325
rect 27617 44316 27629 44319
rect 25976 44288 27629 44316
rect 27617 44285 27629 44288
rect 27663 44285 27675 44319
rect 27617 44279 27675 44285
rect 27706 44276 27712 44328
rect 27764 44316 27770 44328
rect 28629 44319 28687 44325
rect 28629 44316 28641 44319
rect 27764 44288 28641 44316
rect 27764 44276 27770 44288
rect 28629 44285 28641 44288
rect 28675 44285 28687 44319
rect 29472 44316 29500 44347
rect 29638 44344 29644 44356
rect 29696 44344 29702 44396
rect 30742 44384 30748 44396
rect 29748 44356 30748 44384
rect 29748 44316 29776 44356
rect 30742 44344 30748 44356
rect 30800 44344 30806 44396
rect 30926 44316 30932 44328
rect 29472 44288 29776 44316
rect 30887 44288 30932 44316
rect 28629 44279 28687 44285
rect 30926 44276 30932 44288
rect 30984 44276 30990 44328
rect 19058 44208 19064 44260
rect 19116 44248 19122 44260
rect 19153 44251 19211 44257
rect 19153 44248 19165 44251
rect 19116 44220 19165 44248
rect 19116 44208 19122 44220
rect 19153 44217 19165 44220
rect 19199 44217 19211 44251
rect 19153 44211 19211 44217
rect 21450 44208 21456 44260
rect 21508 44248 21514 44260
rect 23842 44248 23848 44260
rect 21508 44220 23704 44248
rect 23803 44220 23848 44248
rect 21508 44208 21514 44220
rect 22370 44180 22376 44192
rect 22331 44152 22376 44180
rect 22370 44140 22376 44152
rect 22428 44140 22434 44192
rect 23676 44180 23704 44220
rect 23842 44208 23848 44220
rect 23900 44208 23906 44260
rect 31036 44248 31064 44424
rect 32582 44412 32588 44424
rect 32640 44412 32646 44464
rect 33689 44455 33747 44461
rect 33689 44421 33701 44455
rect 33735 44452 33747 44455
rect 33778 44452 33784 44464
rect 33735 44424 33784 44452
rect 33735 44421 33747 44424
rect 33689 44415 33747 44421
rect 33778 44412 33784 44424
rect 33836 44452 33842 44464
rect 34333 44455 34391 44461
rect 34333 44452 34345 44455
rect 33836 44424 34345 44452
rect 33836 44412 33842 44424
rect 34333 44421 34345 44424
rect 34379 44421 34391 44455
rect 34333 44415 34391 44421
rect 38470 44412 38476 44464
rect 38528 44452 38534 44464
rect 38528 44424 39160 44452
rect 38528 44412 38534 44424
rect 31113 44387 31171 44393
rect 31113 44353 31125 44387
rect 31159 44384 31171 44387
rect 32398 44384 32404 44396
rect 31159 44356 32404 44384
rect 31159 44353 31171 44356
rect 31113 44347 31171 44353
rect 32398 44344 32404 44356
rect 32456 44344 32462 44396
rect 33042 44344 33048 44396
rect 33100 44344 33106 44396
rect 33962 44344 33968 44396
rect 34020 44384 34026 44396
rect 34149 44387 34207 44393
rect 34149 44384 34161 44387
rect 34020 44356 34161 44384
rect 34020 44344 34026 44356
rect 34149 44353 34161 44356
rect 34195 44353 34207 44387
rect 34514 44384 34520 44396
rect 34475 44356 34520 44384
rect 34149 44347 34207 44353
rect 34514 44344 34520 44356
rect 34572 44344 34578 44396
rect 35713 44387 35771 44393
rect 35713 44353 35725 44387
rect 35759 44384 35771 44387
rect 36538 44384 36544 44396
rect 35759 44356 36544 44384
rect 35759 44353 35771 44356
rect 35713 44347 35771 44353
rect 36538 44344 36544 44356
rect 36596 44344 36602 44396
rect 37458 44384 37464 44396
rect 37419 44356 37464 44384
rect 37458 44344 37464 44356
rect 37516 44344 37522 44396
rect 37642 44384 37648 44396
rect 37603 44356 37648 44384
rect 37642 44344 37648 44356
rect 37700 44344 37706 44396
rect 38105 44387 38163 44393
rect 38105 44353 38117 44387
rect 38151 44384 38163 44387
rect 38378 44384 38384 44396
rect 38151 44356 38384 44384
rect 38151 44353 38163 44356
rect 38105 44347 38163 44353
rect 38378 44344 38384 44356
rect 38436 44344 38442 44396
rect 38562 44344 38568 44396
rect 38620 44384 38626 44396
rect 38841 44387 38899 44393
rect 38841 44384 38853 44387
rect 38620 44356 38853 44384
rect 38620 44344 38626 44356
rect 38841 44353 38853 44356
rect 38887 44353 38899 44387
rect 39022 44384 39028 44396
rect 38983 44356 39028 44384
rect 38841 44347 38899 44353
rect 39022 44344 39028 44356
rect 39080 44344 39086 44396
rect 39132 44393 39160 44424
rect 40034 44412 40040 44464
rect 40092 44452 40098 44464
rect 40681 44455 40739 44461
rect 40681 44452 40693 44455
rect 40092 44424 40693 44452
rect 40092 44412 40098 44424
rect 40681 44421 40693 44424
rect 40727 44421 40739 44455
rect 40681 44415 40739 44421
rect 39117 44387 39175 44393
rect 39117 44353 39129 44387
rect 39163 44384 39175 44387
rect 39577 44387 39635 44393
rect 39577 44384 39589 44387
rect 39163 44356 39589 44384
rect 39163 44353 39175 44356
rect 39117 44347 39175 44353
rect 39577 44353 39589 44356
rect 39623 44353 39635 44387
rect 39577 44347 39635 44353
rect 32858 44316 32864 44328
rect 32819 44288 32864 44316
rect 32858 44276 32864 44288
rect 32916 44276 32922 44328
rect 35805 44319 35863 44325
rect 35805 44285 35817 44319
rect 35851 44316 35863 44319
rect 35894 44316 35900 44328
rect 35851 44288 35900 44316
rect 35851 44285 35863 44288
rect 35805 44279 35863 44285
rect 35894 44276 35900 44288
rect 35952 44276 35958 44328
rect 23952 44220 27108 44248
rect 23952 44180 23980 44220
rect 23676 44152 23980 44180
rect 27080 44180 27108 44220
rect 28736 44220 31064 44248
rect 28736 44180 28764 44220
rect 37550 44180 37556 44192
rect 27080 44152 28764 44180
rect 37511 44152 37556 44180
rect 37550 44140 37556 44152
rect 37608 44140 37614 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 21177 43979 21235 43985
rect 21177 43945 21189 43979
rect 21223 43976 21235 43979
rect 22094 43976 22100 43988
rect 21223 43948 22100 43976
rect 21223 43945 21235 43948
rect 21177 43939 21235 43945
rect 22094 43936 22100 43948
rect 22152 43936 22158 43988
rect 24946 43936 24952 43988
rect 25004 43976 25010 43988
rect 26145 43979 26203 43985
rect 26145 43976 26157 43979
rect 25004 43948 26157 43976
rect 25004 43936 25010 43948
rect 26145 43945 26157 43948
rect 26191 43945 26203 43979
rect 26145 43939 26203 43945
rect 28997 43979 29055 43985
rect 28997 43945 29009 43979
rect 29043 43976 29055 43979
rect 29086 43976 29092 43988
rect 29043 43948 29092 43976
rect 29043 43945 29055 43948
rect 28997 43939 29055 43945
rect 29086 43936 29092 43948
rect 29144 43936 29150 43988
rect 29362 43936 29368 43988
rect 29420 43976 29426 43988
rect 29733 43979 29791 43985
rect 29733 43976 29745 43979
rect 29420 43948 29745 43976
rect 29420 43936 29426 43948
rect 29733 43945 29745 43948
rect 29779 43945 29791 43979
rect 30926 43976 30932 43988
rect 30887 43948 30932 43976
rect 29733 43939 29791 43945
rect 30926 43936 30932 43948
rect 30984 43936 30990 43988
rect 31757 43979 31815 43985
rect 31757 43945 31769 43979
rect 31803 43976 31815 43979
rect 31803 43948 34100 43976
rect 31803 43945 31815 43948
rect 31757 43939 31815 43945
rect 20625 43911 20683 43917
rect 20625 43877 20637 43911
rect 20671 43908 20683 43911
rect 21818 43908 21824 43920
rect 20671 43880 21824 43908
rect 20671 43877 20683 43880
rect 20625 43871 20683 43877
rect 21818 43868 21824 43880
rect 21876 43868 21882 43920
rect 26418 43908 26424 43920
rect 24872 43880 26424 43908
rect 22649 43843 22707 43849
rect 22649 43809 22661 43843
rect 22695 43840 22707 43843
rect 23198 43840 23204 43852
rect 22695 43812 23204 43840
rect 22695 43809 22707 43812
rect 22649 43803 22707 43809
rect 23198 43800 23204 43812
rect 23256 43800 23262 43852
rect 24872 43849 24900 43880
rect 26418 43868 26424 43880
rect 26476 43868 26482 43920
rect 32858 43908 32864 43920
rect 32600 43880 32864 43908
rect 24857 43843 24915 43849
rect 24857 43809 24869 43843
rect 24903 43809 24915 43843
rect 24857 43803 24915 43809
rect 26694 43800 26700 43852
rect 26752 43840 26758 43852
rect 26789 43843 26847 43849
rect 26789 43840 26801 43843
rect 26752 43812 26801 43840
rect 26752 43800 26758 43812
rect 26789 43809 26801 43812
rect 26835 43809 26847 43843
rect 26789 43803 26847 43809
rect 20990 43732 20996 43784
rect 21048 43772 21054 43784
rect 21637 43775 21695 43781
rect 21637 43772 21649 43775
rect 21048 43744 21649 43772
rect 21048 43732 21054 43744
rect 21637 43741 21649 43744
rect 21683 43741 21695 43775
rect 21637 43735 21695 43741
rect 22370 43732 22376 43784
rect 22428 43772 22434 43784
rect 22925 43775 22983 43781
rect 22925 43772 22937 43775
rect 22428 43744 22937 43772
rect 22428 43732 22434 43744
rect 22925 43741 22937 43744
rect 22971 43741 22983 43775
rect 22925 43735 22983 43741
rect 23385 43775 23443 43781
rect 23385 43741 23397 43775
rect 23431 43772 23443 43775
rect 23842 43772 23848 43784
rect 23431 43744 23848 43772
rect 23431 43741 23443 43744
rect 23385 43735 23443 43741
rect 23842 43732 23848 43744
rect 23900 43732 23906 43784
rect 25958 43772 25964 43784
rect 25346 43758 25964 43772
rect 25332 43744 25964 43758
rect 23474 43664 23480 43716
rect 23532 43704 23538 43716
rect 24854 43704 24860 43716
rect 23532 43676 24860 43704
rect 23532 43664 23538 43676
rect 24854 43664 24860 43676
rect 24912 43704 24918 43716
rect 25332 43704 25360 43744
rect 25958 43732 25964 43744
rect 26016 43732 26022 43784
rect 27154 43772 27160 43784
rect 27115 43744 27160 43772
rect 27154 43732 27160 43744
rect 27212 43732 27218 43784
rect 27614 43772 27620 43784
rect 27575 43744 27620 43772
rect 27614 43732 27620 43744
rect 27672 43732 27678 43784
rect 28350 43772 28356 43784
rect 28311 43744 28356 43772
rect 28350 43732 28356 43744
rect 28408 43732 28414 43784
rect 29178 43772 29184 43784
rect 29139 43744 29184 43772
rect 29178 43732 29184 43744
rect 29236 43732 29242 43784
rect 31018 43772 31024 43784
rect 30979 43744 31024 43772
rect 31018 43732 31024 43744
rect 31076 43732 31082 43784
rect 31662 43772 31668 43784
rect 31623 43744 31668 43772
rect 31662 43732 31668 43744
rect 31720 43732 31726 43784
rect 31849 43775 31907 43781
rect 31849 43741 31861 43775
rect 31895 43741 31907 43775
rect 31849 43735 31907 43741
rect 32493 43775 32551 43781
rect 32493 43741 32505 43775
rect 32539 43772 32551 43775
rect 32600 43772 32628 43880
rect 32858 43868 32864 43880
rect 32916 43868 32922 43920
rect 33134 43908 33140 43920
rect 33095 43880 33140 43908
rect 33134 43868 33140 43880
rect 33192 43868 33198 43920
rect 34072 43908 34100 43948
rect 34146 43936 34152 43988
rect 34204 43976 34210 43988
rect 34241 43979 34299 43985
rect 34241 43976 34253 43979
rect 34204 43948 34253 43976
rect 34204 43936 34210 43948
rect 34241 43945 34253 43948
rect 34287 43945 34299 43979
rect 34241 43939 34299 43945
rect 34514 43936 34520 43988
rect 34572 43976 34578 43988
rect 35529 43979 35587 43985
rect 35529 43976 35541 43979
rect 34572 43948 35541 43976
rect 34572 43936 34578 43948
rect 35529 43945 35541 43948
rect 35575 43945 35587 43979
rect 36538 43976 36544 43988
rect 36499 43948 36544 43976
rect 35529 43939 35587 43945
rect 36538 43936 36544 43948
rect 36596 43936 36602 43988
rect 36814 43976 36820 43988
rect 36775 43948 36820 43976
rect 36814 43936 36820 43948
rect 36872 43936 36878 43988
rect 38470 43936 38476 43988
rect 38528 43976 38534 43988
rect 39025 43979 39083 43985
rect 39025 43976 39037 43979
rect 38528 43948 39037 43976
rect 38528 43936 38534 43948
rect 39025 43945 39037 43948
rect 39071 43945 39083 43979
rect 40126 43976 40132 43988
rect 40087 43948 40132 43976
rect 39025 43939 39083 43945
rect 40126 43936 40132 43948
rect 40184 43936 40190 43988
rect 36630 43908 36636 43920
rect 34072 43880 36636 43908
rect 36630 43868 36636 43880
rect 36688 43868 36694 43920
rect 38565 43911 38623 43917
rect 38565 43877 38577 43911
rect 38611 43908 38623 43911
rect 38838 43908 38844 43920
rect 38611 43880 38844 43908
rect 38611 43877 38623 43880
rect 38565 43871 38623 43877
rect 33042 43840 33048 43852
rect 32692 43812 33048 43840
rect 32692 43781 32720 43812
rect 33042 43800 33048 43812
rect 33100 43840 33106 43852
rect 34977 43843 35035 43849
rect 34977 43840 34989 43843
rect 33100 43812 33548 43840
rect 33100 43800 33106 43812
rect 32539 43744 32628 43772
rect 32677 43775 32735 43781
rect 32539 43741 32551 43744
rect 32493 43735 32551 43741
rect 32677 43741 32689 43775
rect 32723 43741 32735 43775
rect 32677 43735 32735 43741
rect 24912 43676 25360 43704
rect 24912 43664 24918 43676
rect 25498 43664 25504 43716
rect 25556 43704 25562 43716
rect 25682 43704 25688 43716
rect 25556 43676 25688 43704
rect 25556 43664 25562 43676
rect 25682 43664 25688 43676
rect 25740 43664 25746 43716
rect 27430 43664 27436 43716
rect 27488 43704 27494 43716
rect 28445 43707 28503 43713
rect 28445 43704 28457 43707
rect 27488 43676 28457 43704
rect 27488 43664 27494 43676
rect 28445 43673 28457 43676
rect 28491 43673 28503 43707
rect 28445 43667 28503 43673
rect 21818 43596 21824 43648
rect 21876 43636 21882 43648
rect 22186 43636 22192 43648
rect 21876 43608 22192 43636
rect 21876 43596 21882 43608
rect 22186 43596 22192 43608
rect 22244 43596 22250 43648
rect 31864 43636 31892 43735
rect 32858 43732 32864 43784
rect 32916 43772 32922 43784
rect 33520 43781 33548 43812
rect 33980 43812 34989 43840
rect 33980 43781 34008 43812
rect 34977 43809 34989 43812
rect 35023 43840 35035 43843
rect 35434 43840 35440 43852
rect 35023 43812 35440 43840
rect 35023 43809 35035 43812
rect 34977 43803 35035 43809
rect 35434 43800 35440 43812
rect 35492 43800 35498 43852
rect 36814 43840 36820 43852
rect 35728 43812 36820 43840
rect 33505 43775 33563 43781
rect 32916 43744 33364 43772
rect 32916 43732 32922 43744
rect 32309 43707 32367 43713
rect 32309 43673 32321 43707
rect 32355 43704 32367 43707
rect 33042 43704 33048 43716
rect 32355 43676 33048 43704
rect 32355 43673 32367 43676
rect 32309 43667 32367 43673
rect 33042 43664 33048 43676
rect 33100 43664 33106 43716
rect 33336 43713 33364 43744
rect 33505 43741 33517 43775
rect 33551 43741 33563 43775
rect 33505 43735 33563 43741
rect 33965 43775 34023 43781
rect 33965 43741 33977 43775
rect 34011 43741 34023 43775
rect 33965 43735 34023 43741
rect 34149 43775 34207 43781
rect 34149 43741 34161 43775
rect 34195 43772 34207 43775
rect 34238 43772 34244 43784
rect 34195 43744 34244 43772
rect 34195 43741 34207 43744
rect 34149 43735 34207 43741
rect 33321 43707 33379 43713
rect 33321 43673 33333 43707
rect 33367 43704 33379 43707
rect 33980 43704 34008 43735
rect 34238 43732 34244 43744
rect 34296 43732 34302 43784
rect 35728 43781 35756 43812
rect 36814 43800 36820 43812
rect 36872 43800 36878 43852
rect 38580 43840 38608 43871
rect 38838 43868 38844 43880
rect 38896 43868 38902 43920
rect 37752 43812 38608 43840
rect 37752 43784 37780 43812
rect 35713 43775 35771 43781
rect 35713 43741 35725 43775
rect 35759 43741 35771 43775
rect 35713 43735 35771 43741
rect 35897 43775 35955 43781
rect 35897 43741 35909 43775
rect 35943 43772 35955 43775
rect 37001 43775 37059 43781
rect 37001 43772 37013 43775
rect 35943 43744 37013 43772
rect 35943 43741 35955 43744
rect 35897 43735 35955 43741
rect 37001 43741 37013 43744
rect 37047 43772 37059 43775
rect 37553 43775 37611 43781
rect 37553 43772 37565 43775
rect 37047 43744 37565 43772
rect 37047 43741 37059 43744
rect 37001 43735 37059 43741
rect 37553 43741 37565 43744
rect 37599 43741 37611 43775
rect 37553 43735 37611 43741
rect 37734 43732 37740 43784
rect 37792 43772 37798 43784
rect 38013 43775 38071 43781
rect 37792 43744 37885 43772
rect 37792 43732 37798 43744
rect 38013 43741 38025 43775
rect 38059 43772 38071 43775
rect 38378 43772 38384 43784
rect 38059 43744 38384 43772
rect 38059 43741 38071 43744
rect 38013 43735 38071 43741
rect 38378 43732 38384 43744
rect 38436 43732 38442 43784
rect 35986 43704 35992 43716
rect 33367 43676 34008 43704
rect 35947 43676 35992 43704
rect 33367 43673 33379 43676
rect 33321 43667 33379 43673
rect 35986 43664 35992 43676
rect 36044 43664 36050 43716
rect 37642 43664 37648 43716
rect 37700 43704 37706 43716
rect 37921 43707 37979 43713
rect 37921 43704 37933 43707
rect 37700 43676 37933 43704
rect 37700 43664 37706 43676
rect 37921 43673 37933 43676
rect 37967 43673 37979 43707
rect 37921 43667 37979 43673
rect 32674 43636 32680 43648
rect 31864 43608 32680 43636
rect 32674 43596 32680 43608
rect 32732 43596 32738 43648
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 22465 43435 22523 43441
rect 22465 43401 22477 43435
rect 22511 43432 22523 43435
rect 22646 43432 22652 43444
rect 22511 43404 22652 43432
rect 22511 43401 22523 43404
rect 22465 43395 22523 43401
rect 22646 43392 22652 43404
rect 22704 43392 22710 43444
rect 23566 43432 23572 43444
rect 23527 43404 23572 43432
rect 23566 43392 23572 43404
rect 23624 43392 23630 43444
rect 26418 43432 26424 43444
rect 25792 43404 26424 43432
rect 24949 43367 25007 43373
rect 24949 43333 24961 43367
rect 24995 43364 25007 43367
rect 25038 43364 25044 43376
rect 24995 43336 25044 43364
rect 24995 43333 25007 43336
rect 24949 43327 25007 43333
rect 25038 43324 25044 43336
rect 25096 43324 25102 43376
rect 25133 43367 25191 43373
rect 25133 43333 25145 43367
rect 25179 43364 25191 43367
rect 25682 43364 25688 43376
rect 25179 43336 25688 43364
rect 25179 43333 25191 43336
rect 25133 43327 25191 43333
rect 25682 43324 25688 43336
rect 25740 43324 25746 43376
rect 25792 43373 25820 43404
rect 26418 43392 26424 43404
rect 26476 43392 26482 43444
rect 27614 43432 27620 43444
rect 27575 43404 27620 43432
rect 27614 43392 27620 43404
rect 27672 43392 27678 43444
rect 33226 43432 33232 43444
rect 33187 43404 33232 43432
rect 33226 43392 33232 43404
rect 33284 43392 33290 43444
rect 35161 43435 35219 43441
rect 35161 43401 35173 43435
rect 35207 43432 35219 43435
rect 35434 43432 35440 43444
rect 35207 43404 35440 43432
rect 35207 43401 35219 43404
rect 35161 43395 35219 43401
rect 35434 43392 35440 43404
rect 35492 43392 35498 43444
rect 35710 43432 35716 43444
rect 35671 43404 35716 43432
rect 35710 43392 35716 43404
rect 35768 43392 35774 43444
rect 36814 43432 36820 43444
rect 36775 43404 36820 43432
rect 36814 43392 36820 43404
rect 36872 43392 36878 43444
rect 37553 43435 37611 43441
rect 37553 43401 37565 43435
rect 37599 43432 37611 43435
rect 37734 43432 37740 43444
rect 37599 43404 37740 43432
rect 37599 43401 37611 43404
rect 37553 43395 37611 43401
rect 37734 43392 37740 43404
rect 37792 43392 37798 43444
rect 38105 43435 38163 43441
rect 38105 43401 38117 43435
rect 38151 43432 38163 43435
rect 38470 43432 38476 43444
rect 38151 43404 38476 43432
rect 38151 43401 38163 43404
rect 38105 43395 38163 43401
rect 38470 43392 38476 43404
rect 38528 43392 38534 43444
rect 38838 43392 38844 43444
rect 38896 43432 38902 43444
rect 39117 43435 39175 43441
rect 39117 43432 39129 43435
rect 38896 43404 39129 43432
rect 38896 43392 38902 43404
rect 39117 43401 39129 43404
rect 39163 43401 39175 43435
rect 39117 43395 39175 43401
rect 25777 43367 25835 43373
rect 25777 43333 25789 43367
rect 25823 43333 25835 43367
rect 25777 43327 25835 43333
rect 23661 43299 23719 43305
rect 23661 43265 23673 43299
rect 23707 43296 23719 43299
rect 24121 43299 24179 43305
rect 24121 43296 24133 43299
rect 23707 43268 24133 43296
rect 23707 43265 23719 43268
rect 23661 43259 23719 43265
rect 24121 43265 24133 43268
rect 24167 43265 24179 43299
rect 24121 43259 24179 43265
rect 24305 43299 24363 43305
rect 24305 43265 24317 43299
rect 24351 43265 24363 43299
rect 24305 43259 24363 43265
rect 24489 43299 24547 43305
rect 24489 43265 24501 43299
rect 24535 43296 24547 43299
rect 24854 43296 24860 43308
rect 24535 43268 24860 43296
rect 24535 43265 24547 43268
rect 24489 43259 24547 43265
rect 23017 43231 23075 43237
rect 23017 43197 23029 43231
rect 23063 43228 23075 43231
rect 23106 43228 23112 43240
rect 23063 43200 23112 43228
rect 23063 43197 23075 43200
rect 23017 43191 23075 43197
rect 23106 43188 23112 43200
rect 23164 43228 23170 43240
rect 24320 43228 24348 43259
rect 24854 43256 24860 43268
rect 24912 43256 24918 43308
rect 25317 43299 25375 43305
rect 25317 43265 25329 43299
rect 25363 43296 25375 43299
rect 25590 43296 25596 43308
rect 25363 43268 25596 43296
rect 25363 43265 25375 43268
rect 25317 43259 25375 43265
rect 25590 43256 25596 43268
rect 25648 43256 25654 43308
rect 25792 43228 25820 43327
rect 26050 43324 26056 43376
rect 26108 43364 26114 43376
rect 26145 43367 26203 43373
rect 26145 43364 26157 43367
rect 26108 43336 26157 43364
rect 26108 43324 26114 43336
rect 26145 43333 26157 43336
rect 26191 43333 26203 43367
rect 29270 43364 29276 43376
rect 29231 43336 29276 43364
rect 26145 43327 26203 43333
rect 29270 43324 29276 43336
rect 29328 43324 29334 43376
rect 32122 43324 32128 43376
rect 32180 43364 32186 43376
rect 32309 43367 32367 43373
rect 32309 43364 32321 43367
rect 32180 43336 32321 43364
rect 32180 43324 32186 43336
rect 32309 43333 32321 43336
rect 32355 43333 32367 43367
rect 32674 43364 32680 43376
rect 32635 43336 32680 43364
rect 32309 43327 32367 43333
rect 32674 43324 32680 43336
rect 32732 43324 32738 43376
rect 33502 43364 33508 43376
rect 32968 43336 33508 43364
rect 25961 43299 26019 43305
rect 25961 43265 25973 43299
rect 26007 43296 26019 43299
rect 26878 43296 26884 43308
rect 26007 43268 26884 43296
rect 26007 43265 26019 43268
rect 25961 43259 26019 43265
rect 26878 43256 26884 43268
rect 26936 43256 26942 43308
rect 27157 43299 27215 43305
rect 27157 43265 27169 43299
rect 27203 43296 27215 43299
rect 27246 43296 27252 43308
rect 27203 43268 27252 43296
rect 27203 43265 27215 43268
rect 27157 43259 27215 43265
rect 27246 43256 27252 43268
rect 27304 43256 27310 43308
rect 31202 43296 31208 43308
rect 31163 43268 31208 43296
rect 31202 43256 31208 43268
rect 31260 43256 31266 43308
rect 31662 43256 31668 43308
rect 31720 43296 31726 43308
rect 31757 43299 31815 43305
rect 31757 43296 31769 43299
rect 31720 43268 31769 43296
rect 31720 43256 31726 43268
rect 31757 43265 31769 43268
rect 31803 43296 31815 43299
rect 32493 43299 32551 43305
rect 32493 43296 32505 43299
rect 31803 43268 32505 43296
rect 31803 43265 31815 43268
rect 31757 43259 31815 43265
rect 32493 43265 32505 43268
rect 32539 43296 32551 43299
rect 32858 43296 32864 43308
rect 32539 43268 32864 43296
rect 32539 43265 32551 43268
rect 32493 43259 32551 43265
rect 32858 43256 32864 43268
rect 32916 43296 32922 43308
rect 32968 43296 32996 43336
rect 33502 43324 33508 43336
rect 33560 43324 33566 43376
rect 35526 43324 35532 43376
rect 35584 43364 35590 43376
rect 36173 43367 36231 43373
rect 36173 43364 36185 43367
rect 35584 43336 36185 43364
rect 35584 43324 35590 43336
rect 36173 43333 36185 43336
rect 36219 43333 36231 43367
rect 36173 43327 36231 43333
rect 38194 43324 38200 43376
rect 38252 43364 38258 43376
rect 38657 43367 38715 43373
rect 38657 43364 38669 43367
rect 38252 43336 38669 43364
rect 38252 43324 38258 43336
rect 38657 43333 38669 43336
rect 38703 43333 38715 43367
rect 38657 43327 38715 43333
rect 32916 43268 32996 43296
rect 32916 43256 32922 43268
rect 33042 43256 33048 43308
rect 33100 43296 33106 43308
rect 33137 43299 33195 43305
rect 33137 43296 33149 43299
rect 33100 43268 33149 43296
rect 33100 43256 33106 43268
rect 33137 43265 33149 43268
rect 33183 43265 33195 43299
rect 33137 43259 33195 43265
rect 33410 43256 33416 43308
rect 33468 43296 33474 43308
rect 33781 43299 33839 43305
rect 33781 43296 33793 43299
rect 33468 43268 33793 43296
rect 33468 43256 33474 43268
rect 33781 43265 33793 43268
rect 33827 43265 33839 43299
rect 33781 43259 33839 43265
rect 33870 43256 33876 43308
rect 33928 43296 33934 43308
rect 34425 43299 34483 43305
rect 34425 43296 34437 43299
rect 33928 43268 34437 43296
rect 33928 43256 33934 43268
rect 34425 43265 34437 43268
rect 34471 43265 34483 43299
rect 34425 43259 34483 43265
rect 36909 43299 36967 43305
rect 36909 43265 36921 43299
rect 36955 43296 36967 43299
rect 37550 43296 37556 43308
rect 36955 43268 37556 43296
rect 36955 43265 36967 43268
rect 36909 43259 36967 43265
rect 37550 43256 37556 43268
rect 37608 43256 37614 43308
rect 23164 43200 25820 43228
rect 28629 43231 28687 43237
rect 23164 43188 23170 43200
rect 28629 43197 28641 43231
rect 28675 43228 28687 43231
rect 29181 43231 29239 43237
rect 29181 43228 29193 43231
rect 28675 43200 29193 43228
rect 28675 43197 28687 43200
rect 28629 43191 28687 43197
rect 29181 43197 29193 43200
rect 29227 43197 29239 43231
rect 29181 43191 29239 43197
rect 29730 43160 29736 43172
rect 29691 43132 29736 43160
rect 29730 43120 29736 43132
rect 29788 43120 29794 43172
rect 27430 43092 27436 43104
rect 27391 43064 27436 43092
rect 27430 43052 27436 43064
rect 27488 43052 27494 43104
rect 30282 43052 30288 43104
rect 30340 43092 30346 43104
rect 30377 43095 30435 43101
rect 30377 43092 30389 43095
rect 30340 43064 30389 43092
rect 30340 43052 30346 43064
rect 30377 43061 30389 43064
rect 30423 43092 30435 43095
rect 30926 43092 30932 43104
rect 30423 43064 30932 43092
rect 30423 43061 30435 43064
rect 30377 43055 30435 43061
rect 30926 43052 30932 43064
rect 30984 43052 30990 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 24673 42891 24731 42897
rect 24673 42857 24685 42891
rect 24719 42888 24731 42891
rect 25777 42891 25835 42897
rect 25777 42888 25789 42891
rect 24719 42860 25789 42888
rect 24719 42857 24731 42860
rect 24673 42851 24731 42857
rect 25777 42857 25789 42860
rect 25823 42888 25835 42891
rect 26237 42891 26295 42897
rect 26237 42888 26249 42891
rect 25823 42860 26249 42888
rect 25823 42857 25835 42860
rect 25777 42851 25835 42857
rect 26237 42857 26249 42860
rect 26283 42888 26295 42891
rect 26418 42888 26424 42900
rect 26283 42860 26424 42888
rect 26283 42857 26295 42860
rect 26237 42851 26295 42857
rect 26418 42848 26424 42860
rect 26476 42848 26482 42900
rect 29178 42848 29184 42900
rect 29236 42888 29242 42900
rect 29733 42891 29791 42897
rect 29733 42888 29745 42891
rect 29236 42860 29745 42888
rect 29236 42848 29242 42860
rect 29733 42857 29745 42860
rect 29779 42857 29791 42891
rect 32858 42888 32864 42900
rect 32819 42860 32864 42888
rect 29733 42851 29791 42857
rect 32858 42848 32864 42860
rect 32916 42848 32922 42900
rect 33413 42891 33471 42897
rect 33413 42857 33425 42891
rect 33459 42888 33471 42891
rect 33965 42891 34023 42897
rect 33965 42888 33977 42891
rect 33459 42860 33977 42888
rect 33459 42857 33471 42860
rect 33413 42851 33471 42857
rect 33965 42857 33977 42860
rect 34011 42888 34023 42891
rect 35434 42888 35440 42900
rect 34011 42860 35440 42888
rect 34011 42857 34023 42860
rect 33965 42851 34023 42857
rect 35434 42848 35440 42860
rect 35492 42848 35498 42900
rect 22646 42780 22652 42832
rect 22704 42820 22710 42832
rect 25133 42823 25191 42829
rect 25133 42820 25145 42823
rect 22704 42792 25145 42820
rect 22704 42780 22710 42792
rect 25133 42789 25145 42792
rect 25179 42789 25191 42823
rect 25133 42783 25191 42789
rect 34977 42823 35035 42829
rect 34977 42789 34989 42823
rect 35023 42820 35035 42823
rect 35526 42820 35532 42832
rect 35023 42792 35532 42820
rect 35023 42789 35035 42792
rect 34977 42783 35035 42789
rect 35526 42780 35532 42792
rect 35584 42820 35590 42832
rect 35986 42820 35992 42832
rect 35584 42792 35992 42820
rect 35584 42780 35590 42792
rect 35986 42780 35992 42792
rect 36044 42780 36050 42832
rect 24029 42755 24087 42761
rect 24029 42721 24041 42755
rect 24075 42752 24087 42755
rect 26326 42752 26332 42764
rect 24075 42724 26332 42752
rect 24075 42721 24087 42724
rect 24029 42715 24087 42721
rect 26326 42712 26332 42724
rect 26384 42712 26390 42764
rect 27249 42755 27307 42761
rect 27249 42721 27261 42755
rect 27295 42752 27307 42755
rect 27338 42752 27344 42764
rect 27295 42724 27344 42752
rect 27295 42721 27307 42724
rect 27249 42715 27307 42721
rect 27338 42712 27344 42724
rect 27396 42712 27402 42764
rect 27522 42712 27528 42764
rect 27580 42752 27586 42764
rect 27709 42755 27767 42761
rect 27709 42752 27721 42755
rect 27580 42724 27721 42752
rect 27580 42712 27586 42724
rect 27709 42721 27721 42724
rect 27755 42752 27767 42755
rect 28445 42755 28503 42761
rect 28445 42752 28457 42755
rect 27755 42724 28457 42752
rect 27755 42721 27767 42724
rect 27709 42715 27767 42721
rect 28445 42721 28457 42724
rect 28491 42721 28503 42755
rect 28445 42715 28503 42721
rect 30377 42755 30435 42761
rect 30377 42721 30389 42755
rect 30423 42752 30435 42755
rect 30742 42752 30748 42764
rect 30423 42724 30748 42752
rect 30423 42721 30435 42724
rect 30377 42715 30435 42721
rect 30742 42712 30748 42724
rect 30800 42712 30806 42764
rect 36633 42755 36691 42761
rect 36633 42721 36645 42755
rect 36679 42752 36691 42755
rect 37274 42752 37280 42764
rect 36679 42724 37280 42752
rect 36679 42721 36691 42724
rect 36633 42715 36691 42721
rect 37274 42712 37280 42724
rect 37332 42752 37338 42764
rect 38194 42752 38200 42764
rect 37332 42724 38200 42752
rect 37332 42712 37338 42724
rect 38194 42712 38200 42724
rect 38252 42712 38258 42764
rect 31941 42687 31999 42693
rect 31941 42684 31953 42687
rect 29012 42656 31953 42684
rect 22186 42508 22192 42560
rect 22244 42548 22250 42560
rect 22925 42551 22983 42557
rect 22925 42548 22937 42551
rect 22244 42520 22937 42548
rect 22244 42508 22250 42520
rect 22925 42517 22937 42520
rect 22971 42517 22983 42551
rect 22925 42511 22983 42517
rect 27246 42508 27252 42560
rect 27304 42548 27310 42560
rect 29012 42557 29040 42656
rect 31941 42653 31953 42656
rect 31987 42653 31999 42687
rect 31941 42647 31999 42653
rect 30926 42616 30932 42628
rect 30887 42588 30932 42616
rect 30926 42576 30932 42588
rect 30984 42576 30990 42628
rect 31754 42616 31760 42628
rect 31496 42588 31760 42616
rect 28997 42551 29055 42557
rect 28997 42548 29009 42551
rect 27304 42520 29009 42548
rect 27304 42508 27310 42520
rect 28997 42517 29009 42520
rect 29043 42517 29055 42551
rect 28997 42511 29055 42517
rect 29270 42508 29276 42560
rect 29328 42548 29334 42560
rect 31496 42557 31524 42588
rect 31754 42576 31760 42588
rect 31812 42576 31818 42628
rect 31481 42551 31539 42557
rect 31481 42548 31493 42551
rect 29328 42520 31493 42548
rect 29328 42508 29334 42520
rect 31481 42517 31493 42520
rect 31527 42517 31539 42551
rect 31481 42511 31539 42517
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 25225 42347 25283 42353
rect 25225 42313 25237 42347
rect 25271 42344 25283 42347
rect 26326 42344 26332 42356
rect 25271 42316 26332 42344
rect 25271 42313 25283 42316
rect 25225 42307 25283 42313
rect 26326 42304 26332 42316
rect 26384 42304 26390 42356
rect 27246 42344 27252 42356
rect 27207 42316 27252 42344
rect 27246 42304 27252 42316
rect 27304 42304 27310 42356
rect 27522 42304 27528 42356
rect 27580 42344 27586 42356
rect 27709 42347 27767 42353
rect 27709 42344 27721 42347
rect 27580 42316 27721 42344
rect 27580 42304 27586 42316
rect 27709 42313 27721 42316
rect 27755 42313 27767 42347
rect 27709 42307 27767 42313
rect 29917 42347 29975 42353
rect 29917 42313 29929 42347
rect 29963 42344 29975 42347
rect 30926 42344 30932 42356
rect 29963 42316 30932 42344
rect 29963 42313 29975 42316
rect 29917 42307 29975 42313
rect 30926 42304 30932 42316
rect 30984 42344 30990 42356
rect 32309 42347 32367 42353
rect 32309 42344 32321 42347
rect 30984 42316 32321 42344
rect 30984 42304 30990 42316
rect 32309 42313 32321 42316
rect 32355 42313 32367 42347
rect 32309 42307 32367 42313
rect 34241 42347 34299 42353
rect 34241 42313 34253 42347
rect 34287 42344 34299 42347
rect 35710 42344 35716 42356
rect 34287 42316 35716 42344
rect 34287 42313 34299 42316
rect 34241 42307 34299 42313
rect 35710 42304 35716 42316
rect 35768 42304 35774 42356
rect 35986 42344 35992 42356
rect 35947 42316 35992 42344
rect 35986 42304 35992 42316
rect 36044 42304 36050 42356
rect 25777 42279 25835 42285
rect 25777 42245 25789 42279
rect 25823 42276 25835 42279
rect 25866 42276 25872 42288
rect 25823 42248 25872 42276
rect 25823 42245 25835 42248
rect 25777 42239 25835 42245
rect 25866 42236 25872 42248
rect 25924 42276 25930 42288
rect 28261 42279 28319 42285
rect 28261 42276 28273 42279
rect 25924 42248 28273 42276
rect 25924 42236 25930 42248
rect 28261 42245 28273 42248
rect 28307 42276 28319 42279
rect 29638 42276 29644 42288
rect 28307 42248 29644 42276
rect 28307 42245 28319 42248
rect 28261 42239 28319 42245
rect 29638 42236 29644 42248
rect 29696 42236 29702 42288
rect 30742 42276 30748 42288
rect 30703 42248 30748 42276
rect 30742 42236 30748 42248
rect 30800 42236 30806 42288
rect 35529 42279 35587 42285
rect 35529 42245 35541 42279
rect 35575 42276 35587 42279
rect 37274 42276 37280 42288
rect 35575 42248 37280 42276
rect 35575 42245 35587 42248
rect 35529 42239 35587 42245
rect 37274 42236 37280 42248
rect 37332 42236 37338 42288
rect 29270 42004 29276 42016
rect 29231 41976 29276 42004
rect 29270 41964 29276 41976
rect 29328 41964 29334 42016
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 25317 41803 25375 41809
rect 25317 41769 25329 41803
rect 25363 41800 25375 41803
rect 29270 41800 29276 41812
rect 25363 41772 29276 41800
rect 25363 41769 25375 41772
rect 25317 41763 25375 41769
rect 29270 41760 29276 41772
rect 29328 41760 29334 41812
rect 29638 41760 29644 41812
rect 29696 41800 29702 41812
rect 29733 41803 29791 41809
rect 29733 41800 29745 41803
rect 29696 41772 29745 41800
rect 29696 41760 29702 41772
rect 29733 41769 29745 41772
rect 29779 41769 29791 41803
rect 29733 41763 29791 41769
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 22925 6783 22983 6789
rect 22925 6749 22937 6783
rect 22971 6780 22983 6783
rect 23014 6780 23020 6792
rect 22971 6752 23020 6780
rect 22971 6749 22983 6752
rect 22925 6743 22983 6749
rect 23014 6740 23020 6752
rect 23072 6740 23078 6792
rect 24394 6740 24400 6792
rect 24452 6780 24458 6792
rect 24581 6783 24639 6789
rect 24581 6780 24593 6783
rect 24452 6752 24593 6780
rect 24452 6740 24458 6752
rect 24581 6749 24593 6752
rect 24627 6749 24639 6783
rect 24581 6743 24639 6749
rect 21913 6647 21971 6653
rect 21913 6613 21925 6647
rect 21959 6644 21971 6647
rect 22186 6644 22192 6656
rect 21959 6616 22192 6644
rect 21959 6613 21971 6616
rect 21913 6607 21971 6613
rect 22186 6604 22192 6616
rect 22244 6644 22250 6656
rect 22373 6647 22431 6653
rect 22373 6644 22385 6647
rect 22244 6616 22385 6644
rect 22244 6604 22250 6616
rect 22373 6613 22385 6616
rect 22419 6613 22431 6647
rect 22373 6607 22431 6613
rect 24673 6647 24731 6653
rect 24673 6613 24685 6647
rect 24719 6644 24731 6647
rect 24762 6644 24768 6656
rect 24719 6616 24768 6644
rect 24719 6613 24731 6616
rect 24673 6607 24731 6613
rect 24762 6604 24768 6616
rect 24820 6604 24826 6656
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 24486 6332 24492 6384
rect 24544 6372 24550 6384
rect 24765 6375 24823 6381
rect 24765 6372 24777 6375
rect 24544 6344 24777 6372
rect 24544 6332 24550 6344
rect 24765 6341 24777 6344
rect 24811 6341 24823 6375
rect 24765 6335 24823 6341
rect 26053 6375 26111 6381
rect 26053 6341 26065 6375
rect 26099 6372 26111 6375
rect 26694 6372 26700 6384
rect 26099 6344 26700 6372
rect 26099 6341 26111 6344
rect 26053 6335 26111 6341
rect 26694 6332 26700 6344
rect 26752 6332 26758 6384
rect 22186 6304 22192 6316
rect 22147 6276 22192 6304
rect 22186 6264 22192 6276
rect 22244 6264 22250 6316
rect 22278 6264 22284 6316
rect 22336 6304 22342 6316
rect 22649 6307 22707 6313
rect 22649 6304 22661 6307
rect 22336 6276 22661 6304
rect 22336 6264 22342 6276
rect 22649 6273 22661 6276
rect 22695 6273 22707 6307
rect 28166 6304 28172 6316
rect 28127 6276 28172 6304
rect 22649 6267 22707 6273
rect 28166 6264 28172 6276
rect 28224 6264 28230 6316
rect 24121 6239 24179 6245
rect 24121 6205 24133 6239
rect 24167 6236 24179 6239
rect 24673 6239 24731 6245
rect 24673 6236 24685 6239
rect 24167 6208 24685 6236
rect 24167 6205 24179 6208
rect 24121 6199 24179 6205
rect 24673 6205 24685 6208
rect 24719 6205 24731 6239
rect 25958 6236 25964 6248
rect 25919 6208 25964 6236
rect 24673 6199 24731 6205
rect 25958 6196 25964 6208
rect 26016 6196 26022 6248
rect 25222 6168 25228 6180
rect 25183 6140 25228 6168
rect 25222 6128 25228 6140
rect 25280 6128 25286 6180
rect 26510 6168 26516 6180
rect 26471 6140 26516 6168
rect 26510 6128 26516 6140
rect 26568 6128 26574 6180
rect 20809 6103 20867 6109
rect 20809 6069 20821 6103
rect 20855 6100 20867 6103
rect 20898 6100 20904 6112
rect 20855 6072 20904 6100
rect 20855 6069 20867 6072
rect 20809 6063 20867 6069
rect 20898 6060 20904 6072
rect 20956 6060 20962 6112
rect 21269 6103 21327 6109
rect 21269 6069 21281 6103
rect 21315 6100 21327 6103
rect 21358 6100 21364 6112
rect 21315 6072 21364 6100
rect 21315 6069 21327 6072
rect 21269 6063 21327 6069
rect 21358 6060 21364 6072
rect 21416 6060 21422 6112
rect 22002 6100 22008 6112
rect 21963 6072 22008 6100
rect 22002 6060 22008 6072
rect 22060 6060 22066 6112
rect 22741 6103 22799 6109
rect 22741 6069 22753 6103
rect 22787 6100 22799 6103
rect 23382 6100 23388 6112
rect 22787 6072 23388 6100
rect 22787 6069 22799 6072
rect 22741 6063 22799 6069
rect 23382 6060 23388 6072
rect 23440 6060 23446 6112
rect 23477 6103 23535 6109
rect 23477 6069 23489 6103
rect 23523 6100 23535 6103
rect 24670 6100 24676 6112
rect 23523 6072 24676 6100
rect 23523 6069 23535 6072
rect 23477 6063 23535 6069
rect 24670 6060 24676 6072
rect 24728 6060 24734 6112
rect 27341 6103 27399 6109
rect 27341 6069 27353 6103
rect 27387 6100 27399 6103
rect 27430 6100 27436 6112
rect 27387 6072 27436 6100
rect 27387 6069 27399 6072
rect 27341 6063 27399 6069
rect 27430 6060 27436 6072
rect 27488 6060 27494 6112
rect 27798 6060 27804 6112
rect 27856 6100 27862 6112
rect 28077 6103 28135 6109
rect 28077 6100 28089 6103
rect 27856 6072 28089 6100
rect 27856 6060 27862 6072
rect 28077 6069 28089 6072
rect 28123 6069 28135 6103
rect 28077 6063 28135 6069
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 25958 5896 25964 5908
rect 25919 5868 25964 5896
rect 25958 5856 25964 5868
rect 26016 5856 26022 5908
rect 26694 5896 26700 5908
rect 26655 5868 26700 5896
rect 26694 5856 26700 5868
rect 26752 5856 26758 5908
rect 21910 5828 21916 5840
rect 21871 5800 21916 5828
rect 21910 5788 21916 5800
rect 21968 5788 21974 5840
rect 23842 5828 23848 5840
rect 23803 5800 23848 5828
rect 23842 5788 23848 5800
rect 23900 5788 23906 5840
rect 27982 5828 27988 5840
rect 27943 5800 27988 5828
rect 27982 5788 27988 5800
rect 28040 5788 28046 5840
rect 21358 5760 21364 5772
rect 21319 5732 21364 5760
rect 21358 5720 21364 5732
rect 21416 5720 21422 5772
rect 22741 5763 22799 5769
rect 22741 5729 22753 5763
rect 22787 5760 22799 5763
rect 23293 5763 23351 5769
rect 23293 5760 23305 5763
rect 22787 5732 23305 5760
rect 22787 5729 22799 5732
rect 22741 5723 22799 5729
rect 23293 5729 23305 5732
rect 23339 5729 23351 5763
rect 24670 5760 24676 5772
rect 24631 5732 24676 5760
rect 23293 5723 23351 5729
rect 24670 5720 24676 5732
rect 24728 5720 24734 5772
rect 24946 5760 24952 5772
rect 24907 5732 24952 5760
rect 24946 5720 24952 5732
rect 25004 5720 25010 5772
rect 27430 5760 27436 5772
rect 27391 5732 27436 5760
rect 27430 5720 27436 5732
rect 27488 5720 27494 5772
rect 20622 5692 20628 5704
rect 20583 5664 20628 5692
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 25682 5652 25688 5704
rect 25740 5692 25746 5704
rect 26605 5695 26663 5701
rect 26605 5692 26617 5695
rect 25740 5664 26617 5692
rect 25740 5652 25746 5664
rect 26605 5661 26617 5664
rect 26651 5661 26663 5695
rect 26605 5655 26663 5661
rect 20717 5627 20775 5633
rect 20717 5593 20729 5627
rect 20763 5624 20775 5627
rect 21453 5627 21511 5633
rect 21453 5624 21465 5627
rect 20763 5596 21465 5624
rect 20763 5593 20775 5596
rect 20717 5587 20775 5593
rect 21453 5593 21465 5596
rect 21499 5593 21511 5627
rect 23382 5624 23388 5636
rect 23343 5596 23388 5624
rect 21453 5587 21511 5593
rect 23382 5584 23388 5596
rect 23440 5584 23446 5636
rect 24762 5624 24768 5636
rect 24723 5596 24768 5624
rect 24762 5584 24768 5596
rect 24820 5584 24826 5636
rect 27522 5584 27528 5636
rect 27580 5624 27586 5636
rect 27580 5596 27625 5624
rect 27580 5584 27586 5596
rect 20165 5559 20223 5565
rect 20165 5525 20177 5559
rect 20211 5556 20223 5559
rect 20806 5556 20812 5568
rect 20211 5528 20812 5556
rect 20211 5525 20223 5528
rect 20165 5519 20223 5525
rect 20806 5516 20812 5528
rect 20864 5516 20870 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 21361 5355 21419 5361
rect 21361 5321 21373 5355
rect 21407 5352 21419 5355
rect 24486 5352 24492 5364
rect 21407 5324 23152 5352
rect 24447 5324 24492 5352
rect 21407 5321 21419 5324
rect 21361 5315 21419 5321
rect 22186 5284 22192 5296
rect 20824 5256 22192 5284
rect 20824 5228 20852 5256
rect 22186 5244 22192 5256
rect 22244 5284 22250 5296
rect 23014 5284 23020 5296
rect 22244 5256 22508 5284
rect 22975 5256 23020 5284
rect 22244 5244 22250 5256
rect 19334 5176 19340 5228
rect 19392 5216 19398 5228
rect 19981 5219 20039 5225
rect 19981 5216 19993 5219
rect 19392 5188 19993 5216
rect 19392 5176 19398 5188
rect 19981 5185 19993 5188
rect 20027 5185 20039 5219
rect 20806 5216 20812 5228
rect 20767 5188 20812 5216
rect 19981 5179 20039 5185
rect 19996 5080 20024 5179
rect 20806 5176 20812 5188
rect 20864 5176 20870 5228
rect 21269 5219 21327 5225
rect 21269 5185 21281 5219
rect 21315 5216 21327 5219
rect 22278 5216 22284 5228
rect 21315 5188 22284 5216
rect 21315 5185 21327 5188
rect 21269 5179 21327 5185
rect 20346 5108 20352 5160
rect 20404 5148 20410 5160
rect 21284 5148 21312 5179
rect 22278 5176 22284 5188
rect 22336 5176 22342 5228
rect 22480 5225 22508 5256
rect 23014 5244 23020 5256
rect 23072 5244 23078 5296
rect 23124 5293 23152 5324
rect 24486 5312 24492 5324
rect 24544 5312 24550 5364
rect 23109 5287 23167 5293
rect 23109 5253 23121 5287
rect 23155 5253 23167 5287
rect 23109 5247 23167 5253
rect 25774 5244 25780 5296
rect 25832 5284 25838 5296
rect 25869 5287 25927 5293
rect 25869 5284 25881 5287
rect 25832 5256 25881 5284
rect 25832 5244 25838 5256
rect 25869 5253 25881 5256
rect 25915 5253 25927 5287
rect 27798 5284 27804 5296
rect 27759 5256 27804 5284
rect 25869 5247 25927 5253
rect 27798 5244 27804 5256
rect 27856 5244 27862 5296
rect 22465 5219 22523 5225
rect 22465 5185 22477 5219
rect 22511 5185 22523 5219
rect 22465 5179 22523 5185
rect 23750 5176 23756 5228
rect 23808 5216 23814 5228
rect 24394 5216 24400 5228
rect 23808 5188 24400 5216
rect 23808 5176 23814 5188
rect 24394 5176 24400 5188
rect 24452 5176 24458 5228
rect 20404 5120 21312 5148
rect 25225 5151 25283 5157
rect 20404 5108 20410 5120
rect 25225 5117 25237 5151
rect 25271 5148 25283 5151
rect 25777 5151 25835 5157
rect 25777 5148 25789 5151
rect 25271 5120 25789 5148
rect 25271 5117 25283 5120
rect 25225 5111 25283 5117
rect 25777 5117 25789 5120
rect 25823 5117 25835 5151
rect 27614 5148 27620 5160
rect 27575 5120 27620 5148
rect 25777 5111 25835 5117
rect 27614 5108 27620 5120
rect 27672 5108 27678 5160
rect 27893 5151 27951 5157
rect 27893 5117 27905 5151
rect 27939 5148 27951 5151
rect 28445 5151 28503 5157
rect 28445 5148 28457 5151
rect 27939 5120 28457 5148
rect 27939 5117 27951 5120
rect 27893 5111 27951 5117
rect 28445 5117 28457 5120
rect 28491 5117 28503 5151
rect 28445 5111 28503 5117
rect 20622 5080 20628 5092
rect 19996 5052 20628 5080
rect 20622 5040 20628 5052
rect 20680 5040 20686 5092
rect 22278 5080 22284 5092
rect 22239 5052 22284 5080
rect 22278 5040 22284 5052
rect 22336 5040 22342 5092
rect 23566 5080 23572 5092
rect 23527 5052 23572 5080
rect 23566 5040 23572 5052
rect 23624 5040 23630 5092
rect 26326 5080 26332 5092
rect 26287 5052 26332 5080
rect 26326 5040 26332 5052
rect 26384 5040 26390 5092
rect 19426 5012 19432 5024
rect 19387 4984 19432 5012
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 20070 5012 20076 5024
rect 20031 4984 20076 5012
rect 20070 4972 20076 4984
rect 20128 4972 20134 5024
rect 29086 5012 29092 5024
rect 29047 4984 29092 5012
rect 29086 4972 29092 4984
rect 29144 4972 29150 5024
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 22097 4811 22155 4817
rect 20088 4780 22048 4808
rect 18877 4675 18935 4681
rect 18877 4641 18889 4675
rect 18923 4672 18935 4675
rect 19978 4672 19984 4684
rect 18923 4644 19984 4672
rect 18923 4641 18935 4644
rect 18877 4635 18935 4641
rect 19978 4632 19984 4644
rect 20036 4632 20042 4684
rect 18046 4604 18052 4616
rect 18007 4576 18052 4604
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4604 19763 4607
rect 20088 4604 20116 4780
rect 22020 4752 22048 4780
rect 22097 4777 22109 4811
rect 22143 4808 22155 4811
rect 23750 4808 23756 4820
rect 22143 4780 23756 4808
rect 22143 4777 22155 4780
rect 22097 4771 22155 4777
rect 23750 4768 23756 4780
rect 23808 4768 23814 4820
rect 25774 4808 25780 4820
rect 25735 4780 25780 4808
rect 25774 4768 25780 4780
rect 25832 4768 25838 4820
rect 27522 4808 27528 4820
rect 27483 4780 27528 4808
rect 27522 4768 27528 4780
rect 27580 4768 27586 4820
rect 20714 4700 20720 4752
rect 20772 4740 20778 4752
rect 22002 4740 22008 4752
rect 20772 4712 21036 4740
rect 21915 4712 22008 4740
rect 20772 4700 20778 4712
rect 20898 4672 20904 4684
rect 20859 4644 20904 4672
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 21008 4672 21036 4712
rect 22002 4700 22008 4712
rect 22060 4740 22066 4752
rect 25041 4743 25099 4749
rect 22060 4712 23520 4740
rect 22060 4700 22066 4712
rect 22833 4675 22891 4681
rect 22833 4672 22845 4675
rect 21008 4644 22845 4672
rect 22833 4641 22845 4644
rect 22879 4641 22891 4675
rect 23290 4672 23296 4684
rect 23251 4644 23296 4672
rect 22833 4635 22891 4641
rect 23290 4632 23296 4644
rect 23348 4632 23354 4684
rect 19751 4576 20116 4604
rect 20165 4607 20223 4613
rect 19751 4573 19763 4576
rect 19705 4567 19763 4573
rect 20165 4573 20177 4607
rect 20211 4604 20223 4607
rect 20346 4604 20352 4616
rect 20211 4576 20352 4604
rect 20211 4573 20223 4576
rect 20165 4567 20223 4573
rect 20346 4564 20352 4576
rect 20404 4564 20410 4616
rect 22002 4564 22008 4616
rect 22060 4604 22066 4616
rect 22281 4607 22339 4613
rect 22281 4604 22293 4607
rect 22060 4576 22293 4604
rect 22060 4564 22066 4576
rect 22281 4573 22293 4576
rect 22327 4573 22339 4607
rect 23492 4604 23520 4712
rect 25041 4709 25053 4743
rect 25087 4740 25099 4743
rect 25682 4740 25688 4752
rect 25087 4712 25688 4740
rect 25087 4709 25099 4712
rect 25041 4703 25099 4709
rect 25682 4700 25688 4712
rect 25740 4700 25746 4752
rect 27540 4712 29776 4740
rect 25240 4644 26234 4672
rect 25240 4613 25268 4644
rect 25225 4607 25283 4613
rect 25225 4604 25237 4607
rect 23492 4576 25237 4604
rect 22281 4567 22339 4573
rect 25225 4573 25237 4576
rect 25271 4573 25283 4607
rect 25682 4604 25688 4616
rect 25643 4576 25688 4604
rect 25225 4567 25283 4573
rect 25682 4564 25688 4576
rect 25740 4564 25746 4616
rect 26206 4604 26234 4644
rect 26973 4607 27031 4613
rect 26973 4604 26985 4607
rect 26206 4576 26985 4604
rect 26973 4573 26985 4576
rect 27019 4604 27031 4607
rect 27540 4604 27568 4712
rect 28810 4672 28816 4684
rect 28771 4644 28816 4672
rect 28810 4632 28816 4644
rect 28868 4632 28874 4684
rect 29086 4672 29092 4684
rect 29047 4644 29092 4672
rect 29086 4632 29092 4644
rect 29144 4632 29150 4684
rect 27019 4576 27568 4604
rect 27617 4607 27675 4613
rect 27019 4573 27031 4576
rect 26973 4567 27031 4573
rect 27617 4573 27629 4607
rect 27663 4604 27675 4607
rect 27890 4604 27896 4616
rect 27663 4576 27896 4604
rect 27663 4573 27675 4576
rect 27617 4567 27675 4573
rect 20070 4496 20076 4548
rect 20128 4536 20134 4548
rect 20993 4539 21051 4545
rect 20993 4536 21005 4539
rect 20128 4508 21005 4536
rect 20128 4496 20134 4508
rect 20993 4505 21005 4508
rect 21039 4505 21051 4539
rect 20993 4499 21051 4505
rect 21545 4539 21603 4545
rect 21545 4505 21557 4539
rect 21591 4536 21603 4539
rect 21634 4536 21640 4548
rect 21591 4508 21640 4536
rect 21591 4505 21603 4508
rect 21545 4499 21603 4505
rect 21634 4496 21640 4508
rect 21692 4496 21698 4548
rect 22925 4539 22983 4545
rect 22066 4508 22784 4536
rect 19613 4471 19671 4477
rect 19613 4437 19625 4471
rect 19659 4468 19671 4471
rect 20162 4468 20168 4480
rect 19659 4440 20168 4468
rect 19659 4437 19671 4440
rect 19613 4431 19671 4437
rect 20162 4428 20168 4440
rect 20220 4428 20226 4480
rect 20257 4471 20315 4477
rect 20257 4437 20269 4471
rect 20303 4468 20315 4471
rect 22066 4468 22094 4508
rect 20303 4440 22094 4468
rect 22756 4468 22784 4508
rect 22925 4505 22937 4539
rect 22971 4505 22983 4539
rect 22925 4499 22983 4505
rect 22940 4468 22968 4499
rect 22756 4440 22968 4468
rect 26789 4471 26847 4477
rect 20303 4437 20315 4440
rect 20257 4431 20315 4437
rect 26789 4437 26801 4471
rect 26835 4468 26847 4471
rect 27632 4468 27660 4567
rect 27890 4564 27896 4576
rect 27948 4604 27954 4616
rect 28166 4604 28172 4616
rect 27948 4576 28172 4604
rect 27948 4564 27954 4576
rect 28166 4564 28172 4576
rect 28224 4564 28230 4616
rect 29748 4613 29776 4712
rect 29733 4607 29791 4613
rect 29733 4573 29745 4607
rect 29779 4573 29791 4607
rect 29733 4567 29791 4573
rect 30561 4607 30619 4613
rect 30561 4573 30573 4607
rect 30607 4573 30619 4607
rect 30561 4567 30619 4573
rect 28997 4539 29055 4545
rect 28997 4505 29009 4539
rect 29043 4536 29055 4539
rect 30469 4539 30527 4545
rect 30469 4536 30481 4539
rect 29043 4508 30481 4536
rect 29043 4505 29055 4508
rect 28997 4499 29055 4505
rect 30469 4505 30481 4508
rect 30515 4505 30527 4539
rect 30469 4499 30527 4505
rect 26835 4440 27660 4468
rect 29917 4471 29975 4477
rect 26835 4437 26847 4440
rect 26789 4431 26847 4437
rect 29917 4437 29929 4471
rect 29963 4468 29975 4471
rect 30374 4468 30380 4480
rect 29963 4440 30380 4468
rect 29963 4437 29975 4440
rect 29917 4431 29975 4437
rect 30374 4428 30380 4440
rect 30432 4468 30438 4480
rect 30576 4468 30604 4567
rect 30432 4440 30604 4468
rect 30432 4428 30438 4440
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 20162 4156 20168 4208
rect 20220 4196 20226 4208
rect 20533 4199 20591 4205
rect 20533 4196 20545 4199
rect 20220 4168 20545 4196
rect 20220 4156 20226 4168
rect 20533 4165 20545 4168
rect 20579 4165 20591 4199
rect 20533 4159 20591 4165
rect 20806 4156 20812 4208
rect 20864 4196 20870 4208
rect 22189 4199 22247 4205
rect 22189 4196 22201 4199
rect 20864 4168 22201 4196
rect 20864 4156 20870 4168
rect 22189 4165 22201 4168
rect 22235 4165 22247 4199
rect 24302 4196 24308 4208
rect 24263 4168 24308 4196
rect 22189 4159 22247 4165
rect 24302 4156 24308 4168
rect 24360 4156 24366 4208
rect 25498 4196 25504 4208
rect 25459 4168 25504 4196
rect 25498 4156 25504 4168
rect 25556 4156 25562 4208
rect 27338 4196 27344 4208
rect 27299 4168 27344 4196
rect 27338 4156 27344 4168
rect 27396 4156 27402 4208
rect 29089 4199 29147 4205
rect 29089 4165 29101 4199
rect 29135 4196 29147 4199
rect 29825 4199 29883 4205
rect 29825 4196 29837 4199
rect 29135 4168 29837 4196
rect 29135 4165 29147 4168
rect 29089 4159 29147 4165
rect 29825 4165 29837 4168
rect 29871 4165 29883 4199
rect 29825 4159 29883 4165
rect 29917 4131 29975 4137
rect 29917 4097 29929 4131
rect 29963 4128 29975 4131
rect 30466 4128 30472 4140
rect 29963 4100 30472 4128
rect 29963 4097 29975 4100
rect 29917 4091 29975 4097
rect 30466 4088 30472 4100
rect 30524 4088 30530 4140
rect 18601 4063 18659 4069
rect 18601 4029 18613 4063
rect 18647 4060 18659 4063
rect 20441 4063 20499 4069
rect 20441 4060 20453 4063
rect 18647 4032 20453 4060
rect 18647 4029 18659 4032
rect 18601 4023 18659 4029
rect 20441 4029 20453 4032
rect 20487 4029 20499 4063
rect 21082 4060 21088 4072
rect 21043 4032 21088 4060
rect 20441 4023 20499 4029
rect 21082 4020 21088 4032
rect 21140 4020 21146 4072
rect 22097 4063 22155 4069
rect 22097 4029 22109 4063
rect 22143 4029 22155 4063
rect 22097 4023 22155 4029
rect 19245 3995 19303 4001
rect 19245 3961 19257 3995
rect 19291 3992 19303 3995
rect 22112 3992 22140 4023
rect 22186 4020 22192 4072
rect 22244 4060 22250 4072
rect 22373 4063 22431 4069
rect 22373 4060 22385 4063
rect 22244 4032 22385 4060
rect 22244 4020 22250 4032
rect 22373 4029 22385 4032
rect 22419 4029 22431 4063
rect 22373 4023 22431 4029
rect 23382 4020 23388 4072
rect 23440 4060 23446 4072
rect 24213 4063 24271 4069
rect 24213 4060 24225 4063
rect 23440 4032 24225 4060
rect 23440 4020 23446 4032
rect 24213 4029 24225 4032
rect 24259 4029 24271 4063
rect 25409 4063 25467 4069
rect 25409 4060 25421 4063
rect 24213 4023 24271 4029
rect 24504 4032 25421 4060
rect 19291 3964 22140 3992
rect 23661 3995 23719 4001
rect 19291 3961 19303 3964
rect 19245 3955 19303 3961
rect 23661 3961 23673 3995
rect 23707 3992 23719 3995
rect 24504 3992 24532 4032
rect 25409 4029 25421 4032
rect 25455 4029 25467 4063
rect 26050 4060 26056 4072
rect 26011 4032 26056 4060
rect 25409 4023 25467 4029
rect 26050 4020 26056 4032
rect 26108 4020 26114 4072
rect 26602 4020 26608 4072
rect 26660 4060 26666 4072
rect 27249 4063 27307 4069
rect 27249 4060 27261 4063
rect 26660 4032 27261 4060
rect 26660 4020 26666 4032
rect 27249 4029 27261 4032
rect 27295 4029 27307 4063
rect 27249 4023 27307 4029
rect 27430 4020 27436 4072
rect 27488 4060 27494 4072
rect 27525 4063 27583 4069
rect 27525 4060 27537 4063
rect 27488 4032 27537 4060
rect 27488 4020 27494 4032
rect 27525 4029 27537 4032
rect 27571 4029 27583 4063
rect 27525 4023 27583 4029
rect 28905 4063 28963 4069
rect 28905 4029 28917 4063
rect 28951 4060 28963 4063
rect 29086 4060 29092 4072
rect 28951 4032 29092 4060
rect 28951 4029 28963 4032
rect 28905 4023 28963 4029
rect 29086 4020 29092 4032
rect 29144 4020 29150 4072
rect 29181 4063 29239 4069
rect 29181 4029 29193 4063
rect 29227 4060 29239 4063
rect 30377 4063 30435 4069
rect 30377 4060 30389 4063
rect 29227 4032 30389 4060
rect 29227 4029 29239 4032
rect 29181 4023 29239 4029
rect 30377 4029 30389 4032
rect 30423 4029 30435 4063
rect 30377 4023 30435 4029
rect 23707 3964 24532 3992
rect 23707 3961 23719 3964
rect 23661 3955 23719 3961
rect 24670 3952 24676 4004
rect 24728 3992 24734 4004
rect 24765 3995 24823 4001
rect 24765 3992 24777 3995
rect 24728 3964 24777 3992
rect 24728 3952 24734 3964
rect 24765 3961 24777 3964
rect 24811 3961 24823 3995
rect 24765 3955 24823 3961
rect 15010 3924 15016 3936
rect 14971 3896 15016 3924
rect 15010 3884 15016 3896
rect 15068 3884 15074 3936
rect 16114 3924 16120 3936
rect 16075 3896 16120 3924
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 17218 3924 17224 3936
rect 17179 3896 17224 3924
rect 17218 3884 17224 3896
rect 17276 3884 17282 3936
rect 17957 3927 18015 3933
rect 17957 3893 17969 3927
rect 18003 3924 18015 3927
rect 18874 3924 18880 3936
rect 18003 3896 18880 3924
rect 18003 3893 18015 3896
rect 17957 3887 18015 3893
rect 18874 3884 18880 3896
rect 18932 3884 18938 3936
rect 19889 3927 19947 3933
rect 19889 3893 19901 3927
rect 19935 3924 19947 3927
rect 20714 3924 20720 3936
rect 19935 3896 20720 3924
rect 19935 3893 19947 3896
rect 19889 3887 19947 3893
rect 20714 3884 20720 3896
rect 20772 3884 20778 3936
rect 20898 3884 20904 3936
rect 20956 3924 20962 3936
rect 23750 3924 23756 3936
rect 20956 3896 23756 3924
rect 20956 3884 20962 3896
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 18138 3680 18144 3732
rect 18196 3720 18202 3732
rect 21726 3720 21732 3732
rect 18196 3692 21732 3720
rect 18196 3680 18202 3692
rect 21726 3680 21732 3692
rect 21784 3680 21790 3732
rect 23382 3720 23388 3732
rect 23343 3692 23388 3720
rect 23382 3680 23388 3692
rect 23440 3680 23446 3732
rect 23937 3723 23995 3729
rect 23937 3689 23949 3723
rect 23983 3720 23995 3723
rect 24302 3720 24308 3732
rect 23983 3692 24308 3720
rect 23983 3689 23995 3692
rect 23937 3683 23995 3689
rect 24302 3680 24308 3692
rect 24360 3680 24366 3732
rect 25498 3680 25504 3732
rect 25556 3720 25562 3732
rect 25869 3723 25927 3729
rect 25869 3720 25881 3723
rect 25556 3692 25881 3720
rect 25556 3680 25562 3692
rect 25869 3689 25881 3692
rect 25915 3689 25927 3723
rect 25869 3683 25927 3689
rect 16301 3655 16359 3661
rect 16301 3621 16313 3655
rect 16347 3652 16359 3655
rect 16942 3652 16948 3664
rect 16347 3624 16948 3652
rect 16347 3621 16359 3624
rect 16301 3615 16359 3621
rect 16942 3612 16948 3624
rect 17000 3612 17006 3664
rect 20162 3612 20168 3664
rect 20220 3652 20226 3664
rect 30466 3652 30472 3664
rect 20220 3624 23980 3652
rect 20220 3612 20226 3624
rect 15013 3587 15071 3593
rect 15013 3553 15025 3587
rect 15059 3584 15071 3587
rect 15838 3584 15844 3596
rect 15059 3556 15844 3584
rect 15059 3553 15071 3556
rect 15013 3547 15071 3553
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 17589 3587 17647 3593
rect 17589 3553 17601 3587
rect 17635 3584 17647 3587
rect 20254 3584 20260 3596
rect 17635 3556 20260 3584
rect 17635 3553 17647 3556
rect 17589 3547 17647 3553
rect 20254 3544 20260 3556
rect 20312 3544 20318 3596
rect 20349 3587 20407 3593
rect 20349 3553 20361 3587
rect 20395 3584 20407 3587
rect 20395 3556 22600 3584
rect 20395 3553 20407 3556
rect 20349 3547 20407 3553
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 4249 3519 4307 3525
rect 4249 3516 4261 3519
rect 4212 3488 4261 3516
rect 4212 3476 4218 3488
rect 4249 3485 4261 3488
rect 4295 3485 4307 3519
rect 5166 3516 5172 3528
rect 5127 3488 5172 3516
rect 4249 3479 4307 3485
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 5994 3516 6000 3528
rect 5955 3488 6000 3516
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 6822 3516 6828 3528
rect 6783 3488 6828 3516
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 7650 3516 7656 3528
rect 7611 3488 7656 3516
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 8478 3516 8484 3528
rect 8439 3488 8484 3516
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 9306 3516 9312 3528
rect 9267 3488 9312 3516
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 10134 3516 10140 3528
rect 10095 3488 10140 3516
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 10962 3516 10968 3528
rect 10923 3488 10968 3516
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3516 11759 3519
rect 11790 3516 11796 3528
rect 11747 3488 11796 3516
rect 11747 3485 11759 3488
rect 11701 3479 11759 3485
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 12345 3519 12403 3525
rect 12345 3485 12357 3519
rect 12391 3516 12403 3519
rect 12526 3516 12532 3528
rect 12391 3488 12532 3516
rect 12391 3485 12403 3488
rect 12345 3479 12403 3485
rect 12526 3476 12532 3488
rect 12584 3476 12590 3528
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3516 13047 3519
rect 13078 3516 13084 3528
rect 13035 3488 13084 3516
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 13630 3516 13636 3528
rect 13591 3488 13636 3516
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 15657 3519 15715 3525
rect 15657 3485 15669 3519
rect 15703 3516 15715 3519
rect 16390 3516 16396 3528
rect 15703 3488 16396 3516
rect 15703 3485 15715 3488
rect 15657 3479 15715 3485
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 16945 3519 17003 3525
rect 16945 3485 16957 3519
rect 16991 3485 17003 3519
rect 16945 3479 17003 3485
rect 18233 3519 18291 3525
rect 18233 3485 18245 3519
rect 18279 3516 18291 3519
rect 18598 3516 18604 3528
rect 18279 3488 18604 3516
rect 18279 3485 18291 3488
rect 18233 3479 18291 3485
rect 16960 3448 16988 3479
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 18690 3476 18696 3528
rect 18748 3516 18754 3528
rect 19334 3516 19340 3528
rect 18748 3488 19340 3516
rect 18748 3476 18754 3488
rect 19334 3476 19340 3488
rect 19392 3516 19398 3528
rect 19613 3519 19671 3525
rect 19613 3516 19625 3519
rect 19392 3488 19625 3516
rect 19392 3476 19398 3488
rect 19613 3485 19625 3488
rect 19659 3485 19671 3519
rect 19613 3479 19671 3485
rect 20441 3519 20499 3525
rect 20441 3485 20453 3519
rect 20487 3516 20499 3519
rect 20898 3516 20904 3528
rect 20487 3488 20904 3516
rect 20487 3485 20499 3488
rect 20441 3479 20499 3485
rect 20898 3476 20904 3488
rect 20956 3476 20962 3528
rect 18506 3448 18512 3460
rect 16960 3420 18512 3448
rect 18506 3408 18512 3420
rect 18564 3408 18570 3460
rect 20346 3448 20352 3460
rect 19352 3420 20352 3448
rect 19352 3392 19380 3420
rect 20346 3408 20352 3420
rect 20404 3408 20410 3460
rect 20622 3408 20628 3460
rect 20680 3448 20686 3460
rect 21637 3451 21695 3457
rect 21637 3448 21649 3451
rect 20680 3420 21649 3448
rect 20680 3408 20686 3420
rect 21637 3417 21649 3420
rect 21683 3417 21695 3451
rect 21637 3411 21695 3417
rect 21726 3408 21732 3460
rect 21784 3448 21790 3460
rect 22281 3451 22339 3457
rect 21784 3420 21829 3448
rect 21784 3408 21790 3420
rect 22281 3417 22293 3451
rect 22327 3448 22339 3451
rect 22462 3448 22468 3460
rect 22327 3420 22468 3448
rect 22327 3417 22339 3420
rect 22281 3411 22339 3417
rect 22462 3408 22468 3420
rect 22520 3408 22526 3460
rect 22572 3448 22600 3556
rect 23750 3476 23756 3528
rect 23808 3516 23814 3528
rect 23845 3519 23903 3525
rect 23845 3516 23857 3519
rect 23808 3488 23857 3516
rect 23808 3476 23814 3488
rect 23845 3485 23857 3488
rect 23891 3485 23903 3519
rect 23952 3516 23980 3624
rect 29932 3624 30472 3652
rect 24210 3544 24216 3596
rect 24268 3584 24274 3596
rect 24949 3587 25007 3593
rect 24949 3584 24961 3587
rect 24268 3556 24961 3584
rect 24268 3544 24274 3556
rect 24949 3553 24961 3556
rect 24995 3553 25007 3587
rect 24949 3547 25007 3553
rect 27065 3587 27123 3593
rect 27065 3553 27077 3587
rect 27111 3584 27123 3587
rect 27154 3584 27160 3596
rect 27111 3556 27160 3584
rect 27111 3553 27123 3556
rect 27065 3547 27123 3553
rect 27154 3544 27160 3556
rect 27212 3544 27218 3596
rect 28258 3584 28264 3596
rect 28219 3556 28264 3584
rect 28258 3544 28264 3556
rect 28316 3544 28322 3596
rect 23952 3488 24532 3516
rect 23845 3479 23903 3485
rect 24504 3448 24532 3488
rect 25682 3476 25688 3528
rect 25740 3516 25746 3528
rect 29932 3525 29960 3624
rect 30466 3612 30472 3624
rect 30524 3652 30530 3664
rect 31386 3652 31392 3664
rect 30524 3624 31392 3652
rect 30524 3612 30530 3624
rect 31386 3612 31392 3624
rect 31444 3612 31450 3664
rect 32950 3612 32956 3664
rect 33008 3652 33014 3664
rect 33597 3655 33655 3661
rect 33597 3652 33609 3655
rect 33008 3624 33609 3652
rect 33008 3612 33014 3624
rect 33597 3621 33609 3624
rect 33643 3621 33655 3655
rect 33597 3615 33655 3621
rect 36814 3612 36820 3664
rect 36872 3652 36878 3664
rect 37461 3655 37519 3661
rect 37461 3652 37473 3655
rect 36872 3624 37473 3652
rect 36872 3612 36878 3624
rect 37461 3621 37473 3624
rect 37507 3621 37519 3655
rect 37461 3615 37519 3621
rect 30190 3544 30196 3596
rect 30248 3584 30254 3596
rect 31021 3587 31079 3593
rect 31021 3584 31033 3587
rect 30248 3556 31033 3584
rect 30248 3544 30254 3556
rect 31021 3553 31033 3556
rect 31067 3553 31079 3587
rect 31021 3547 31079 3553
rect 34790 3544 34796 3596
rect 34848 3584 34854 3596
rect 35529 3587 35587 3593
rect 35529 3584 35541 3587
rect 34848 3556 35541 3584
rect 34848 3544 34854 3556
rect 35529 3553 35541 3556
rect 35575 3553 35587 3587
rect 35529 3547 35587 3553
rect 25961 3519 26019 3525
rect 25961 3516 25973 3519
rect 25740 3488 25973 3516
rect 25740 3476 25746 3488
rect 25961 3485 25973 3488
rect 26007 3485 26019 3519
rect 25961 3479 26019 3485
rect 29917 3519 29975 3525
rect 29917 3485 29929 3519
rect 29963 3485 29975 3519
rect 29917 3479 29975 3485
rect 30006 3476 30012 3528
rect 30064 3516 30070 3528
rect 30377 3519 30435 3525
rect 30377 3516 30389 3519
rect 30064 3488 30389 3516
rect 30064 3476 30070 3488
rect 30377 3485 30389 3488
rect 30423 3485 30435 3519
rect 30377 3479 30435 3485
rect 31110 3476 31116 3528
rect 31168 3516 31174 3528
rect 31665 3519 31723 3525
rect 31665 3516 31677 3519
rect 31168 3488 31677 3516
rect 31168 3476 31174 3488
rect 31665 3485 31677 3488
rect 31711 3485 31723 3519
rect 31665 3479 31723 3485
rect 31846 3476 31852 3528
rect 31904 3516 31910 3528
rect 32309 3519 32367 3525
rect 32309 3516 32321 3519
rect 31904 3488 32321 3516
rect 31904 3476 31910 3488
rect 32309 3485 32321 3488
rect 32355 3485 32367 3519
rect 32309 3479 32367 3485
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 32953 3519 33011 3525
rect 32953 3516 32965 3519
rect 32456 3488 32965 3516
rect 32456 3476 32462 3488
rect 32953 3485 32965 3488
rect 32999 3485 33011 3519
rect 32953 3479 33011 3485
rect 34330 3476 34336 3528
rect 34388 3516 34394 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34388 3488 34897 3516
rect 34388 3476 34394 3488
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 34885 3479 34943 3485
rect 35710 3476 35716 3528
rect 35768 3516 35774 3528
rect 36173 3519 36231 3525
rect 36173 3516 36185 3519
rect 35768 3488 36185 3516
rect 35768 3476 35774 3488
rect 36173 3485 36185 3488
rect 36219 3485 36231 3519
rect 36173 3479 36231 3485
rect 36262 3476 36268 3528
rect 36320 3516 36326 3528
rect 36817 3519 36875 3525
rect 36817 3516 36829 3519
rect 36320 3488 36829 3516
rect 36320 3476 36326 3488
rect 36817 3485 36829 3488
rect 36863 3485 36875 3519
rect 36817 3479 36875 3485
rect 37642 3476 37648 3528
rect 37700 3516 37706 3528
rect 38105 3519 38163 3525
rect 38105 3516 38117 3519
rect 37700 3488 38117 3516
rect 37700 3476 37706 3488
rect 38105 3485 38117 3488
rect 38151 3485 38163 3519
rect 38105 3479 38163 3485
rect 38194 3476 38200 3528
rect 38252 3516 38258 3528
rect 38749 3519 38807 3525
rect 38749 3516 38761 3519
rect 38252 3488 38761 3516
rect 38252 3476 38258 3488
rect 38749 3485 38761 3488
rect 38795 3485 38807 3519
rect 38749 3479 38807 3485
rect 39574 3476 39580 3528
rect 39632 3516 39638 3528
rect 40037 3519 40095 3525
rect 40037 3516 40049 3519
rect 39632 3488 40049 3516
rect 39632 3476 39638 3488
rect 40037 3485 40049 3488
rect 40083 3485 40095 3519
rect 40037 3479 40095 3485
rect 40402 3476 40408 3528
rect 40460 3516 40466 3528
rect 40681 3519 40739 3525
rect 40681 3516 40693 3519
rect 40460 3488 40693 3516
rect 40460 3476 40466 3488
rect 40681 3485 40693 3488
rect 40727 3485 40739 3519
rect 40681 3479 40739 3485
rect 40954 3476 40960 3528
rect 41012 3516 41018 3528
rect 41325 3519 41383 3525
rect 41325 3516 41337 3519
rect 41012 3488 41337 3516
rect 41012 3476 41018 3488
rect 41325 3485 41337 3488
rect 41371 3485 41383 3519
rect 41325 3479 41383 3485
rect 41506 3476 41512 3528
rect 41564 3516 41570 3528
rect 41969 3519 42027 3525
rect 41969 3516 41981 3519
rect 41564 3488 41981 3516
rect 41564 3476 41570 3488
rect 41969 3485 41981 3488
rect 42015 3485 42027 3519
rect 42886 3516 42892 3528
rect 42847 3488 42892 3516
rect 41969 3479 42027 3485
rect 42886 3476 42892 3488
rect 42944 3476 42950 3528
rect 43162 3476 43168 3528
rect 43220 3516 43226 3528
rect 43349 3519 43407 3525
rect 43349 3516 43361 3519
rect 43220 3488 43361 3516
rect 43220 3476 43226 3488
rect 43349 3485 43361 3488
rect 43395 3485 43407 3519
rect 43349 3479 43407 3485
rect 44818 3476 44824 3528
rect 44876 3516 44882 3528
rect 45189 3519 45247 3525
rect 45189 3516 45201 3519
rect 44876 3488 45201 3516
rect 44876 3476 44882 3488
rect 45189 3485 45201 3488
rect 45235 3485 45247 3519
rect 45189 3479 45247 3485
rect 45646 3476 45652 3528
rect 45704 3516 45710 3528
rect 45833 3519 45891 3525
rect 45833 3516 45845 3519
rect 45704 3488 45845 3516
rect 45704 3476 45710 3488
rect 45833 3485 45845 3488
rect 45879 3485 45891 3519
rect 46474 3516 46480 3528
rect 46435 3488 46480 3516
rect 45833 3479 45891 3485
rect 46474 3476 46480 3488
rect 46532 3476 46538 3528
rect 46750 3476 46756 3528
rect 46808 3516 46814 3528
rect 47121 3519 47179 3525
rect 47121 3516 47133 3519
rect 46808 3488 47133 3516
rect 46808 3476 46814 3488
rect 47121 3485 47133 3488
rect 47167 3485 47179 3519
rect 47121 3479 47179 3485
rect 47302 3476 47308 3528
rect 47360 3516 47366 3528
rect 47765 3519 47823 3525
rect 47765 3516 47777 3519
rect 47360 3488 47777 3516
rect 47360 3476 47366 3488
rect 47765 3485 47777 3488
rect 47811 3485 47823 3519
rect 47765 3479 47823 3485
rect 24673 3451 24731 3457
rect 24673 3448 24685 3451
rect 22572 3420 24440 3448
rect 24504 3420 24685 3448
rect 18782 3380 18788 3392
rect 18743 3352 18788 3380
rect 18782 3340 18788 3352
rect 18840 3340 18846 3392
rect 19334 3340 19340 3392
rect 19392 3340 19398 3392
rect 19705 3383 19763 3389
rect 19705 3349 19717 3383
rect 19751 3380 19763 3383
rect 20806 3380 20812 3392
rect 19751 3352 20812 3380
rect 19751 3349 19763 3352
rect 19705 3343 19763 3349
rect 20806 3340 20812 3352
rect 20864 3340 20870 3392
rect 20993 3383 21051 3389
rect 20993 3349 21005 3383
rect 21039 3380 21051 3383
rect 24118 3380 24124 3392
rect 21039 3352 24124 3380
rect 21039 3349 21051 3352
rect 20993 3343 21051 3349
rect 24118 3340 24124 3352
rect 24176 3340 24182 3392
rect 24412 3380 24440 3420
rect 24673 3417 24685 3420
rect 24719 3417 24731 3451
rect 24673 3411 24731 3417
rect 24765 3451 24823 3457
rect 24765 3417 24777 3451
rect 24811 3417 24823 3451
rect 24765 3411 24823 3417
rect 24780 3380 24808 3411
rect 25038 3408 25044 3460
rect 25096 3448 25102 3460
rect 25700 3448 25728 3476
rect 25096 3420 25728 3448
rect 27249 3451 27307 3457
rect 25096 3408 25102 3420
rect 27249 3417 27261 3451
rect 27295 3417 27307 3451
rect 27249 3411 27307 3417
rect 27341 3451 27399 3457
rect 27341 3417 27353 3451
rect 27387 3448 27399 3451
rect 28166 3448 28172 3460
rect 27387 3420 28172 3448
rect 27387 3417 27399 3420
rect 27341 3411 27399 3417
rect 24412 3352 24808 3380
rect 27264 3380 27292 3411
rect 28166 3408 28172 3420
rect 28224 3408 28230 3460
rect 28445 3451 28503 3457
rect 28445 3417 28457 3451
rect 28491 3417 28503 3451
rect 28445 3411 28503 3417
rect 28537 3451 28595 3457
rect 28537 3417 28549 3451
rect 28583 3448 28595 3451
rect 30742 3448 30748 3460
rect 28583 3420 30748 3448
rect 28583 3417 28595 3420
rect 28537 3411 28595 3417
rect 28350 3380 28356 3392
rect 27264 3352 28356 3380
rect 28350 3340 28356 3352
rect 28408 3340 28414 3392
rect 28460 3380 28488 3411
rect 30742 3408 30748 3420
rect 30800 3408 30806 3460
rect 29825 3383 29883 3389
rect 29825 3380 29837 3383
rect 28460 3352 29837 3380
rect 29825 3349 29837 3352
rect 29871 3349 29883 3383
rect 29825 3343 29883 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 18138 3176 18144 3188
rect 18099 3148 18144 3176
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 19429 3179 19487 3185
rect 19429 3145 19441 3179
rect 19475 3176 19487 3179
rect 22002 3176 22008 3188
rect 19475 3148 22008 3176
rect 19475 3145 19487 3148
rect 19429 3139 19487 3145
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 30282 3176 30288 3188
rect 28920 3148 30288 3176
rect 18782 3068 18788 3120
rect 18840 3108 18846 3120
rect 20809 3111 20867 3117
rect 20809 3108 20821 3111
rect 18840 3080 20821 3108
rect 18840 3068 18846 3080
rect 20809 3077 20821 3080
rect 20855 3077 20867 3111
rect 20809 3071 20867 3077
rect 20898 3068 20904 3120
rect 20956 3108 20962 3120
rect 22741 3111 22799 3117
rect 22741 3108 22753 3111
rect 20956 3080 22753 3108
rect 20956 3068 20962 3080
rect 22741 3077 22753 3080
rect 22787 3077 22799 3111
rect 24118 3108 24124 3120
rect 24079 3080 24124 3108
rect 22741 3071 22799 3077
rect 24118 3068 24124 3080
rect 24176 3068 24182 3120
rect 24854 3068 24860 3120
rect 24912 3108 24918 3120
rect 25317 3111 25375 3117
rect 25317 3108 25329 3111
rect 24912 3080 25329 3108
rect 24912 3068 24918 3080
rect 25317 3077 25329 3080
rect 25363 3077 25375 3111
rect 27706 3108 27712 3120
rect 27667 3080 27712 3108
rect 25317 3071 25375 3077
rect 27706 3068 27712 3080
rect 27764 3068 27770 3120
rect 28920 3117 28948 3148
rect 30282 3136 30288 3148
rect 30340 3136 30346 3188
rect 28905 3111 28963 3117
rect 28905 3077 28917 3111
rect 28951 3077 28963 3111
rect 28905 3071 28963 3077
rect 28997 3111 29055 3117
rect 28997 3077 29009 3111
rect 29043 3108 29055 3111
rect 30006 3108 30012 3120
rect 29043 3080 30012 3108
rect 29043 3077 29055 3080
rect 28997 3071 29055 3077
rect 30006 3068 30012 3080
rect 30064 3068 30070 3120
rect 30101 3111 30159 3117
rect 30101 3077 30113 3111
rect 30147 3108 30159 3111
rect 31481 3111 31539 3117
rect 31481 3108 31493 3111
rect 30147 3080 31493 3108
rect 30147 3077 30159 3080
rect 30101 3071 30159 3077
rect 31481 3077 31493 3080
rect 31527 3077 31539 3111
rect 31481 3071 31539 3077
rect 18233 3043 18291 3049
rect 18233 3009 18245 3043
rect 18279 3040 18291 3043
rect 18690 3040 18696 3052
rect 18279 3012 18696 3040
rect 18279 3009 18291 3012
rect 18233 3003 18291 3009
rect 18690 3000 18696 3012
rect 18748 3000 18754 3052
rect 19334 3000 19340 3052
rect 19392 3040 19398 3052
rect 19521 3043 19579 3049
rect 19521 3040 19533 3043
rect 19392 3012 19533 3040
rect 19392 3000 19398 3012
rect 19521 3009 19533 3012
rect 19567 3009 19579 3043
rect 20162 3040 20168 3052
rect 20123 3012 20168 3040
rect 19521 3003 19579 3009
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 26602 3040 26608 3052
rect 26563 3012 26608 3040
rect 26602 3000 26608 3012
rect 26660 3000 26666 3052
rect 30742 3040 30748 3052
rect 30703 3012 30748 3040
rect 30742 3000 30748 3012
rect 30800 3000 30806 3052
rect 31386 3040 31392 3052
rect 31347 3012 31392 3040
rect 31386 3000 31392 3012
rect 31444 3000 31450 3052
rect 32674 3000 32680 3052
rect 32732 3040 32738 3052
rect 34241 3043 34299 3049
rect 34241 3040 34253 3043
rect 32732 3012 34253 3040
rect 32732 3000 32738 3012
rect 34241 3009 34253 3012
rect 34287 3009 34299 3043
rect 34241 3003 34299 3009
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2972 4767 2975
rect 5442 2972 5448 2984
rect 4755 2944 5448 2972
rect 4755 2941 4767 2944
rect 4709 2935 4767 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 7285 2975 7343 2981
rect 7285 2941 7297 2975
rect 7331 2972 7343 2975
rect 7926 2972 7932 2984
rect 7331 2944 7932 2972
rect 7331 2941 7343 2944
rect 7285 2935 7343 2941
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 9858 2972 9864 2984
rect 9263 2944 9864 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 14369 2975 14427 2981
rect 14369 2941 14381 2975
rect 14415 2972 14427 2975
rect 15286 2972 15292 2984
rect 14415 2944 15292 2972
rect 14415 2941 14427 2944
rect 14369 2935 14427 2941
rect 15286 2932 15292 2944
rect 15344 2932 15350 2984
rect 15657 2975 15715 2981
rect 15657 2941 15669 2975
rect 15703 2972 15715 2975
rect 17494 2972 17500 2984
rect 15703 2944 17500 2972
rect 15703 2941 15715 2944
rect 15657 2935 15715 2941
rect 17494 2932 17500 2944
rect 17552 2932 17558 2984
rect 18598 2932 18604 2984
rect 18656 2972 18662 2984
rect 20717 2975 20775 2981
rect 20717 2972 20729 2975
rect 18656 2944 20729 2972
rect 18656 2932 18662 2944
rect 20717 2941 20729 2944
rect 20763 2941 20775 2975
rect 21358 2972 21364 2984
rect 21319 2944 21364 2972
rect 20717 2935 20775 2941
rect 21358 2932 21364 2944
rect 21416 2932 21422 2984
rect 22649 2975 22707 2981
rect 22649 2941 22661 2975
rect 22695 2941 22707 2975
rect 22649 2935 22707 2941
rect 4065 2907 4123 2913
rect 4065 2873 4077 2907
rect 4111 2904 4123 2907
rect 4890 2904 4896 2916
rect 4111 2876 4896 2904
rect 4111 2873 4123 2876
rect 4065 2867 4123 2873
rect 4890 2864 4896 2876
rect 4948 2864 4954 2916
rect 5353 2907 5411 2913
rect 5353 2873 5365 2907
rect 5399 2904 5411 2907
rect 6270 2904 6276 2916
rect 5399 2876 6276 2904
rect 5399 2873 5411 2876
rect 5353 2867 5411 2873
rect 6270 2864 6276 2876
rect 6328 2864 6334 2916
rect 8754 2904 8760 2916
rect 7944 2876 8760 2904
rect 2777 2839 2835 2845
rect 2777 2805 2789 2839
rect 2823 2836 2835 2839
rect 3142 2836 3148 2848
rect 2823 2808 3148 2836
rect 2823 2805 2835 2808
rect 2777 2799 2835 2805
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 3421 2839 3479 2845
rect 3421 2805 3433 2839
rect 3467 2836 3479 2839
rect 3878 2836 3884 2848
rect 3467 2808 3884 2836
rect 3467 2805 3479 2808
rect 3421 2799 3479 2805
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 5997 2839 6055 2845
rect 5997 2805 6009 2839
rect 6043 2836 6055 2839
rect 6546 2836 6552 2848
rect 6043 2808 6552 2836
rect 6043 2805 6055 2808
rect 5997 2799 6055 2805
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 7944 2845 7972 2876
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 10505 2907 10563 2913
rect 10505 2873 10517 2907
rect 10551 2904 10563 2907
rect 11238 2904 11244 2916
rect 10551 2876 11244 2904
rect 10551 2873 10563 2876
rect 10505 2867 10563 2873
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 12437 2907 12495 2913
rect 12437 2873 12449 2907
rect 12483 2904 12495 2907
rect 13354 2904 13360 2916
rect 12483 2876 13360 2904
rect 12483 2873 12495 2876
rect 12437 2867 12495 2873
rect 13354 2864 13360 2876
rect 13412 2864 13418 2916
rect 13725 2907 13783 2913
rect 13725 2873 13737 2907
rect 13771 2904 13783 2907
rect 14458 2904 14464 2916
rect 13771 2876 14464 2904
rect 13771 2873 13783 2876
rect 13725 2867 13783 2873
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 15013 2907 15071 2913
rect 15013 2873 15025 2907
rect 15059 2904 15071 2907
rect 16666 2904 16672 2916
rect 15059 2876 16672 2904
rect 15059 2873 15071 2876
rect 15013 2867 15071 2873
rect 16666 2864 16672 2876
rect 16724 2864 16730 2916
rect 18322 2904 18328 2916
rect 17512 2876 18328 2904
rect 7929 2839 7987 2845
rect 7929 2805 7941 2839
rect 7975 2805 7987 2839
rect 7929 2799 7987 2805
rect 8573 2839 8631 2845
rect 8573 2805 8585 2839
rect 8619 2836 8631 2839
rect 9030 2836 9036 2848
rect 8619 2808 9036 2836
rect 8619 2805 8631 2808
rect 8573 2799 8631 2805
rect 9030 2796 9036 2808
rect 9088 2796 9094 2848
rect 9861 2839 9919 2845
rect 9861 2805 9873 2839
rect 9907 2836 9919 2839
rect 10686 2836 10692 2848
rect 9907 2808 10692 2836
rect 9907 2805 9919 2808
rect 9861 2799 9919 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2836 11207 2839
rect 12066 2836 12072 2848
rect 11195 2808 12072 2836
rect 11195 2805 11207 2808
rect 11149 2799 11207 2805
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 13081 2839 13139 2845
rect 13081 2805 13093 2839
rect 13127 2836 13139 2839
rect 13906 2836 13912 2848
rect 13127 2808 13912 2836
rect 13127 2805 13139 2808
rect 13081 2799 13139 2805
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 16301 2839 16359 2845
rect 16301 2805 16313 2839
rect 16347 2836 16359 2839
rect 17512 2836 17540 2876
rect 18322 2864 18328 2876
rect 18380 2864 18386 2916
rect 18877 2907 18935 2913
rect 18877 2873 18889 2907
rect 18923 2904 18935 2907
rect 22664 2904 22692 2935
rect 22738 2932 22744 2984
rect 22796 2972 22802 2984
rect 22925 2975 22983 2981
rect 22925 2972 22937 2975
rect 22796 2944 22937 2972
rect 22796 2932 22802 2944
rect 22925 2941 22937 2944
rect 22971 2941 22983 2975
rect 22925 2935 22983 2941
rect 24029 2975 24087 2981
rect 24029 2941 24041 2975
rect 24075 2941 24087 2975
rect 24394 2972 24400 2984
rect 24355 2944 24400 2972
rect 24029 2935 24087 2941
rect 18923 2876 22692 2904
rect 18923 2873 18935 2876
rect 18877 2867 18935 2873
rect 16347 2808 17540 2836
rect 17589 2839 17647 2845
rect 16347 2805 16359 2808
rect 16301 2799 16359 2805
rect 17589 2805 17601 2839
rect 17635 2836 17647 2839
rect 20530 2836 20536 2848
rect 17635 2808 20536 2836
rect 17635 2805 17647 2808
rect 17589 2799 17647 2805
rect 20530 2796 20536 2808
rect 20588 2796 20594 2848
rect 22094 2796 22100 2848
rect 22152 2836 22158 2848
rect 24044 2836 24072 2935
rect 24394 2932 24400 2944
rect 24452 2932 24458 2984
rect 24486 2932 24492 2984
rect 24544 2972 24550 2984
rect 25225 2975 25283 2981
rect 25225 2972 25237 2975
rect 24544 2944 25237 2972
rect 24544 2932 24550 2944
rect 25225 2941 25237 2944
rect 25271 2941 25283 2975
rect 25498 2972 25504 2984
rect 25459 2944 25504 2972
rect 25225 2935 25283 2941
rect 25498 2932 25504 2944
rect 25556 2932 25562 2984
rect 26878 2932 26884 2984
rect 26936 2972 26942 2984
rect 27157 2975 27215 2981
rect 27157 2972 27169 2975
rect 26936 2944 27169 2972
rect 26936 2932 26942 2944
rect 27157 2941 27169 2944
rect 27203 2941 27215 2975
rect 27798 2972 27804 2984
rect 27759 2944 27804 2972
rect 27157 2935 27215 2941
rect 27798 2932 27804 2944
rect 27856 2932 27862 2984
rect 28534 2972 28540 2984
rect 28495 2944 28540 2972
rect 28534 2932 28540 2944
rect 28592 2932 28598 2984
rect 29362 2932 29368 2984
rect 29420 2972 29426 2984
rect 29549 2975 29607 2981
rect 29549 2972 29561 2975
rect 29420 2944 29561 2972
rect 29420 2932 29426 2944
rect 29549 2941 29561 2944
rect 29595 2941 29607 2975
rect 29549 2935 29607 2941
rect 30193 2975 30251 2981
rect 30193 2941 30205 2975
rect 30239 2972 30251 2975
rect 31018 2972 31024 2984
rect 30239 2944 31024 2972
rect 30239 2941 30251 2944
rect 30193 2935 30251 2941
rect 31018 2932 31024 2944
rect 31076 2932 31082 2984
rect 32122 2932 32128 2984
rect 32180 2972 32186 2984
rect 33597 2975 33655 2981
rect 33597 2972 33609 2975
rect 32180 2944 33609 2972
rect 32180 2932 32186 2944
rect 33597 2941 33609 2944
rect 33643 2941 33655 2975
rect 33597 2935 33655 2941
rect 34054 2932 34060 2984
rect 34112 2972 34118 2984
rect 35529 2975 35587 2981
rect 35529 2972 35541 2975
rect 34112 2944 35541 2972
rect 34112 2932 34118 2944
rect 35529 2941 35541 2944
rect 35575 2941 35587 2975
rect 35529 2935 35587 2941
rect 37090 2932 37096 2984
rect 37148 2972 37154 2984
rect 38105 2975 38163 2981
rect 38105 2972 38117 2975
rect 37148 2944 38117 2972
rect 37148 2932 37154 2944
rect 38105 2941 38117 2944
rect 38151 2941 38163 2975
rect 38105 2935 38163 2941
rect 38746 2932 38752 2984
rect 38804 2972 38810 2984
rect 39393 2975 39451 2981
rect 39393 2972 39405 2975
rect 38804 2944 39405 2972
rect 38804 2932 38810 2944
rect 39393 2941 39405 2944
rect 39439 2941 39451 2975
rect 39393 2935 39451 2941
rect 40678 2932 40684 2984
rect 40736 2972 40742 2984
rect 41325 2975 41383 2981
rect 41325 2972 41337 2975
rect 40736 2944 41337 2972
rect 40736 2932 40742 2944
rect 41325 2941 41337 2944
rect 41371 2941 41383 2975
rect 41325 2935 41383 2941
rect 42610 2932 42616 2984
rect 42668 2972 42674 2984
rect 43257 2975 43315 2981
rect 43257 2972 43269 2975
rect 42668 2944 43269 2972
rect 42668 2932 42674 2944
rect 43257 2941 43269 2944
rect 43303 2941 43315 2975
rect 43257 2935 43315 2941
rect 44542 2932 44548 2984
rect 44600 2972 44606 2984
rect 45189 2975 45247 2981
rect 45189 2972 45201 2975
rect 44600 2944 45201 2972
rect 44600 2932 44606 2944
rect 45189 2941 45201 2944
rect 45235 2941 45247 2975
rect 45189 2935 45247 2941
rect 31570 2864 31576 2916
rect 31628 2904 31634 2916
rect 32953 2907 33011 2913
rect 32953 2904 32965 2907
rect 31628 2876 32965 2904
rect 31628 2864 31634 2876
rect 32953 2873 32965 2876
rect 32999 2873 33011 2907
rect 32953 2867 33011 2873
rect 33502 2864 33508 2916
rect 33560 2904 33566 2916
rect 34885 2907 34943 2913
rect 34885 2904 34897 2907
rect 33560 2876 34897 2904
rect 33560 2864 33566 2876
rect 34885 2873 34897 2876
rect 34931 2873 34943 2907
rect 34885 2867 34943 2873
rect 35342 2864 35348 2916
rect 35400 2904 35406 2916
rect 36173 2907 36231 2913
rect 36173 2904 36185 2907
rect 35400 2876 36185 2904
rect 35400 2864 35406 2876
rect 36173 2873 36185 2876
rect 36219 2873 36231 2907
rect 36173 2867 36231 2873
rect 37918 2864 37924 2916
rect 37976 2904 37982 2916
rect 37976 2876 38792 2904
rect 37976 2864 37982 2876
rect 22152 2808 24072 2836
rect 22152 2796 22158 2808
rect 30742 2796 30748 2848
rect 30800 2836 30806 2848
rect 32309 2839 32367 2845
rect 32309 2836 32321 2839
rect 30800 2808 32321 2836
rect 30800 2796 30806 2808
rect 32309 2805 32321 2808
rect 32355 2805 32367 2839
rect 32309 2799 32367 2805
rect 35986 2796 35992 2848
rect 36044 2836 36050 2848
rect 38764 2845 38792 2876
rect 37461 2839 37519 2845
rect 37461 2836 37473 2839
rect 36044 2808 37473 2836
rect 36044 2796 36050 2808
rect 37461 2805 37473 2808
rect 37507 2805 37519 2839
rect 37461 2799 37519 2805
rect 38749 2839 38807 2845
rect 38749 2805 38761 2839
rect 38795 2805 38807 2839
rect 38749 2799 38807 2805
rect 39022 2796 39028 2848
rect 39080 2836 39086 2848
rect 40037 2839 40095 2845
rect 40037 2836 40049 2839
rect 39080 2808 40049 2836
rect 39080 2796 39086 2808
rect 40037 2805 40049 2808
rect 40083 2805 40095 2839
rect 40037 2799 40095 2805
rect 40126 2796 40132 2848
rect 40184 2836 40190 2848
rect 40681 2839 40739 2845
rect 40681 2836 40693 2839
rect 40184 2808 40693 2836
rect 40184 2796 40190 2808
rect 40681 2805 40693 2808
rect 40727 2805 40739 2839
rect 40681 2799 40739 2805
rect 42058 2796 42064 2848
rect 42116 2836 42122 2848
rect 42613 2839 42671 2845
rect 42613 2836 42625 2839
rect 42116 2808 42625 2836
rect 42116 2796 42122 2808
rect 42613 2805 42625 2808
rect 42659 2805 42671 2839
rect 42613 2799 42671 2805
rect 43438 2796 43444 2848
rect 43496 2836 43502 2848
rect 43901 2839 43959 2845
rect 43901 2836 43913 2839
rect 43496 2808 43913 2836
rect 43496 2796 43502 2808
rect 43901 2805 43913 2808
rect 43947 2805 43959 2839
rect 43901 2799 43959 2805
rect 43990 2796 43996 2848
rect 44048 2836 44054 2848
rect 44545 2839 44603 2845
rect 44545 2836 44557 2839
rect 44048 2808 44557 2836
rect 44048 2796 44054 2808
rect 44545 2805 44557 2808
rect 44591 2805 44603 2839
rect 44545 2799 44603 2805
rect 45370 2796 45376 2848
rect 45428 2836 45434 2848
rect 45833 2839 45891 2845
rect 45833 2836 45845 2839
rect 45428 2808 45845 2836
rect 45428 2796 45434 2808
rect 45833 2805 45845 2808
rect 45879 2805 45891 2839
rect 45833 2799 45891 2805
rect 45922 2796 45928 2848
rect 45980 2836 45986 2848
rect 46477 2839 46535 2845
rect 46477 2836 46489 2839
rect 45980 2808 46489 2836
rect 45980 2796 45986 2808
rect 46477 2805 46489 2808
rect 46523 2805 46535 2839
rect 46477 2799 46535 2805
rect 47026 2796 47032 2848
rect 47084 2836 47090 2848
rect 47765 2839 47823 2845
rect 47765 2836 47777 2839
rect 47084 2808 47777 2836
rect 47084 2796 47090 2808
rect 47765 2805 47777 2808
rect 47811 2805 47823 2839
rect 47765 2799 47823 2805
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 15657 2635 15715 2641
rect 15657 2601 15669 2635
rect 15703 2632 15715 2635
rect 19150 2632 19156 2644
rect 15703 2604 19156 2632
rect 15703 2601 15715 2604
rect 15657 2595 15715 2601
rect 19150 2592 19156 2604
rect 19208 2592 19214 2644
rect 20622 2632 20628 2644
rect 19904 2604 20628 2632
rect 5353 2567 5411 2573
rect 5353 2533 5365 2567
rect 5399 2564 5411 2567
rect 7098 2564 7104 2576
rect 5399 2536 7104 2564
rect 5399 2533 5411 2536
rect 5353 2527 5411 2533
rect 7098 2524 7104 2536
rect 7156 2524 7162 2576
rect 7929 2567 7987 2573
rect 7929 2533 7941 2567
rect 7975 2564 7987 2567
rect 9582 2564 9588 2576
rect 7975 2536 9588 2564
rect 7975 2533 7987 2536
rect 7929 2527 7987 2533
rect 9582 2524 9588 2536
rect 9640 2524 9646 2576
rect 9861 2567 9919 2573
rect 9861 2533 9873 2567
rect 9907 2564 9919 2567
rect 11514 2564 11520 2576
rect 9907 2536 11520 2564
rect 9907 2533 9919 2536
rect 9861 2527 9919 2533
rect 11514 2524 11520 2536
rect 11572 2524 11578 2576
rect 12437 2567 12495 2573
rect 12437 2533 12449 2567
rect 12483 2564 12495 2567
rect 14182 2564 14188 2576
rect 12483 2536 14188 2564
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 14182 2524 14188 2536
rect 14240 2524 14246 2576
rect 18233 2567 18291 2573
rect 18233 2533 18245 2567
rect 18279 2564 18291 2567
rect 19904 2564 19932 2604
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 20809 2635 20867 2641
rect 20809 2601 20821 2635
rect 20855 2632 20867 2635
rect 22094 2632 22100 2644
rect 20855 2604 22100 2632
rect 20855 2601 20867 2604
rect 20809 2595 20867 2601
rect 22094 2592 22100 2604
rect 22152 2592 22158 2644
rect 22189 2635 22247 2641
rect 22189 2601 22201 2635
rect 22235 2632 22247 2635
rect 24486 2632 24492 2644
rect 22235 2604 24492 2632
rect 22235 2601 22247 2604
rect 22189 2595 22247 2601
rect 24486 2592 24492 2604
rect 24544 2592 24550 2644
rect 27249 2635 27307 2641
rect 27249 2601 27261 2635
rect 27295 2632 27307 2635
rect 27338 2632 27344 2644
rect 27295 2604 27344 2632
rect 27295 2601 27307 2604
rect 27249 2595 27307 2601
rect 27338 2592 27344 2604
rect 27396 2592 27402 2644
rect 27798 2632 27804 2644
rect 27759 2604 27804 2632
rect 27798 2592 27804 2604
rect 27856 2592 27862 2644
rect 28350 2592 28356 2644
rect 28408 2632 28414 2644
rect 28537 2635 28595 2641
rect 28537 2632 28549 2635
rect 28408 2604 28549 2632
rect 28408 2592 28414 2604
rect 28537 2601 28549 2604
rect 28583 2601 28595 2635
rect 28537 2595 28595 2601
rect 30282 2592 30288 2644
rect 30340 2632 30346 2644
rect 30469 2635 30527 2641
rect 30469 2632 30481 2635
rect 30340 2604 30481 2632
rect 30340 2592 30346 2604
rect 30469 2601 30481 2604
rect 30515 2601 30527 2635
rect 31018 2632 31024 2644
rect 30979 2604 31024 2632
rect 30469 2595 30527 2601
rect 31018 2592 31024 2604
rect 31076 2592 31082 2644
rect 18279 2536 19932 2564
rect 20073 2567 20131 2573
rect 18279 2533 18291 2536
rect 18233 2527 18291 2533
rect 20073 2533 20085 2567
rect 20119 2564 20131 2567
rect 20898 2564 20904 2576
rect 20119 2536 20904 2564
rect 20119 2533 20131 2536
rect 20073 2527 20131 2533
rect 20898 2524 20904 2536
rect 20956 2524 20962 2576
rect 21453 2567 21511 2573
rect 21453 2533 21465 2567
rect 21499 2564 21511 2567
rect 26513 2567 26571 2573
rect 21499 2536 25360 2564
rect 21499 2533 21511 2536
rect 21453 2527 21511 2533
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 3510 2496 3516 2508
rect 2823 2468 3516 2496
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 3510 2456 3516 2468
rect 3568 2456 3574 2508
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2496 7343 2499
rect 8202 2496 8208 2508
rect 7331 2468 8208 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 10410 2496 10416 2508
rect 8619 2468 10416 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 10410 2456 10416 2468
rect 10468 2456 10474 2508
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2496 11207 2499
rect 12802 2496 12808 2508
rect 11195 2468 12808 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 12802 2456 12808 2468
rect 12860 2456 12866 2508
rect 13081 2499 13139 2505
rect 13081 2465 13093 2499
rect 13127 2496 13139 2499
rect 14734 2496 14740 2508
rect 13127 2468 14740 2496
rect 13127 2465 13139 2468
rect 13081 2459 13139 2465
rect 14734 2456 14740 2468
rect 14792 2456 14798 2508
rect 15013 2499 15071 2505
rect 15013 2465 15025 2499
rect 15059 2496 15071 2499
rect 17770 2496 17776 2508
rect 15059 2468 17776 2496
rect 15059 2465 15071 2468
rect 15013 2459 15071 2465
rect 17770 2456 17776 2468
rect 17828 2456 17834 2508
rect 18877 2499 18935 2505
rect 18877 2465 18889 2499
rect 18923 2496 18935 2499
rect 22741 2499 22799 2505
rect 22741 2496 22753 2499
rect 18923 2468 22753 2496
rect 18923 2465 18935 2468
rect 18877 2459 18935 2465
rect 22741 2465 22753 2468
rect 22787 2465 22799 2499
rect 23014 2496 23020 2508
rect 22975 2468 23020 2496
rect 22741 2459 22799 2465
rect 23014 2456 23020 2468
rect 23072 2456 23078 2508
rect 23937 2499 23995 2505
rect 23937 2465 23949 2499
rect 23983 2496 23995 2499
rect 24854 2496 24860 2508
rect 23983 2468 24860 2496
rect 23983 2465 23995 2468
rect 23937 2459 23995 2465
rect 24854 2456 24860 2468
rect 24912 2456 24918 2508
rect 25332 2505 25360 2536
rect 26513 2533 26525 2567
rect 26559 2564 26571 2567
rect 27706 2564 27712 2576
rect 26559 2536 27712 2564
rect 26559 2533 26571 2536
rect 26513 2527 26571 2533
rect 27706 2524 27712 2536
rect 27764 2524 27770 2576
rect 28166 2524 28172 2576
rect 28224 2564 28230 2576
rect 29733 2567 29791 2573
rect 29733 2564 29745 2567
rect 28224 2536 29745 2564
rect 28224 2524 28230 2536
rect 29733 2533 29745 2536
rect 29779 2533 29791 2567
rect 29733 2527 29791 2533
rect 29914 2524 29920 2576
rect 29972 2564 29978 2576
rect 32309 2567 32367 2573
rect 32309 2564 32321 2567
rect 29972 2536 32321 2564
rect 29972 2524 29978 2536
rect 32309 2533 32321 2536
rect 32355 2533 32367 2567
rect 32309 2527 32367 2533
rect 33226 2524 33232 2576
rect 33284 2564 33290 2576
rect 34885 2567 34943 2573
rect 34885 2564 34897 2567
rect 33284 2536 34897 2564
rect 33284 2524 33290 2536
rect 34885 2533 34897 2536
rect 34931 2533 34943 2567
rect 34885 2527 34943 2533
rect 35434 2524 35440 2576
rect 35492 2564 35498 2576
rect 37461 2567 37519 2573
rect 37461 2564 37473 2567
rect 35492 2536 37473 2564
rect 35492 2524 35498 2536
rect 37461 2533 37473 2536
rect 37507 2533 37519 2567
rect 37461 2527 37519 2533
rect 38470 2524 38476 2576
rect 38528 2564 38534 2576
rect 40037 2567 40095 2573
rect 40037 2564 40049 2567
rect 38528 2536 40049 2564
rect 38528 2524 38534 2536
rect 40037 2533 40049 2536
rect 40083 2533 40095 2567
rect 40037 2527 40095 2533
rect 42334 2524 42340 2576
rect 42392 2564 42398 2576
rect 43901 2567 43959 2573
rect 43901 2564 43913 2567
rect 42392 2536 43913 2564
rect 42392 2524 42398 2536
rect 43901 2533 43913 2536
rect 43947 2533 43959 2567
rect 43901 2527 43959 2533
rect 45094 2524 45100 2576
rect 45152 2564 45158 2576
rect 46477 2567 46535 2573
rect 46477 2564 46489 2567
rect 45152 2536 46489 2564
rect 45152 2524 45158 2536
rect 46477 2533 46489 2536
rect 46523 2533 46535 2567
rect 46477 2527 46535 2533
rect 25317 2499 25375 2505
rect 25317 2465 25329 2499
rect 25363 2465 25375 2499
rect 25774 2496 25780 2508
rect 25735 2468 25780 2496
rect 25317 2459 25375 2465
rect 25774 2456 25780 2468
rect 25832 2456 25838 2508
rect 31294 2456 31300 2508
rect 31352 2496 31358 2508
rect 33597 2499 33655 2505
rect 33597 2496 33609 2499
rect 31352 2468 33609 2496
rect 31352 2456 31358 2468
rect 33597 2465 33609 2468
rect 33643 2465 33655 2499
rect 33597 2459 33655 2465
rect 34606 2456 34612 2508
rect 34664 2496 34670 2508
rect 36173 2499 36231 2505
rect 36173 2496 36185 2499
rect 34664 2468 36185 2496
rect 34664 2456 34670 2468
rect 36173 2465 36185 2468
rect 36219 2465 36231 2499
rect 36173 2459 36231 2465
rect 37366 2456 37372 2508
rect 37424 2496 37430 2508
rect 38749 2499 38807 2505
rect 38749 2496 38761 2499
rect 37424 2468 38761 2496
rect 37424 2456 37430 2468
rect 38749 2465 38761 2468
rect 38795 2465 38807 2499
rect 38749 2459 38807 2465
rect 39298 2456 39304 2508
rect 39356 2496 39362 2508
rect 40681 2499 40739 2505
rect 40681 2496 40693 2499
rect 39356 2468 40693 2496
rect 39356 2456 39362 2468
rect 40681 2465 40693 2468
rect 40727 2465 40739 2499
rect 40681 2459 40739 2465
rect 41230 2456 41236 2508
rect 41288 2496 41294 2508
rect 42613 2499 42671 2505
rect 42613 2496 42625 2499
rect 41288 2468 42625 2496
rect 41288 2456 41294 2468
rect 42613 2465 42625 2468
rect 42659 2465 42671 2499
rect 42613 2459 42671 2465
rect 43714 2456 43720 2508
rect 43772 2496 43778 2508
rect 45189 2499 45247 2505
rect 45189 2496 45201 2499
rect 43772 2468 45201 2496
rect 43772 2456 43778 2468
rect 45189 2465 45201 2468
rect 45235 2465 45247 2499
rect 45189 2459 45247 2465
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2590 2428 2596 2440
rect 2179 2400 2596 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 4614 2428 4620 2440
rect 3467 2400 4620 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 5718 2428 5724 2440
rect 4755 2400 5724 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 10505 2431 10563 2437
rect 6043 2400 6914 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6886 2360 6914 2400
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 12250 2428 12256 2440
rect 10551 2400 12256 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 12250 2388 12256 2400
rect 12308 2388 12314 2440
rect 13725 2431 13783 2437
rect 13725 2397 13737 2431
rect 13771 2428 13783 2431
rect 15562 2428 15568 2440
rect 13771 2400 15568 2428
rect 13771 2397 13783 2400
rect 13725 2391 13783 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 16301 2431 16359 2437
rect 16301 2397 16313 2431
rect 16347 2428 16359 2431
rect 17589 2431 17647 2437
rect 16347 2400 16574 2428
rect 16347 2397 16359 2400
rect 16301 2391 16359 2397
rect 7374 2360 7380 2372
rect 6886 2332 7380 2360
rect 7374 2320 7380 2332
rect 7432 2320 7438 2372
rect 16546 2360 16574 2400
rect 17589 2397 17601 2431
rect 17635 2428 17647 2431
rect 17635 2400 19196 2428
rect 17635 2397 17647 2400
rect 17589 2391 17647 2397
rect 17402 2360 17408 2372
rect 16546 2332 17408 2360
rect 17402 2320 17408 2332
rect 17460 2320 17466 2372
rect 19168 2292 19196 2400
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19981 2431 20039 2437
rect 19981 2428 19993 2431
rect 19392 2400 19993 2428
rect 19392 2388 19398 2400
rect 19981 2397 19993 2400
rect 20027 2397 20039 2431
rect 19981 2391 20039 2397
rect 24029 2431 24087 2437
rect 24029 2397 24041 2431
rect 24075 2428 24087 2431
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 24075 2400 24593 2428
rect 24075 2397 24087 2400
rect 24029 2391 24087 2397
rect 24581 2397 24593 2400
rect 24627 2428 24639 2431
rect 25038 2428 25044 2440
rect 24627 2400 25044 2428
rect 24627 2397 24639 2400
rect 24581 2391 24639 2397
rect 25038 2388 25044 2400
rect 25096 2388 25102 2440
rect 26605 2431 26663 2437
rect 26605 2397 26617 2431
rect 26651 2428 26663 2431
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 26651 2400 27169 2428
rect 26651 2397 26663 2400
rect 26605 2391 26663 2397
rect 27157 2397 27169 2400
rect 27203 2428 27215 2431
rect 27890 2428 27896 2440
rect 27203 2400 27896 2428
rect 27203 2397 27215 2400
rect 27157 2391 27215 2397
rect 27890 2388 27896 2400
rect 27948 2428 27954 2440
rect 28445 2431 28503 2437
rect 28445 2428 28457 2431
rect 27948 2400 28457 2428
rect 27948 2388 27954 2400
rect 28445 2397 28457 2400
rect 28491 2397 28503 2431
rect 28445 2391 28503 2397
rect 30561 2431 30619 2437
rect 30561 2397 30573 2431
rect 30607 2428 30619 2431
rect 31386 2428 31392 2440
rect 30607 2400 31392 2428
rect 30607 2397 30619 2400
rect 30561 2391 30619 2397
rect 31386 2388 31392 2400
rect 31444 2388 31450 2440
rect 32953 2431 33011 2437
rect 32953 2397 32965 2431
rect 32999 2397 33011 2431
rect 32953 2391 33011 2397
rect 22002 2320 22008 2372
rect 22060 2360 22066 2372
rect 22833 2363 22891 2369
rect 22833 2360 22845 2363
rect 22060 2332 22845 2360
rect 22060 2320 22066 2332
rect 22833 2329 22845 2332
rect 22879 2329 22891 2363
rect 22833 2323 22891 2329
rect 25409 2363 25467 2369
rect 25409 2329 25421 2363
rect 25455 2329 25467 2363
rect 25409 2323 25467 2329
rect 20806 2292 20812 2304
rect 19168 2264 20812 2292
rect 20806 2252 20812 2264
rect 20864 2252 20870 2304
rect 24673 2295 24731 2301
rect 24673 2261 24685 2295
rect 24719 2292 24731 2295
rect 25424 2292 25452 2323
rect 30466 2320 30472 2372
rect 30524 2360 30530 2372
rect 32968 2360 32996 2391
rect 33778 2388 33784 2440
rect 33836 2428 33842 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 33836 2400 35541 2428
rect 33836 2388 33842 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 36538 2388 36544 2440
rect 36596 2428 36602 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 36596 2400 38117 2428
rect 36596 2388 36602 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 39850 2388 39856 2440
rect 39908 2428 39914 2440
rect 41325 2431 41383 2437
rect 41325 2428 41337 2431
rect 39908 2400 41337 2428
rect 39908 2388 39914 2400
rect 41325 2397 41337 2400
rect 41371 2397 41383 2431
rect 41325 2391 41383 2397
rect 41782 2388 41788 2440
rect 41840 2428 41846 2440
rect 43257 2431 43315 2437
rect 43257 2428 43269 2431
rect 41840 2400 43269 2428
rect 41840 2388 41846 2400
rect 43257 2397 43269 2400
rect 43303 2397 43315 2431
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 43257 2391 43315 2397
rect 45526 2400 45845 2428
rect 30524 2332 32996 2360
rect 30524 2320 30530 2332
rect 44266 2320 44272 2372
rect 44324 2360 44330 2372
rect 45526 2360 45554 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 46198 2388 46204 2440
rect 46256 2428 46262 2440
rect 47765 2431 47823 2437
rect 47765 2428 47777 2431
rect 46256 2400 47777 2428
rect 46256 2388 46262 2400
rect 47765 2397 47777 2400
rect 47811 2397 47823 2431
rect 47765 2391 47823 2397
rect 44324 2332 45554 2360
rect 44324 2320 44330 2332
rect 24719 2264 25452 2292
rect 24719 2261 24731 2264
rect 24673 2255 24731 2261
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 17402 1844 17408 1896
rect 17460 1884 17466 1896
rect 19978 1884 19984 1896
rect 17460 1856 19984 1884
rect 17460 1844 17466 1856
rect 19978 1844 19984 1856
rect 20036 1844 20042 1896
<< via1 >>
rect 19432 47744 19484 47796
rect 23940 47744 23992 47796
rect 16948 47676 17000 47728
rect 23756 47676 23808 47728
rect 18880 47608 18932 47660
rect 24584 47608 24636 47660
rect 5080 47540 5132 47592
rect 22100 47540 22152 47592
rect 29000 47540 29052 47592
rect 34704 47540 34756 47592
rect 36452 47540 36504 47592
rect 41236 47540 41288 47592
rect 17592 47472 17644 47524
rect 21272 47472 21324 47524
rect 23756 47472 23808 47524
rect 24768 47472 24820 47524
rect 27528 47472 27580 47524
rect 33600 47472 33652 47524
rect 36360 47472 36412 47524
rect 11704 47404 11756 47456
rect 20076 47404 20128 47456
rect 22192 47404 22244 47456
rect 29644 47404 29696 47456
rect 31576 47404 31628 47456
rect 36544 47404 36596 47456
rect 41972 47404 42024 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 4712 47243 4764 47252
rect 4712 47209 4721 47243
rect 4721 47209 4755 47243
rect 4755 47209 4764 47243
rect 4712 47200 4764 47209
rect 5816 47200 5868 47252
rect 6000 47243 6052 47252
rect 6000 47209 6009 47243
rect 6009 47209 6043 47243
rect 6043 47209 6052 47243
rect 6000 47200 6052 47209
rect 7104 47243 7156 47252
rect 7104 47209 7113 47243
rect 7113 47209 7147 47243
rect 7147 47209 7156 47243
rect 7104 47200 7156 47209
rect 7748 47243 7800 47252
rect 7748 47209 7757 47243
rect 7757 47209 7791 47243
rect 7791 47209 7800 47243
rect 7748 47200 7800 47209
rect 8392 47243 8444 47252
rect 8392 47209 8401 47243
rect 8401 47209 8435 47243
rect 8435 47209 8444 47243
rect 8392 47200 8444 47209
rect 9128 47243 9180 47252
rect 9128 47209 9137 47243
rect 9137 47209 9171 47243
rect 9171 47209 9180 47243
rect 9128 47200 9180 47209
rect 10232 47243 10284 47252
rect 10232 47209 10241 47243
rect 10241 47209 10275 47243
rect 10275 47209 10284 47243
rect 10232 47200 10284 47209
rect 11152 47243 11204 47252
rect 11152 47209 11161 47243
rect 11161 47209 11195 47243
rect 11195 47209 11204 47243
rect 11152 47200 11204 47209
rect 12440 47243 12492 47252
rect 12440 47209 12449 47243
rect 12449 47209 12483 47243
rect 12483 47209 12492 47243
rect 13544 47243 13596 47252
rect 12440 47200 12492 47209
rect 13544 47209 13553 47243
rect 13553 47209 13587 47243
rect 13587 47209 13596 47243
rect 13544 47200 13596 47209
rect 15752 47200 15804 47252
rect 19064 47200 19116 47252
rect 20076 47243 20128 47252
rect 20076 47209 20085 47243
rect 20085 47209 20119 47243
rect 20119 47209 20128 47243
rect 20076 47200 20128 47209
rect 22100 47243 22152 47252
rect 22100 47209 22109 47243
rect 22109 47209 22143 47243
rect 22143 47209 22152 47243
rect 22100 47200 22152 47209
rect 26792 47200 26844 47252
rect 32680 47200 32732 47252
rect 39304 47200 39356 47252
rect 43352 47200 43404 47252
rect 44088 47200 44140 47252
rect 44824 47200 44876 47252
rect 45836 47243 45888 47252
rect 45836 47209 45845 47243
rect 45845 47209 45879 47243
rect 45879 47209 45888 47243
rect 45836 47200 45888 47209
rect 45928 47200 45980 47252
rect 16856 47132 16908 47184
rect 16948 47175 17000 47184
rect 16948 47141 16957 47175
rect 16957 47141 16991 47175
rect 16991 47141 17000 47175
rect 17592 47175 17644 47184
rect 16948 47132 17000 47141
rect 17592 47141 17601 47175
rect 17601 47141 17635 47175
rect 17635 47141 17644 47175
rect 17592 47132 17644 47141
rect 18880 47175 18932 47184
rect 18880 47141 18889 47175
rect 18889 47141 18923 47175
rect 18923 47141 18932 47175
rect 18880 47132 18932 47141
rect 19340 47132 19392 47184
rect 19984 47132 20036 47184
rect 22376 47132 22428 47184
rect 28264 47132 28316 47184
rect 30472 47132 30524 47184
rect 36820 47132 36872 47184
rect 41880 47132 41932 47184
rect 41972 47175 42024 47184
rect 41972 47141 41981 47175
rect 41981 47141 42015 47175
rect 42015 47141 42024 47175
rect 41972 47132 42024 47141
rect 16120 46860 16172 46912
rect 19064 46996 19116 47048
rect 21364 47064 21416 47116
rect 17960 46928 18012 46980
rect 21272 47039 21324 47048
rect 21272 47005 21281 47039
rect 21281 47005 21315 47039
rect 21315 47005 21324 47039
rect 21272 46996 21324 47005
rect 22192 46996 22244 47048
rect 22376 47039 22428 47048
rect 22376 47005 22385 47039
rect 22385 47005 22419 47039
rect 22419 47005 22428 47039
rect 23388 47064 23440 47116
rect 25780 47064 25832 47116
rect 28724 47107 28776 47116
rect 22376 46996 22428 47005
rect 23572 46996 23624 47048
rect 23756 46996 23808 47048
rect 21824 46928 21876 46980
rect 22928 46928 22980 46980
rect 24584 46928 24636 46980
rect 25872 47039 25924 47048
rect 25136 46971 25188 46980
rect 18512 46860 18564 46912
rect 19800 46860 19852 46912
rect 20076 46860 20128 46912
rect 22744 46860 22796 46912
rect 23664 46860 23716 46912
rect 25136 46937 25145 46971
rect 25145 46937 25179 46971
rect 25179 46937 25188 46971
rect 25136 46928 25188 46937
rect 25872 47005 25881 47039
rect 25881 47005 25915 47039
rect 25915 47005 25924 47039
rect 25872 46996 25924 47005
rect 26516 46996 26568 47048
rect 27344 47039 27396 47048
rect 27344 47005 27353 47039
rect 27353 47005 27387 47039
rect 27387 47005 27396 47039
rect 27344 46996 27396 47005
rect 26608 46928 26660 46980
rect 28724 47073 28733 47107
rect 28733 47073 28767 47107
rect 28767 47073 28776 47107
rect 28724 47064 28776 47073
rect 29276 47064 29328 47116
rect 28816 47039 28868 47048
rect 28816 47005 28825 47039
rect 28825 47005 28859 47039
rect 28859 47005 28868 47039
rect 28816 46996 28868 47005
rect 29092 47039 29144 47048
rect 29092 47005 29101 47039
rect 29101 47005 29135 47039
rect 29135 47005 29144 47039
rect 29092 46996 29144 47005
rect 30656 46996 30708 47048
rect 30564 46971 30616 46980
rect 25044 46903 25096 46912
rect 25044 46869 25053 46903
rect 25053 46869 25087 46903
rect 25087 46869 25096 46903
rect 25044 46860 25096 46869
rect 25688 46903 25740 46912
rect 25688 46869 25697 46903
rect 25697 46869 25731 46903
rect 25731 46869 25740 46903
rect 25688 46860 25740 46869
rect 26056 46860 26108 46912
rect 30564 46937 30573 46971
rect 30573 46937 30607 46971
rect 30607 46937 30616 46971
rect 30564 46928 30616 46937
rect 32036 46996 32088 47048
rect 31024 46971 31076 46980
rect 27252 46860 27304 46912
rect 31024 46937 31033 46971
rect 31033 46937 31067 46971
rect 31067 46937 31076 46971
rect 31024 46928 31076 46937
rect 30932 46903 30984 46912
rect 30932 46869 30941 46903
rect 30941 46869 30975 46903
rect 30975 46869 30984 46903
rect 30932 46860 30984 46869
rect 31484 46860 31536 46912
rect 31760 46860 31812 46912
rect 33324 46996 33376 47048
rect 33232 46928 33284 46980
rect 34244 47064 34296 47116
rect 34520 47064 34572 47116
rect 33600 47039 33652 47048
rect 33600 47005 33609 47039
rect 33609 47005 33643 47039
rect 33643 47005 33652 47039
rect 33876 47039 33928 47048
rect 33600 46996 33652 47005
rect 33876 47005 33885 47039
rect 33885 47005 33919 47039
rect 33919 47005 33928 47039
rect 33876 46996 33928 47005
rect 34704 46996 34756 47048
rect 37740 47064 37792 47116
rect 35900 46996 35952 47048
rect 36820 47039 36872 47048
rect 36820 47005 36829 47039
rect 36829 47005 36863 47039
rect 36863 47005 36872 47039
rect 36820 46996 36872 47005
rect 37648 46996 37700 47048
rect 39488 47064 39540 47116
rect 38016 47039 38068 47048
rect 38016 47005 38025 47039
rect 38025 47005 38059 47039
rect 38059 47005 38068 47039
rect 38016 46996 38068 47005
rect 40132 46996 40184 47048
rect 40684 47039 40736 47048
rect 40684 47005 40693 47039
rect 40693 47005 40727 47039
rect 40727 47005 40736 47039
rect 40684 46996 40736 47005
rect 32772 46860 32824 46912
rect 37740 46860 37792 46912
rect 38384 46860 38436 46912
rect 39672 46860 39724 46912
rect 40224 46860 40276 46912
rect 43260 47039 43312 47048
rect 41236 46928 41288 46980
rect 43260 47005 43269 47039
rect 43269 47005 43303 47039
rect 43303 47005 43312 47039
rect 43260 46996 43312 47005
rect 44088 46928 44140 46980
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 19340 46656 19392 46708
rect 19432 46656 19484 46708
rect 19892 46656 19944 46708
rect 18328 46588 18380 46640
rect 6920 46563 6972 46572
rect 6920 46529 6929 46563
rect 6929 46529 6963 46563
rect 6963 46529 6972 46563
rect 14648 46563 14700 46572
rect 6920 46520 6972 46529
rect 14648 46529 14657 46563
rect 14657 46529 14691 46563
rect 14691 46529 14700 46563
rect 14648 46520 14700 46529
rect 17960 46563 18012 46572
rect 17960 46529 17969 46563
rect 17969 46529 18003 46563
rect 18003 46529 18012 46563
rect 17960 46520 18012 46529
rect 18972 46520 19024 46572
rect 20444 46588 20496 46640
rect 21272 46656 21324 46708
rect 21456 46588 21508 46640
rect 18052 46452 18104 46504
rect 19892 46563 19944 46572
rect 19892 46529 19901 46563
rect 19901 46529 19935 46563
rect 19935 46529 19944 46563
rect 19892 46520 19944 46529
rect 20260 46520 20312 46572
rect 20536 46520 20588 46572
rect 21180 46563 21232 46572
rect 21180 46529 21191 46563
rect 21191 46529 21225 46563
rect 21225 46529 21232 46563
rect 21180 46520 21232 46529
rect 15016 46384 15068 46436
rect 19708 46495 19760 46504
rect 19708 46461 19717 46495
rect 19717 46461 19751 46495
rect 19751 46461 19760 46495
rect 19708 46452 19760 46461
rect 23480 46588 23532 46640
rect 23848 46631 23900 46640
rect 23848 46597 23857 46631
rect 23857 46597 23891 46631
rect 23891 46597 23900 46631
rect 23848 46588 23900 46597
rect 24308 46631 24360 46640
rect 24308 46597 24317 46631
rect 24317 46597 24351 46631
rect 24351 46597 24360 46631
rect 24308 46588 24360 46597
rect 22744 46520 22796 46572
rect 22928 46520 22980 46572
rect 23296 46563 23348 46572
rect 23296 46529 23304 46563
rect 23304 46529 23338 46563
rect 23338 46529 23348 46563
rect 23296 46520 23348 46529
rect 23388 46563 23440 46572
rect 23388 46529 23397 46563
rect 23397 46529 23431 46563
rect 23431 46529 23440 46563
rect 23664 46563 23716 46572
rect 23388 46520 23440 46529
rect 23664 46529 23673 46563
rect 23673 46529 23707 46563
rect 23707 46529 23716 46563
rect 24860 46588 24912 46640
rect 25228 46699 25280 46708
rect 25228 46665 25237 46699
rect 25237 46665 25271 46699
rect 25271 46665 25280 46699
rect 25228 46656 25280 46665
rect 25872 46656 25924 46708
rect 25688 46588 25740 46640
rect 28632 46656 28684 46708
rect 28264 46631 28316 46640
rect 23664 46520 23716 46529
rect 23204 46452 23256 46504
rect 24308 46452 24360 46504
rect 25780 46520 25832 46572
rect 26608 46563 26660 46572
rect 25228 46452 25280 46504
rect 26608 46529 26617 46563
rect 26617 46529 26651 46563
rect 26651 46529 26660 46563
rect 26608 46520 26660 46529
rect 26884 46520 26936 46572
rect 27528 46563 27580 46572
rect 27528 46529 27537 46563
rect 27537 46529 27571 46563
rect 27571 46529 27580 46563
rect 27528 46520 27580 46529
rect 26516 46452 26568 46504
rect 27804 46563 27856 46572
rect 27804 46529 27813 46563
rect 27813 46529 27847 46563
rect 27847 46529 27856 46563
rect 27804 46520 27856 46529
rect 28264 46597 28273 46631
rect 28273 46597 28307 46631
rect 28307 46597 28316 46631
rect 28264 46588 28316 46597
rect 29644 46699 29696 46708
rect 29644 46665 29653 46699
rect 29653 46665 29687 46699
rect 29687 46665 29696 46699
rect 29644 46656 29696 46665
rect 30104 46656 30156 46708
rect 34520 46656 34572 46708
rect 34980 46656 35032 46708
rect 30288 46588 30340 46640
rect 29276 46563 29328 46572
rect 29276 46529 29285 46563
rect 29285 46529 29319 46563
rect 29319 46529 29328 46563
rect 29276 46520 29328 46529
rect 29460 46563 29512 46572
rect 29460 46529 29469 46563
rect 29469 46529 29503 46563
rect 29503 46529 29512 46563
rect 29460 46520 29512 46529
rect 29828 46520 29880 46572
rect 30656 46588 30708 46640
rect 33140 46588 33192 46640
rect 30932 46520 30984 46572
rect 31668 46563 31720 46572
rect 31024 46495 31076 46504
rect 13912 46316 13964 46368
rect 19294 46316 19346 46368
rect 22376 46427 22428 46436
rect 20076 46316 20128 46368
rect 22376 46393 22385 46427
rect 22385 46393 22419 46427
rect 22419 46393 22428 46427
rect 22376 46384 22428 46393
rect 23940 46384 23992 46436
rect 22836 46316 22888 46368
rect 22928 46316 22980 46368
rect 23756 46316 23808 46368
rect 27068 46316 27120 46368
rect 27252 46359 27304 46368
rect 27252 46325 27261 46359
rect 27261 46325 27295 46359
rect 27295 46325 27304 46359
rect 27252 46316 27304 46325
rect 31024 46461 31033 46495
rect 31033 46461 31067 46495
rect 31067 46461 31076 46495
rect 31024 46452 31076 46461
rect 31668 46529 31677 46563
rect 31677 46529 31711 46563
rect 31711 46529 31720 46563
rect 31668 46520 31720 46529
rect 32496 46563 32548 46572
rect 32496 46529 32505 46563
rect 32505 46529 32539 46563
rect 32539 46529 32548 46563
rect 32496 46520 32548 46529
rect 33232 46520 33284 46572
rect 34244 46520 34296 46572
rect 35532 46588 35584 46640
rect 36728 46656 36780 46708
rect 39948 46656 40000 46708
rect 40040 46656 40092 46708
rect 43260 46656 43312 46708
rect 37096 46588 37148 46640
rect 34612 46563 34664 46572
rect 34612 46529 34641 46563
rect 34641 46529 34664 46563
rect 34612 46520 34664 46529
rect 34796 46520 34848 46572
rect 34980 46520 35032 46572
rect 35624 46563 35676 46572
rect 35624 46529 35631 46563
rect 35631 46529 35665 46563
rect 35665 46529 35676 46563
rect 35624 46520 35676 46529
rect 35992 46520 36044 46572
rect 37188 46520 37240 46572
rect 37740 46520 37792 46572
rect 38016 46520 38068 46572
rect 33876 46452 33928 46504
rect 34336 46495 34388 46504
rect 34336 46461 34345 46495
rect 34345 46461 34379 46495
rect 34379 46461 34388 46495
rect 34336 46452 34388 46461
rect 36728 46452 36780 46504
rect 37464 46452 37516 46504
rect 34888 46384 34940 46436
rect 31668 46316 31720 46368
rect 35348 46316 35400 46368
rect 35992 46359 36044 46368
rect 35992 46325 36001 46359
rect 36001 46325 36035 46359
rect 36035 46325 36044 46359
rect 35992 46316 36044 46325
rect 36544 46359 36596 46368
rect 36544 46325 36553 46359
rect 36553 46325 36587 46359
rect 36587 46325 36596 46359
rect 36544 46316 36596 46325
rect 37648 46359 37700 46368
rect 37648 46325 37657 46359
rect 37657 46325 37691 46359
rect 37691 46325 37700 46359
rect 37648 46316 37700 46325
rect 39028 46520 39080 46572
rect 38476 46452 38528 46504
rect 38844 46452 38896 46504
rect 38292 46384 38344 46436
rect 42616 46520 42668 46572
rect 43904 46563 43956 46572
rect 43904 46529 43913 46563
rect 43913 46529 43947 46563
rect 43947 46529 43956 46563
rect 43904 46520 43956 46529
rect 44548 46563 44600 46572
rect 44548 46529 44557 46563
rect 44557 46529 44591 46563
rect 44591 46529 44600 46563
rect 44548 46520 44600 46529
rect 42708 46452 42760 46504
rect 45192 46452 45244 46504
rect 39120 46427 39172 46436
rect 39120 46393 39129 46427
rect 39129 46393 39163 46427
rect 39163 46393 39172 46427
rect 39120 46384 39172 46393
rect 40040 46384 40092 46436
rect 41144 46384 41196 46436
rect 41696 46359 41748 46368
rect 41696 46325 41705 46359
rect 41705 46325 41739 46359
rect 41739 46325 41748 46359
rect 41696 46316 41748 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 18512 46112 18564 46164
rect 19708 46112 19760 46164
rect 12808 46044 12860 46096
rect 19294 46044 19346 46096
rect 19892 46044 19944 46096
rect 20076 46087 20128 46096
rect 20076 46053 20085 46087
rect 20085 46053 20119 46087
rect 20119 46053 20128 46087
rect 20076 46044 20128 46053
rect 20444 46112 20496 46164
rect 26424 46112 26476 46164
rect 27068 46112 27120 46164
rect 21640 46044 21692 46096
rect 18420 45908 18472 45960
rect 20168 45976 20220 46028
rect 23388 46044 23440 46096
rect 25136 46087 25188 46096
rect 25136 46053 25145 46087
rect 25145 46053 25179 46087
rect 25179 46053 25188 46087
rect 25136 46044 25188 46053
rect 18880 45951 18932 45960
rect 18880 45917 18889 45951
rect 18889 45917 18923 45951
rect 18923 45917 18932 45951
rect 18880 45908 18932 45917
rect 18696 45840 18748 45892
rect 19432 45917 19448 45926
rect 19448 45917 19482 45926
rect 19482 45917 19484 45926
rect 19432 45874 19484 45917
rect 19616 45908 19668 45960
rect 20444 45908 20496 45960
rect 21180 45908 21232 45960
rect 22652 45976 22704 46028
rect 23664 46019 23716 46028
rect 23664 45985 23673 46019
rect 23673 45985 23707 46019
rect 23707 45985 23716 46019
rect 23664 45976 23716 45985
rect 23848 45976 23900 46028
rect 25596 46044 25648 46096
rect 27804 46112 27856 46164
rect 27896 46112 27948 46164
rect 34796 46112 34848 46164
rect 37372 46155 37424 46164
rect 37372 46121 37381 46155
rect 37381 46121 37415 46155
rect 37415 46121 37424 46155
rect 37372 46112 37424 46121
rect 38016 46112 38068 46164
rect 38936 46112 38988 46164
rect 41512 46112 41564 46164
rect 42248 46112 42300 46164
rect 44088 46112 44140 46164
rect 26332 45976 26384 46028
rect 27252 45976 27304 46028
rect 28816 46044 28868 46096
rect 29460 46044 29512 46096
rect 35992 46044 36044 46096
rect 27528 45976 27580 46028
rect 21916 45951 21968 45960
rect 21916 45917 21925 45951
rect 21925 45917 21959 45951
rect 21959 45917 21968 45951
rect 21916 45908 21968 45917
rect 22376 45951 22428 45960
rect 22376 45917 22385 45951
rect 22385 45917 22419 45951
rect 22419 45917 22428 45951
rect 22376 45908 22428 45917
rect 22836 45908 22888 45960
rect 20720 45883 20772 45892
rect 20720 45849 20729 45883
rect 20729 45849 20763 45883
rect 20763 45849 20772 45883
rect 20720 45840 20772 45849
rect 22652 45840 22704 45892
rect 17868 45772 17920 45824
rect 19708 45772 19760 45824
rect 20352 45772 20404 45824
rect 23940 45951 23992 45960
rect 23940 45917 23949 45951
rect 23949 45917 23983 45951
rect 23983 45917 23992 45951
rect 23940 45908 23992 45917
rect 24768 45908 24820 45960
rect 25044 45908 25096 45960
rect 26700 45951 26752 45960
rect 23020 45840 23072 45892
rect 26700 45917 26709 45951
rect 26709 45917 26743 45951
rect 26743 45917 26752 45951
rect 26700 45908 26752 45917
rect 26792 45951 26844 45960
rect 26792 45917 26801 45951
rect 26801 45917 26835 45951
rect 26835 45917 26844 45951
rect 26792 45908 26844 45917
rect 27436 45908 27488 45960
rect 28724 45976 28776 46028
rect 28908 45908 28960 45960
rect 30564 45976 30616 46028
rect 31484 46019 31536 46028
rect 31484 45985 31493 46019
rect 31493 45985 31527 46019
rect 31527 45985 31536 46019
rect 31484 45976 31536 45985
rect 30196 45951 30248 45960
rect 30196 45917 30205 45951
rect 30205 45917 30239 45951
rect 30239 45917 30248 45951
rect 30196 45908 30248 45917
rect 30288 45951 30340 45960
rect 30288 45917 30297 45951
rect 30297 45917 30331 45951
rect 30331 45917 30340 45951
rect 31760 45976 31812 46028
rect 32036 46019 32088 46028
rect 32036 45985 32045 46019
rect 32045 45985 32079 46019
rect 32079 45985 32088 46019
rect 32036 45976 32088 45985
rect 35348 46019 35400 46028
rect 35348 45985 35357 46019
rect 35357 45985 35391 46019
rect 35391 45985 35400 46019
rect 35348 45976 35400 45985
rect 35532 46019 35584 46028
rect 35532 45985 35541 46019
rect 35541 45985 35575 46019
rect 35575 45985 35584 46019
rect 35532 45976 35584 45985
rect 37740 46087 37792 46096
rect 37740 46053 37749 46087
rect 37749 46053 37783 46087
rect 37783 46053 37792 46087
rect 37740 46044 37792 46053
rect 38200 46044 38252 46096
rect 30288 45908 30340 45917
rect 28540 45840 28592 45892
rect 23296 45772 23348 45824
rect 24860 45772 24912 45824
rect 26792 45772 26844 45824
rect 29000 45772 29052 45824
rect 29644 45772 29696 45824
rect 33876 45951 33928 45960
rect 33876 45917 33885 45951
rect 33885 45917 33919 45951
rect 33919 45917 33928 45951
rect 35624 45951 35676 45960
rect 33876 45908 33928 45917
rect 35624 45917 35633 45951
rect 35633 45917 35667 45951
rect 35667 45917 35676 45951
rect 35624 45908 35676 45917
rect 36176 45908 36228 45960
rect 36452 45951 36504 45960
rect 36452 45917 36461 45951
rect 36461 45917 36495 45951
rect 36495 45917 36504 45951
rect 36452 45908 36504 45917
rect 36544 45951 36596 45960
rect 36544 45917 36553 45951
rect 36553 45917 36587 45951
rect 36587 45917 36596 45951
rect 36728 45951 36780 45960
rect 36544 45908 36596 45917
rect 36728 45917 36737 45951
rect 36737 45917 36771 45951
rect 36771 45917 36780 45951
rect 36728 45908 36780 45917
rect 36820 45951 36872 45960
rect 36820 45917 36829 45951
rect 36829 45917 36863 45951
rect 36863 45917 36872 45951
rect 36820 45908 36872 45917
rect 38108 45908 38160 45960
rect 39120 45976 39172 46028
rect 39948 45976 40000 46028
rect 39488 45951 39540 45960
rect 37648 45840 37700 45892
rect 39488 45917 39497 45951
rect 39497 45917 39531 45951
rect 39531 45917 39540 45951
rect 39488 45908 39540 45917
rect 40776 45908 40828 45960
rect 40316 45840 40368 45892
rect 32680 45772 32732 45824
rect 34152 45772 34204 45824
rect 35808 45772 35860 45824
rect 36544 45772 36596 45824
rect 37004 45772 37056 45824
rect 39028 45772 39080 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 17224 45568 17276 45620
rect 19432 45568 19484 45620
rect 17868 45500 17920 45552
rect 18420 45500 18472 45552
rect 18328 45475 18380 45484
rect 18328 45441 18337 45475
rect 18337 45441 18371 45475
rect 18371 45441 18380 45475
rect 18328 45432 18380 45441
rect 20720 45500 20772 45552
rect 20168 45475 20220 45484
rect 9680 45364 9732 45416
rect 20168 45441 20177 45475
rect 20177 45441 20211 45475
rect 20211 45441 20220 45475
rect 20168 45432 20220 45441
rect 20444 45475 20496 45484
rect 20444 45441 20453 45475
rect 20453 45441 20487 45475
rect 20487 45441 20496 45475
rect 23020 45568 23072 45620
rect 20444 45432 20496 45441
rect 21364 45432 21416 45484
rect 23848 45500 23900 45552
rect 24860 45568 24912 45620
rect 26332 45568 26384 45620
rect 26884 45568 26936 45620
rect 27988 45568 28040 45620
rect 22284 45364 22336 45416
rect 22744 45475 22796 45484
rect 22744 45441 22753 45475
rect 22753 45441 22787 45475
rect 22787 45441 22796 45475
rect 22744 45432 22796 45441
rect 22468 45364 22520 45416
rect 23572 45432 23624 45484
rect 23756 45364 23808 45416
rect 29000 45500 29052 45552
rect 29276 45568 29328 45620
rect 29828 45568 29880 45620
rect 31668 45568 31720 45620
rect 33324 45568 33376 45620
rect 34612 45568 34664 45620
rect 30564 45543 30616 45552
rect 30564 45509 30573 45543
rect 30573 45509 30607 45543
rect 30607 45509 30616 45543
rect 30564 45500 30616 45509
rect 33140 45500 33192 45552
rect 24860 45475 24912 45484
rect 24860 45441 24869 45475
rect 24869 45441 24903 45475
rect 24903 45441 24912 45475
rect 24860 45432 24912 45441
rect 27344 45432 27396 45484
rect 27620 45432 27672 45484
rect 27988 45475 28040 45484
rect 27988 45441 27997 45475
rect 27997 45441 28031 45475
rect 28031 45441 28040 45475
rect 27988 45432 28040 45441
rect 28724 45432 28776 45484
rect 29184 45475 29236 45484
rect 29184 45441 29193 45475
rect 29193 45441 29236 45475
rect 29184 45432 29236 45441
rect 26516 45364 26568 45416
rect 30288 45475 30340 45484
rect 30288 45441 30297 45475
rect 30297 45441 30331 45475
rect 30331 45441 30340 45475
rect 30288 45432 30340 45441
rect 30748 45432 30800 45484
rect 32312 45432 32364 45484
rect 34520 45500 34572 45552
rect 36452 45568 36504 45620
rect 37832 45568 37884 45620
rect 39212 45568 39264 45620
rect 42708 45611 42760 45620
rect 42708 45577 42717 45611
rect 42717 45577 42751 45611
rect 42751 45577 42760 45611
rect 42708 45568 42760 45577
rect 33600 45475 33652 45484
rect 31760 45364 31812 45416
rect 32128 45364 32180 45416
rect 33600 45441 33609 45475
rect 33609 45441 33643 45475
rect 33643 45441 33652 45475
rect 33600 45432 33652 45441
rect 33232 45364 33284 45416
rect 33968 45364 34020 45416
rect 34152 45407 34204 45416
rect 34152 45373 34161 45407
rect 34161 45373 34195 45407
rect 34195 45373 34204 45407
rect 34152 45364 34204 45373
rect 34244 45364 34296 45416
rect 35440 45500 35492 45552
rect 36176 45475 36228 45484
rect 36176 45441 36185 45475
rect 36185 45441 36219 45475
rect 36219 45441 36228 45475
rect 36636 45475 36688 45484
rect 36176 45432 36228 45441
rect 36636 45441 36645 45475
rect 36645 45441 36679 45475
rect 36679 45441 36688 45475
rect 36636 45432 36688 45441
rect 38016 45432 38068 45484
rect 38292 45475 38344 45484
rect 38292 45441 38300 45475
rect 38300 45441 38334 45475
rect 38334 45441 38344 45475
rect 38292 45432 38344 45441
rect 38568 45432 38620 45484
rect 38660 45432 38712 45484
rect 40132 45432 40184 45484
rect 40316 45432 40368 45484
rect 35624 45364 35676 45416
rect 35900 45364 35952 45416
rect 37464 45364 37516 45416
rect 37924 45407 37976 45416
rect 37924 45373 37933 45407
rect 37933 45373 37967 45407
rect 37967 45373 37976 45407
rect 37924 45364 37976 45373
rect 38108 45364 38160 45416
rect 25872 45296 25924 45348
rect 27344 45296 27396 45348
rect 27620 45296 27672 45348
rect 29092 45296 29144 45348
rect 30196 45339 30248 45348
rect 30196 45305 30205 45339
rect 30205 45305 30239 45339
rect 30239 45305 30248 45339
rect 30196 45296 30248 45305
rect 36728 45339 36780 45348
rect 36728 45305 36737 45339
rect 36737 45305 36771 45339
rect 36771 45305 36780 45339
rect 36728 45296 36780 45305
rect 37188 45296 37240 45348
rect 40408 45296 40460 45348
rect 18972 45228 19024 45280
rect 25780 45228 25832 45280
rect 26332 45228 26384 45280
rect 26516 45271 26568 45280
rect 26516 45237 26525 45271
rect 26525 45237 26559 45271
rect 26559 45237 26568 45271
rect 26516 45228 26568 45237
rect 27804 45228 27856 45280
rect 28632 45228 28684 45280
rect 29184 45228 29236 45280
rect 29736 45228 29788 45280
rect 31024 45228 31076 45280
rect 32404 45271 32456 45280
rect 32404 45237 32413 45271
rect 32413 45237 32447 45271
rect 32447 45237 32456 45271
rect 32404 45228 32456 45237
rect 32588 45228 32640 45280
rect 35532 45228 35584 45280
rect 38384 45271 38436 45280
rect 38384 45237 38393 45271
rect 38393 45237 38427 45271
rect 38427 45237 38436 45271
rect 38384 45228 38436 45237
rect 39028 45228 39080 45280
rect 41144 45228 41196 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 20536 45024 20588 45076
rect 23572 45024 23624 45076
rect 20168 44956 20220 45008
rect 23664 44956 23716 45008
rect 18696 44863 18748 44872
rect 18696 44829 18705 44863
rect 18705 44829 18739 44863
rect 18739 44829 18748 44863
rect 18696 44820 18748 44829
rect 19984 44863 20036 44872
rect 19984 44829 19993 44863
rect 19993 44829 20027 44863
rect 20027 44829 20036 44863
rect 19984 44820 20036 44829
rect 20996 44820 21048 44872
rect 21456 44863 21508 44872
rect 21456 44829 21465 44863
rect 21465 44829 21499 44863
rect 21499 44829 21508 44863
rect 21456 44820 21508 44829
rect 22376 44863 22428 44872
rect 22376 44829 22385 44863
rect 22385 44829 22419 44863
rect 22419 44829 22428 44863
rect 22376 44820 22428 44829
rect 25044 44888 25096 44940
rect 20812 44752 20864 44804
rect 22468 44752 22520 44804
rect 23756 44863 23808 44872
rect 23756 44829 23765 44863
rect 23765 44829 23799 44863
rect 23799 44829 23808 44863
rect 23756 44820 23808 44829
rect 24032 44863 24084 44872
rect 24032 44829 24041 44863
rect 24041 44829 24075 44863
rect 24075 44829 24084 44863
rect 24584 44863 24636 44872
rect 24032 44820 24084 44829
rect 24584 44829 24593 44863
rect 24593 44829 24627 44863
rect 24627 44829 24636 44863
rect 24584 44820 24636 44829
rect 25596 44820 25648 44872
rect 26056 44863 26108 44872
rect 26056 44829 26065 44863
rect 26065 44829 26099 44863
rect 26099 44829 26108 44863
rect 26056 44820 26108 44829
rect 26424 44820 26476 44872
rect 27344 44820 27396 44872
rect 27436 44820 27488 44872
rect 28356 44888 28408 44940
rect 27804 44863 27856 44872
rect 27804 44829 27813 44863
rect 27813 44829 27847 44863
rect 27847 44829 27856 44863
rect 27804 44820 27856 44829
rect 28632 44863 28684 44872
rect 28632 44829 28641 44863
rect 28641 44829 28675 44863
rect 28675 44829 28684 44863
rect 28632 44820 28684 44829
rect 31484 45024 31536 45076
rect 35624 45024 35676 45076
rect 30564 44931 30616 44940
rect 30564 44897 30573 44931
rect 30573 44897 30607 44931
rect 30607 44897 30616 44931
rect 30564 44888 30616 44897
rect 29000 44820 29052 44872
rect 31760 44820 31812 44872
rect 31944 44820 31996 44872
rect 33140 44888 33192 44940
rect 33600 44956 33652 45008
rect 32312 44863 32364 44872
rect 32312 44829 32321 44863
rect 32321 44829 32355 44863
rect 32355 44829 32364 44863
rect 32312 44820 32364 44829
rect 33232 44820 33284 44872
rect 33324 44820 33376 44872
rect 33784 44863 33836 44872
rect 33784 44829 33793 44863
rect 33793 44829 33827 44863
rect 33827 44829 33836 44863
rect 33784 44820 33836 44829
rect 34520 44820 34572 44872
rect 38108 45024 38160 45076
rect 38384 45024 38436 45076
rect 39212 45067 39264 45076
rect 39212 45033 39221 45067
rect 39221 45033 39255 45067
rect 39255 45033 39264 45067
rect 39212 45024 39264 45033
rect 40040 45067 40092 45076
rect 40040 45033 40049 45067
rect 40049 45033 40083 45067
rect 40083 45033 40092 45067
rect 40040 45024 40092 45033
rect 40132 45024 40184 45076
rect 40776 45024 40828 45076
rect 42708 45024 42760 45076
rect 35808 44956 35860 45008
rect 37464 44956 37516 45008
rect 38844 44956 38896 45008
rect 37004 44863 37056 44872
rect 18972 44684 19024 44736
rect 21180 44684 21232 44736
rect 25504 44795 25556 44804
rect 25504 44761 25513 44795
rect 25513 44761 25547 44795
rect 25547 44761 25556 44795
rect 25504 44752 25556 44761
rect 26884 44752 26936 44804
rect 24860 44684 24912 44736
rect 25872 44727 25924 44736
rect 25872 44693 25881 44727
rect 25881 44693 25915 44727
rect 25915 44693 25924 44727
rect 25872 44684 25924 44693
rect 25964 44684 26016 44736
rect 27712 44752 27764 44804
rect 27252 44684 27304 44736
rect 29184 44752 29236 44804
rect 33048 44684 33100 44736
rect 37004 44829 37013 44863
rect 37013 44829 37047 44863
rect 37047 44829 37056 44863
rect 37004 44820 37056 44829
rect 37188 44863 37240 44872
rect 37188 44829 37197 44863
rect 37197 44829 37231 44863
rect 37231 44829 37240 44863
rect 37188 44820 37240 44829
rect 38016 44888 38068 44940
rect 38568 44888 38620 44940
rect 38292 44863 38344 44872
rect 38292 44829 38302 44863
rect 38302 44829 38336 44863
rect 38336 44829 38344 44863
rect 38292 44820 38344 44829
rect 41144 44863 41196 44872
rect 37648 44795 37700 44804
rect 37648 44761 37657 44795
rect 37657 44761 37691 44795
rect 37691 44761 37700 44795
rect 37648 44752 37700 44761
rect 37924 44752 37976 44804
rect 38476 44752 38528 44804
rect 41144 44829 41153 44863
rect 41153 44829 41187 44863
rect 41187 44829 41196 44863
rect 41144 44820 41196 44829
rect 38660 44684 38712 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 18328 44480 18380 44532
rect 19984 44480 20036 44532
rect 22744 44480 22796 44532
rect 25504 44523 25556 44532
rect 23756 44412 23808 44464
rect 24860 44455 24912 44464
rect 18972 44387 19024 44396
rect 18972 44353 18981 44387
rect 18981 44353 19015 44387
rect 19015 44353 19024 44387
rect 18972 44344 19024 44353
rect 20076 44344 20128 44396
rect 20812 44387 20864 44396
rect 20812 44353 20821 44387
rect 20821 44353 20855 44387
rect 20855 44353 20864 44387
rect 20812 44344 20864 44353
rect 20996 44344 21048 44396
rect 22468 44387 22520 44396
rect 22468 44353 22477 44387
rect 22477 44353 22511 44387
rect 22511 44353 22520 44387
rect 22468 44344 22520 44353
rect 23112 44387 23164 44396
rect 23112 44353 23121 44387
rect 23121 44353 23155 44387
rect 23155 44353 23164 44387
rect 23112 44344 23164 44353
rect 23480 44344 23532 44396
rect 24860 44421 24869 44455
rect 24869 44421 24903 44455
rect 24903 44421 24912 44455
rect 24860 44412 24912 44421
rect 25504 44489 25513 44523
rect 25513 44489 25547 44523
rect 25547 44489 25556 44523
rect 25504 44480 25556 44489
rect 27252 44523 27304 44532
rect 27252 44489 27261 44523
rect 27261 44489 27295 44523
rect 27295 44489 27304 44523
rect 27252 44480 27304 44489
rect 27344 44480 27396 44532
rect 25504 44387 25556 44396
rect 25504 44353 25513 44387
rect 25513 44353 25547 44387
rect 25547 44353 25556 44387
rect 25504 44344 25556 44353
rect 23572 44276 23624 44328
rect 24032 44276 24084 44328
rect 25044 44276 25096 44328
rect 25872 44319 25924 44328
rect 25872 44285 25881 44319
rect 25881 44285 25915 44319
rect 25915 44285 25924 44319
rect 25872 44276 25924 44285
rect 26240 44344 26292 44396
rect 26516 44412 26568 44464
rect 27160 44455 27212 44464
rect 27160 44421 27169 44455
rect 27169 44421 27203 44455
rect 27203 44421 27212 44455
rect 27160 44412 27212 44421
rect 29276 44412 29328 44464
rect 27436 44387 27488 44396
rect 27436 44353 27445 44387
rect 27445 44353 27479 44387
rect 27479 44353 27488 44387
rect 30932 44480 30984 44532
rect 37740 44480 37792 44532
rect 38660 44523 38712 44532
rect 38660 44489 38669 44523
rect 38669 44489 38703 44523
rect 38703 44489 38712 44523
rect 38660 44480 38712 44489
rect 40132 44523 40184 44532
rect 40132 44489 40141 44523
rect 40141 44489 40175 44523
rect 40175 44489 40184 44523
rect 40132 44480 40184 44489
rect 42708 44480 42760 44532
rect 27436 44344 27488 44353
rect 29644 44387 29696 44396
rect 27712 44276 27764 44328
rect 29644 44353 29653 44387
rect 29653 44353 29687 44387
rect 29687 44353 29696 44387
rect 29644 44344 29696 44353
rect 30748 44344 30800 44396
rect 30932 44319 30984 44328
rect 30932 44285 30941 44319
rect 30941 44285 30975 44319
rect 30975 44285 30984 44319
rect 30932 44276 30984 44285
rect 19064 44208 19116 44260
rect 21456 44208 21508 44260
rect 23848 44251 23900 44260
rect 22376 44183 22428 44192
rect 22376 44149 22385 44183
rect 22385 44149 22419 44183
rect 22419 44149 22428 44183
rect 22376 44140 22428 44149
rect 23848 44217 23857 44251
rect 23857 44217 23891 44251
rect 23891 44217 23900 44251
rect 23848 44208 23900 44217
rect 32588 44412 32640 44464
rect 33784 44412 33836 44464
rect 38476 44412 38528 44464
rect 32404 44344 32456 44396
rect 33048 44344 33100 44396
rect 33968 44344 34020 44396
rect 34520 44387 34572 44396
rect 34520 44353 34529 44387
rect 34529 44353 34563 44387
rect 34563 44353 34572 44387
rect 34520 44344 34572 44353
rect 36544 44344 36596 44396
rect 37464 44387 37516 44396
rect 37464 44353 37473 44387
rect 37473 44353 37507 44387
rect 37507 44353 37516 44387
rect 37464 44344 37516 44353
rect 37648 44387 37700 44396
rect 37648 44353 37657 44387
rect 37657 44353 37691 44387
rect 37691 44353 37700 44387
rect 37648 44344 37700 44353
rect 38384 44344 38436 44396
rect 38568 44344 38620 44396
rect 39028 44387 39080 44396
rect 39028 44353 39037 44387
rect 39037 44353 39071 44387
rect 39071 44353 39080 44387
rect 39028 44344 39080 44353
rect 40040 44412 40092 44464
rect 32864 44319 32916 44328
rect 32864 44285 32873 44319
rect 32873 44285 32907 44319
rect 32907 44285 32916 44319
rect 32864 44276 32916 44285
rect 35900 44276 35952 44328
rect 37556 44183 37608 44192
rect 37556 44149 37565 44183
rect 37565 44149 37599 44183
rect 37599 44149 37608 44183
rect 37556 44140 37608 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 22100 43936 22152 43988
rect 24952 43936 25004 43988
rect 29092 43936 29144 43988
rect 29368 43936 29420 43988
rect 30932 43979 30984 43988
rect 30932 43945 30941 43979
rect 30941 43945 30975 43979
rect 30975 43945 30984 43979
rect 30932 43936 30984 43945
rect 21824 43911 21876 43920
rect 21824 43877 21833 43911
rect 21833 43877 21867 43911
rect 21867 43877 21876 43911
rect 21824 43868 21876 43877
rect 23204 43800 23256 43852
rect 26424 43868 26476 43920
rect 26700 43800 26752 43852
rect 20996 43732 21048 43784
rect 22376 43732 22428 43784
rect 23848 43732 23900 43784
rect 23480 43664 23532 43716
rect 24860 43664 24912 43716
rect 25964 43732 26016 43784
rect 27160 43775 27212 43784
rect 27160 43741 27169 43775
rect 27169 43741 27203 43775
rect 27203 43741 27212 43775
rect 27160 43732 27212 43741
rect 27620 43775 27672 43784
rect 27620 43741 27629 43775
rect 27629 43741 27663 43775
rect 27663 43741 27672 43775
rect 27620 43732 27672 43741
rect 28356 43775 28408 43784
rect 28356 43741 28365 43775
rect 28365 43741 28399 43775
rect 28399 43741 28408 43775
rect 28356 43732 28408 43741
rect 29184 43775 29236 43784
rect 29184 43741 29193 43775
rect 29193 43741 29227 43775
rect 29227 43741 29236 43775
rect 29184 43732 29236 43741
rect 31024 43775 31076 43784
rect 31024 43741 31033 43775
rect 31033 43741 31067 43775
rect 31067 43741 31076 43775
rect 31024 43732 31076 43741
rect 31668 43775 31720 43784
rect 31668 43741 31677 43775
rect 31677 43741 31711 43775
rect 31711 43741 31720 43775
rect 31668 43732 31720 43741
rect 32864 43868 32916 43920
rect 33140 43911 33192 43920
rect 33140 43877 33149 43911
rect 33149 43877 33183 43911
rect 33183 43877 33192 43911
rect 33140 43868 33192 43877
rect 34152 43936 34204 43988
rect 34520 43936 34572 43988
rect 36544 43979 36596 43988
rect 36544 43945 36553 43979
rect 36553 43945 36587 43979
rect 36587 43945 36596 43979
rect 36544 43936 36596 43945
rect 36820 43979 36872 43988
rect 36820 43945 36829 43979
rect 36829 43945 36863 43979
rect 36863 43945 36872 43979
rect 36820 43936 36872 43945
rect 38476 43936 38528 43988
rect 40132 43979 40184 43988
rect 40132 43945 40141 43979
rect 40141 43945 40175 43979
rect 40175 43945 40184 43979
rect 40132 43936 40184 43945
rect 36636 43868 36688 43920
rect 33048 43800 33100 43852
rect 25504 43664 25556 43716
rect 25688 43707 25740 43716
rect 25688 43673 25697 43707
rect 25697 43673 25731 43707
rect 25731 43673 25740 43707
rect 25688 43664 25740 43673
rect 27436 43664 27488 43716
rect 21824 43596 21876 43648
rect 22192 43596 22244 43648
rect 32864 43732 32916 43784
rect 35440 43800 35492 43852
rect 33048 43664 33100 43716
rect 34244 43732 34296 43784
rect 36820 43800 36872 43852
rect 38844 43868 38896 43920
rect 37740 43775 37792 43784
rect 37740 43741 37749 43775
rect 37749 43741 37783 43775
rect 37783 43741 37792 43775
rect 37740 43732 37792 43741
rect 38384 43732 38436 43784
rect 35992 43707 36044 43716
rect 35992 43673 36001 43707
rect 36001 43673 36035 43707
rect 36035 43673 36044 43707
rect 35992 43664 36044 43673
rect 37648 43664 37700 43716
rect 32680 43596 32732 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 22652 43392 22704 43444
rect 23572 43435 23624 43444
rect 23572 43401 23581 43435
rect 23581 43401 23615 43435
rect 23615 43401 23624 43435
rect 23572 43392 23624 43401
rect 25044 43324 25096 43376
rect 25688 43324 25740 43376
rect 26424 43392 26476 43444
rect 27620 43435 27672 43444
rect 27620 43401 27629 43435
rect 27629 43401 27663 43435
rect 27663 43401 27672 43435
rect 27620 43392 27672 43401
rect 33232 43435 33284 43444
rect 33232 43401 33241 43435
rect 33241 43401 33275 43435
rect 33275 43401 33284 43435
rect 33232 43392 33284 43401
rect 35440 43392 35492 43444
rect 35716 43435 35768 43444
rect 35716 43401 35725 43435
rect 35725 43401 35759 43435
rect 35759 43401 35768 43435
rect 35716 43392 35768 43401
rect 36820 43435 36872 43444
rect 36820 43401 36829 43435
rect 36829 43401 36863 43435
rect 36863 43401 36872 43435
rect 36820 43392 36872 43401
rect 37740 43392 37792 43444
rect 38476 43392 38528 43444
rect 38844 43392 38896 43444
rect 23112 43188 23164 43240
rect 24860 43256 24912 43308
rect 25596 43256 25648 43308
rect 26056 43324 26108 43376
rect 29276 43367 29328 43376
rect 29276 43333 29285 43367
rect 29285 43333 29319 43367
rect 29319 43333 29328 43367
rect 29276 43324 29328 43333
rect 32128 43324 32180 43376
rect 32680 43367 32732 43376
rect 32680 43333 32689 43367
rect 32689 43333 32723 43367
rect 32723 43333 32732 43367
rect 32680 43324 32732 43333
rect 26884 43256 26936 43308
rect 27252 43256 27304 43308
rect 31208 43299 31260 43308
rect 31208 43265 31217 43299
rect 31217 43265 31251 43299
rect 31251 43265 31260 43299
rect 31208 43256 31260 43265
rect 31668 43256 31720 43308
rect 32864 43256 32916 43308
rect 33508 43324 33560 43376
rect 35532 43324 35584 43376
rect 38200 43324 38252 43376
rect 33048 43256 33100 43308
rect 33416 43256 33468 43308
rect 33876 43256 33928 43308
rect 37556 43256 37608 43308
rect 29736 43163 29788 43172
rect 29736 43129 29745 43163
rect 29745 43129 29779 43163
rect 29779 43129 29788 43163
rect 29736 43120 29788 43129
rect 27436 43095 27488 43104
rect 27436 43061 27445 43095
rect 27445 43061 27479 43095
rect 27479 43061 27488 43095
rect 27436 43052 27488 43061
rect 30288 43052 30340 43104
rect 30932 43052 30984 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 26424 42848 26476 42900
rect 29184 42848 29236 42900
rect 32864 42891 32916 42900
rect 32864 42857 32873 42891
rect 32873 42857 32907 42891
rect 32907 42857 32916 42891
rect 32864 42848 32916 42857
rect 35440 42891 35492 42900
rect 35440 42857 35449 42891
rect 35449 42857 35483 42891
rect 35483 42857 35492 42891
rect 35440 42848 35492 42857
rect 22652 42780 22704 42832
rect 35532 42780 35584 42832
rect 35992 42823 36044 42832
rect 35992 42789 36001 42823
rect 36001 42789 36035 42823
rect 36035 42789 36044 42823
rect 35992 42780 36044 42789
rect 26332 42712 26384 42764
rect 27344 42712 27396 42764
rect 27528 42712 27580 42764
rect 30748 42712 30800 42764
rect 37280 42712 37332 42764
rect 38200 42712 38252 42764
rect 22192 42508 22244 42560
rect 27252 42508 27304 42560
rect 30932 42619 30984 42628
rect 30932 42585 30941 42619
rect 30941 42585 30975 42619
rect 30975 42585 30984 42619
rect 30932 42576 30984 42585
rect 29276 42508 29328 42560
rect 31760 42576 31812 42628
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 26332 42347 26384 42356
rect 26332 42313 26341 42347
rect 26341 42313 26375 42347
rect 26375 42313 26384 42347
rect 26332 42304 26384 42313
rect 27252 42347 27304 42356
rect 27252 42313 27261 42347
rect 27261 42313 27295 42347
rect 27295 42313 27304 42347
rect 27252 42304 27304 42313
rect 27528 42304 27580 42356
rect 30932 42304 30984 42356
rect 35716 42304 35768 42356
rect 35992 42347 36044 42356
rect 35992 42313 36001 42347
rect 36001 42313 36035 42347
rect 36035 42313 36044 42347
rect 35992 42304 36044 42313
rect 25872 42236 25924 42288
rect 29644 42236 29696 42288
rect 30748 42279 30800 42288
rect 30748 42245 30757 42279
rect 30757 42245 30791 42279
rect 30791 42245 30800 42279
rect 30748 42236 30800 42245
rect 37280 42236 37332 42288
rect 29276 42007 29328 42016
rect 29276 41973 29285 42007
rect 29285 41973 29319 42007
rect 29319 41973 29328 42007
rect 29276 41964 29328 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 29276 41760 29328 41812
rect 29644 41760 29696 41812
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 23020 6740 23072 6792
rect 24400 6740 24452 6792
rect 22192 6604 22244 6656
rect 24768 6604 24820 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 24492 6332 24544 6384
rect 26700 6332 26752 6384
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 22192 6264 22244 6273
rect 22284 6264 22336 6316
rect 28172 6307 28224 6316
rect 28172 6273 28181 6307
rect 28181 6273 28215 6307
rect 28215 6273 28224 6307
rect 28172 6264 28224 6273
rect 25964 6239 26016 6248
rect 25964 6205 25973 6239
rect 25973 6205 26007 6239
rect 26007 6205 26016 6239
rect 25964 6196 26016 6205
rect 25228 6171 25280 6180
rect 25228 6137 25237 6171
rect 25237 6137 25271 6171
rect 25271 6137 25280 6171
rect 25228 6128 25280 6137
rect 26516 6171 26568 6180
rect 26516 6137 26525 6171
rect 26525 6137 26559 6171
rect 26559 6137 26568 6171
rect 26516 6128 26568 6137
rect 20904 6060 20956 6112
rect 21364 6060 21416 6112
rect 22008 6103 22060 6112
rect 22008 6069 22017 6103
rect 22017 6069 22051 6103
rect 22051 6069 22060 6103
rect 22008 6060 22060 6069
rect 23388 6060 23440 6112
rect 24676 6060 24728 6112
rect 27436 6060 27488 6112
rect 27804 6060 27856 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 25964 5899 26016 5908
rect 25964 5865 25973 5899
rect 25973 5865 26007 5899
rect 26007 5865 26016 5899
rect 25964 5856 26016 5865
rect 26700 5899 26752 5908
rect 26700 5865 26709 5899
rect 26709 5865 26743 5899
rect 26743 5865 26752 5899
rect 26700 5856 26752 5865
rect 21916 5831 21968 5840
rect 21916 5797 21925 5831
rect 21925 5797 21959 5831
rect 21959 5797 21968 5831
rect 21916 5788 21968 5797
rect 23848 5831 23900 5840
rect 23848 5797 23857 5831
rect 23857 5797 23891 5831
rect 23891 5797 23900 5831
rect 23848 5788 23900 5797
rect 27988 5831 28040 5840
rect 27988 5797 27997 5831
rect 27997 5797 28031 5831
rect 28031 5797 28040 5831
rect 27988 5788 28040 5797
rect 21364 5763 21416 5772
rect 21364 5729 21373 5763
rect 21373 5729 21407 5763
rect 21407 5729 21416 5763
rect 21364 5720 21416 5729
rect 24676 5763 24728 5772
rect 24676 5729 24685 5763
rect 24685 5729 24719 5763
rect 24719 5729 24728 5763
rect 24676 5720 24728 5729
rect 24952 5763 25004 5772
rect 24952 5729 24961 5763
rect 24961 5729 24995 5763
rect 24995 5729 25004 5763
rect 24952 5720 25004 5729
rect 27436 5763 27488 5772
rect 27436 5729 27445 5763
rect 27445 5729 27479 5763
rect 27479 5729 27488 5763
rect 27436 5720 27488 5729
rect 20628 5695 20680 5704
rect 20628 5661 20637 5695
rect 20637 5661 20671 5695
rect 20671 5661 20680 5695
rect 20628 5652 20680 5661
rect 25688 5652 25740 5704
rect 23388 5627 23440 5636
rect 23388 5593 23397 5627
rect 23397 5593 23431 5627
rect 23431 5593 23440 5627
rect 23388 5584 23440 5593
rect 24768 5627 24820 5636
rect 24768 5593 24777 5627
rect 24777 5593 24811 5627
rect 24811 5593 24820 5627
rect 24768 5584 24820 5593
rect 27528 5627 27580 5636
rect 27528 5593 27537 5627
rect 27537 5593 27571 5627
rect 27571 5593 27580 5627
rect 27528 5584 27580 5593
rect 20812 5516 20864 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 24492 5355 24544 5364
rect 22192 5244 22244 5296
rect 23020 5287 23072 5296
rect 19340 5176 19392 5228
rect 20812 5219 20864 5228
rect 20812 5185 20821 5219
rect 20821 5185 20855 5219
rect 20855 5185 20864 5219
rect 20812 5176 20864 5185
rect 20352 5108 20404 5160
rect 22284 5176 22336 5228
rect 23020 5253 23029 5287
rect 23029 5253 23063 5287
rect 23063 5253 23072 5287
rect 23020 5244 23072 5253
rect 24492 5321 24501 5355
rect 24501 5321 24535 5355
rect 24535 5321 24544 5355
rect 24492 5312 24544 5321
rect 25780 5244 25832 5296
rect 27804 5287 27856 5296
rect 27804 5253 27813 5287
rect 27813 5253 27847 5287
rect 27847 5253 27856 5287
rect 27804 5244 27856 5253
rect 23756 5176 23808 5228
rect 24400 5219 24452 5228
rect 24400 5185 24409 5219
rect 24409 5185 24443 5219
rect 24443 5185 24452 5219
rect 24400 5176 24452 5185
rect 27620 5151 27672 5160
rect 27620 5117 27629 5151
rect 27629 5117 27663 5151
rect 27663 5117 27672 5151
rect 27620 5108 27672 5117
rect 20628 5083 20680 5092
rect 20628 5049 20637 5083
rect 20637 5049 20671 5083
rect 20671 5049 20680 5083
rect 20628 5040 20680 5049
rect 22284 5083 22336 5092
rect 22284 5049 22293 5083
rect 22293 5049 22327 5083
rect 22327 5049 22336 5083
rect 22284 5040 22336 5049
rect 23572 5083 23624 5092
rect 23572 5049 23581 5083
rect 23581 5049 23615 5083
rect 23615 5049 23624 5083
rect 23572 5040 23624 5049
rect 26332 5083 26384 5092
rect 26332 5049 26341 5083
rect 26341 5049 26375 5083
rect 26375 5049 26384 5083
rect 26332 5040 26384 5049
rect 19432 5015 19484 5024
rect 19432 4981 19441 5015
rect 19441 4981 19475 5015
rect 19475 4981 19484 5015
rect 19432 4972 19484 4981
rect 20076 5015 20128 5024
rect 20076 4981 20085 5015
rect 20085 4981 20119 5015
rect 20119 4981 20128 5015
rect 20076 4972 20128 4981
rect 29092 5015 29144 5024
rect 29092 4981 29101 5015
rect 29101 4981 29135 5015
rect 29135 4981 29144 5015
rect 29092 4972 29144 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19984 4632 20036 4684
rect 18052 4607 18104 4616
rect 18052 4573 18061 4607
rect 18061 4573 18095 4607
rect 18095 4573 18104 4607
rect 18052 4564 18104 4573
rect 23756 4768 23808 4820
rect 25780 4811 25832 4820
rect 25780 4777 25789 4811
rect 25789 4777 25823 4811
rect 25823 4777 25832 4811
rect 25780 4768 25832 4777
rect 27528 4811 27580 4820
rect 27528 4777 27537 4811
rect 27537 4777 27571 4811
rect 27571 4777 27580 4811
rect 27528 4768 27580 4777
rect 20720 4700 20772 4752
rect 20904 4675 20956 4684
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 20904 4632 20956 4641
rect 22008 4700 22060 4752
rect 23296 4675 23348 4684
rect 23296 4641 23305 4675
rect 23305 4641 23339 4675
rect 23339 4641 23348 4675
rect 23296 4632 23348 4641
rect 20352 4564 20404 4616
rect 22008 4564 22060 4616
rect 25688 4700 25740 4752
rect 25688 4607 25740 4616
rect 25688 4573 25697 4607
rect 25697 4573 25731 4607
rect 25731 4573 25740 4607
rect 25688 4564 25740 4573
rect 28816 4675 28868 4684
rect 28816 4641 28825 4675
rect 28825 4641 28859 4675
rect 28859 4641 28868 4675
rect 28816 4632 28868 4641
rect 29092 4675 29144 4684
rect 29092 4641 29101 4675
rect 29101 4641 29135 4675
rect 29135 4641 29144 4675
rect 29092 4632 29144 4641
rect 20076 4496 20128 4548
rect 21640 4496 21692 4548
rect 20168 4428 20220 4480
rect 27896 4564 27948 4616
rect 28172 4564 28224 4616
rect 30380 4428 30432 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 20168 4156 20220 4208
rect 20812 4156 20864 4208
rect 24308 4199 24360 4208
rect 24308 4165 24317 4199
rect 24317 4165 24351 4199
rect 24351 4165 24360 4199
rect 24308 4156 24360 4165
rect 25504 4199 25556 4208
rect 25504 4165 25513 4199
rect 25513 4165 25547 4199
rect 25547 4165 25556 4199
rect 25504 4156 25556 4165
rect 27344 4199 27396 4208
rect 27344 4165 27353 4199
rect 27353 4165 27387 4199
rect 27387 4165 27396 4199
rect 27344 4156 27396 4165
rect 30472 4088 30524 4140
rect 21088 4063 21140 4072
rect 21088 4029 21097 4063
rect 21097 4029 21131 4063
rect 21131 4029 21140 4063
rect 21088 4020 21140 4029
rect 22192 4020 22244 4072
rect 23388 4020 23440 4072
rect 26056 4063 26108 4072
rect 26056 4029 26065 4063
rect 26065 4029 26099 4063
rect 26099 4029 26108 4063
rect 26056 4020 26108 4029
rect 26608 4020 26660 4072
rect 27436 4020 27488 4072
rect 29092 4020 29144 4072
rect 24676 3952 24728 4004
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 16120 3927 16172 3936
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 17224 3927 17276 3936
rect 17224 3893 17233 3927
rect 17233 3893 17267 3927
rect 17267 3893 17276 3927
rect 17224 3884 17276 3893
rect 18880 3884 18932 3936
rect 20720 3884 20772 3936
rect 20904 3884 20956 3936
rect 23756 3884 23808 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 18144 3680 18196 3732
rect 21732 3680 21784 3732
rect 23388 3723 23440 3732
rect 23388 3689 23397 3723
rect 23397 3689 23431 3723
rect 23431 3689 23440 3723
rect 23388 3680 23440 3689
rect 24308 3680 24360 3732
rect 25504 3680 25556 3732
rect 16948 3612 17000 3664
rect 20168 3612 20220 3664
rect 15844 3544 15896 3596
rect 20260 3544 20312 3596
rect 4160 3476 4212 3528
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 11796 3476 11848 3528
rect 12532 3476 12584 3528
rect 13084 3476 13136 3528
rect 13636 3519 13688 3528
rect 13636 3485 13645 3519
rect 13645 3485 13679 3519
rect 13679 3485 13688 3519
rect 13636 3476 13688 3485
rect 16396 3476 16448 3528
rect 18604 3476 18656 3528
rect 18696 3519 18748 3528
rect 18696 3485 18705 3519
rect 18705 3485 18739 3519
rect 18739 3485 18748 3519
rect 18696 3476 18748 3485
rect 19340 3476 19392 3528
rect 20904 3519 20956 3528
rect 20904 3485 20913 3519
rect 20913 3485 20947 3519
rect 20947 3485 20956 3519
rect 20904 3476 20956 3485
rect 18512 3408 18564 3460
rect 20352 3408 20404 3460
rect 20628 3408 20680 3460
rect 21732 3451 21784 3460
rect 21732 3417 21741 3451
rect 21741 3417 21775 3451
rect 21775 3417 21784 3451
rect 21732 3408 21784 3417
rect 22468 3408 22520 3460
rect 23756 3476 23808 3528
rect 24216 3544 24268 3596
rect 27160 3544 27212 3596
rect 28264 3587 28316 3596
rect 28264 3553 28273 3587
rect 28273 3553 28307 3587
rect 28307 3553 28316 3587
rect 28264 3544 28316 3553
rect 25688 3476 25740 3528
rect 30472 3612 30524 3664
rect 31392 3612 31444 3664
rect 32956 3612 33008 3664
rect 36820 3612 36872 3664
rect 30196 3544 30248 3596
rect 34796 3544 34848 3596
rect 30012 3476 30064 3528
rect 31116 3476 31168 3528
rect 31852 3476 31904 3528
rect 32404 3476 32456 3528
rect 34336 3476 34388 3528
rect 35716 3476 35768 3528
rect 36268 3476 36320 3528
rect 37648 3476 37700 3528
rect 38200 3476 38252 3528
rect 39580 3476 39632 3528
rect 40408 3476 40460 3528
rect 40960 3476 41012 3528
rect 41512 3476 41564 3528
rect 42892 3519 42944 3528
rect 42892 3485 42901 3519
rect 42901 3485 42935 3519
rect 42935 3485 42944 3519
rect 42892 3476 42944 3485
rect 43168 3476 43220 3528
rect 44824 3476 44876 3528
rect 45652 3476 45704 3528
rect 46480 3519 46532 3528
rect 46480 3485 46489 3519
rect 46489 3485 46523 3519
rect 46523 3485 46532 3519
rect 46480 3476 46532 3485
rect 46756 3476 46808 3528
rect 47308 3476 47360 3528
rect 18788 3383 18840 3392
rect 18788 3349 18797 3383
rect 18797 3349 18831 3383
rect 18831 3349 18840 3383
rect 18788 3340 18840 3349
rect 19340 3340 19392 3392
rect 20812 3340 20864 3392
rect 24124 3340 24176 3392
rect 25044 3408 25096 3460
rect 28172 3408 28224 3460
rect 28356 3340 28408 3392
rect 30748 3408 30800 3460
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 18144 3179 18196 3188
rect 18144 3145 18153 3179
rect 18153 3145 18187 3179
rect 18187 3145 18196 3179
rect 18144 3136 18196 3145
rect 22008 3136 22060 3188
rect 18788 3068 18840 3120
rect 20904 3068 20956 3120
rect 24124 3111 24176 3120
rect 24124 3077 24133 3111
rect 24133 3077 24167 3111
rect 24167 3077 24176 3111
rect 24124 3068 24176 3077
rect 24860 3068 24912 3120
rect 27712 3111 27764 3120
rect 27712 3077 27721 3111
rect 27721 3077 27755 3111
rect 27755 3077 27764 3111
rect 27712 3068 27764 3077
rect 30288 3136 30340 3188
rect 30012 3068 30064 3120
rect 18696 3000 18748 3052
rect 19340 3000 19392 3052
rect 20168 3043 20220 3052
rect 20168 3009 20177 3043
rect 20177 3009 20211 3043
rect 20211 3009 20220 3043
rect 20168 3000 20220 3009
rect 26608 3043 26660 3052
rect 26608 3009 26617 3043
rect 26617 3009 26651 3043
rect 26651 3009 26660 3043
rect 26608 3000 26660 3009
rect 30748 3043 30800 3052
rect 30748 3009 30757 3043
rect 30757 3009 30791 3043
rect 30791 3009 30800 3043
rect 30748 3000 30800 3009
rect 31392 3043 31444 3052
rect 31392 3009 31401 3043
rect 31401 3009 31435 3043
rect 31435 3009 31444 3043
rect 31392 3000 31444 3009
rect 32680 3000 32732 3052
rect 5448 2932 5500 2984
rect 7932 2932 7984 2984
rect 9864 2932 9916 2984
rect 15292 2932 15344 2984
rect 17500 2932 17552 2984
rect 18604 2932 18656 2984
rect 21364 2975 21416 2984
rect 21364 2941 21373 2975
rect 21373 2941 21407 2975
rect 21407 2941 21416 2975
rect 21364 2932 21416 2941
rect 4896 2864 4948 2916
rect 6276 2864 6328 2916
rect 3148 2796 3200 2848
rect 3884 2796 3936 2848
rect 6552 2796 6604 2848
rect 8760 2864 8812 2916
rect 11244 2864 11296 2916
rect 13360 2864 13412 2916
rect 14464 2864 14516 2916
rect 16672 2864 16724 2916
rect 9036 2796 9088 2848
rect 10692 2796 10744 2848
rect 12072 2796 12124 2848
rect 13912 2796 13964 2848
rect 18328 2864 18380 2916
rect 22744 2932 22796 2984
rect 24400 2975 24452 2984
rect 20536 2796 20588 2848
rect 22100 2796 22152 2848
rect 24400 2941 24409 2975
rect 24409 2941 24443 2975
rect 24443 2941 24452 2975
rect 24400 2932 24452 2941
rect 24492 2932 24544 2984
rect 25504 2975 25556 2984
rect 25504 2941 25513 2975
rect 25513 2941 25547 2975
rect 25547 2941 25556 2975
rect 25504 2932 25556 2941
rect 26884 2932 26936 2984
rect 27804 2975 27856 2984
rect 27804 2941 27813 2975
rect 27813 2941 27847 2975
rect 27847 2941 27856 2975
rect 27804 2932 27856 2941
rect 28540 2975 28592 2984
rect 28540 2941 28549 2975
rect 28549 2941 28583 2975
rect 28583 2941 28592 2975
rect 28540 2932 28592 2941
rect 29368 2932 29420 2984
rect 31024 2932 31076 2984
rect 32128 2932 32180 2984
rect 34060 2932 34112 2984
rect 37096 2932 37148 2984
rect 38752 2932 38804 2984
rect 40684 2932 40736 2984
rect 42616 2932 42668 2984
rect 44548 2932 44600 2984
rect 31576 2864 31628 2916
rect 33508 2864 33560 2916
rect 35348 2864 35400 2916
rect 37924 2864 37976 2916
rect 30748 2796 30800 2848
rect 35992 2796 36044 2848
rect 39028 2796 39080 2848
rect 40132 2796 40184 2848
rect 42064 2796 42116 2848
rect 43444 2796 43496 2848
rect 43996 2796 44048 2848
rect 45376 2796 45428 2848
rect 45928 2796 45980 2848
rect 47032 2796 47084 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 19156 2592 19208 2644
rect 7104 2524 7156 2576
rect 9588 2524 9640 2576
rect 11520 2524 11572 2576
rect 14188 2524 14240 2576
rect 20628 2592 20680 2644
rect 22100 2592 22152 2644
rect 24492 2592 24544 2644
rect 27344 2592 27396 2644
rect 27804 2635 27856 2644
rect 27804 2601 27813 2635
rect 27813 2601 27847 2635
rect 27847 2601 27856 2635
rect 27804 2592 27856 2601
rect 28356 2592 28408 2644
rect 30288 2592 30340 2644
rect 31024 2635 31076 2644
rect 31024 2601 31033 2635
rect 31033 2601 31067 2635
rect 31067 2601 31076 2635
rect 31024 2592 31076 2601
rect 20904 2524 20956 2576
rect 3516 2456 3568 2508
rect 8208 2456 8260 2508
rect 10416 2456 10468 2508
rect 12808 2456 12860 2508
rect 14740 2456 14792 2508
rect 17776 2456 17828 2508
rect 23020 2499 23072 2508
rect 23020 2465 23029 2499
rect 23029 2465 23063 2499
rect 23063 2465 23072 2499
rect 23020 2456 23072 2465
rect 24860 2456 24912 2508
rect 27712 2524 27764 2576
rect 28172 2524 28224 2576
rect 29920 2524 29972 2576
rect 33232 2524 33284 2576
rect 35440 2524 35492 2576
rect 38476 2524 38528 2576
rect 42340 2524 42392 2576
rect 45100 2524 45152 2576
rect 25780 2499 25832 2508
rect 25780 2465 25789 2499
rect 25789 2465 25823 2499
rect 25823 2465 25832 2499
rect 25780 2456 25832 2465
rect 31300 2456 31352 2508
rect 34612 2456 34664 2508
rect 37372 2456 37424 2508
rect 39304 2456 39356 2508
rect 41236 2456 41288 2508
rect 43720 2456 43772 2508
rect 2596 2388 2648 2440
rect 4620 2388 4672 2440
rect 5724 2388 5776 2440
rect 12256 2388 12308 2440
rect 15568 2388 15620 2440
rect 7380 2320 7432 2372
rect 17408 2320 17460 2372
rect 19340 2388 19392 2440
rect 25044 2388 25096 2440
rect 27896 2388 27948 2440
rect 31392 2388 31444 2440
rect 22008 2320 22060 2372
rect 20812 2252 20864 2304
rect 30472 2320 30524 2372
rect 33784 2388 33836 2440
rect 36544 2388 36596 2440
rect 39856 2388 39908 2440
rect 41788 2388 41840 2440
rect 44272 2320 44324 2372
rect 46204 2388 46256 2440
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 17408 1844 17460 1896
rect 19984 1844 20036 1896
<< metal2 >>
rect 3974 49200 4030 50000
rect 4342 49200 4398 50000
rect 4710 49200 4766 50000
rect 5078 49200 5134 50000
rect 5446 49200 5502 50000
rect 5814 49200 5870 50000
rect 6182 49314 6238 50000
rect 6012 49286 6238 49314
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4724 47258 4752 49200
rect 5092 47598 5120 49200
rect 5080 47592 5132 47598
rect 5080 47534 5132 47540
rect 5828 47258 5856 49200
rect 6012 47258 6040 49286
rect 6182 49200 6238 49286
rect 6550 49200 6606 50000
rect 6918 49200 6974 50000
rect 7286 49314 7342 50000
rect 7116 49286 7342 49314
rect 4712 47252 4764 47258
rect 4712 47194 4764 47200
rect 5816 47252 5868 47258
rect 5816 47194 5868 47200
rect 6000 47252 6052 47258
rect 6000 47194 6052 47200
rect 6932 46578 6960 49200
rect 7116 47258 7144 49286
rect 7286 49200 7342 49286
rect 7654 49200 7710 50000
rect 8022 49314 8078 50000
rect 7760 49286 8078 49314
rect 7760 47258 7788 49286
rect 8022 49200 8078 49286
rect 8390 49200 8446 50000
rect 8758 49200 8814 50000
rect 9126 49200 9182 50000
rect 9494 49200 9550 50000
rect 9862 49200 9918 50000
rect 10230 49200 10286 50000
rect 10598 49314 10654 50000
rect 10336 49286 10654 49314
rect 8404 47258 8432 49200
rect 9140 47258 9168 49200
rect 7104 47252 7156 47258
rect 7104 47194 7156 47200
rect 7748 47252 7800 47258
rect 7748 47194 7800 47200
rect 8392 47252 8444 47258
rect 8392 47194 8444 47200
rect 9128 47252 9180 47258
rect 9128 47194 9180 47200
rect 6920 46572 6972 46578
rect 6920 46514 6972 46520
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 9508 46209 9536 49200
rect 10244 47258 10272 49200
rect 10232 47252 10284 47258
rect 10232 47194 10284 47200
rect 9494 46200 9550 46209
rect 9494 46135 9550 46144
rect 10336 45554 10364 49286
rect 10598 49200 10654 49286
rect 10966 49200 11022 50000
rect 11334 49314 11390 50000
rect 11164 49286 11390 49314
rect 11164 47258 11192 49286
rect 11334 49200 11390 49286
rect 11702 49200 11758 50000
rect 12070 49200 12126 50000
rect 12438 49200 12494 50000
rect 12806 49200 12862 50000
rect 13174 49200 13230 50000
rect 13542 49200 13598 50000
rect 13910 49200 13966 50000
rect 14278 49200 14334 50000
rect 14646 49200 14702 50000
rect 15014 49200 15070 50000
rect 15382 49200 15438 50000
rect 15750 49200 15806 50000
rect 16118 49200 16174 50000
rect 16486 49200 16542 50000
rect 16854 49200 16910 50000
rect 17222 49200 17278 50000
rect 17590 49200 17646 50000
rect 17958 49200 18014 50000
rect 18326 49200 18382 50000
rect 18694 49200 18750 50000
rect 19062 49200 19118 50000
rect 19430 49200 19486 50000
rect 19798 49200 19854 50000
rect 20166 49314 20222 50000
rect 20534 49314 20590 50000
rect 19904 49286 20222 49314
rect 11716 47462 11744 49200
rect 11704 47456 11756 47462
rect 11704 47398 11756 47404
rect 12452 47258 12480 49200
rect 11152 47252 11204 47258
rect 11152 47194 11204 47200
rect 12440 47252 12492 47258
rect 12440 47194 12492 47200
rect 12820 46102 12848 49200
rect 13556 47258 13584 49200
rect 13544 47252 13596 47258
rect 13544 47194 13596 47200
rect 13924 46374 13952 49200
rect 14660 46578 14688 49200
rect 14648 46572 14700 46578
rect 14648 46514 14700 46520
rect 15028 46442 15056 49200
rect 15764 47258 15792 49200
rect 15752 47252 15804 47258
rect 15752 47194 15804 47200
rect 16132 46918 16160 49200
rect 16868 47190 16896 49200
rect 16948 47728 17000 47734
rect 16948 47670 17000 47676
rect 16960 47190 16988 47670
rect 16856 47184 16908 47190
rect 16856 47126 16908 47132
rect 16948 47184 17000 47190
rect 16948 47126 17000 47132
rect 16120 46912 16172 46918
rect 16120 46854 16172 46860
rect 15016 46436 15068 46442
rect 15016 46378 15068 46384
rect 13912 46368 13964 46374
rect 13912 46310 13964 46316
rect 12808 46096 12860 46102
rect 12808 46038 12860 46044
rect 17236 45626 17264 49200
rect 17592 47524 17644 47530
rect 17592 47466 17644 47472
rect 17604 47190 17632 47466
rect 17972 47274 18000 49200
rect 17972 47246 18092 47274
rect 17592 47184 17644 47190
rect 17592 47126 17644 47132
rect 17960 46980 18012 46986
rect 17960 46922 18012 46928
rect 17972 46578 18000 46922
rect 17960 46572 18012 46578
rect 17960 46514 18012 46520
rect 18064 46510 18092 47246
rect 18340 46646 18368 49200
rect 18880 47660 18932 47666
rect 18880 47602 18932 47608
rect 18892 47190 18920 47602
rect 19076 47258 19104 49200
rect 19444 47802 19472 49200
rect 19432 47796 19484 47802
rect 19432 47738 19484 47744
rect 19064 47252 19116 47258
rect 19064 47194 19116 47200
rect 18880 47184 18932 47190
rect 18880 47126 18932 47132
rect 19340 47184 19392 47190
rect 19340 47126 19392 47132
rect 19064 47048 19116 47054
rect 19064 46990 19116 46996
rect 18512 46912 18564 46918
rect 18512 46854 18564 46860
rect 18328 46640 18380 46646
rect 18328 46582 18380 46588
rect 18052 46504 18104 46510
rect 18052 46446 18104 46452
rect 18524 46170 18552 46854
rect 18972 46572 19024 46578
rect 18972 46514 19024 46520
rect 18878 46472 18934 46481
rect 18878 46407 18934 46416
rect 18512 46164 18564 46170
rect 18512 46106 18564 46112
rect 18892 45966 18920 46407
rect 18420 45960 18472 45966
rect 17866 45928 17922 45937
rect 18420 45902 18472 45908
rect 18880 45960 18932 45966
rect 18880 45902 18932 45908
rect 17866 45863 17922 45872
rect 17880 45830 17908 45863
rect 17868 45824 17920 45830
rect 17868 45766 17920 45772
rect 17224 45620 17276 45626
rect 17224 45562 17276 45568
rect 17880 45558 17908 45766
rect 18432 45558 18460 45902
rect 18696 45892 18748 45898
rect 18696 45834 18748 45840
rect 9692 45526 10364 45554
rect 17868 45552 17920 45558
rect 9692 45422 9720 45526
rect 17868 45494 17920 45500
rect 18420 45552 18472 45558
rect 18420 45494 18472 45500
rect 18328 45484 18380 45490
rect 18328 45426 18380 45432
rect 9680 45416 9732 45422
rect 9680 45358 9732 45364
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 18340 44538 18368 45426
rect 18708 44878 18736 45834
rect 18984 45286 19012 46514
rect 18972 45280 19024 45286
rect 18972 45222 19024 45228
rect 18696 44872 18748 44878
rect 18696 44814 18748 44820
rect 18972 44736 19024 44742
rect 18972 44678 19024 44684
rect 18328 44532 18380 44538
rect 18328 44474 18380 44480
rect 18984 44402 19012 44678
rect 18972 44396 19024 44402
rect 18972 44338 19024 44344
rect 19076 44266 19104 46990
rect 19352 46714 19380 47126
rect 19800 46912 19852 46918
rect 19904 46900 19932 49286
rect 20166 49200 20222 49286
rect 20272 49286 20590 49314
rect 20272 48314 20300 49286
rect 20534 49200 20590 49286
rect 20902 49200 20958 50000
rect 21270 49200 21326 50000
rect 21638 49200 21694 50000
rect 22006 49200 22062 50000
rect 22374 49200 22430 50000
rect 22742 49314 22798 50000
rect 22742 49286 22876 49314
rect 22742 49200 22798 49286
rect 19996 48286 20300 48314
rect 19996 47190 20024 48286
rect 21284 47530 21312 49200
rect 21272 47524 21324 47530
rect 21272 47466 21324 47472
rect 20076 47456 20128 47462
rect 20076 47398 20128 47404
rect 20088 47258 20116 47398
rect 20076 47252 20128 47258
rect 20076 47194 20128 47200
rect 19984 47184 20036 47190
rect 19984 47126 20036 47132
rect 21364 47116 21416 47122
rect 21364 47058 21416 47064
rect 21272 47048 21324 47054
rect 21272 46990 21324 46996
rect 19852 46872 19932 46900
rect 20076 46912 20128 46918
rect 19800 46854 19852 46860
rect 20076 46854 20128 46860
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19340 46708 19392 46714
rect 19340 46650 19392 46656
rect 19432 46708 19484 46714
rect 19892 46708 19944 46714
rect 19484 46668 19892 46696
rect 19432 46650 19484 46656
rect 19892 46650 19944 46656
rect 20088 46617 20116 46854
rect 21284 46714 21312 46990
rect 21272 46708 21324 46714
rect 21272 46650 21324 46656
rect 20444 46640 20496 46646
rect 20074 46608 20130 46617
rect 19892 46572 19944 46578
rect 20074 46543 20130 46552
rect 20258 46608 20314 46617
rect 20444 46582 20496 46588
rect 20314 46552 20392 46560
rect 20258 46543 20260 46552
rect 19892 46514 19944 46520
rect 20312 46532 20392 46552
rect 20260 46514 20312 46520
rect 19708 46504 19760 46510
rect 19760 46452 19840 46458
rect 19708 46446 19840 46452
rect 19720 46430 19840 46446
rect 19294 46368 19346 46374
rect 19346 46336 19394 46345
rect 19294 46310 19338 46316
rect 19306 46294 19338 46310
rect 19338 46271 19394 46280
rect 19708 46164 19760 46170
rect 19708 46106 19760 46112
rect 19294 46096 19346 46102
rect 19346 46064 19394 46073
rect 19294 46038 19338 46044
rect 19306 46022 19338 46038
rect 19338 45999 19394 46008
rect 19616 45960 19668 45966
rect 19432 45926 19484 45932
rect 19720 45948 19748 46106
rect 19668 45920 19748 45948
rect 19616 45902 19668 45908
rect 19432 45868 19484 45874
rect 19444 45626 19472 45868
rect 19720 45830 19748 45920
rect 19708 45824 19760 45830
rect 19812 45812 19840 46430
rect 19904 46102 19932 46514
rect 20076 46368 20128 46374
rect 20074 46336 20076 46345
rect 20128 46336 20130 46345
rect 20074 46271 20130 46280
rect 19892 46096 19944 46102
rect 20076 46096 20128 46102
rect 19892 46038 19944 46044
rect 20074 46064 20076 46073
rect 20128 46064 20130 46073
rect 20074 45999 20130 46008
rect 20168 46028 20220 46034
rect 20168 45970 20220 45976
rect 19812 45784 20116 45812
rect 19708 45766 19760 45772
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19432 45620 19484 45626
rect 19432 45562 19484 45568
rect 19984 44872 20036 44878
rect 19984 44814 20036 44820
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19996 44538 20024 44814
rect 19984 44532 20036 44538
rect 19984 44474 20036 44480
rect 20088 44402 20116 45784
rect 20180 45490 20208 45970
rect 20364 45937 20392 46532
rect 20456 46170 20484 46582
rect 20536 46572 20588 46578
rect 20536 46514 20588 46520
rect 21180 46572 21232 46578
rect 21180 46514 21232 46520
rect 20444 46164 20496 46170
rect 20444 46106 20496 46112
rect 20444 45960 20496 45966
rect 20350 45928 20406 45937
rect 20444 45902 20496 45908
rect 20350 45863 20406 45872
rect 20364 45830 20392 45863
rect 20352 45824 20404 45830
rect 20352 45766 20404 45772
rect 20456 45490 20484 45902
rect 20168 45484 20220 45490
rect 20168 45426 20220 45432
rect 20444 45484 20496 45490
rect 20444 45426 20496 45432
rect 20180 45014 20208 45426
rect 20548 45082 20576 46514
rect 21192 45966 21220 46514
rect 21180 45960 21232 45966
rect 21180 45902 21232 45908
rect 20720 45892 20772 45898
rect 20720 45834 20772 45840
rect 20732 45558 20760 45834
rect 20720 45552 20772 45558
rect 20720 45494 20772 45500
rect 20536 45076 20588 45082
rect 20536 45018 20588 45024
rect 20168 45008 20220 45014
rect 20168 44950 20220 44956
rect 20996 44872 21048 44878
rect 20996 44814 21048 44820
rect 20812 44804 20864 44810
rect 20812 44746 20864 44752
rect 20824 44402 20852 44746
rect 21008 44402 21036 44814
rect 21192 44742 21220 45902
rect 21376 45490 21404 47058
rect 21456 46640 21508 46646
rect 21456 46582 21508 46588
rect 21364 45484 21416 45490
rect 21364 45426 21416 45432
rect 21468 44878 21496 46582
rect 21652 46102 21680 49200
rect 22100 47592 22152 47598
rect 22100 47534 22152 47540
rect 22112 47258 22140 47534
rect 22192 47456 22244 47462
rect 22192 47398 22244 47404
rect 22100 47252 22152 47258
rect 22100 47194 22152 47200
rect 22204 47054 22232 47398
rect 22388 47190 22416 49200
rect 22376 47184 22428 47190
rect 22376 47126 22428 47132
rect 22192 47048 22244 47054
rect 22112 47008 22192 47036
rect 21824 46980 21876 46986
rect 21824 46922 21876 46928
rect 21640 46096 21692 46102
rect 21640 46038 21692 46044
rect 21456 44872 21508 44878
rect 21456 44814 21508 44820
rect 21180 44736 21232 44742
rect 21180 44678 21232 44684
rect 20076 44396 20128 44402
rect 20076 44338 20128 44344
rect 20812 44396 20864 44402
rect 20812 44338 20864 44344
rect 20996 44396 21048 44402
rect 20996 44338 21048 44344
rect 19064 44260 19116 44266
rect 19064 44202 19116 44208
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 21008 43790 21036 44338
rect 21468 44266 21496 44814
rect 21456 44260 21508 44266
rect 21456 44202 21508 44208
rect 21836 43926 21864 46922
rect 22112 46209 22140 47008
rect 22376 47048 22428 47054
rect 22192 46990 22244 46996
rect 22296 47008 22376 47036
rect 22098 46200 22154 46209
rect 22098 46135 22154 46144
rect 21916 45960 21968 45966
rect 21916 45902 21968 45908
rect 21928 45801 21956 45902
rect 21914 45792 21970 45801
rect 21914 45727 21970 45736
rect 22112 43994 22140 46135
rect 22296 45422 22324 47008
rect 22376 46990 22428 46996
rect 22744 46912 22796 46918
rect 22744 46854 22796 46860
rect 22756 46578 22784 46854
rect 22744 46572 22796 46578
rect 22744 46514 22796 46520
rect 22376 46436 22428 46442
rect 22376 46378 22428 46384
rect 22388 46050 22416 46378
rect 22848 46374 22876 49286
rect 23110 49200 23166 50000
rect 23478 49200 23534 50000
rect 23846 49200 23902 50000
rect 24214 49314 24270 50000
rect 24214 49286 24348 49314
rect 24214 49200 24270 49286
rect 23388 47116 23440 47122
rect 23388 47058 23440 47064
rect 22928 46980 22980 46986
rect 22928 46922 22980 46928
rect 22940 46578 22968 46922
rect 23400 46578 23428 47058
rect 23492 46646 23520 49200
rect 23756 47728 23808 47734
rect 23756 47670 23808 47676
rect 23768 47530 23796 47670
rect 23756 47524 23808 47530
rect 23756 47466 23808 47472
rect 23768 47054 23796 47466
rect 23572 47048 23624 47054
rect 23572 46990 23624 46996
rect 23756 47048 23808 47054
rect 23756 46990 23808 46996
rect 23480 46640 23532 46646
rect 23480 46582 23532 46588
rect 22928 46572 22980 46578
rect 22928 46514 22980 46520
rect 23296 46572 23348 46578
rect 23296 46514 23348 46520
rect 23388 46572 23440 46578
rect 23388 46514 23440 46520
rect 23204 46504 23256 46510
rect 23204 46446 23256 46452
rect 22836 46368 22888 46374
rect 22836 46310 22888 46316
rect 22928 46368 22980 46374
rect 22928 46310 22980 46316
rect 22388 46034 22692 46050
rect 22388 46028 22704 46034
rect 22388 46022 22652 46028
rect 22652 45970 22704 45976
rect 22376 45960 22428 45966
rect 22836 45960 22888 45966
rect 22376 45902 22428 45908
rect 22834 45928 22836 45937
rect 22888 45928 22890 45937
rect 22284 45416 22336 45422
rect 22284 45358 22336 45364
rect 22388 45404 22416 45902
rect 22652 45892 22704 45898
rect 22704 45852 22784 45880
rect 22834 45863 22890 45872
rect 22652 45834 22704 45840
rect 22468 45416 22520 45422
rect 22388 45376 22468 45404
rect 22388 44878 22416 45376
rect 22468 45358 22520 45364
rect 22376 44872 22428 44878
rect 22376 44814 22428 44820
rect 22468 44804 22520 44810
rect 22468 44746 22520 44752
rect 22480 44402 22508 44746
rect 22468 44396 22520 44402
rect 22468 44338 22520 44344
rect 22376 44192 22428 44198
rect 22376 44134 22428 44140
rect 22100 43988 22152 43994
rect 22100 43930 22152 43936
rect 21824 43920 21876 43926
rect 21824 43862 21876 43868
rect 20996 43784 21048 43790
rect 20996 43726 21048 43732
rect 21836 43654 21864 43862
rect 22388 43790 22416 44134
rect 22376 43784 22428 43790
rect 22376 43726 22428 43732
rect 21824 43648 21876 43654
rect 21824 43590 21876 43596
rect 22192 43648 22244 43654
rect 22192 43590 22244 43596
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 22204 42566 22232 43590
rect 22664 43450 22692 45834
rect 22756 45812 22784 45852
rect 22940 45812 22968 46310
rect 23020 45892 23072 45898
rect 23020 45834 23072 45840
rect 22756 45784 22968 45812
rect 23032 45626 23060 45834
rect 23020 45620 23072 45626
rect 23020 45562 23072 45568
rect 22744 45484 22796 45490
rect 22744 45426 22796 45432
rect 22756 44538 22784 45426
rect 22744 44532 22796 44538
rect 22744 44474 22796 44480
rect 23112 44396 23164 44402
rect 23112 44338 23164 44344
rect 22652 43444 22704 43450
rect 22652 43386 22704 43392
rect 22664 42838 22692 43386
rect 23124 43246 23152 44338
rect 23216 43858 23244 46446
rect 23308 45830 23336 46514
rect 23400 46102 23428 46514
rect 23388 46096 23440 46102
rect 23388 46038 23440 46044
rect 23584 45937 23612 46990
rect 23664 46912 23716 46918
rect 23664 46854 23716 46860
rect 23676 46578 23704 46854
rect 23664 46572 23716 46578
rect 23664 46514 23716 46520
rect 23768 46374 23796 46990
rect 23860 46646 23888 49200
rect 23940 47796 23992 47802
rect 23940 47738 23992 47744
rect 23848 46640 23900 46646
rect 23848 46582 23900 46588
rect 23756 46368 23808 46374
rect 23756 46310 23808 46316
rect 23662 46200 23718 46209
rect 23662 46135 23718 46144
rect 23676 46034 23704 46135
rect 23860 46034 23888 46582
rect 23952 46442 23980 47738
rect 24320 46646 24348 49286
rect 24582 49200 24638 50000
rect 24950 49200 25006 50000
rect 25318 49314 25374 50000
rect 25686 49314 25742 50000
rect 25318 49286 25636 49314
rect 25318 49200 25374 49286
rect 24596 47666 24624 49200
rect 24584 47660 24636 47666
rect 24584 47602 24636 47608
rect 24768 47524 24820 47530
rect 24768 47466 24820 47472
rect 24584 46980 24636 46986
rect 24584 46922 24636 46928
rect 24308 46640 24360 46646
rect 24308 46582 24360 46588
rect 24320 46510 24348 46582
rect 24308 46504 24360 46510
rect 24308 46446 24360 46452
rect 23940 46436 23992 46442
rect 23940 46378 23992 46384
rect 23664 46028 23716 46034
rect 23664 45970 23716 45976
rect 23848 46028 23900 46034
rect 23848 45970 23900 45976
rect 23952 45966 23980 46378
rect 23940 45960 23992 45966
rect 23570 45928 23626 45937
rect 23626 45886 23704 45914
rect 23940 45902 23992 45908
rect 23570 45863 23626 45872
rect 23296 45824 23348 45830
rect 23294 45792 23296 45801
rect 23584 45803 23612 45863
rect 23348 45792 23350 45801
rect 23294 45727 23350 45736
rect 23572 45484 23624 45490
rect 23572 45426 23624 45432
rect 23584 45082 23612 45426
rect 23572 45076 23624 45082
rect 23572 45018 23624 45024
rect 23676 45014 23704 45886
rect 23848 45552 23900 45558
rect 23768 45512 23848 45540
rect 23768 45422 23796 45512
rect 23848 45494 23900 45500
rect 23756 45416 23808 45422
rect 23756 45358 23808 45364
rect 23664 45008 23716 45014
rect 23664 44950 23716 44956
rect 24596 44878 24624 46922
rect 24780 45966 24808 47466
rect 24860 46640 24912 46646
rect 24860 46582 24912 46588
rect 24768 45960 24820 45966
rect 24768 45902 24820 45908
rect 24872 45830 24900 46582
rect 24860 45824 24912 45830
rect 24860 45766 24912 45772
rect 24872 45626 24900 45766
rect 24860 45620 24912 45626
rect 24860 45562 24912 45568
rect 24872 45490 24900 45562
rect 24860 45484 24912 45490
rect 24860 45426 24912 45432
rect 23756 44872 23808 44878
rect 23756 44814 23808 44820
rect 24032 44872 24084 44878
rect 24032 44814 24084 44820
rect 24584 44872 24636 44878
rect 24584 44814 24636 44820
rect 23768 44470 23796 44814
rect 23756 44464 23808 44470
rect 23756 44406 23808 44412
rect 23480 44396 23532 44402
rect 23480 44338 23532 44344
rect 23204 43852 23256 43858
rect 23204 43794 23256 43800
rect 23492 43722 23520 44338
rect 24044 44334 24072 44814
rect 24860 44736 24912 44742
rect 24860 44678 24912 44684
rect 24872 44470 24900 44678
rect 24860 44464 24912 44470
rect 24860 44406 24912 44412
rect 23572 44328 23624 44334
rect 23572 44270 23624 44276
rect 24032 44328 24084 44334
rect 24032 44270 24084 44276
rect 23480 43716 23532 43722
rect 23480 43658 23532 43664
rect 23584 43450 23612 44270
rect 23848 44260 23900 44266
rect 23848 44202 23900 44208
rect 23860 43790 23888 44202
rect 24964 43994 24992 49200
rect 25136 46980 25188 46986
rect 25136 46922 25188 46928
rect 25044 46912 25096 46918
rect 25044 46854 25096 46860
rect 25056 45966 25084 46854
rect 25148 46102 25176 46922
rect 25228 46708 25280 46714
rect 25228 46650 25280 46656
rect 25240 46510 25268 46650
rect 25228 46504 25280 46510
rect 25228 46446 25280 46452
rect 25608 46102 25636 49286
rect 25686 49286 26004 49314
rect 25686 49200 25742 49286
rect 25780 47116 25832 47122
rect 25780 47058 25832 47064
rect 25688 46912 25740 46918
rect 25688 46854 25740 46860
rect 25700 46646 25728 46854
rect 25688 46640 25740 46646
rect 25688 46582 25740 46588
rect 25792 46578 25820 47058
rect 25872 47048 25924 47054
rect 25872 46990 25924 46996
rect 25884 46714 25912 46990
rect 25872 46708 25924 46714
rect 25872 46650 25924 46656
rect 25780 46572 25832 46578
rect 25780 46514 25832 46520
rect 25136 46096 25188 46102
rect 25136 46038 25188 46044
rect 25596 46096 25648 46102
rect 25596 46038 25648 46044
rect 25044 45960 25096 45966
rect 25044 45902 25096 45908
rect 25792 45286 25820 46514
rect 25976 46322 26004 49286
rect 26054 49200 26110 50000
rect 26422 49200 26478 50000
rect 26790 49200 26846 50000
rect 27158 49200 27214 50000
rect 27526 49200 27582 50000
rect 27894 49200 27950 50000
rect 28262 49314 28318 50000
rect 28262 49286 28580 49314
rect 28262 49200 28318 49286
rect 26068 46918 26096 49200
rect 26056 46912 26108 46918
rect 26056 46854 26108 46860
rect 25976 46294 26280 46322
rect 25872 45348 25924 45354
rect 25872 45290 25924 45296
rect 25780 45280 25832 45286
rect 25780 45222 25832 45228
rect 25044 44940 25096 44946
rect 25044 44882 25096 44888
rect 25056 44334 25084 44882
rect 25596 44872 25648 44878
rect 25596 44814 25648 44820
rect 25504 44804 25556 44810
rect 25504 44746 25556 44752
rect 25516 44538 25544 44746
rect 25504 44532 25556 44538
rect 25504 44474 25556 44480
rect 25504 44396 25556 44402
rect 25504 44338 25556 44344
rect 25044 44328 25096 44334
rect 25044 44270 25096 44276
rect 24952 43988 25004 43994
rect 24952 43930 25004 43936
rect 23848 43784 23900 43790
rect 23848 43726 23900 43732
rect 24860 43716 24912 43722
rect 24860 43658 24912 43664
rect 23572 43444 23624 43450
rect 23572 43386 23624 43392
rect 24872 43314 24900 43658
rect 25056 43382 25084 44270
rect 25516 43722 25544 44338
rect 25504 43716 25556 43722
rect 25504 43658 25556 43664
rect 25044 43376 25096 43382
rect 25044 43318 25096 43324
rect 25608 43314 25636 44814
rect 25884 44742 25912 45290
rect 26056 44872 26108 44878
rect 26056 44814 26108 44820
rect 25872 44736 25924 44742
rect 25872 44678 25924 44684
rect 25964 44736 26016 44742
rect 25964 44678 26016 44684
rect 25884 44334 25912 44678
rect 25872 44328 25924 44334
rect 25872 44270 25924 44276
rect 25688 43716 25740 43722
rect 25688 43658 25740 43664
rect 25700 43382 25728 43658
rect 25688 43376 25740 43382
rect 25688 43318 25740 43324
rect 24860 43308 24912 43314
rect 24860 43250 24912 43256
rect 25596 43308 25648 43314
rect 25596 43250 25648 43256
rect 23112 43240 23164 43246
rect 23112 43182 23164 43188
rect 22652 42832 22704 42838
rect 22652 42774 22704 42780
rect 22192 42560 22244 42566
rect 22192 42502 22244 42508
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 22204 6662 22232 42502
rect 25884 42294 25912 44270
rect 25976 43790 26004 44678
rect 25964 43784 26016 43790
rect 25964 43726 26016 43732
rect 26068 43382 26096 44814
rect 26252 44402 26280 46294
rect 26436 46170 26464 49200
rect 26804 47258 26832 49200
rect 26792 47252 26844 47258
rect 26792 47194 26844 47200
rect 26516 47048 26568 47054
rect 26516 46990 26568 46996
rect 26528 46510 26556 46990
rect 26608 46980 26660 46986
rect 26608 46922 26660 46928
rect 26620 46578 26648 46922
rect 27172 46900 27200 49200
rect 27540 47530 27568 49200
rect 27528 47524 27580 47530
rect 27528 47466 27580 47472
rect 27344 47048 27396 47054
rect 27344 46990 27396 46996
rect 27252 46912 27304 46918
rect 27172 46872 27252 46900
rect 27252 46854 27304 46860
rect 26608 46572 26660 46578
rect 26608 46514 26660 46520
rect 26884 46572 26936 46578
rect 26884 46514 26936 46520
rect 26516 46504 26568 46510
rect 26516 46446 26568 46452
rect 26424 46164 26476 46170
rect 26424 46106 26476 46112
rect 26332 46028 26384 46034
rect 26332 45970 26384 45976
rect 26344 45626 26372 45970
rect 26332 45620 26384 45626
rect 26332 45562 26384 45568
rect 26332 45280 26384 45286
rect 26332 45222 26384 45228
rect 26240 44396 26292 44402
rect 26240 44338 26292 44344
rect 26056 43376 26108 43382
rect 26056 43318 26108 43324
rect 26344 42770 26372 45222
rect 26436 44878 26464 46106
rect 26528 45422 26556 46446
rect 26700 45960 26752 45966
rect 26700 45902 26752 45908
rect 26792 45960 26844 45966
rect 26792 45902 26844 45908
rect 26516 45416 26568 45422
rect 26516 45358 26568 45364
rect 26516 45280 26568 45286
rect 26516 45222 26568 45228
rect 26424 44872 26476 44878
rect 26424 44814 26476 44820
rect 26436 43926 26464 44814
rect 26528 44470 26556 45222
rect 26516 44464 26568 44470
rect 26516 44406 26568 44412
rect 26424 43920 26476 43926
rect 26424 43862 26476 43868
rect 26436 43450 26464 43862
rect 26712 43858 26740 45902
rect 26804 45830 26832 45902
rect 26792 45824 26844 45830
rect 26792 45766 26844 45772
rect 26896 45626 26924 46514
rect 27068 46368 27120 46374
rect 27068 46310 27120 46316
rect 27252 46368 27304 46374
rect 27252 46310 27304 46316
rect 27080 46170 27108 46310
rect 27068 46164 27120 46170
rect 27068 46106 27120 46112
rect 26884 45620 26936 45626
rect 26884 45562 26936 45568
rect 26896 44810 26924 45562
rect 26884 44804 26936 44810
rect 26884 44746 26936 44752
rect 26700 43852 26752 43858
rect 26700 43794 26752 43800
rect 26424 43444 26476 43450
rect 26424 43386 26476 43392
rect 26436 42906 26464 43386
rect 26896 43314 26924 44746
rect 26884 43308 26936 43314
rect 26884 43250 26936 43256
rect 27080 43194 27108 46106
rect 27264 46034 27292 46310
rect 27252 46028 27304 46034
rect 27252 45970 27304 45976
rect 27356 45490 27384 46990
rect 27528 46572 27580 46578
rect 27528 46514 27580 46520
rect 27804 46572 27856 46578
rect 27804 46514 27856 46520
rect 27540 46034 27568 46514
rect 27816 46170 27844 46514
rect 27908 46170 27936 49200
rect 28264 47184 28316 47190
rect 28264 47126 28316 47132
rect 28276 46646 28304 47126
rect 28264 46640 28316 46646
rect 28264 46582 28316 46588
rect 27804 46164 27856 46170
rect 27804 46106 27856 46112
rect 27896 46164 27948 46170
rect 27896 46106 27948 46112
rect 27528 46028 27580 46034
rect 27580 45988 27660 46016
rect 27528 45970 27580 45976
rect 27436 45960 27488 45966
rect 27436 45902 27488 45908
rect 27344 45484 27396 45490
rect 27344 45426 27396 45432
rect 27356 45354 27384 45426
rect 27344 45348 27396 45354
rect 27344 45290 27396 45296
rect 27448 44878 27476 45902
rect 27632 45490 27660 45988
rect 28552 45898 28580 49286
rect 28630 49200 28686 50000
rect 28998 49200 29054 50000
rect 29366 49200 29422 50000
rect 29734 49200 29790 50000
rect 30102 49200 30158 50000
rect 30470 49200 30526 50000
rect 30838 49314 30894 50000
rect 30760 49286 30894 49314
rect 28644 46714 28672 49200
rect 29012 47598 29040 49200
rect 29000 47592 29052 47598
rect 29000 47534 29052 47540
rect 28724 47116 28776 47122
rect 28724 47058 28776 47064
rect 29276 47116 29328 47122
rect 29276 47058 29328 47064
rect 28632 46708 28684 46714
rect 28632 46650 28684 46656
rect 28736 46034 28764 47058
rect 28816 47048 28868 47054
rect 28816 46990 28868 46996
rect 29092 47048 29144 47054
rect 29092 46990 29144 46996
rect 28828 46753 28856 46990
rect 28814 46744 28870 46753
rect 28814 46679 28870 46688
rect 28828 46102 28856 46679
rect 28816 46096 28868 46102
rect 28816 46038 28868 46044
rect 28724 46028 28776 46034
rect 28724 45970 28776 45976
rect 28540 45892 28592 45898
rect 28540 45834 28592 45840
rect 27988 45620 28040 45626
rect 27988 45562 28040 45568
rect 28000 45490 28028 45562
rect 28736 45490 28764 45970
rect 28908 45960 28960 45966
rect 29104 45937 29132 46990
rect 29288 46578 29316 47058
rect 29276 46572 29328 46578
rect 29276 46514 29328 46520
rect 28908 45902 28960 45908
rect 29090 45928 29146 45937
rect 27620 45484 27672 45490
rect 27620 45426 27672 45432
rect 27988 45484 28040 45490
rect 27988 45426 28040 45432
rect 28724 45484 28776 45490
rect 28724 45426 28776 45432
rect 27632 45354 27660 45426
rect 27620 45348 27672 45354
rect 27620 45290 27672 45296
rect 27804 45280 27856 45286
rect 27804 45222 27856 45228
rect 28632 45280 28684 45286
rect 28632 45222 28684 45228
rect 28920 45234 28948 45902
rect 29090 45863 29146 45872
rect 29000 45824 29052 45830
rect 29000 45766 29052 45772
rect 29012 45558 29040 45766
rect 29276 45620 29328 45626
rect 29276 45562 29328 45568
rect 29000 45552 29052 45558
rect 29000 45494 29052 45500
rect 29184 45484 29236 45490
rect 29184 45426 29236 45432
rect 29092 45348 29144 45354
rect 29092 45290 29144 45296
rect 27816 44878 27844 45222
rect 28356 44940 28408 44946
rect 28356 44882 28408 44888
rect 27344 44872 27396 44878
rect 27344 44814 27396 44820
rect 27436 44872 27488 44878
rect 27804 44872 27856 44878
rect 27488 44832 27568 44860
rect 27436 44814 27488 44820
rect 27252 44736 27304 44742
rect 27252 44678 27304 44684
rect 27264 44538 27292 44678
rect 27356 44538 27384 44814
rect 27252 44532 27304 44538
rect 27252 44474 27304 44480
rect 27344 44532 27396 44538
rect 27344 44474 27396 44480
rect 27160 44464 27212 44470
rect 27160 44406 27212 44412
rect 27172 43790 27200 44406
rect 27160 43784 27212 43790
rect 27160 43726 27212 43732
rect 27264 43314 27292 44474
rect 27252 43308 27304 43314
rect 27252 43250 27304 43256
rect 27080 43166 27292 43194
rect 26424 42900 26476 42906
rect 26424 42842 26476 42848
rect 26332 42764 26384 42770
rect 26332 42706 26384 42712
rect 26344 42362 26372 42706
rect 27264 42566 27292 43166
rect 27356 42770 27384 44474
rect 27436 44396 27488 44402
rect 27436 44338 27488 44344
rect 27448 43722 27476 44338
rect 27436 43716 27488 43722
rect 27436 43658 27488 43664
rect 27448 43110 27476 43658
rect 27436 43104 27488 43110
rect 27436 43046 27488 43052
rect 27540 42770 27568 44832
rect 27804 44814 27856 44820
rect 27712 44804 27764 44810
rect 27712 44746 27764 44752
rect 27724 44334 27752 44746
rect 27712 44328 27764 44334
rect 27712 44270 27764 44276
rect 28368 43790 28396 44882
rect 28644 44878 28672 45222
rect 28920 45206 29040 45234
rect 29012 44878 29040 45206
rect 28632 44872 28684 44878
rect 28632 44814 28684 44820
rect 29000 44872 29052 44878
rect 29000 44814 29052 44820
rect 29104 43994 29132 45290
rect 29196 45286 29224 45426
rect 29184 45280 29236 45286
rect 29184 45222 29236 45228
rect 29196 44810 29224 45222
rect 29184 44804 29236 44810
rect 29184 44746 29236 44752
rect 29092 43988 29144 43994
rect 29092 43930 29144 43936
rect 29196 43790 29224 44746
rect 29288 44470 29316 45562
rect 29276 44464 29328 44470
rect 29276 44406 29328 44412
rect 27620 43784 27672 43790
rect 27620 43726 27672 43732
rect 28356 43784 28408 43790
rect 28356 43726 28408 43732
rect 29184 43784 29236 43790
rect 29184 43726 29236 43732
rect 27632 43450 27660 43726
rect 27620 43444 27672 43450
rect 27620 43386 27672 43392
rect 29196 42906 29224 43726
rect 29288 43382 29316 44406
rect 29380 43994 29408 49200
rect 29644 47456 29696 47462
rect 29644 47398 29696 47404
rect 29656 46714 29684 47398
rect 29644 46708 29696 46714
rect 29644 46650 29696 46656
rect 29460 46572 29512 46578
rect 29460 46514 29512 46520
rect 29472 46102 29500 46514
rect 29460 46096 29512 46102
rect 29460 46038 29512 46044
rect 29644 45824 29696 45830
rect 29644 45766 29696 45772
rect 29656 44402 29684 45766
rect 29748 45286 29776 49200
rect 30116 46714 30144 49200
rect 30484 47190 30512 49200
rect 30472 47184 30524 47190
rect 30472 47126 30524 47132
rect 30656 47048 30708 47054
rect 30656 46990 30708 46996
rect 30564 46980 30616 46986
rect 30564 46922 30616 46928
rect 30104 46708 30156 46714
rect 30104 46650 30156 46656
rect 30288 46640 30340 46646
rect 30288 46582 30340 46588
rect 29828 46572 29880 46578
rect 29828 46514 29880 46520
rect 29840 45626 29868 46514
rect 30300 46345 30328 46582
rect 30286 46336 30342 46345
rect 30286 46271 30342 46280
rect 30300 45966 30328 46271
rect 30576 46209 30604 46922
rect 30668 46646 30696 46990
rect 30656 46640 30708 46646
rect 30656 46582 30708 46588
rect 30562 46200 30618 46209
rect 30562 46135 30618 46144
rect 30564 46028 30616 46034
rect 30564 45970 30616 45976
rect 30196 45960 30248 45966
rect 30196 45902 30248 45908
rect 30288 45960 30340 45966
rect 30288 45902 30340 45908
rect 29828 45620 29880 45626
rect 29828 45562 29880 45568
rect 30208 45354 30236 45902
rect 30300 45490 30328 45902
rect 30576 45558 30604 45970
rect 30564 45552 30616 45558
rect 30564 45494 30616 45500
rect 30288 45484 30340 45490
rect 30288 45426 30340 45432
rect 30196 45348 30248 45354
rect 30196 45290 30248 45296
rect 29736 45280 29788 45286
rect 29736 45222 29788 45228
rect 29644 44396 29696 44402
rect 29644 44338 29696 44344
rect 29368 43988 29420 43994
rect 29368 43930 29420 43936
rect 29276 43376 29328 43382
rect 29276 43318 29328 43324
rect 29736 43172 29788 43178
rect 29736 43114 29788 43120
rect 29184 42900 29236 42906
rect 29184 42842 29236 42848
rect 27344 42764 27396 42770
rect 27344 42706 27396 42712
rect 27528 42764 27580 42770
rect 27528 42706 27580 42712
rect 27252 42560 27304 42566
rect 27252 42502 27304 42508
rect 27264 42362 27292 42502
rect 27540 42362 27568 42706
rect 29276 42560 29328 42566
rect 29276 42502 29328 42508
rect 26332 42356 26384 42362
rect 26332 42298 26384 42304
rect 27252 42356 27304 42362
rect 27252 42298 27304 42304
rect 27528 42356 27580 42362
rect 27528 42298 27580 42304
rect 25872 42288 25924 42294
rect 25872 42230 25924 42236
rect 29288 42022 29316 42502
rect 29644 42288 29696 42294
rect 29644 42230 29696 42236
rect 29276 42016 29328 42022
rect 29276 41958 29328 41964
rect 29288 41818 29316 41958
rect 29656 41818 29684 42230
rect 29276 41812 29328 41818
rect 29276 41754 29328 41760
rect 29644 41812 29696 41818
rect 29644 41754 29696 41760
rect 29748 6914 29776 43114
rect 30300 43110 30328 45426
rect 30576 44946 30604 45494
rect 30760 45490 30788 49286
rect 30838 49200 30894 49286
rect 31206 49200 31262 50000
rect 31574 49200 31630 50000
rect 31942 49200 31998 50000
rect 32310 49314 32366 50000
rect 32310 49286 32628 49314
rect 32310 49200 32366 49286
rect 31024 46980 31076 46986
rect 31024 46922 31076 46928
rect 30932 46912 30984 46918
rect 30932 46854 30984 46860
rect 30944 46578 30972 46854
rect 30932 46572 30984 46578
rect 30932 46514 30984 46520
rect 31036 46510 31064 46922
rect 31024 46504 31076 46510
rect 31024 46446 31076 46452
rect 31036 45812 31064 46446
rect 30944 45784 31064 45812
rect 30748 45484 30800 45490
rect 30748 45426 30800 45432
rect 30564 44940 30616 44946
rect 30564 44882 30616 44888
rect 30760 44402 30788 45426
rect 30944 44538 30972 45784
rect 31024 45280 31076 45286
rect 31024 45222 31076 45228
rect 30932 44532 30984 44538
rect 30932 44474 30984 44480
rect 30748 44396 30800 44402
rect 30748 44338 30800 44344
rect 30288 43104 30340 43110
rect 30288 43046 30340 43052
rect 30760 42770 30788 44338
rect 30932 44328 30984 44334
rect 30932 44270 30984 44276
rect 30944 43994 30972 44270
rect 30932 43988 30984 43994
rect 30932 43930 30984 43936
rect 31036 43790 31064 45222
rect 31024 43784 31076 43790
rect 31024 43726 31076 43732
rect 31220 43314 31248 49200
rect 31588 47462 31616 49200
rect 31576 47456 31628 47462
rect 31576 47398 31628 47404
rect 31484 46912 31536 46918
rect 31484 46854 31536 46860
rect 31760 46912 31812 46918
rect 31760 46854 31812 46860
rect 31496 46034 31524 46854
rect 31666 46744 31722 46753
rect 31666 46679 31722 46688
rect 31680 46578 31708 46679
rect 31668 46572 31720 46578
rect 31668 46514 31720 46520
rect 31668 46368 31720 46374
rect 31668 46310 31720 46316
rect 31484 46028 31536 46034
rect 31484 45970 31536 45976
rect 31496 45082 31524 45970
rect 31680 45626 31708 46310
rect 31772 46034 31800 46854
rect 31760 46028 31812 46034
rect 31760 45970 31812 45976
rect 31668 45620 31720 45626
rect 31668 45562 31720 45568
rect 31772 45422 31800 45970
rect 31760 45416 31812 45422
rect 31760 45358 31812 45364
rect 31484 45076 31536 45082
rect 31484 45018 31536 45024
rect 31956 44878 31984 49200
rect 32036 47048 32088 47054
rect 32036 46990 32088 46996
rect 32048 46034 32076 46990
rect 32600 46866 32628 49286
rect 32678 49200 32734 50000
rect 33046 49200 33102 50000
rect 33414 49200 33470 50000
rect 33782 49200 33838 50000
rect 34150 49200 34206 50000
rect 34518 49200 34574 50000
rect 34886 49200 34942 50000
rect 35254 49314 35310 50000
rect 35254 49286 35480 49314
rect 35254 49200 35310 49286
rect 32692 47258 32720 49200
rect 32680 47252 32732 47258
rect 32680 47194 32732 47200
rect 32772 46912 32824 46918
rect 32600 46860 32772 46866
rect 32600 46854 32824 46860
rect 32600 46838 32812 46854
rect 33060 46628 33088 49200
rect 33324 47048 33376 47054
rect 33324 46990 33376 46996
rect 33232 46980 33284 46986
rect 33232 46922 33284 46928
rect 33140 46640 33192 46646
rect 33060 46600 33140 46628
rect 33140 46582 33192 46588
rect 33244 46578 33272 46922
rect 32496 46572 32548 46578
rect 32496 46514 32548 46520
rect 33232 46572 33284 46578
rect 33232 46514 33284 46520
rect 32508 46345 32536 46514
rect 32494 46336 32550 46345
rect 32494 46271 32550 46280
rect 32036 46028 32088 46034
rect 32036 45970 32088 45976
rect 32680 45824 32732 45830
rect 32680 45766 32732 45772
rect 32312 45484 32364 45490
rect 32312 45426 32364 45432
rect 32128 45416 32180 45422
rect 32128 45358 32180 45364
rect 31760 44872 31812 44878
rect 31760 44814 31812 44820
rect 31944 44872 31996 44878
rect 31944 44814 31996 44820
rect 31668 43784 31720 43790
rect 31668 43726 31720 43732
rect 31680 43314 31708 43726
rect 31208 43308 31260 43314
rect 31208 43250 31260 43256
rect 31668 43308 31720 43314
rect 31668 43250 31720 43256
rect 30932 43104 30984 43110
rect 30932 43046 30984 43052
rect 30748 42764 30800 42770
rect 30748 42706 30800 42712
rect 30760 42294 30788 42706
rect 30944 42634 30972 43046
rect 31772 42634 31800 44814
rect 32140 43382 32168 45358
rect 32324 44985 32352 45426
rect 32404 45280 32456 45286
rect 32404 45222 32456 45228
rect 32588 45280 32640 45286
rect 32588 45222 32640 45228
rect 32310 44976 32366 44985
rect 32310 44911 32366 44920
rect 32324 44878 32352 44911
rect 32312 44872 32364 44878
rect 32312 44814 32364 44820
rect 32416 44402 32444 45222
rect 32600 44470 32628 45222
rect 32588 44464 32640 44470
rect 32588 44406 32640 44412
rect 32404 44396 32456 44402
rect 32404 44338 32456 44344
rect 32692 43654 32720 45766
rect 33336 45626 33364 46990
rect 33324 45620 33376 45626
rect 33324 45562 33376 45568
rect 33140 45552 33192 45558
rect 33140 45494 33192 45500
rect 33152 44946 33180 45494
rect 33232 45416 33284 45422
rect 33232 45358 33284 45364
rect 33140 44940 33192 44946
rect 33140 44882 33192 44888
rect 33048 44736 33100 44742
rect 33048 44678 33100 44684
rect 33060 44402 33088 44678
rect 33048 44396 33100 44402
rect 33048 44338 33100 44344
rect 32864 44328 32916 44334
rect 32864 44270 32916 44276
rect 32876 43926 32904 44270
rect 32864 43920 32916 43926
rect 32864 43862 32916 43868
rect 32876 43790 32904 43862
rect 33060 43858 33088 44338
rect 33152 43926 33180 44882
rect 33244 44878 33272 45358
rect 33336 44878 33364 45562
rect 33232 44872 33284 44878
rect 33232 44814 33284 44820
rect 33324 44872 33376 44878
rect 33324 44814 33376 44820
rect 33140 43920 33192 43926
rect 33140 43862 33192 43868
rect 33048 43852 33100 43858
rect 33048 43794 33100 43800
rect 32864 43784 32916 43790
rect 32864 43726 32916 43732
rect 33048 43716 33100 43722
rect 33048 43658 33100 43664
rect 32680 43648 32732 43654
rect 32680 43590 32732 43596
rect 32692 43382 32720 43590
rect 32128 43376 32180 43382
rect 32128 43318 32180 43324
rect 32680 43376 32732 43382
rect 32680 43318 32732 43324
rect 33060 43314 33088 43658
rect 33244 43450 33272 44814
rect 33232 43444 33284 43450
rect 33232 43386 33284 43392
rect 33428 43314 33456 49200
rect 33600 47524 33652 47530
rect 33600 47466 33652 47472
rect 33612 47054 33640 47466
rect 33600 47048 33652 47054
rect 33520 47008 33600 47036
rect 33520 43382 33548 47008
rect 33600 46990 33652 46996
rect 33600 45484 33652 45490
rect 33600 45426 33652 45432
rect 33612 45014 33640 45426
rect 33600 45008 33652 45014
rect 33600 44950 33652 44956
rect 33796 44962 33824 49200
rect 33874 47152 33930 47161
rect 33874 47087 33930 47096
rect 33888 47054 33916 47087
rect 33876 47048 33928 47054
rect 33876 46990 33928 46996
rect 33888 46510 33916 46990
rect 33876 46504 33928 46510
rect 33876 46446 33928 46452
rect 33888 45966 33916 46446
rect 33876 45960 33928 45966
rect 33876 45902 33928 45908
rect 34164 45830 34192 49200
rect 34532 47274 34560 49200
rect 34704 47592 34756 47598
rect 34900 47546 34928 49200
rect 34704 47534 34756 47540
rect 34532 47246 34652 47274
rect 34244 47116 34296 47122
rect 34244 47058 34296 47064
rect 34520 47116 34572 47122
rect 34520 47058 34572 47064
rect 34256 46578 34284 47058
rect 34532 46714 34560 47058
rect 34624 46753 34652 47246
rect 34716 47054 34744 47534
rect 34808 47518 34928 47546
rect 34704 47048 34756 47054
rect 34704 46990 34756 46996
rect 34610 46744 34666 46753
rect 34520 46708 34572 46714
rect 34808 46730 34836 47518
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34808 46702 34928 46730
rect 34610 46679 34666 46688
rect 34520 46650 34572 46656
rect 34244 46572 34296 46578
rect 34244 46514 34296 46520
rect 34612 46572 34664 46578
rect 34612 46514 34664 46520
rect 34796 46572 34848 46578
rect 34796 46514 34848 46520
rect 34152 45824 34204 45830
rect 34152 45766 34204 45772
rect 34256 45422 34284 46514
rect 34336 46504 34388 46510
rect 34334 46472 34336 46481
rect 34388 46472 34390 46481
rect 34334 46407 34390 46416
rect 34624 45801 34652 46514
rect 34808 46170 34836 46514
rect 34900 46442 34928 46702
rect 34980 46708 35032 46714
rect 34980 46650 35032 46656
rect 34992 46578 35020 46650
rect 34980 46572 35032 46578
rect 34980 46514 35032 46520
rect 34888 46436 34940 46442
rect 34888 46378 34940 46384
rect 35348 46368 35400 46374
rect 35348 46310 35400 46316
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34796 46164 34848 46170
rect 34796 46106 34848 46112
rect 35360 46034 35388 46310
rect 35348 46028 35400 46034
rect 35348 45970 35400 45976
rect 34610 45792 34666 45801
rect 34610 45727 34666 45736
rect 34624 45626 34652 45727
rect 34612 45620 34664 45626
rect 34612 45562 34664 45568
rect 35452 45558 35480 49286
rect 35622 49200 35678 50000
rect 35990 49200 36046 50000
rect 36358 49200 36414 50000
rect 36726 49200 36782 50000
rect 37094 49200 37150 50000
rect 37462 49200 37518 50000
rect 37830 49200 37886 50000
rect 38198 49200 38254 50000
rect 38566 49200 38622 50000
rect 38934 49200 38990 50000
rect 39302 49200 39358 50000
rect 39670 49200 39726 50000
rect 40038 49200 40094 50000
rect 40406 49200 40462 50000
rect 40774 49200 40830 50000
rect 41142 49200 41198 50000
rect 41510 49200 41566 50000
rect 41878 49200 41934 50000
rect 42246 49200 42302 50000
rect 42614 49200 42670 50000
rect 42982 49200 43038 50000
rect 43350 49200 43406 50000
rect 43718 49314 43774 50000
rect 43718 49286 43944 49314
rect 43718 49200 43774 49286
rect 35636 46889 35664 49200
rect 35714 47152 35770 47161
rect 35714 47087 35770 47096
rect 35622 46880 35678 46889
rect 35622 46815 35678 46824
rect 35532 46640 35584 46646
rect 35532 46582 35584 46588
rect 35544 46034 35572 46582
rect 35624 46572 35676 46578
rect 35624 46514 35676 46520
rect 35532 46028 35584 46034
rect 35532 45970 35584 45976
rect 34520 45552 34572 45558
rect 34520 45494 34572 45500
rect 35440 45552 35492 45558
rect 35440 45494 35492 45500
rect 33968 45416 34020 45422
rect 33968 45358 34020 45364
rect 34152 45416 34204 45422
rect 34152 45358 34204 45364
rect 34244 45416 34296 45422
rect 34244 45358 34296 45364
rect 33796 44934 33916 44962
rect 33784 44872 33836 44878
rect 33784 44814 33836 44820
rect 33796 44470 33824 44814
rect 33784 44464 33836 44470
rect 33784 44406 33836 44412
rect 33508 43376 33560 43382
rect 33508 43318 33560 43324
rect 33888 43314 33916 44934
rect 33980 44402 34008 45358
rect 33968 44396 34020 44402
rect 33968 44338 34020 44344
rect 34164 43994 34192 45358
rect 34152 43988 34204 43994
rect 34152 43930 34204 43936
rect 34256 43790 34284 45358
rect 34532 44878 34560 45494
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34520 44872 34572 44878
rect 34520 44814 34572 44820
rect 34532 44402 34560 44814
rect 34520 44396 34572 44402
rect 34520 44338 34572 44344
rect 34532 43994 34560 44338
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34520 43988 34572 43994
rect 34520 43930 34572 43936
rect 35452 43858 35480 45494
rect 35544 45286 35572 45970
rect 35636 45966 35664 46514
rect 35624 45960 35676 45966
rect 35624 45902 35676 45908
rect 35624 45416 35676 45422
rect 35624 45358 35676 45364
rect 35532 45280 35584 45286
rect 35532 45222 35584 45228
rect 35440 43852 35492 43858
rect 35440 43794 35492 43800
rect 34244 43784 34296 43790
rect 34244 43726 34296 43732
rect 35452 43450 35480 43794
rect 35440 43444 35492 43450
rect 35440 43386 35492 43392
rect 32864 43308 32916 43314
rect 32864 43250 32916 43256
rect 33048 43308 33100 43314
rect 33048 43250 33100 43256
rect 33416 43308 33468 43314
rect 33416 43250 33468 43256
rect 33876 43308 33928 43314
rect 33876 43250 33928 43256
rect 32876 42906 32904 43250
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 35452 42906 35480 43386
rect 35544 43382 35572 45222
rect 35636 45082 35664 45358
rect 35624 45076 35676 45082
rect 35624 45018 35676 45024
rect 35728 43450 35756 47087
rect 35900 47048 35952 47054
rect 35898 47016 35900 47025
rect 35952 47016 35954 47025
rect 35898 46951 35954 46960
rect 36004 46578 36032 49200
rect 36372 47530 36400 49200
rect 36452 47592 36504 47598
rect 36452 47534 36504 47540
rect 36360 47524 36412 47530
rect 36360 47466 36412 47472
rect 35992 46572 36044 46578
rect 35992 46514 36044 46520
rect 35992 46368 36044 46374
rect 35992 46310 36044 46316
rect 36004 46102 36032 46310
rect 35992 46096 36044 46102
rect 35992 46038 36044 46044
rect 36464 45966 36492 47534
rect 36544 47456 36596 47462
rect 36544 47398 36596 47404
rect 36556 46374 36584 47398
rect 36740 46714 36768 49200
rect 36820 47184 36872 47190
rect 36820 47126 36872 47132
rect 36832 47054 36860 47126
rect 36820 47048 36872 47054
rect 36820 46990 36872 46996
rect 36728 46708 36780 46714
rect 36728 46650 36780 46656
rect 37108 46646 37136 49200
rect 37096 46640 37148 46646
rect 37096 46582 37148 46588
rect 37370 46608 37426 46617
rect 37188 46572 37240 46578
rect 37370 46543 37426 46552
rect 37188 46514 37240 46520
rect 36728 46504 36780 46510
rect 37200 46481 37228 46514
rect 36728 46446 36780 46452
rect 37186 46472 37242 46481
rect 36544 46368 36596 46374
rect 36544 46310 36596 46316
rect 36740 46073 36768 46446
rect 37186 46407 37242 46416
rect 36818 46336 36874 46345
rect 36818 46271 36874 46280
rect 36726 46064 36782 46073
rect 36726 45999 36782 46008
rect 36740 45966 36768 45999
rect 36832 45966 36860 46271
rect 37384 46170 37412 46543
rect 37476 46510 37504 49200
rect 37738 47152 37794 47161
rect 37738 47087 37740 47096
rect 37792 47087 37794 47096
rect 37740 47058 37792 47064
rect 37648 47048 37700 47054
rect 37648 46990 37700 46996
rect 37464 46504 37516 46510
rect 37464 46446 37516 46452
rect 37372 46164 37424 46170
rect 37372 46106 37424 46112
rect 36176 45960 36228 45966
rect 36176 45902 36228 45908
rect 36452 45960 36504 45966
rect 36452 45902 36504 45908
rect 36544 45960 36596 45966
rect 36544 45902 36596 45908
rect 36728 45960 36780 45966
rect 36728 45902 36780 45908
rect 36820 45960 36872 45966
rect 36820 45902 36872 45908
rect 35808 45824 35860 45830
rect 35808 45766 35860 45772
rect 35820 45014 35848 45766
rect 36188 45490 36216 45902
rect 36464 45626 36492 45902
rect 36556 45830 36584 45902
rect 36544 45824 36596 45830
rect 36544 45766 36596 45772
rect 37004 45824 37056 45830
rect 37004 45766 37056 45772
rect 36452 45620 36504 45626
rect 36452 45562 36504 45568
rect 36176 45484 36228 45490
rect 36176 45426 36228 45432
rect 36636 45484 36688 45490
rect 36636 45426 36688 45432
rect 35900 45416 35952 45422
rect 35900 45358 35952 45364
rect 35808 45008 35860 45014
rect 35808 44950 35860 44956
rect 35912 44334 35940 45358
rect 36544 44396 36596 44402
rect 36544 44338 36596 44344
rect 35900 44328 35952 44334
rect 35900 44270 35952 44276
rect 35912 43738 35940 44270
rect 36556 43994 36584 44338
rect 36544 43988 36596 43994
rect 36544 43930 36596 43936
rect 36648 43926 36676 45426
rect 36728 45348 36780 45354
rect 36728 45290 36780 45296
rect 36740 44985 36768 45290
rect 36726 44976 36782 44985
rect 36726 44911 36782 44920
rect 37016 44878 37044 45766
rect 37476 45422 37504 46446
rect 37660 46374 37688 46990
rect 37740 46912 37792 46918
rect 37740 46854 37792 46860
rect 37752 46578 37780 46854
rect 37740 46572 37792 46578
rect 37740 46514 37792 46520
rect 37648 46368 37700 46374
rect 37648 46310 37700 46316
rect 37660 45898 37688 46310
rect 37740 46096 37792 46102
rect 37740 46038 37792 46044
rect 37648 45892 37700 45898
rect 37648 45834 37700 45840
rect 37464 45416 37516 45422
rect 37464 45358 37516 45364
rect 37188 45348 37240 45354
rect 37188 45290 37240 45296
rect 37200 44878 37228 45290
rect 37464 45008 37516 45014
rect 37464 44950 37516 44956
rect 37004 44872 37056 44878
rect 37004 44814 37056 44820
rect 37188 44872 37240 44878
rect 37188 44814 37240 44820
rect 37476 44402 37504 44950
rect 37648 44804 37700 44810
rect 37648 44746 37700 44752
rect 37660 44402 37688 44746
rect 37752 44538 37780 46038
rect 37844 45626 37872 49200
rect 38016 47048 38068 47054
rect 38016 46990 38068 46996
rect 38028 46578 38056 46990
rect 38016 46572 38068 46578
rect 38016 46514 38068 46520
rect 38028 46170 38056 46514
rect 38016 46164 38068 46170
rect 38016 46106 38068 46112
rect 37832 45620 37884 45626
rect 37832 45562 37884 45568
rect 38028 45490 38056 46106
rect 38212 46102 38240 49200
rect 38384 46912 38436 46918
rect 38384 46854 38436 46860
rect 38290 46472 38346 46481
rect 38290 46407 38292 46416
rect 38344 46407 38346 46416
rect 38292 46378 38344 46384
rect 38200 46096 38252 46102
rect 38200 46038 38252 46044
rect 38108 45960 38160 45966
rect 38108 45902 38160 45908
rect 38120 45801 38148 45902
rect 38106 45792 38162 45801
rect 38106 45727 38162 45736
rect 38016 45484 38068 45490
rect 38016 45426 38068 45432
rect 37924 45416 37976 45422
rect 37924 45358 37976 45364
rect 37936 44810 37964 45358
rect 38028 44946 38056 45426
rect 38120 45422 38148 45727
rect 38396 45642 38424 46854
rect 38476 46504 38528 46510
rect 38476 46446 38528 46452
rect 38488 46345 38516 46446
rect 38474 46336 38530 46345
rect 38474 46271 38530 46280
rect 38212 45614 38424 45642
rect 38108 45416 38160 45422
rect 38108 45358 38160 45364
rect 38108 45076 38160 45082
rect 38212 45064 38240 45614
rect 38580 45490 38608 49200
rect 38844 46504 38896 46510
rect 38844 46446 38896 46452
rect 38292 45484 38344 45490
rect 38292 45426 38344 45432
rect 38568 45484 38620 45490
rect 38568 45426 38620 45432
rect 38660 45484 38712 45490
rect 38660 45426 38712 45432
rect 38160 45036 38240 45064
rect 38108 45018 38160 45024
rect 38016 44940 38068 44946
rect 38016 44882 38068 44888
rect 37924 44804 37976 44810
rect 37924 44746 37976 44752
rect 37740 44532 37792 44538
rect 37740 44474 37792 44480
rect 37464 44396 37516 44402
rect 37464 44338 37516 44344
rect 37648 44396 37700 44402
rect 37648 44338 37700 44344
rect 37556 44192 37608 44198
rect 37556 44134 37608 44140
rect 36820 43988 36872 43994
rect 36820 43930 36872 43936
rect 36636 43920 36688 43926
rect 36636 43862 36688 43868
rect 36832 43858 36860 43930
rect 36820 43852 36872 43858
rect 36820 43794 36872 43800
rect 35912 43722 36032 43738
rect 35912 43716 36044 43722
rect 35912 43710 35992 43716
rect 35992 43658 36044 43664
rect 36832 43450 36860 43794
rect 35716 43444 35768 43450
rect 35716 43386 35768 43392
rect 36820 43444 36872 43450
rect 36820 43386 36872 43392
rect 35532 43376 35584 43382
rect 35532 43318 35584 43324
rect 32864 42900 32916 42906
rect 32864 42842 32916 42848
rect 35440 42900 35492 42906
rect 35440 42842 35492 42848
rect 35544 42838 35572 43318
rect 35532 42832 35584 42838
rect 35532 42774 35584 42780
rect 30932 42628 30984 42634
rect 30932 42570 30984 42576
rect 31760 42628 31812 42634
rect 31760 42570 31812 42576
rect 30944 42362 30972 42570
rect 35728 42362 35756 43386
rect 37568 43314 37596 44134
rect 37660 43722 37688 44338
rect 37740 43784 37792 43790
rect 37740 43726 37792 43732
rect 37648 43716 37700 43722
rect 37648 43658 37700 43664
rect 37752 43450 37780 43726
rect 37740 43444 37792 43450
rect 37740 43386 37792 43392
rect 38212 43382 38240 45036
rect 38304 44878 38332 45426
rect 38672 45370 38700 45426
rect 38488 45342 38700 45370
rect 38384 45280 38436 45286
rect 38384 45222 38436 45228
rect 38396 45082 38424 45222
rect 38384 45076 38436 45082
rect 38384 45018 38436 45024
rect 38292 44872 38344 44878
rect 38292 44814 38344 44820
rect 38396 44402 38424 45018
rect 38488 44810 38516 45342
rect 38856 45014 38884 46446
rect 38948 46170 38976 49200
rect 39316 47258 39344 49200
rect 39304 47252 39356 47258
rect 39304 47194 39356 47200
rect 39488 47116 39540 47122
rect 39488 47058 39540 47064
rect 39028 46572 39080 46578
rect 39028 46514 39080 46520
rect 38936 46164 38988 46170
rect 38936 46106 38988 46112
rect 39040 45830 39068 46514
rect 39120 46436 39172 46442
rect 39120 46378 39172 46384
rect 39132 46034 39160 46378
rect 39120 46028 39172 46034
rect 39120 45970 39172 45976
rect 39500 45966 39528 47058
rect 39684 46918 39712 49200
rect 39672 46912 39724 46918
rect 39672 46854 39724 46860
rect 40052 46714 40080 49200
rect 40132 47048 40184 47054
rect 40132 46990 40184 46996
rect 40144 46753 40172 46990
rect 40224 46912 40276 46918
rect 40224 46854 40276 46860
rect 40130 46744 40186 46753
rect 39948 46708 40000 46714
rect 39948 46650 40000 46656
rect 40040 46708 40092 46714
rect 40130 46679 40186 46688
rect 40040 46650 40092 46656
rect 39960 46034 39988 46650
rect 40236 46594 40264 46854
rect 40052 46566 40264 46594
rect 40052 46442 40080 46566
rect 40040 46436 40092 46442
rect 40040 46378 40092 46384
rect 39948 46028 40000 46034
rect 39948 45970 40000 45976
rect 39488 45960 39540 45966
rect 39488 45902 39540 45908
rect 39028 45824 39080 45830
rect 39028 45766 39080 45772
rect 39040 45286 39068 45766
rect 39212 45620 39264 45626
rect 39212 45562 39264 45568
rect 39028 45280 39080 45286
rect 39028 45222 39080 45228
rect 38844 45008 38896 45014
rect 38844 44950 38896 44956
rect 38568 44940 38620 44946
rect 38568 44882 38620 44888
rect 38476 44804 38528 44810
rect 38476 44746 38528 44752
rect 38488 44470 38516 44746
rect 38476 44464 38528 44470
rect 38476 44406 38528 44412
rect 38384 44396 38436 44402
rect 38384 44338 38436 44344
rect 38396 43790 38424 44338
rect 38488 43994 38516 44406
rect 38580 44402 38608 44882
rect 38660 44736 38712 44742
rect 38660 44678 38712 44684
rect 38672 44538 38700 44678
rect 38660 44532 38712 44538
rect 38660 44474 38712 44480
rect 38568 44396 38620 44402
rect 38568 44338 38620 44344
rect 38476 43988 38528 43994
rect 38476 43930 38528 43936
rect 38384 43784 38436 43790
rect 38384 43726 38436 43732
rect 38488 43450 38516 43930
rect 38856 43926 38884 44950
rect 39040 44402 39068 45222
rect 39224 45082 39252 45562
rect 40052 45082 40080 46378
rect 40316 45892 40368 45898
rect 40316 45834 40368 45840
rect 40328 45490 40356 45834
rect 40132 45484 40184 45490
rect 40132 45426 40184 45432
rect 40316 45484 40368 45490
rect 40316 45426 40368 45432
rect 40144 45082 40172 45426
rect 40420 45354 40448 49200
rect 40684 47048 40736 47054
rect 40684 46990 40736 46996
rect 40696 46889 40724 46990
rect 40682 46880 40738 46889
rect 40682 46815 40738 46824
rect 40788 45966 40816 49200
rect 41156 46442 41184 49200
rect 41236 47592 41288 47598
rect 41236 47534 41288 47540
rect 41248 46986 41276 47534
rect 41236 46980 41288 46986
rect 41236 46922 41288 46928
rect 41144 46436 41196 46442
rect 41144 46378 41196 46384
rect 41524 46170 41552 49200
rect 41892 47190 41920 49200
rect 41972 47456 42024 47462
rect 41972 47398 42024 47404
rect 41984 47190 42012 47398
rect 41880 47184 41932 47190
rect 41880 47126 41932 47132
rect 41972 47184 42024 47190
rect 41972 47126 42024 47132
rect 41696 46368 41748 46374
rect 41696 46310 41748 46316
rect 41512 46164 41564 46170
rect 41512 46106 41564 46112
rect 41708 46073 41736 46310
rect 42260 46170 42288 49200
rect 42628 46578 42656 49200
rect 42616 46572 42668 46578
rect 42616 46514 42668 46520
rect 42708 46504 42760 46510
rect 42708 46446 42760 46452
rect 42248 46164 42300 46170
rect 42248 46106 42300 46112
rect 41694 46064 41750 46073
rect 41694 45999 41750 46008
rect 40776 45960 40828 45966
rect 40776 45902 40828 45908
rect 40408 45348 40460 45354
rect 40408 45290 40460 45296
rect 40788 45082 40816 45902
rect 42720 45626 42748 46446
rect 42996 45937 43024 49200
rect 43364 47258 43392 49200
rect 43352 47252 43404 47258
rect 43352 47194 43404 47200
rect 43260 47048 43312 47054
rect 43260 46990 43312 46996
rect 43272 46714 43300 46990
rect 43260 46708 43312 46714
rect 43260 46650 43312 46656
rect 43916 46578 43944 49286
rect 44086 49200 44142 50000
rect 44454 49314 44510 50000
rect 44454 49286 44588 49314
rect 44454 49200 44510 49286
rect 44100 47258 44128 49200
rect 44088 47252 44140 47258
rect 44088 47194 44140 47200
rect 44100 46986 44128 47194
rect 44088 46980 44140 46986
rect 44088 46922 44140 46928
rect 43904 46572 43956 46578
rect 43904 46514 43956 46520
rect 44100 46170 44128 46922
rect 44560 46578 44588 49286
rect 44822 49200 44878 50000
rect 45190 49200 45246 50000
rect 45558 49314 45614 50000
rect 45558 49286 45876 49314
rect 45558 49200 45614 49286
rect 44836 47258 44864 49200
rect 44824 47252 44876 47258
rect 44824 47194 44876 47200
rect 44548 46572 44600 46578
rect 44548 46514 44600 46520
rect 45204 46510 45232 49200
rect 45848 47258 45876 49286
rect 45926 49200 45982 50000
rect 45940 47258 45968 49200
rect 45836 47252 45888 47258
rect 45836 47194 45888 47200
rect 45928 47252 45980 47258
rect 45928 47194 45980 47200
rect 45192 46504 45244 46510
rect 45192 46446 45244 46452
rect 44088 46164 44140 46170
rect 44088 46106 44140 46112
rect 42982 45928 43038 45937
rect 42982 45863 43038 45872
rect 42708 45620 42760 45626
rect 42708 45562 42760 45568
rect 41144 45280 41196 45286
rect 41144 45222 41196 45228
rect 39212 45076 39264 45082
rect 39212 45018 39264 45024
rect 40040 45076 40092 45082
rect 40040 45018 40092 45024
rect 40132 45076 40184 45082
rect 40132 45018 40184 45024
rect 40776 45076 40828 45082
rect 40776 45018 40828 45024
rect 40052 44470 40080 45018
rect 40144 44538 40172 45018
rect 41156 44878 41184 45222
rect 42720 45082 42748 45562
rect 42708 45076 42760 45082
rect 42708 45018 42760 45024
rect 41144 44872 41196 44878
rect 41144 44814 41196 44820
rect 42720 44538 42748 45018
rect 40132 44532 40184 44538
rect 40132 44474 40184 44480
rect 42708 44532 42760 44538
rect 42708 44474 42760 44480
rect 40040 44464 40092 44470
rect 40040 44406 40092 44412
rect 39028 44396 39080 44402
rect 39028 44338 39080 44344
rect 40144 43994 40172 44474
rect 40132 43988 40184 43994
rect 40132 43930 40184 43936
rect 38844 43920 38896 43926
rect 38844 43862 38896 43868
rect 38856 43450 38884 43862
rect 38476 43444 38528 43450
rect 38476 43386 38528 43392
rect 38844 43444 38896 43450
rect 38844 43386 38896 43392
rect 38200 43376 38252 43382
rect 38200 43318 38252 43324
rect 37556 43308 37608 43314
rect 37556 43250 37608 43256
rect 35992 42832 36044 42838
rect 35992 42774 36044 42780
rect 36004 42362 36032 42774
rect 38212 42770 38240 43318
rect 37280 42764 37332 42770
rect 37280 42706 37332 42712
rect 38200 42764 38252 42770
rect 38200 42706 38252 42712
rect 30932 42356 30984 42362
rect 30932 42298 30984 42304
rect 35716 42356 35768 42362
rect 35716 42298 35768 42304
rect 35992 42356 36044 42362
rect 35992 42298 36044 42304
rect 37292 42294 37320 42706
rect 30748 42288 30800 42294
rect 30748 42230 30800 42236
rect 37280 42288 37332 42294
rect 37280 42230 37332 42236
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 29656 6886 29776 6914
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 24400 6792 24452 6798
rect 24400 6734 24452 6740
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 22204 6322 22232 6598
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 4172 2938 4200 3470
rect 4080 2910 4200 2938
rect 4896 2916 4948 2922
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2608 800 2636 2382
rect 3160 800 3188 2790
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 3528 800 3556 2450
rect 3896 800 3924 2790
rect 4080 2564 4108 2910
rect 4896 2858 4948 2864
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4080 2536 4292 2564
rect 4264 800 4292 2536
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4632 800 4660 2382
rect 4908 800 4936 2858
rect 5184 800 5212 3470
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5460 800 5488 2926
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5736 800 5764 2382
rect 6012 800 6040 3470
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 6288 800 6316 2858
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6564 800 6592 2790
rect 6840 800 6868 3470
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7116 800 7144 2518
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 7392 800 7420 2314
rect 7668 800 7696 3470
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7944 800 7972 2926
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8220 800 8248 2450
rect 8496 800 8524 3470
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8772 800 8800 2858
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 9048 800 9076 2790
rect 9324 800 9352 3470
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9588 2576 9640 2582
rect 9588 2518 9640 2524
rect 9600 800 9628 2518
rect 9876 800 9904 2926
rect 10152 800 10180 3470
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10416 2508 10468 2514
rect 10416 2450 10468 2456
rect 10428 800 10456 2450
rect 10704 800 10732 2790
rect 10980 800 11008 3470
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11256 800 11284 2858
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 11532 800 11560 2518
rect 11808 800 11836 3470
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12084 800 12112 2790
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12268 800 12296 2382
rect 12544 800 12572 3470
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 12820 800 12848 2450
rect 13096 800 13124 3470
rect 13360 2916 13412 2922
rect 13360 2858 13412 2864
rect 13372 800 13400 2858
rect 13648 800 13676 3470
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13924 800 13952 2790
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 14200 800 14228 2518
rect 14476 800 14504 2858
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 14752 800 14780 2450
rect 15028 800 15056 3878
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 15304 800 15332 2926
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15580 800 15608 2382
rect 15856 800 15884 3538
rect 16132 800 16160 3878
rect 16948 3664 17000 3670
rect 16948 3606 17000 3612
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16408 800 16436 3470
rect 16672 2916 16724 2922
rect 16672 2858 16724 2864
rect 16684 800 16712 2858
rect 16960 800 16988 3606
rect 17236 800 17264 3878
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17408 2372 17460 2378
rect 17408 2314 17460 2320
rect 17420 1902 17448 2314
rect 17408 1896 17460 1902
rect 17408 1838 17460 1844
rect 17512 800 17540 2926
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 17788 800 17816 2450
rect 18064 800 18092 4558
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 18156 3194 18184 3674
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18512 3460 18564 3466
rect 18512 3402 18564 3408
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18328 2916 18380 2922
rect 18328 2858 18380 2864
rect 18340 800 18368 2858
rect 18524 1850 18552 3402
rect 18616 2990 18644 3470
rect 18708 3058 18736 3470
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18800 3126 18828 3334
rect 18788 3120 18840 3126
rect 18788 3062 18840 3068
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 18524 1822 18644 1850
rect 18616 800 18644 1822
rect 18892 800 18920 3878
rect 19352 3534 19380 5170
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19352 3058 19380 3334
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 19168 800 19196 2586
rect 19352 2446 19380 2994
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19444 800 19472 4966
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 1986 20024 4626
rect 20088 4554 20116 4966
rect 20364 4622 20392 5102
rect 20640 5098 20668 5646
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20824 5234 20852 5510
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20628 5092 20680 5098
rect 20628 5034 20680 5040
rect 20720 4752 20772 4758
rect 20720 4694 20772 4700
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20076 4548 20128 4554
rect 20076 4490 20128 4496
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 20180 4214 20208 4422
rect 20168 4208 20220 4214
rect 20168 4150 20220 4156
rect 20168 3664 20220 3670
rect 20168 3606 20220 3612
rect 20180 3058 20208 3606
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 19720 1958 20024 1986
rect 19720 800 19748 1958
rect 19984 1896 20036 1902
rect 19984 1838 20036 1844
rect 19996 800 20024 1838
rect 20272 800 20300 3538
rect 20364 3466 20392 4558
rect 20732 3942 20760 4694
rect 20916 4690 20944 6054
rect 21376 5778 21404 6054
rect 21916 5840 21968 5846
rect 21916 5782 21968 5788
rect 21364 5772 21416 5778
rect 21364 5714 21416 5720
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 21640 4548 21692 4554
rect 21640 4490 21692 4496
rect 20812 4208 20864 4214
rect 20812 4150 20864 4156
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20352 3460 20404 3466
rect 20352 3402 20404 3408
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 20548 800 20576 2790
rect 20640 2650 20668 3402
rect 20824 3398 20852 4150
rect 21088 4072 21140 4078
rect 21088 4014 21140 4020
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 20916 3534 20944 3878
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20904 3120 20956 3126
rect 20904 3062 20956 3068
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20916 2582 20944 3062
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20824 800 20852 2246
rect 21100 800 21128 4014
rect 21364 2984 21416 2990
rect 21364 2926 21416 2932
rect 21376 800 21404 2926
rect 21652 800 21680 4490
rect 21732 3732 21784 3738
rect 21732 3674 21784 3680
rect 21744 3466 21772 3674
rect 21732 3460 21784 3466
rect 21732 3402 21784 3408
rect 21928 800 21956 5782
rect 22020 4758 22048 6054
rect 22204 5302 22232 6258
rect 22192 5296 22244 5302
rect 22192 5238 22244 5244
rect 22296 5234 22324 6258
rect 23032 5302 23060 6734
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 23400 5642 23428 6054
rect 23848 5840 23900 5846
rect 23848 5782 23900 5788
rect 23388 5636 23440 5642
rect 23388 5578 23440 5584
rect 23020 5296 23072 5302
rect 23020 5238 23072 5244
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 22296 5098 22324 5170
rect 22284 5092 22336 5098
rect 22284 5034 22336 5040
rect 23572 5092 23624 5098
rect 23572 5034 23624 5040
rect 22008 4752 22060 4758
rect 22008 4694 22060 4700
rect 22020 4622 22048 4694
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22020 2378 22048 3130
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 22112 2650 22140 2790
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 22008 2372 22060 2378
rect 22008 2314 22060 2320
rect 22204 800 22232 4014
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 22480 800 22508 3402
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 22756 800 22784 2926
rect 23020 2508 23072 2514
rect 23020 2450 23072 2456
rect 23032 800 23060 2450
rect 23308 800 23336 4626
rect 23388 4072 23440 4078
rect 23388 4014 23440 4020
rect 23400 3738 23428 4014
rect 23388 3732 23440 3738
rect 23388 3674 23440 3680
rect 23584 800 23612 5034
rect 23768 4826 23796 5170
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 23768 3942 23796 4762
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23768 3534 23796 3878
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 23860 800 23888 5782
rect 24412 5234 24440 6734
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 24492 6384 24544 6390
rect 24492 6326 24544 6332
rect 24504 5370 24532 6326
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24688 5778 24716 6054
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24780 5642 24808 6598
rect 26700 6384 26752 6390
rect 26700 6326 26752 6332
rect 25964 6248 26016 6254
rect 25964 6190 26016 6196
rect 25228 6180 25280 6186
rect 25228 6122 25280 6128
rect 24952 5772 25004 5778
rect 24952 5714 25004 5720
rect 24768 5636 24820 5642
rect 24768 5578 24820 5584
rect 24492 5364 24544 5370
rect 24492 5306 24544 5312
rect 24400 5228 24452 5234
rect 24400 5170 24452 5176
rect 24308 4208 24360 4214
rect 24308 4150 24360 4156
rect 24320 3738 24348 4150
rect 24676 4004 24728 4010
rect 24676 3946 24728 3952
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 24136 3126 24164 3334
rect 24124 3120 24176 3126
rect 24124 3062 24176 3068
rect 24228 1714 24256 3538
rect 24400 2984 24452 2990
rect 24400 2926 24452 2932
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 24136 1686 24256 1714
rect 24136 800 24164 1686
rect 24412 800 24440 2926
rect 24504 2650 24532 2926
rect 24492 2644 24544 2650
rect 24492 2586 24544 2592
rect 24688 800 24716 3946
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 24872 2514 24900 3062
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 24964 800 24992 5714
rect 25044 3460 25096 3466
rect 25044 3402 25096 3408
rect 25056 2446 25084 3402
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 25240 800 25268 6122
rect 25976 5914 26004 6190
rect 26516 6180 26568 6186
rect 26516 6122 26568 6128
rect 25964 5908 26016 5914
rect 25964 5850 26016 5856
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25700 4758 25728 5646
rect 25780 5296 25832 5302
rect 25780 5238 25832 5244
rect 25792 4826 25820 5238
rect 26332 5092 26384 5098
rect 26332 5034 26384 5040
rect 25780 4820 25832 4826
rect 25780 4762 25832 4768
rect 25688 4752 25740 4758
rect 25688 4694 25740 4700
rect 25700 4622 25728 4694
rect 25688 4616 25740 4622
rect 25688 4558 25740 4564
rect 25504 4208 25556 4214
rect 25504 4150 25556 4156
rect 25516 3738 25544 4150
rect 25504 3732 25556 3738
rect 25504 3674 25556 3680
rect 25700 3534 25728 4558
rect 26056 4072 26108 4078
rect 26056 4014 26108 4020
rect 25688 3528 25740 3534
rect 25688 3470 25740 3476
rect 25504 2984 25556 2990
rect 25504 2926 25556 2932
rect 25516 800 25544 2926
rect 25780 2508 25832 2514
rect 25780 2450 25832 2456
rect 25792 800 25820 2450
rect 26068 800 26096 4014
rect 26344 800 26372 5034
rect 26528 2938 26556 6122
rect 26712 5914 26740 6326
rect 28172 6316 28224 6322
rect 28172 6258 28224 6264
rect 27436 6112 27488 6118
rect 27436 6054 27488 6060
rect 27804 6112 27856 6118
rect 27804 6054 27856 6060
rect 26700 5908 26752 5914
rect 26700 5850 26752 5856
rect 27448 5778 27476 6054
rect 27436 5772 27488 5778
rect 27436 5714 27488 5720
rect 27528 5636 27580 5642
rect 27528 5578 27580 5584
rect 27540 4826 27568 5578
rect 27816 5302 27844 6054
rect 27988 5840 28040 5846
rect 27988 5782 28040 5788
rect 27804 5296 27856 5302
rect 27804 5238 27856 5244
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 27528 4820 27580 4826
rect 27528 4762 27580 4768
rect 27344 4208 27396 4214
rect 27344 4150 27396 4156
rect 26608 4072 26660 4078
rect 26608 4014 26660 4020
rect 26620 3058 26648 4014
rect 27160 3596 27212 3602
rect 27160 3538 27212 3544
rect 26608 3052 26660 3058
rect 26608 2994 26660 3000
rect 26884 2984 26936 2990
rect 26528 2910 26648 2938
rect 26884 2926 26936 2932
rect 26620 800 26648 2910
rect 26896 800 26924 2926
rect 27172 800 27200 3538
rect 27356 2650 27384 4150
rect 27436 4072 27488 4078
rect 27436 4014 27488 4020
rect 27344 2644 27396 2650
rect 27344 2586 27396 2592
rect 27448 800 27476 4014
rect 27632 2394 27660 5102
rect 27896 4616 27948 4622
rect 27896 4558 27948 4564
rect 27712 3120 27764 3126
rect 27712 3062 27764 3068
rect 27724 2582 27752 3062
rect 27804 2984 27856 2990
rect 27804 2926 27856 2932
rect 27816 2650 27844 2926
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 27712 2576 27764 2582
rect 27712 2518 27764 2524
rect 27908 2446 27936 4558
rect 27896 2440 27948 2446
rect 27632 2366 27752 2394
rect 27896 2382 27948 2388
rect 27724 800 27752 2366
rect 28000 800 28028 5782
rect 28184 4622 28212 6258
rect 29092 5024 29144 5030
rect 29092 4966 29144 4972
rect 29104 4690 29132 4966
rect 28816 4684 28868 4690
rect 28816 4626 28868 4632
rect 29092 4684 29144 4690
rect 29092 4626 29144 4632
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 28264 3596 28316 3602
rect 28264 3538 28316 3544
rect 28172 3460 28224 3466
rect 28172 3402 28224 3408
rect 28184 2582 28212 3402
rect 28172 2576 28224 2582
rect 28172 2518 28224 2524
rect 28276 800 28304 3538
rect 28356 3392 28408 3398
rect 28356 3334 28408 3340
rect 28368 2650 28396 3334
rect 28540 2984 28592 2990
rect 28540 2926 28592 2932
rect 28356 2644 28408 2650
rect 28356 2586 28408 2592
rect 28552 800 28580 2926
rect 28828 800 28856 4626
rect 29092 4072 29144 4078
rect 29092 4014 29144 4020
rect 29104 800 29132 4014
rect 29368 2984 29420 2990
rect 29368 2926 29420 2932
rect 29380 800 29408 2926
rect 29656 800 29684 6886
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 30380 4480 30432 4486
rect 30432 4428 30512 4434
rect 30380 4422 30512 4428
rect 30392 4406 30512 4422
rect 30484 4146 30512 4406
rect 30472 4140 30524 4146
rect 30472 4082 30524 4088
rect 30484 3670 30512 4082
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 30472 3664 30524 3670
rect 30472 3606 30524 3612
rect 31392 3664 31444 3670
rect 31392 3606 31444 3612
rect 32956 3664 33008 3670
rect 32956 3606 33008 3612
rect 36820 3664 36872 3670
rect 36820 3606 36872 3612
rect 30196 3596 30248 3602
rect 30196 3538 30248 3544
rect 30012 3528 30064 3534
rect 30012 3470 30064 3476
rect 30024 3126 30052 3470
rect 30012 3120 30064 3126
rect 30012 3062 30064 3068
rect 29920 2576 29972 2582
rect 29920 2518 29972 2524
rect 29932 800 29960 2518
rect 30208 800 30236 3538
rect 31116 3528 31168 3534
rect 31116 3470 31168 3476
rect 30748 3460 30800 3466
rect 30748 3402 30800 3408
rect 30288 3188 30340 3194
rect 30288 3130 30340 3136
rect 30300 2650 30328 3130
rect 30760 3058 30788 3402
rect 30748 3052 30800 3058
rect 30748 2994 30800 3000
rect 31024 2984 31076 2990
rect 31024 2926 31076 2932
rect 30748 2848 30800 2854
rect 30748 2790 30800 2796
rect 30288 2644 30340 2650
rect 30288 2586 30340 2592
rect 30472 2372 30524 2378
rect 30472 2314 30524 2320
rect 30484 800 30512 2314
rect 30760 800 30788 2790
rect 31036 2650 31064 2926
rect 31024 2644 31076 2650
rect 31024 2586 31076 2592
rect 31128 1850 31156 3470
rect 31404 3058 31432 3606
rect 31852 3528 31904 3534
rect 31852 3470 31904 3476
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 31392 3052 31444 3058
rect 31392 2994 31444 3000
rect 31300 2508 31352 2514
rect 31300 2450 31352 2456
rect 31036 1822 31156 1850
rect 31036 800 31064 1822
rect 31312 800 31340 2450
rect 31404 2446 31432 2994
rect 31576 2916 31628 2922
rect 31576 2858 31628 2864
rect 31392 2440 31444 2446
rect 31392 2382 31444 2388
rect 31588 800 31616 2858
rect 31864 800 31892 3470
rect 32128 2984 32180 2990
rect 32128 2926 32180 2932
rect 32140 800 32168 2926
rect 32416 800 32444 3470
rect 32680 3052 32732 3058
rect 32680 2994 32732 3000
rect 32692 800 32720 2994
rect 32968 800 32996 3606
rect 34796 3596 34848 3602
rect 34796 3538 34848 3544
rect 34336 3528 34388 3534
rect 34336 3470 34388 3476
rect 34060 2984 34112 2990
rect 34060 2926 34112 2932
rect 33508 2916 33560 2922
rect 33508 2858 33560 2864
rect 33232 2576 33284 2582
rect 33232 2518 33284 2524
rect 33244 800 33272 2518
rect 33520 800 33548 2858
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 33796 800 33824 2382
rect 34072 800 34100 2926
rect 34348 800 34376 3470
rect 34612 2508 34664 2514
rect 34612 2450 34664 2456
rect 34624 800 34652 2450
rect 34808 1850 34836 3538
rect 35716 3528 35768 3534
rect 35716 3470 35768 3476
rect 36268 3528 36320 3534
rect 36268 3470 36320 3476
rect 35348 2916 35400 2922
rect 35348 2858 35400 2864
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34808 1822 34928 1850
rect 34900 800 34928 1822
rect 35360 1442 35388 2858
rect 35440 2576 35492 2582
rect 35440 2518 35492 2524
rect 35176 1414 35388 1442
rect 35176 800 35204 1414
rect 35452 800 35480 2518
rect 35728 800 35756 3470
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36004 800 36032 2790
rect 36280 800 36308 3470
rect 36544 2440 36596 2446
rect 36544 2382 36596 2388
rect 36556 800 36584 2382
rect 36832 800 36860 3606
rect 37648 3528 37700 3534
rect 37648 3470 37700 3476
rect 38200 3528 38252 3534
rect 38200 3470 38252 3476
rect 39580 3528 39632 3534
rect 39580 3470 39632 3476
rect 40408 3528 40460 3534
rect 40408 3470 40460 3476
rect 40960 3528 41012 3534
rect 40960 3470 41012 3476
rect 41512 3528 41564 3534
rect 41512 3470 41564 3476
rect 42892 3528 42944 3534
rect 42892 3470 42944 3476
rect 43168 3528 43220 3534
rect 43168 3470 43220 3476
rect 44824 3528 44876 3534
rect 44824 3470 44876 3476
rect 45652 3528 45704 3534
rect 45652 3470 45704 3476
rect 46480 3528 46532 3534
rect 46480 3470 46532 3476
rect 46756 3528 46808 3534
rect 46756 3470 46808 3476
rect 47308 3528 47360 3534
rect 47308 3470 47360 3476
rect 37096 2984 37148 2990
rect 37096 2926 37148 2932
rect 37108 800 37136 2926
rect 37372 2508 37424 2514
rect 37372 2450 37424 2456
rect 37384 800 37412 2450
rect 37660 800 37688 3470
rect 37924 2916 37976 2922
rect 37924 2858 37976 2864
rect 37936 800 37964 2858
rect 38212 800 38240 3470
rect 38752 2984 38804 2990
rect 38752 2926 38804 2932
rect 38476 2576 38528 2582
rect 38476 2518 38528 2524
rect 38488 800 38516 2518
rect 38764 800 38792 2926
rect 39028 2848 39080 2854
rect 39028 2790 39080 2796
rect 39040 800 39068 2790
rect 39304 2508 39356 2514
rect 39304 2450 39356 2456
rect 39316 800 39344 2450
rect 39592 800 39620 3470
rect 40132 2848 40184 2854
rect 40132 2790 40184 2796
rect 39856 2440 39908 2446
rect 39856 2382 39908 2388
rect 39868 800 39896 2382
rect 40144 800 40172 2790
rect 40420 800 40448 3470
rect 40684 2984 40736 2990
rect 40684 2926 40736 2932
rect 40696 800 40724 2926
rect 40972 800 41000 3470
rect 41236 2508 41288 2514
rect 41236 2450 41288 2456
rect 41248 800 41276 2450
rect 41524 800 41552 3470
rect 42616 2984 42668 2990
rect 42616 2926 42668 2932
rect 42064 2848 42116 2854
rect 42064 2790 42116 2796
rect 41788 2440 41840 2446
rect 41788 2382 41840 2388
rect 41800 800 41828 2382
rect 42076 800 42104 2790
rect 42340 2576 42392 2582
rect 42340 2518 42392 2524
rect 42352 800 42380 2518
rect 42628 800 42656 2926
rect 42904 800 42932 3470
rect 43180 800 43208 3470
rect 44548 2984 44600 2990
rect 44548 2926 44600 2932
rect 43444 2848 43496 2854
rect 43444 2790 43496 2796
rect 43996 2848 44048 2854
rect 43996 2790 44048 2796
rect 43456 800 43484 2790
rect 43720 2508 43772 2514
rect 43720 2450 43772 2456
rect 43732 800 43760 2450
rect 44008 800 44036 2790
rect 44272 2372 44324 2378
rect 44272 2314 44324 2320
rect 44284 800 44312 2314
rect 44560 800 44588 2926
rect 44836 800 44864 3470
rect 45376 2848 45428 2854
rect 45376 2790 45428 2796
rect 45100 2576 45152 2582
rect 45100 2518 45152 2524
rect 45112 800 45140 2518
rect 45388 800 45416 2790
rect 45664 800 45692 3470
rect 45928 2848 45980 2854
rect 45928 2790 45980 2796
rect 45940 800 45968 2790
rect 46204 2440 46256 2446
rect 46204 2382 46256 2388
rect 46216 800 46244 2382
rect 46492 800 46520 3470
rect 46768 800 46796 3470
rect 47032 2848 47084 2854
rect 47032 2790 47084 2796
rect 47044 800 47072 2790
rect 47320 800 47348 3470
rect 2410 0 2466 800
rect 2502 0 2558 800
rect 2594 0 2650 800
rect 2686 0 2742 800
rect 2778 0 2834 800
rect 2870 0 2926 800
rect 2962 0 3018 800
rect 3054 0 3110 800
rect 3146 0 3202 800
rect 3238 0 3294 800
rect 3330 0 3386 800
rect 3422 0 3478 800
rect 3514 0 3570 800
rect 3606 0 3662 800
rect 3698 0 3754 800
rect 3790 0 3846 800
rect 3882 0 3938 800
rect 3974 0 4030 800
rect 4066 0 4122 800
rect 4158 0 4214 800
rect 4250 0 4306 800
rect 4342 0 4398 800
rect 4434 0 4490 800
rect 4526 0 4582 800
rect 4618 0 4674 800
rect 4710 0 4766 800
rect 4802 0 4858 800
rect 4894 0 4950 800
rect 4986 0 5042 800
rect 5078 0 5134 800
rect 5170 0 5226 800
rect 5262 0 5318 800
rect 5354 0 5410 800
rect 5446 0 5502 800
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5722 0 5778 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6366 0 6422 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6642 0 6698 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7010 0 7066 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
<< via2 >>
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 9494 46144 9550 46200
rect 18878 46416 18934 46472
rect 17866 45872 17922 45928
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 20074 46552 20130 46608
rect 20258 46572 20314 46608
rect 20258 46552 20260 46572
rect 20260 46552 20312 46572
rect 20312 46552 20314 46572
rect 19338 46316 19346 46336
rect 19346 46316 19394 46336
rect 19338 46280 19394 46316
rect 19338 46044 19346 46064
rect 19346 46044 19394 46064
rect 19338 46008 19394 46044
rect 20074 46316 20076 46336
rect 20076 46316 20128 46336
rect 20128 46316 20130 46336
rect 20074 46280 20130 46316
rect 20074 46044 20076 46064
rect 20076 46044 20128 46064
rect 20128 46044 20130 46064
rect 20074 46008 20130 46044
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 20350 45872 20406 45928
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 22098 46144 22154 46200
rect 21914 45736 21970 45792
rect 22834 45908 22836 45928
rect 22836 45908 22888 45928
rect 22888 45908 22890 45928
rect 22834 45872 22890 45908
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 23662 46144 23718 46200
rect 23570 45872 23626 45928
rect 23294 45772 23296 45792
rect 23296 45772 23348 45792
rect 23348 45772 23350 45792
rect 23294 45736 23350 45772
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 28814 46688 28870 46744
rect 29090 45872 29146 45928
rect 30286 46280 30342 46336
rect 30562 46144 30618 46200
rect 31666 46688 31722 46744
rect 32494 46280 32550 46336
rect 32310 44920 32366 44976
rect 33874 47096 33930 47152
rect 34610 46688 34666 46744
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34334 46452 34336 46472
rect 34336 46452 34388 46472
rect 34388 46452 34390 46472
rect 34334 46416 34390 46452
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34610 45736 34666 45792
rect 35714 47096 35770 47152
rect 35622 46824 35678 46880
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 35898 46996 35900 47016
rect 35900 46996 35952 47016
rect 35952 46996 35954 47016
rect 35898 46960 35954 46996
rect 37370 46552 37426 46608
rect 37186 46416 37242 46472
rect 36818 46280 36874 46336
rect 36726 46008 36782 46064
rect 37738 47116 37794 47152
rect 37738 47096 37740 47116
rect 37740 47096 37792 47116
rect 37792 47096 37794 47116
rect 36726 44920 36782 44976
rect 38290 46436 38346 46472
rect 38290 46416 38292 46436
rect 38292 46416 38344 46436
rect 38344 46416 38346 46436
rect 38106 45736 38162 45792
rect 38474 46280 38530 46336
rect 40130 46688 40186 46744
rect 40682 46824 40738 46880
rect 41694 46008 41750 46064
rect 42982 45872 43038 45928
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
<< metal3 >>
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 33869 47154 33935 47157
rect 35709 47154 35775 47157
rect 37733 47154 37799 47157
rect 33869 47152 37799 47154
rect 33869 47096 33874 47152
rect 33930 47096 35714 47152
rect 35770 47096 37738 47152
rect 37794 47096 37799 47152
rect 33869 47094 37799 47096
rect 33869 47091 33935 47094
rect 35709 47091 35775 47094
rect 37733 47091 37799 47094
rect 35893 47018 35959 47021
rect 35390 47016 35959 47018
rect 35390 46960 35898 47016
rect 35954 46960 35959 47016
rect 35390 46958 35959 46960
rect 35390 46882 35450 46958
rect 35893 46955 35959 46958
rect 34470 46822 35450 46882
rect 35617 46882 35683 46885
rect 40677 46882 40743 46885
rect 35617 46880 40743 46882
rect 35617 46824 35622 46880
rect 35678 46824 40682 46880
rect 40738 46824 40743 46880
rect 35617 46822 40743 46824
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 28809 46746 28875 46749
rect 31661 46746 31727 46749
rect 34470 46746 34530 46822
rect 35617 46819 35683 46822
rect 40677 46819 40743 46822
rect 28809 46744 34530 46746
rect 28809 46688 28814 46744
rect 28870 46688 31666 46744
rect 31722 46688 34530 46744
rect 28809 46686 34530 46688
rect 34605 46746 34671 46749
rect 40125 46746 40191 46749
rect 34605 46744 40191 46746
rect 34605 46688 34610 46744
rect 34666 46688 40130 46744
rect 40186 46688 40191 46744
rect 34605 46686 40191 46688
rect 28809 46683 28875 46686
rect 31661 46683 31727 46686
rect 34605 46683 34671 46686
rect 40125 46683 40191 46686
rect 20069 46610 20135 46613
rect 20253 46610 20319 46613
rect 37365 46610 37431 46613
rect 20069 46608 20178 46610
rect 20069 46552 20074 46608
rect 20130 46552 20178 46608
rect 20069 46547 20178 46552
rect 20253 46608 37431 46610
rect 20253 46552 20258 46608
rect 20314 46552 37370 46608
rect 37426 46552 37431 46608
rect 20253 46550 37431 46552
rect 20253 46547 20319 46550
rect 37365 46547 37431 46550
rect 18873 46474 18939 46477
rect 20118 46474 20178 46547
rect 34329 46474 34395 46477
rect 18873 46472 34395 46474
rect 18873 46416 18878 46472
rect 18934 46416 34334 46472
rect 34390 46416 34395 46472
rect 18873 46414 34395 46416
rect 18873 46411 18939 46414
rect 34329 46411 34395 46414
rect 37181 46474 37247 46477
rect 38285 46474 38351 46477
rect 37181 46472 38351 46474
rect 37181 46416 37186 46472
rect 37242 46416 38290 46472
rect 38346 46416 38351 46472
rect 37181 46414 38351 46416
rect 37181 46411 37247 46414
rect 38285 46411 38351 46414
rect 19333 46338 19399 46341
rect 20069 46338 20135 46341
rect 19333 46336 20135 46338
rect 19333 46280 19338 46336
rect 19394 46280 20074 46336
rect 20130 46280 20135 46336
rect 19333 46278 20135 46280
rect 19333 46275 19399 46278
rect 20069 46275 20135 46278
rect 30281 46338 30347 46341
rect 32489 46338 32555 46341
rect 30281 46336 32555 46338
rect 30281 46280 30286 46336
rect 30342 46280 32494 46336
rect 32550 46280 32555 46336
rect 30281 46278 32555 46280
rect 30281 46275 30347 46278
rect 32489 46275 32555 46278
rect 36813 46338 36879 46341
rect 38469 46338 38535 46341
rect 36813 46336 38535 46338
rect 36813 46280 36818 46336
rect 36874 46280 38474 46336
rect 38530 46280 38535 46336
rect 36813 46278 38535 46280
rect 36813 46275 36879 46278
rect 38469 46275 38535 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 9489 46202 9555 46205
rect 22093 46202 22159 46205
rect 9489 46200 22159 46202
rect 9489 46144 9494 46200
rect 9550 46144 22098 46200
rect 22154 46144 22159 46200
rect 9489 46142 22159 46144
rect 9489 46139 9555 46142
rect 22093 46139 22159 46142
rect 23657 46202 23723 46205
rect 30557 46202 30623 46205
rect 23657 46200 30623 46202
rect 23657 46144 23662 46200
rect 23718 46144 30562 46200
rect 30618 46144 30623 46200
rect 23657 46142 30623 46144
rect 23657 46139 23723 46142
rect 30557 46139 30623 46142
rect 19333 46066 19399 46069
rect 20069 46066 20135 46069
rect 19333 46064 20135 46066
rect 19333 46008 19338 46064
rect 19394 46008 20074 46064
rect 20130 46008 20135 46064
rect 19333 46006 20135 46008
rect 19333 46003 19399 46006
rect 20069 46003 20135 46006
rect 36721 46066 36787 46069
rect 41689 46066 41755 46069
rect 36721 46064 41755 46066
rect 36721 46008 36726 46064
rect 36782 46008 41694 46064
rect 41750 46008 41755 46064
rect 36721 46006 41755 46008
rect 36721 46003 36787 46006
rect 41689 46003 41755 46006
rect 17861 45930 17927 45933
rect 20345 45930 20411 45933
rect 17861 45928 20411 45930
rect 17861 45872 17866 45928
rect 17922 45872 20350 45928
rect 20406 45872 20411 45928
rect 17861 45870 20411 45872
rect 17861 45867 17927 45870
rect 20345 45867 20411 45870
rect 22829 45930 22895 45933
rect 23565 45930 23631 45933
rect 22829 45928 23631 45930
rect 22829 45872 22834 45928
rect 22890 45872 23570 45928
rect 23626 45872 23631 45928
rect 22829 45870 23631 45872
rect 22829 45867 22895 45870
rect 23565 45867 23631 45870
rect 29085 45930 29151 45933
rect 42977 45930 43043 45933
rect 29085 45928 43043 45930
rect 29085 45872 29090 45928
rect 29146 45872 42982 45928
rect 43038 45872 43043 45928
rect 29085 45870 43043 45872
rect 29085 45867 29151 45870
rect 42977 45867 43043 45870
rect 21909 45794 21975 45797
rect 23289 45794 23355 45797
rect 21909 45792 23355 45794
rect 21909 45736 21914 45792
rect 21970 45736 23294 45792
rect 23350 45736 23355 45792
rect 21909 45734 23355 45736
rect 21909 45731 21975 45734
rect 23289 45731 23355 45734
rect 34605 45794 34671 45797
rect 38101 45794 38167 45797
rect 34605 45792 38167 45794
rect 34605 45736 34610 45792
rect 34666 45736 38106 45792
rect 38162 45736 38167 45792
rect 34605 45734 38167 45736
rect 34605 45731 34671 45734
rect 38101 45731 38167 45734
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 32305 44978 32371 44981
rect 36721 44978 36787 44981
rect 32305 44976 36787 44978
rect 32305 44920 32310 44976
rect 32366 44920 36726 44976
rect 36782 44920 36787 44976
rect 32305 44918 36787 44920
rect 32305 44915 32371 44918
rect 36721 44915 36787 44918
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 21804 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A
timestamp 1666199351
transform 1 0 22356 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A
timestamp 1666199351
transform -1 0 20240 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A
timestamp 1666199351
transform -1 0 29900 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A_N
timestamp 1666199351
transform -1 0 29900 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__B
timestamp 1666199351
transform 1 0 36800 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A1
timestamp 1666199351
transform -1 0 30912 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A2
timestamp 1666199351
transform -1 0 29992 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A
timestamp 1666199351
transform 1 0 31372 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A
timestamp 1666199351
transform 1 0 22356 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A1
timestamp 1666199351
transform 1 0 30820 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1666199351
transform 1 0 30268 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1666199351
transform -1 0 23092 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A
timestamp 1666199351
transform -1 0 32476 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A1
timestamp 1666199351
transform 1 0 30268 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__B1_N
timestamp 1666199351
transform -1 0 33028 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__B1
timestamp 1666199351
transform 1 0 28428 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A
timestamp 1666199351
transform 1 0 24288 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A
timestamp 1666199351
transform 1 0 27692 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A
timestamp 1666199351
transform -1 0 17020 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A
timestamp 1666199351
transform -1 0 24748 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A1
timestamp 1666199351
transform 1 0 29256 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A
timestamp 1666199351
transform 1 0 25668 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1666199351
transform -1 0 40204 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A_N
timestamp 1666199351
transform 1 0 42596 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__B
timestamp 1666199351
transform -1 0 40848 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A1
timestamp 1666199351
transform 1 0 38548 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A2
timestamp 1666199351
transform -1 0 41676 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A
timestamp 1666199351
transform 1 0 39376 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1666199351
transform -1 0 32936 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A1
timestamp 1666199351
transform 1 0 39008 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A
timestamp 1666199351
transform 1 0 36524 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A
timestamp 1666199351
transform 1 0 34868 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1666199351
transform 1 0 41124 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A1
timestamp 1666199351
transform 1 0 39560 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__B1_N
timestamp 1666199351
transform -1 0 40756 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A1
timestamp 1666199351
transform -1 0 38180 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__B1_N
timestamp 1666199351
transform 1 0 40112 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__B1
timestamp 1666199351
transform -1 0 37628 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A
timestamp 1666199351
transform 1 0 35972 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A
timestamp 1666199351
transform 1 0 38456 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A
timestamp 1666199351
transform -1 0 31832 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A
timestamp 1666199351
transform -1 0 33488 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A1
timestamp 1666199351
transform -1 0 41860 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1666199351
transform -1 0 41400 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__B1
timestamp 1666199351
transform -1 0 21252 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A
timestamp 1666199351
transform 1 0 28244 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A2_N
timestamp 1666199351
transform -1 0 26404 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__B2
timestamp 1666199351
transform -1 0 27324 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A2
timestamp 1666199351
transform -1 0 25300 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A3
timestamp 1666199351
transform -1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A
timestamp 1666199351
transform 1 0 42228 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A2_N
timestamp 1666199351
transform -1 0 36156 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__B2
timestamp 1666199351
transform 1 0 40020 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A2
timestamp 1666199351
transform -1 0 36340 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__A3
timestamp 1666199351
transform 1 0 34868 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1666199351
transform 1 0 20516 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1666199351
transform 1 0 31924 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A2
timestamp 1666199351
transform 1 0 28980 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__B1
timestamp 1666199351
transform -1 0 27876 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A
timestamp 1666199351
transform -1 0 44712 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A2
timestamp 1666199351
transform 1 0 43240 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__B1
timestamp 1666199351
transform -1 0 39284 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__B
timestamp 1666199351
transform -1 0 16836 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A2_N
timestamp 1666199351
transform -1 0 17756 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__A2
timestamp 1666199351
transform 1 0 25668 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__B1
timestamp 1666199351
transform 1 0 27140 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__B
timestamp 1666199351
transform -1 0 26404 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__A
timestamp 1666199351
transform -1 0 25852 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__B1
timestamp 1666199351
transform -1 0 24932 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__A1
timestamp 1666199351
transform 1 0 27140 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A2
timestamp 1666199351
transform -1 0 35604 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__B1
timestamp 1666199351
transform -1 0 35604 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__B
timestamp 1666199351
transform 1 0 35052 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A
timestamp 1666199351
transform -1 0 34040 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__A1
timestamp 1666199351
transform -1 0 23276 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__B1
timestamp 1666199351
transform -1 0 25300 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A1
timestamp 1666199351
transform -1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__A1
timestamp 1666199351
transform -1 0 34316 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__B1
timestamp 1666199351
transform -1 0 42136 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A1
timestamp 1666199351
transform 1 0 35604 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__C1
timestamp 1666199351
transform 1 0 22908 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19
timestamp 1666199351
transform 1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40
timestamp 1666199351
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47
timestamp 1666199351
transform 1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1666199351
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1666199351
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1666199351
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1666199351
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1666199351
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1666199351
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1666199351
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1666199351
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1666199351
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1666199351
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124
timestamp 1666199351
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 1666199351
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1666199351
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1666199351
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152
timestamp 1666199351
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_159
timestamp 1666199351
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1666199351
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1666199351
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_180
timestamp 1666199351
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1666199351
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1666199351
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1666199351
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_208
timestamp 1666199351
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_215
timestamp 1666199351
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1666199351
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1666199351
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1666199351
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1666199351
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1666199351
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1666199351
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1666199351
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_271
timestamp 1666199351
transform 1 0 26036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1666199351
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1666199351
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1666199351
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_293
timestamp 1666199351
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_300
timestamp 1666199351
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1666199351
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 1666199351
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1666199351
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 1666199351
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666199351
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_342
timestamp 1666199351
transform 1 0 32568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1666199351
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1666199351
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1666199351
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_370
timestamp 1666199351
transform 1 0 35144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1666199351
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1666199351
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1666199351
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_398
timestamp 1666199351
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_405
timestamp 1666199351
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1666199351
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1666199351
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_426
timestamp 1666199351
transform 1 0 40296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_433
timestamp 1666199351
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_440
timestamp 1666199351
transform 1 0 41584 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1666199351
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_454
timestamp 1666199351
transform 1 0 42872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1666199351
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_468
timestamp 1666199351
transform 1 0 44160 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1666199351
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_482
timestamp 1666199351
transform 1 0 45448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1666199351
transform 1 0 46092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_496
timestamp 1666199351
transform 1 0 46736 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1666199351
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_510
timestamp 1666199351
transform 1 0 48024 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_15 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_19
timestamp 1666199351
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1666199351
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_33
timestamp 1666199351
transform 1 0 4140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1666199351
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_47
timestamp 1666199351
transform 1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1666199351
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1666199351
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_68
timestamp 1666199351
transform 1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1666199351
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1666199351
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_89
timestamp 1666199351
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1666199351
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1666199351
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1666199351
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1666199351
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_124
timestamp 1666199351
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_131
timestamp 1666199351
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_138
timestamp 1666199351
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1666199351
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_152
timestamp 1666199351
transform 1 0 15088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_159
timestamp 1666199351
transform 1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1666199351
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_169
timestamp 1666199351
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1666199351
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1666199351
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_194
timestamp 1666199351
transform 1 0 18952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1666199351
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1666199351
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1666199351
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_242
timestamp 1666199351
transform 1 0 23368 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_257
timestamp 1666199351
transform 1 0 24748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_270
timestamp 1666199351
transform 1 0 25944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_274
timestamp 1666199351
transform 1 0 26312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1666199351
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1666199351
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_292
timestamp 1666199351
transform 1 0 27968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_305
timestamp 1666199351
transform 1 0 29164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_318
timestamp 1666199351
transform 1 0 30360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_325
timestamp 1666199351
transform 1 0 31004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1666199351
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1666199351
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_342
timestamp 1666199351
transform 1 0 32568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_349
timestamp 1666199351
transform 1 0 33212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_356
timestamp 1666199351
transform 1 0 33856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_363
timestamp 1666199351
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_370
timestamp 1666199351
transform 1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_377
timestamp 1666199351
transform 1 0 35788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_384
timestamp 1666199351
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1666199351
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_398
timestamp 1666199351
transform 1 0 37720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_405
timestamp 1666199351
transform 1 0 38364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_412
timestamp 1666199351
transform 1 0 39008 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_419
timestamp 1666199351
transform 1 0 39652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_426
timestamp 1666199351
transform 1 0 40296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_433
timestamp 1666199351
transform 1 0 40940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_440
timestamp 1666199351
transform 1 0 41584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1666199351
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_454
timestamp 1666199351
transform 1 0 42872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1666199351
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_468
timestamp 1666199351
transform 1 0 44160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_475
timestamp 1666199351
transform 1 0 44804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_482
timestamp 1666199351
transform 1 0 45448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_489
timestamp 1666199351
transform 1 0 46092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_496
timestamp 1666199351
transform 1 0 46736 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1666199351
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_510
timestamp 1666199351
transform 1 0 48024 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666199351
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666199351
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666199351
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp 1666199351
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_35
timestamp 1666199351
transform 1 0 4324 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1666199351
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_45
timestamp 1666199351
transform 1 0 5244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_54
timestamp 1666199351
transform 1 0 6072 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_63
timestamp 1666199351
transform 1 0 6900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_72
timestamp 1666199351
transform 1 0 7728 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1666199351
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1666199351
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_90
timestamp 1666199351
transform 1 0 9384 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_99
timestamp 1666199351
transform 1 0 10212 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1666199351
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_112
timestamp 1666199351
transform 1 0 11408 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_116
timestamp 1666199351
transform 1 0 11776 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_123
timestamp 1666199351
transform 1 0 12420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_130
timestamp 1666199351
transform 1 0 13064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1666199351
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1666199351
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_152
timestamp 1666199351
transform 1 0 15088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1666199351
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1666199351
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1666199351
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1666199351
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_187
timestamp 1666199351
transform 1 0 18308 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1666199351
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1666199351
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_204
timestamp 1666199351
transform 1 0 19872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_211
timestamp 1666199351
transform 1 0 20516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_218
timestamp 1666199351
transform 1 0 21160 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_231
timestamp 1666199351
transform 1 0 22356 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_239
timestamp 1666199351
transform 1 0 23092 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_243
timestamp 1666199351
transform 1 0 23460 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1666199351
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1666199351
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_264
timestamp 1666199351
transform 1 0 25392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_271
timestamp 1666199351
transform 1 0 26036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_277
timestamp 1666199351
transform 1 0 26588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_287
timestamp 1666199351
transform 1 0 27508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp 1666199351
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1666199351
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_314
timestamp 1666199351
transform 1 0 29992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1666199351
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_328
timestamp 1666199351
transform 1 0 31280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_335
timestamp 1666199351
transform 1 0 31924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_342
timestamp 1666199351
transform 1 0 32568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_349
timestamp 1666199351
transform 1 0 33212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp 1666199351
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1666199351
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_370
timestamp 1666199351
transform 1 0 35144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_377
timestamp 1666199351
transform 1 0 35788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_384
timestamp 1666199351
transform 1 0 36432 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_391
timestamp 1666199351
transform 1 0 37076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_398
timestamp 1666199351
transform 1 0 37720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_405
timestamp 1666199351
transform 1 0 38364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_412
timestamp 1666199351
transform 1 0 39008 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1666199351
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_426
timestamp 1666199351
transform 1 0 40296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_433
timestamp 1666199351
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_440
timestamp 1666199351
transform 1 0 41584 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_447
timestamp 1666199351
transform 1 0 42228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_451
timestamp 1666199351
transform 1 0 42596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_455
timestamp 1666199351
transform 1 0 42964 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_462
timestamp 1666199351
transform 1 0 43608 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1666199351
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1666199351
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_482
timestamp 1666199351
transform 1 0 45448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_489
timestamp 1666199351
transform 1 0 46092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_496
timestamp 1666199351
transform 1 0 46736 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_503
timestamp 1666199351
transform 1 0 47380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_510
timestamp 1666199351
transform 1 0 48024 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666199351
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666199351
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666199351
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666199351
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1666199351
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666199351
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666199351
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666199351
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666199351
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666199351
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666199351
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666199351
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666199351
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666199351
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666199351
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_152
timestamp 1666199351
transform 1 0 15088 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_160
timestamp 1666199351
transform 1 0 15824 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1666199351
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1666199351
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_176
timestamp 1666199351
transform 1 0 17296 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_180
timestamp 1666199351
transform 1 0 17664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_184
timestamp 1666199351
transform 1 0 18032 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_191
timestamp 1666199351
transform 1 0 18676 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_198
timestamp 1666199351
transform 1 0 19320 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_205
timestamp 1666199351
transform 1 0 19964 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1666199351
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1666199351
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_236
timestamp 1666199351
transform 1 0 22816 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_242
timestamp 1666199351
transform 1 0 23368 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_246
timestamp 1666199351
transform 1 0 23736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_259
timestamp 1666199351
transform 1 0 24932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_272
timestamp 1666199351
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1666199351
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_292
timestamp 1666199351
transform 1 0 27968 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_307
timestamp 1666199351
transform 1 0 29348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_314
timestamp 1666199351
transform 1 0 29992 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_321
timestamp 1666199351
transform 1 0 30636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_333
timestamp 1666199351
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1666199351
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1666199351
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1666199351
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1666199351
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1666199351
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1666199351
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1666199351
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1666199351
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1666199351
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1666199351
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1666199351
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1666199351
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1666199351
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1666199351
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1666199351
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1666199351
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1666199351
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1666199351
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_505
timestamp 1666199351
transform 1 0 47564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_513
timestamp 1666199351
transform 1 0 48300 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666199351
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666199351
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666199351
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666199351
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666199351
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666199351
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666199351
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666199351
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666199351
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666199351
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666199351
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666199351
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666199351
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666199351
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666199351
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666199351
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666199351
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666199351
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_177
timestamp 1666199351
transform 1 0 17388 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_181
timestamp 1666199351
transform 1 0 17756 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_185
timestamp 1666199351
transform 1 0 18124 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1666199351
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1666199351
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_203
timestamp 1666199351
transform 1 0 19780 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1666199351
transform 1 0 20424 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_223
timestamp 1666199351
transform 1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_227
timestamp 1666199351
transform 1 0 21988 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_231
timestamp 1666199351
transform 1 0 22356 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp 1666199351
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_253
timestamp 1666199351
transform 1 0 24380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_259
timestamp 1666199351
transform 1 0 24932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_263
timestamp 1666199351
transform 1 0 25300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_270
timestamp 1666199351
transform 1 0 25944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_278
timestamp 1666199351
transform 1 0 26680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_282
timestamp 1666199351
transform 1 0 27048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_289
timestamp 1666199351
transform 1 0 27692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1666199351
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1666199351
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_314
timestamp 1666199351
transform 1 0 29992 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1666199351
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1666199351
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1666199351
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1666199351
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1666199351
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1666199351
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1666199351
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1666199351
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1666199351
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1666199351
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1666199351
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1666199351
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1666199351
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1666199351
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1666199351
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1666199351
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1666199351
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1666199351
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1666199351
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1666199351
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_513
timestamp 1666199351
transform 1 0 48300 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666199351
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666199351
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666199351
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1666199351
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666199351
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666199351
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666199351
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666199351
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666199351
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666199351
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666199351
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666199351
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666199351
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666199351
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666199351
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666199351
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666199351
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666199351
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666199351
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666199351
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_193
timestamp 1666199351
transform 1 0 18860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_200
timestamp 1666199351
transform 1 0 19504 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_204
timestamp 1666199351
transform 1 0 19872 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_208
timestamp 1666199351
transform 1 0 20240 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1666199351
transform 1 0 20884 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1666199351
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_225
timestamp 1666199351
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_229
timestamp 1666199351
transform 1 0 22172 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_233
timestamp 1666199351
transform 1 0 22540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_246
timestamp 1666199351
transform 1 0 23736 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_252
timestamp 1666199351
transform 1 0 24288 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_256
timestamp 1666199351
transform 1 0 24656 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_263
timestamp 1666199351
transform 1 0 25300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1666199351
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp 1666199351
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_293
timestamp 1666199351
transform 1 0 28060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_300
timestamp 1666199351
transform 1 0 28704 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_307
timestamp 1666199351
transform 1 0 29348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_319
timestamp 1666199351
transform 1 0 30452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 1666199351
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1666199351
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1666199351
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1666199351
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1666199351
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1666199351
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1666199351
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1666199351
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1666199351
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1666199351
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1666199351
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1666199351
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1666199351
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1666199351
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1666199351
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1666199351
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1666199351
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1666199351
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1666199351
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1666199351
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_505
timestamp 1666199351
transform 1 0 47564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_513
timestamp 1666199351
transform 1 0 48300 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666199351
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666199351
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666199351
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666199351
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666199351
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666199351
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666199351
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666199351
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666199351
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666199351
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666199351
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666199351
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666199351
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666199351
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666199351
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666199351
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666199351
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666199351
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666199351
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666199351
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666199351
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1666199351
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_205
timestamp 1666199351
transform 1 0 19964 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_208
timestamp 1666199351
transform 1 0 20240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1666199351
transform 1 0 20884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_228
timestamp 1666199351
transform 1 0 22080 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_232
timestamp 1666199351
transform 1 0 22448 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_236
timestamp 1666199351
transform 1 0 22816 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1666199351
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1666199351
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_264
timestamp 1666199351
transform 1 0 25392 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_273
timestamp 1666199351
transform 1 0 26220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_280
timestamp 1666199351
transform 1 0 26864 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_284
timestamp 1666199351
transform 1 0 27232 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_294
timestamp 1666199351
transform 1 0 28152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1666199351
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1666199351
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1666199351
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1666199351
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1666199351
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1666199351
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1666199351
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1666199351
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1666199351
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1666199351
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1666199351
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1666199351
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1666199351
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1666199351
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1666199351
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1666199351
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1666199351
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1666199351
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1666199351
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1666199351
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1666199351
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1666199351
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_513
timestamp 1666199351
transform 1 0 48300 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666199351
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666199351
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666199351
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666199351
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666199351
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666199351
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666199351
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666199351
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666199351
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666199351
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666199351
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666199351
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666199351
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666199351
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666199351
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666199351
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666199351
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666199351
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666199351
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666199351
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666199351
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_205
timestamp 1666199351
transform 1 0 19964 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_211
timestamp 1666199351
transform 1 0 20516 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1666199351
transform 1 0 20884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1666199351
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1666199351
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_230
timestamp 1666199351
transform 1 0 22264 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_237
timestamp 1666199351
transform 1 0 22908 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1666199351
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_251
timestamp 1666199351
transform 1 0 24196 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_264
timestamp 1666199351
transform 1 0 25392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_268
timestamp 1666199351
transform 1 0 25760 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1666199351
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_281
timestamp 1666199351
transform 1 0 26956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_288
timestamp 1666199351
transform 1 0 27600 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_295
timestamp 1666199351
transform 1 0 28244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_307
timestamp 1666199351
transform 1 0 29348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_319
timestamp 1666199351
transform 1 0 30452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_331
timestamp 1666199351
transform 1 0 31556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1666199351
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1666199351
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1666199351
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1666199351
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1666199351
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1666199351
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1666199351
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1666199351
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1666199351
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1666199351
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1666199351
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1666199351
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1666199351
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1666199351
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1666199351
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1666199351
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1666199351
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1666199351
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1666199351
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1666199351
transform 1 0 47564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_513
timestamp 1666199351
transform 1 0 48300 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666199351
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666199351
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666199351
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666199351
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666199351
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666199351
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666199351
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666199351
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666199351
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666199351
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666199351
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666199351
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666199351
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666199351
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666199351
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666199351
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666199351
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666199351
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666199351
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666199351
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666199351
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666199351
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666199351
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_221
timestamp 1666199351
transform 1 0 21436 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_227
timestamp 1666199351
transform 1 0 21988 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_233
timestamp 1666199351
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_240
timestamp 1666199351
transform 1 0 23184 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1666199351
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_258
timestamp 1666199351
transform 1 0 24840 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_270
timestamp 1666199351
transform 1 0 25944 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_282
timestamp 1666199351
transform 1 0 27048 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_294
timestamp 1666199351
transform 1 0 28152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1666199351
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1666199351
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1666199351
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1666199351
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1666199351
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1666199351
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1666199351
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1666199351
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1666199351
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1666199351
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1666199351
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1666199351
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1666199351
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1666199351
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1666199351
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1666199351
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1666199351
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1666199351
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1666199351
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1666199351
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1666199351
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1666199351
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_513
timestamp 1666199351
transform 1 0 48300 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666199351
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666199351
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666199351
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1666199351
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1666199351
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666199351
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666199351
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666199351
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666199351
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666199351
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666199351
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666199351
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666199351
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666199351
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666199351
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666199351
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666199351
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666199351
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666199351
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666199351
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666199351
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666199351
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666199351
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666199351
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666199351
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1666199351
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1666199351
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1666199351
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1666199351
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1666199351
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666199351
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1666199351
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1666199351
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1666199351
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1666199351
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1666199351
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1666199351
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1666199351
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1666199351
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1666199351
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1666199351
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1666199351
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1666199351
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1666199351
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1666199351
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1666199351
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1666199351
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1666199351
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1666199351
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1666199351
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1666199351
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1666199351
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1666199351
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1666199351
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_505
timestamp 1666199351
transform 1 0 47564 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_513
timestamp 1666199351
transform 1 0 48300 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666199351
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666199351
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666199351
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666199351
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666199351
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666199351
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666199351
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666199351
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666199351
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666199351
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666199351
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666199351
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666199351
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666199351
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666199351
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666199351
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666199351
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666199351
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666199351
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666199351
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666199351
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666199351
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666199351
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666199351
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1666199351
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1666199351
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666199351
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1666199351
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1666199351
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1666199351
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1666199351
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1666199351
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1666199351
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1666199351
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1666199351
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1666199351
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1666199351
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1666199351
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1666199351
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1666199351
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1666199351
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1666199351
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1666199351
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1666199351
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1666199351
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1666199351
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1666199351
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1666199351
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1666199351
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1666199351
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1666199351
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1666199351
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1666199351
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1666199351
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_513
timestamp 1666199351
transform 1 0 48300 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666199351
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666199351
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666199351
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666199351
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666199351
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666199351
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666199351
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666199351
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666199351
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666199351
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666199351
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666199351
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666199351
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666199351
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666199351
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666199351
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666199351
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666199351
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666199351
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666199351
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666199351
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666199351
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666199351
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666199351
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1666199351
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1666199351
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1666199351
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1666199351
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1666199351
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666199351
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666199351
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1666199351
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1666199351
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1666199351
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1666199351
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1666199351
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1666199351
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1666199351
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1666199351
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1666199351
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1666199351
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1666199351
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1666199351
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1666199351
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1666199351
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1666199351
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1666199351
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1666199351
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1666199351
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1666199351
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1666199351
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1666199351
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1666199351
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1666199351
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1666199351
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1666199351
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666199351
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666199351
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666199351
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666199351
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666199351
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666199351
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666199351
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666199351
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666199351
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666199351
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666199351
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666199351
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666199351
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666199351
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666199351
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666199351
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666199351
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666199351
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666199351
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666199351
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666199351
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666199351
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666199351
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1666199351
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1666199351
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1666199351
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1666199351
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1666199351
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1666199351
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1666199351
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1666199351
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1666199351
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1666199351
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1666199351
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1666199351
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1666199351
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1666199351
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1666199351
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1666199351
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1666199351
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1666199351
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1666199351
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1666199351
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1666199351
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1666199351
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1666199351
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1666199351
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1666199351
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1666199351
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1666199351
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1666199351
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1666199351
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1666199351
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1666199351
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_513
timestamp 1666199351
transform 1 0 48300 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666199351
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666199351
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1666199351
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1666199351
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1666199351
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666199351
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666199351
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666199351
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666199351
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666199351
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666199351
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666199351
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666199351
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666199351
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666199351
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666199351
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666199351
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666199351
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666199351
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666199351
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666199351
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666199351
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666199351
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666199351
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666199351
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666199351
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666199351
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666199351
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666199351
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666199351
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1666199351
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1666199351
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1666199351
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1666199351
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1666199351
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1666199351
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1666199351
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1666199351
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1666199351
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1666199351
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1666199351
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1666199351
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1666199351
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1666199351
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1666199351
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1666199351
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1666199351
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1666199351
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1666199351
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1666199351
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1666199351
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1666199351
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1666199351
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1666199351
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1666199351
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1666199351
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666199351
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1666199351
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666199351
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666199351
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666199351
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666199351
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666199351
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666199351
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666199351
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666199351
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666199351
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666199351
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666199351
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666199351
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666199351
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666199351
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666199351
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666199351
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666199351
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666199351
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666199351
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666199351
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666199351
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1666199351
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1666199351
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1666199351
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666199351
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1666199351
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1666199351
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1666199351
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1666199351
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1666199351
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1666199351
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1666199351
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1666199351
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1666199351
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1666199351
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1666199351
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1666199351
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1666199351
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1666199351
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1666199351
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1666199351
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1666199351
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1666199351
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1666199351
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1666199351
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1666199351
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1666199351
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1666199351
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1666199351
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1666199351
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1666199351
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1666199351
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_513
timestamp 1666199351
transform 1 0 48300 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666199351
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666199351
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666199351
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666199351
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1666199351
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666199351
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666199351
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666199351
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666199351
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666199351
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666199351
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666199351
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666199351
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666199351
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666199351
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666199351
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666199351
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666199351
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666199351
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666199351
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666199351
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666199351
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666199351
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666199351
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666199351
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666199351
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1666199351
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666199351
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1666199351
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666199351
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1666199351
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1666199351
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1666199351
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1666199351
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1666199351
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1666199351
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1666199351
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1666199351
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1666199351
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1666199351
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1666199351
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1666199351
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1666199351
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1666199351
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1666199351
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1666199351
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1666199351
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1666199351
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1666199351
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1666199351
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1666199351
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1666199351
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1666199351
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1666199351
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1666199351
transform 1 0 47564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_513
timestamp 1666199351
transform 1 0 48300 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666199351
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666199351
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666199351
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666199351
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666199351
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666199351
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666199351
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666199351
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666199351
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666199351
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666199351
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666199351
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666199351
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666199351
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666199351
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666199351
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666199351
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666199351
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666199351
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666199351
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666199351
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666199351
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666199351
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666199351
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1666199351
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1666199351
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666199351
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666199351
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1666199351
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1666199351
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1666199351
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1666199351
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1666199351
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1666199351
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1666199351
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1666199351
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1666199351
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1666199351
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1666199351
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1666199351
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1666199351
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1666199351
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1666199351
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1666199351
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1666199351
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1666199351
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1666199351
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1666199351
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1666199351
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1666199351
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1666199351
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1666199351
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1666199351
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1666199351
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_513
timestamp 1666199351
transform 1 0 48300 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666199351
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666199351
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1666199351
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1666199351
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1666199351
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666199351
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666199351
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666199351
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666199351
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666199351
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666199351
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666199351
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666199351
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666199351
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666199351
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666199351
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666199351
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666199351
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666199351
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666199351
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666199351
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666199351
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666199351
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666199351
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1666199351
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1666199351
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1666199351
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1666199351
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666199351
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666199351
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1666199351
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1666199351
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1666199351
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1666199351
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1666199351
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1666199351
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1666199351
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1666199351
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1666199351
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1666199351
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1666199351
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1666199351
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1666199351
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1666199351
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1666199351
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1666199351
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1666199351
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1666199351
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1666199351
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1666199351
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1666199351
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1666199351
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1666199351
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1666199351
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1666199351
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_513
timestamp 1666199351
transform 1 0 48300 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666199351
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1666199351
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666199351
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666199351
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666199351
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666199351
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666199351
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666199351
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666199351
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666199351
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666199351
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666199351
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666199351
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666199351
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666199351
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666199351
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666199351
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666199351
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666199351
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666199351
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666199351
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666199351
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666199351
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1666199351
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1666199351
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1666199351
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666199351
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1666199351
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1666199351
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1666199351
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1666199351
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1666199351
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1666199351
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1666199351
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1666199351
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1666199351
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1666199351
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1666199351
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1666199351
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1666199351
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1666199351
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1666199351
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1666199351
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1666199351
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1666199351
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1666199351
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1666199351
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1666199351
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1666199351
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1666199351
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1666199351
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1666199351
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1666199351
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1666199351
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1666199351
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666199351
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666199351
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666199351
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666199351
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666199351
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666199351
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666199351
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666199351
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666199351
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666199351
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666199351
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666199351
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666199351
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666199351
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666199351
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666199351
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666199351
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666199351
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666199351
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666199351
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666199351
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666199351
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666199351
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666199351
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666199351
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1666199351
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1666199351
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1666199351
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1666199351
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666199351
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1666199351
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1666199351
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1666199351
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1666199351
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1666199351
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1666199351
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1666199351
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1666199351
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1666199351
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1666199351
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1666199351
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1666199351
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1666199351
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1666199351
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1666199351
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1666199351
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1666199351
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1666199351
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1666199351
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1666199351
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1666199351
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1666199351
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1666199351
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1666199351
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1666199351
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1666199351
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1666199351
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1666199351
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666199351
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666199351
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666199351
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666199351
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666199351
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666199351
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666199351
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666199351
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666199351
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666199351
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666199351
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666199351
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666199351
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666199351
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666199351
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666199351
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666199351
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666199351
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666199351
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666199351
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666199351
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666199351
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1666199351
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1666199351
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1666199351
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1666199351
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1666199351
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1666199351
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1666199351
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1666199351
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1666199351
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1666199351
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1666199351
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1666199351
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1666199351
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1666199351
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1666199351
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1666199351
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1666199351
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1666199351
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1666199351
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1666199351
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1666199351
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1666199351
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1666199351
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1666199351
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1666199351
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1666199351
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1666199351
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1666199351
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1666199351
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1666199351
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_513
timestamp 1666199351
transform 1 0 48300 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666199351
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666199351
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666199351
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666199351
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666199351
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666199351
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666199351
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666199351
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666199351
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666199351
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666199351
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666199351
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666199351
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666199351
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666199351
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666199351
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666199351
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666199351
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666199351
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666199351
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666199351
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666199351
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666199351
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666199351
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1666199351
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1666199351
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1666199351
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1666199351
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1666199351
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666199351
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1666199351
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1666199351
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1666199351
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1666199351
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1666199351
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1666199351
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1666199351
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1666199351
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1666199351
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1666199351
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1666199351
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1666199351
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1666199351
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1666199351
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1666199351
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1666199351
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1666199351
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1666199351
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1666199351
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1666199351
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1666199351
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1666199351
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1666199351
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1666199351
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1666199351
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_513
timestamp 1666199351
transform 1 0 48300 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666199351
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1666199351
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666199351
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666199351
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666199351
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666199351
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666199351
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666199351
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666199351
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666199351
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666199351
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666199351
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666199351
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666199351
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666199351
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666199351
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666199351
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666199351
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666199351
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666199351
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666199351
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666199351
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666199351
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666199351
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1666199351
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1666199351
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1666199351
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1666199351
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1666199351
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1666199351
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1666199351
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1666199351
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1666199351
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1666199351
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1666199351
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1666199351
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1666199351
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1666199351
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1666199351
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1666199351
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1666199351
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1666199351
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1666199351
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1666199351
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1666199351
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1666199351
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1666199351
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1666199351
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1666199351
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1666199351
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1666199351
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1666199351
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1666199351
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1666199351
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1666199351
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666199351
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666199351
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666199351
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666199351
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666199351
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666199351
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666199351
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666199351
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666199351
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666199351
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666199351
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666199351
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666199351
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666199351
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666199351
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666199351
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666199351
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666199351
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666199351
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666199351
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666199351
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666199351
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666199351
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666199351
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1666199351
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1666199351
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1666199351
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1666199351
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1666199351
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1666199351
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1666199351
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1666199351
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1666199351
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1666199351
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1666199351
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1666199351
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1666199351
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1666199351
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1666199351
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1666199351
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1666199351
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1666199351
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1666199351
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1666199351
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1666199351
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1666199351
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1666199351
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1666199351
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1666199351
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1666199351
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1666199351
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1666199351
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1666199351
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1666199351
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1666199351
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1666199351
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666199351
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1666199351
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666199351
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666199351
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666199351
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666199351
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666199351
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666199351
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666199351
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666199351
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666199351
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666199351
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666199351
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666199351
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666199351
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666199351
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666199351
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666199351
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666199351
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666199351
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666199351
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666199351
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666199351
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1666199351
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1666199351
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1666199351
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1666199351
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1666199351
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1666199351
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1666199351
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1666199351
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1666199351
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1666199351
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1666199351
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1666199351
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1666199351
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1666199351
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1666199351
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1666199351
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1666199351
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1666199351
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1666199351
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1666199351
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1666199351
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1666199351
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1666199351
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1666199351
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1666199351
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1666199351
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1666199351
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1666199351
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1666199351
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1666199351
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1666199351
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_513
timestamp 1666199351
transform 1 0 48300 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666199351
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666199351
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666199351
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1666199351
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1666199351
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666199351
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666199351
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666199351
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666199351
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666199351
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666199351
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666199351
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666199351
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666199351
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666199351
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666199351
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666199351
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666199351
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666199351
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666199351
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666199351
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666199351
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666199351
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666199351
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1666199351
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1666199351
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1666199351
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1666199351
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1666199351
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1666199351
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1666199351
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1666199351
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1666199351
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1666199351
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1666199351
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1666199351
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1666199351
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1666199351
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1666199351
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1666199351
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1666199351
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1666199351
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1666199351
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1666199351
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1666199351
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1666199351
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1666199351
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1666199351
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1666199351
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1666199351
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1666199351
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1666199351
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1666199351
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1666199351
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_505
timestamp 1666199351
transform 1 0 47564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_513
timestamp 1666199351
transform 1 0 48300 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666199351
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666199351
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666199351
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666199351
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666199351
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666199351
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666199351
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666199351
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666199351
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666199351
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666199351
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666199351
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666199351
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666199351
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666199351
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666199351
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666199351
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666199351
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666199351
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666199351
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666199351
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666199351
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666199351
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1666199351
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1666199351
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1666199351
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1666199351
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1666199351
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1666199351
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1666199351
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1666199351
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1666199351
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1666199351
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1666199351
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1666199351
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1666199351
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1666199351
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1666199351
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1666199351
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1666199351
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1666199351
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1666199351
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1666199351
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1666199351
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1666199351
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1666199351
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1666199351
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1666199351
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1666199351
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1666199351
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1666199351
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1666199351
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1666199351
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1666199351
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_513
timestamp 1666199351
transform 1 0 48300 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666199351
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666199351
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666199351
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666199351
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666199351
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666199351
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666199351
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666199351
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666199351
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666199351
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666199351
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666199351
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666199351
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666199351
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666199351
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666199351
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666199351
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666199351
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666199351
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666199351
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666199351
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666199351
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666199351
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666199351
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1666199351
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1666199351
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1666199351
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1666199351
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1666199351
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1666199351
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1666199351
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1666199351
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1666199351
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1666199351
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1666199351
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1666199351
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1666199351
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1666199351
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1666199351
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1666199351
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1666199351
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1666199351
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1666199351
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1666199351
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1666199351
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1666199351
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1666199351
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1666199351
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1666199351
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1666199351
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1666199351
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1666199351
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1666199351
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1666199351
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1666199351
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_513
timestamp 1666199351
transform 1 0 48300 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666199351
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1666199351
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666199351
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666199351
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666199351
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666199351
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666199351
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666199351
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666199351
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666199351
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666199351
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666199351
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666199351
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666199351
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666199351
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666199351
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666199351
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666199351
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666199351
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666199351
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666199351
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666199351
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666199351
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666199351
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1666199351
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1666199351
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1666199351
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1666199351
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1666199351
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1666199351
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1666199351
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1666199351
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1666199351
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1666199351
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1666199351
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1666199351
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1666199351
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1666199351
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1666199351
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1666199351
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1666199351
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1666199351
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1666199351
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1666199351
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1666199351
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1666199351
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1666199351
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1666199351
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1666199351
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1666199351
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1666199351
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1666199351
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1666199351
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1666199351
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_513
timestamp 1666199351
transform 1 0 48300 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666199351
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1666199351
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1666199351
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1666199351
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1666199351
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1666199351
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666199351
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666199351
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666199351
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666199351
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666199351
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666199351
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666199351
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666199351
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666199351
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666199351
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666199351
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666199351
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666199351
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666199351
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666199351
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666199351
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666199351
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666199351
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1666199351
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1666199351
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1666199351
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1666199351
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1666199351
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1666199351
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1666199351
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1666199351
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1666199351
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1666199351
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1666199351
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1666199351
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1666199351
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1666199351
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1666199351
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1666199351
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1666199351
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1666199351
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1666199351
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1666199351
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1666199351
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1666199351
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1666199351
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1666199351
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1666199351
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1666199351
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1666199351
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1666199351
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1666199351
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1666199351
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1666199351
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_513
timestamp 1666199351
transform 1 0 48300 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666199351
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666199351
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666199351
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666199351
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666199351
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666199351
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666199351
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666199351
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666199351
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666199351
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666199351
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666199351
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666199351
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666199351
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666199351
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666199351
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666199351
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666199351
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666199351
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666199351
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666199351
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666199351
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666199351
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1666199351
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1666199351
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1666199351
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1666199351
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1666199351
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1666199351
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1666199351
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1666199351
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1666199351
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1666199351
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1666199351
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1666199351
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1666199351
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1666199351
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1666199351
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1666199351
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1666199351
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1666199351
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1666199351
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1666199351
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1666199351
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1666199351
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1666199351
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1666199351
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1666199351
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1666199351
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1666199351
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1666199351
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1666199351
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1666199351
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1666199351
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_513
timestamp 1666199351
transform 1 0 48300 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666199351
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666199351
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666199351
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666199351
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666199351
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666199351
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666199351
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666199351
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666199351
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666199351
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666199351
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666199351
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666199351
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666199351
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666199351
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666199351
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666199351
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666199351
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666199351
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666199351
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666199351
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666199351
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666199351
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666199351
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1666199351
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1666199351
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1666199351
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1666199351
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1666199351
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1666199351
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1666199351
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1666199351
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1666199351
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1666199351
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1666199351
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1666199351
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1666199351
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1666199351
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1666199351
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1666199351
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1666199351
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1666199351
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1666199351
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1666199351
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1666199351
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1666199351
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1666199351
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1666199351
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1666199351
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1666199351
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1666199351
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1666199351
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1666199351
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1666199351
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_505
timestamp 1666199351
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_513
timestamp 1666199351
transform 1 0 48300 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666199351
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666199351
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666199351
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666199351
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666199351
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666199351
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666199351
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666199351
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666199351
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666199351
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666199351
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666199351
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666199351
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666199351
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666199351
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666199351
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666199351
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666199351
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666199351
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666199351
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666199351
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666199351
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1666199351
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1666199351
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1666199351
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1666199351
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1666199351
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1666199351
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1666199351
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1666199351
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1666199351
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1666199351
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1666199351
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1666199351
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1666199351
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1666199351
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1666199351
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1666199351
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1666199351
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1666199351
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1666199351
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1666199351
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1666199351
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1666199351
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1666199351
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1666199351
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1666199351
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1666199351
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1666199351
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1666199351
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1666199351
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1666199351
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1666199351
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1666199351
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_513
timestamp 1666199351
transform 1 0 48300 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666199351
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666199351
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1666199351
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666199351
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666199351
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666199351
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666199351
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666199351
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666199351
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666199351
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666199351
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666199351
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666199351
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666199351
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666199351
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666199351
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666199351
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666199351
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666199351
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666199351
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666199351
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1666199351
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666199351
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666199351
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1666199351
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1666199351
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1666199351
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1666199351
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1666199351
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1666199351
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1666199351
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1666199351
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1666199351
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1666199351
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1666199351
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1666199351
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1666199351
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1666199351
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1666199351
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1666199351
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1666199351
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1666199351
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1666199351
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1666199351
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1666199351
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1666199351
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1666199351
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1666199351
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1666199351
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1666199351
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1666199351
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1666199351
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1666199351
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1666199351
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1666199351
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_513
timestamp 1666199351
transform 1 0 48300 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666199351
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666199351
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666199351
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666199351
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666199351
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666199351
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666199351
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666199351
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666199351
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666199351
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666199351
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666199351
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666199351
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666199351
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666199351
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666199351
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666199351
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666199351
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666199351
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666199351
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666199351
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666199351
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666199351
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666199351
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1666199351
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1666199351
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1666199351
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1666199351
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1666199351
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1666199351
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1666199351
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1666199351
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1666199351
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1666199351
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1666199351
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1666199351
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1666199351
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1666199351
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1666199351
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1666199351
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1666199351
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1666199351
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1666199351
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1666199351
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1666199351
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1666199351
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1666199351
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1666199351
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1666199351
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1666199351
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1666199351
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1666199351
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1666199351
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1666199351
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_513
timestamp 1666199351
transform 1 0 48300 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666199351
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666199351
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1666199351
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1666199351
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1666199351
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666199351
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666199351
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666199351
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666199351
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666199351
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666199351
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666199351
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666199351
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666199351
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666199351
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666199351
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666199351
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666199351
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666199351
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666199351
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1666199351
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1666199351
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1666199351
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1666199351
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1666199351
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1666199351
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1666199351
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1666199351
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1666199351
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1666199351
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1666199351
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1666199351
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1666199351
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1666199351
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1666199351
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1666199351
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1666199351
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1666199351
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1666199351
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1666199351
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1666199351
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1666199351
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1666199351
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1666199351
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1666199351
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1666199351
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1666199351
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1666199351
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1666199351
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1666199351
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1666199351
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1666199351
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1666199351
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1666199351
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1666199351
transform 1 0 47564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_513
timestamp 1666199351
transform 1 0 48300 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666199351
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666199351
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666199351
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666199351
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666199351
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666199351
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666199351
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666199351
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666199351
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666199351
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666199351
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666199351
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666199351
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666199351
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666199351
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666199351
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666199351
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666199351
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1666199351
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1666199351
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1666199351
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1666199351
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1666199351
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1666199351
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1666199351
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1666199351
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666199351
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1666199351
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1666199351
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1666199351
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1666199351
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1666199351
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1666199351
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1666199351
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1666199351
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1666199351
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1666199351
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1666199351
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1666199351
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1666199351
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1666199351
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1666199351
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1666199351
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1666199351
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1666199351
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1666199351
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1666199351
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1666199351
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1666199351
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1666199351
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1666199351
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1666199351
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1666199351
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1666199351
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_513
timestamp 1666199351
transform 1 0 48300 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666199351
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666199351
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1666199351
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1666199351
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1666199351
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1666199351
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666199351
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666199351
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666199351
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666199351
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666199351
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666199351
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666199351
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666199351
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666199351
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666199351
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666199351
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666199351
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1666199351
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1666199351
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1666199351
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1666199351
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1666199351
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666199351
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1666199351
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1666199351
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1666199351
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1666199351
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1666199351
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666199351
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1666199351
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1666199351
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1666199351
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1666199351
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1666199351
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1666199351
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1666199351
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1666199351
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1666199351
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1666199351
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1666199351
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1666199351
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1666199351
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1666199351
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1666199351
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1666199351
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1666199351
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1666199351
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1666199351
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1666199351
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1666199351
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1666199351
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1666199351
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1666199351
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1666199351
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_513
timestamp 1666199351
transform 1 0 48300 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666199351
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666199351
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666199351
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666199351
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666199351
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666199351
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666199351
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666199351
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666199351
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666199351
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666199351
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666199351
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666199351
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666199351
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666199351
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666199351
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1666199351
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1666199351
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1666199351
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1666199351
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666199351
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1666199351
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1666199351
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1666199351
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1666199351
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1666199351
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1666199351
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1666199351
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1666199351
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1666199351
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1666199351
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1666199351
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1666199351
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1666199351
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1666199351
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1666199351
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1666199351
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1666199351
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1666199351
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1666199351
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1666199351
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1666199351
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1666199351
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1666199351
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1666199351
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1666199351
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1666199351
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1666199351
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1666199351
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1666199351
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1666199351
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1666199351
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1666199351
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1666199351
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_513
timestamp 1666199351
transform 1 0 48300 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1666199351
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666199351
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1666199351
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1666199351
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1666199351
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1666199351
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666199351
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666199351
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666199351
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666199351
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666199351
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666199351
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666199351
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666199351
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666199351
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1666199351
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666199351
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666199351
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666199351
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1666199351
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1666199351
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1666199351
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1666199351
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666199351
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1666199351
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1666199351
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1666199351
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1666199351
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1666199351
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1666199351
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1666199351
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1666199351
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1666199351
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1666199351
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1666199351
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1666199351
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1666199351
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1666199351
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1666199351
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1666199351
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1666199351
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1666199351
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1666199351
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1666199351
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1666199351
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1666199351
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1666199351
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1666199351
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1666199351
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1666199351
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1666199351
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1666199351
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1666199351
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1666199351
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1666199351
transform 1 0 47564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_513
timestamp 1666199351
transform 1 0 48300 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666199351
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1666199351
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666199351
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666199351
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666199351
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666199351
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666199351
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666199351
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666199351
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666199351
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666199351
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666199351
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666199351
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666199351
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666199351
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666199351
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1666199351
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1666199351
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1666199351
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1666199351
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1666199351
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666199351
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1666199351
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1666199351
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1666199351
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1666199351
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1666199351
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1666199351
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1666199351
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1666199351
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1666199351
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1666199351
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1666199351
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1666199351
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1666199351
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1666199351
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1666199351
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1666199351
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1666199351
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1666199351
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1666199351
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1666199351
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1666199351
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1666199351
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1666199351
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1666199351
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1666199351
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1666199351
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1666199351
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1666199351
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1666199351
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1666199351
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1666199351
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1666199351
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_513
timestamp 1666199351
transform 1 0 48300 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666199351
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666199351
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666199351
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666199351
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666199351
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666199351
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666199351
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666199351
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666199351
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666199351
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666199351
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666199351
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666199351
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666199351
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666199351
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1666199351
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1666199351
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1666199351
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666199351
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1666199351
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1666199351
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1666199351
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1666199351
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1666199351
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1666199351
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1666199351
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1666199351
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1666199351
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1666199351
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1666199351
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666199351
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1666199351
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1666199351
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1666199351
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1666199351
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1666199351
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1666199351
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1666199351
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1666199351
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1666199351
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1666199351
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1666199351
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1666199351
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1666199351
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1666199351
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1666199351
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1666199351
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1666199351
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1666199351
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1666199351
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1666199351
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1666199351
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1666199351
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1666199351
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_505
timestamp 1666199351
transform 1 0 47564 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_513
timestamp 1666199351
transform 1 0 48300 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666199351
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1666199351
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666199351
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666199351
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666199351
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666199351
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666199351
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666199351
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666199351
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666199351
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666199351
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1666199351
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1666199351
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1666199351
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666199351
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666199351
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1666199351
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1666199351
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1666199351
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1666199351
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1666199351
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1666199351
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1666199351
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1666199351
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1666199351
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1666199351
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666199351
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1666199351
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1666199351
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1666199351
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1666199351
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1666199351
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1666199351
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1666199351
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1666199351
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1666199351
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1666199351
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1666199351
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1666199351
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1666199351
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1666199351
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1666199351
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1666199351
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1666199351
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1666199351
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1666199351
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1666199351
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1666199351
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1666199351
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1666199351
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1666199351
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1666199351
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1666199351
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1666199351
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_513
timestamp 1666199351
transform 1 0 48300 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666199351
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666199351
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1666199351
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1666199351
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1666199351
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666199351
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666199351
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666199351
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666199351
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1666199351
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666199351
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666199351
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666199351
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1666199351
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1666199351
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1666199351
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1666199351
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1666199351
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1666199351
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1666199351
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1666199351
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1666199351
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1666199351
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1666199351
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666199351
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666199351
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1666199351
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1666199351
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1666199351
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1666199351
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1666199351
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1666199351
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1666199351
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1666199351
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1666199351
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1666199351
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1666199351
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1666199351
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1666199351
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1666199351
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1666199351
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1666199351
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1666199351
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1666199351
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1666199351
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1666199351
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1666199351
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1666199351
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1666199351
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1666199351
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1666199351
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1666199351
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1666199351
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1666199351
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_505
timestamp 1666199351
transform 1 0 47564 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_513
timestamp 1666199351
transform 1 0 48300 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666199351
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1666199351
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666199351
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666199351
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666199351
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666199351
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666199351
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666199351
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666199351
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1666199351
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1666199351
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1666199351
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1666199351
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1666199351
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666199351
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666199351
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666199351
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1666199351
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1666199351
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1666199351
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1666199351
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1666199351
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1666199351
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1666199351
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1666199351
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1666199351
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666199351
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1666199351
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1666199351
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1666199351
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1666199351
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1666199351
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1666199351
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1666199351
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1666199351
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1666199351
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1666199351
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1666199351
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1666199351
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1666199351
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1666199351
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1666199351
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1666199351
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1666199351
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1666199351
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1666199351
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1666199351
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1666199351
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1666199351
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1666199351
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1666199351
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1666199351
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1666199351
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1666199351
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_513
timestamp 1666199351
transform 1 0 48300 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666199351
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666199351
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666199351
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666199351
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666199351
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666199351
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666199351
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666199351
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1666199351
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1666199351
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1666199351
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666199351
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1666199351
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1666199351
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1666199351
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1666199351
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666199351
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666199351
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666199351
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1666199351
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1666199351
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1666199351
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1666199351
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666199351
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1666199351
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1666199351
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1666199351
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1666199351
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1666199351
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1666199351
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1666199351
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1666199351
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1666199351
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1666199351
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1666199351
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1666199351
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1666199351
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1666199351
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1666199351
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1666199351
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1666199351
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1666199351
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1666199351
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1666199351
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1666199351
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1666199351
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1666199351
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1666199351
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1666199351
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1666199351
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1666199351
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1666199351
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1666199351
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1666199351
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1666199351
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1666199351
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666199351
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666199351
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666199351
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666199351
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666199351
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666199351
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666199351
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1666199351
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666199351
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1666199351
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1666199351
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1666199351
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1666199351
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1666199351
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666199351
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1666199351
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1666199351
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1666199351
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1666199351
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1666199351
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666199351
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666199351
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1666199351
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1666199351
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1666199351
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1666199351
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1666199351
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1666199351
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1666199351
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1666199351
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1666199351
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1666199351
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1666199351
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1666199351
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1666199351
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1666199351
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1666199351
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1666199351
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1666199351
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1666199351
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1666199351
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1666199351
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1666199351
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1666199351
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1666199351
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1666199351
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1666199351
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1666199351
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1666199351
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1666199351
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1666199351
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1666199351
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1666199351
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1666199351
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_513
timestamp 1666199351
transform 1 0 48300 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666199351
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666199351
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666199351
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1666199351
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1666199351
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666199351
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666199351
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1666199351
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1666199351
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1666199351
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1666199351
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666199351
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1666199351
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1666199351
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666199351
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1666199351
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1666199351
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1666199351
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1666199351
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1666199351
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1666199351
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1666199351
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1666199351
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1666199351
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1666199351
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1666199351
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1666199351
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1666199351
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1666199351
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1666199351
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1666199351
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1666199351
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1666199351
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1666199351
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1666199351
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1666199351
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1666199351
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1666199351
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1666199351
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1666199351
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1666199351
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1666199351
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1666199351
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1666199351
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1666199351
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1666199351
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1666199351
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1666199351
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1666199351
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1666199351
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1666199351
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1666199351
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1666199351
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1666199351
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_505
timestamp 1666199351
transform 1 0 47564 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_513
timestamp 1666199351
transform 1 0 48300 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666199351
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1666199351
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666199351
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666199351
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666199351
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666199351
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666199351
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666199351
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666199351
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1666199351
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1666199351
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1666199351
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1666199351
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1666199351
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666199351
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1666199351
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1666199351
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1666199351
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1666199351
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1666199351
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1666199351
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1666199351
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1666199351
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1666199351
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1666199351
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1666199351
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1666199351
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1666199351
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1666199351
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1666199351
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1666199351
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1666199351
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1666199351
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1666199351
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1666199351
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1666199351
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1666199351
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1666199351
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1666199351
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1666199351
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1666199351
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1666199351
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1666199351
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1666199351
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1666199351
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1666199351
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1666199351
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1666199351
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1666199351
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1666199351
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1666199351
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1666199351
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1666199351
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1666199351
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_513
timestamp 1666199351
transform 1 0 48300 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666199351
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666199351
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666199351
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666199351
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666199351
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666199351
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666199351
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1666199351
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1666199351
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1666199351
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1666199351
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1666199351
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1666199351
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1666199351
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1666199351
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1666199351
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1666199351
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666199351
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1666199351
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1666199351
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1666199351
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1666199351
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1666199351
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1666199351
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1666199351
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1666199351
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1666199351
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1666199351
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1666199351
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1666199351
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1666199351
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1666199351
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1666199351
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1666199351
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1666199351
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1666199351
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1666199351
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1666199351
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1666199351
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1666199351
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1666199351
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1666199351
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1666199351
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1666199351
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1666199351
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1666199351
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1666199351
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1666199351
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1666199351
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1666199351
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1666199351
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1666199351
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1666199351
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1666199351
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1666199351
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1666199351
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666199351
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666199351
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666199351
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666199351
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666199351
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666199351
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666199351
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666199351
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666199351
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1666199351
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1666199351
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1666199351
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1666199351
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1666199351
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1666199351
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1666199351
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1666199351
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1666199351
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1666199351
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1666199351
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666199351
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1666199351
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1666199351
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1666199351
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1666199351
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1666199351
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1666199351
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1666199351
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1666199351
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1666199351
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1666199351
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1666199351
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666199351
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1666199351
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1666199351
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1666199351
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1666199351
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1666199351
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1666199351
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1666199351
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1666199351
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1666199351
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1666199351
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1666199351
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1666199351
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1666199351
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1666199351
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1666199351
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1666199351
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1666199351
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1666199351
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1666199351
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1666199351
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1666199351
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_513
timestamp 1666199351
transform 1 0 48300 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666199351
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666199351
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666199351
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666199351
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666199351
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666199351
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666199351
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666199351
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666199351
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666199351
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666199351
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666199351
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666199351
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1666199351
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1666199351
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1666199351
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1666199351
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666199351
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1666199351
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1666199351
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1666199351
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1666199351
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1666199351
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666199351
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1666199351
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1666199351
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1666199351
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1666199351
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1666199351
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666199351
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1666199351
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1666199351
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1666199351
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1666199351
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1666199351
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1666199351
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1666199351
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1666199351
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1666199351
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1666199351
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1666199351
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1666199351
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1666199351
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1666199351
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1666199351
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1666199351
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1666199351
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1666199351
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1666199351
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1666199351
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1666199351
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1666199351
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1666199351
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1666199351
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1666199351
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1666199351
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666199351
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666199351
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666199351
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666199351
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666199351
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666199351
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666199351
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666199351
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666199351
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1666199351
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1666199351
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1666199351
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1666199351
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1666199351
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666199351
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1666199351
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1666199351
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1666199351
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1666199351
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1666199351
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1666199351
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1666199351
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1666199351
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1666199351
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1666199351
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1666199351
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1666199351
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1666199351
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1666199351
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1666199351
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1666199351
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1666199351
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666199351
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1666199351
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1666199351
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1666199351
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1666199351
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1666199351
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1666199351
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1666199351
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1666199351
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1666199351
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1666199351
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1666199351
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1666199351
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1666199351
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1666199351
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1666199351
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1666199351
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1666199351
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1666199351
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1666199351
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1666199351
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1666199351
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1666199351
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666199351
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666199351
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666199351
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1666199351
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1666199351
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1666199351
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666199351
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666199351
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666199351
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1666199351
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1666199351
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666199351
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666199351
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1666199351
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1666199351
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1666199351
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1666199351
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666199351
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1666199351
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1666199351
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1666199351
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1666199351
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1666199351
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1666199351
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1666199351
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1666199351
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1666199351
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1666199351
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1666199351
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1666199351
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1666199351
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1666199351
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1666199351
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1666199351
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1666199351
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1666199351
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1666199351
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1666199351
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1666199351
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1666199351
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1666199351
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1666199351
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1666199351
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1666199351
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1666199351
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1666199351
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1666199351
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1666199351
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1666199351
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1666199351
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1666199351
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1666199351
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1666199351
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1666199351
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1666199351
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1666199351
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666199351
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1666199351
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666199351
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666199351
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666199351
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666199351
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666199351
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666199351
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666199351
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666199351
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666199351
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1666199351
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1666199351
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1666199351
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666199351
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1666199351
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1666199351
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1666199351
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1666199351
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1666199351
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1666199351
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1666199351
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1666199351
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1666199351
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1666199351
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1666199351
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1666199351
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1666199351
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1666199351
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1666199351
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1666199351
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1666199351
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1666199351
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1666199351
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1666199351
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1666199351
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1666199351
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1666199351
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1666199351
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1666199351
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1666199351
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1666199351
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1666199351
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1666199351
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1666199351
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1666199351
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1666199351
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1666199351
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1666199351
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1666199351
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1666199351
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1666199351
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1666199351
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1666199351
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_513
timestamp 1666199351
transform 1 0 48300 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666199351
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666199351
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666199351
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666199351
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666199351
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666199351
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666199351
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666199351
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1666199351
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666199351
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666199351
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666199351
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1666199351
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1666199351
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666199351
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666199351
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666199351
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666199351
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1666199351
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1666199351
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1666199351
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1666199351
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1666199351
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1666199351
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1666199351
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1666199351
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1666199351
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1666199351
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1666199351
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1666199351
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1666199351
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1666199351
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1666199351
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1666199351
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1666199351
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1666199351
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1666199351
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1666199351
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1666199351
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1666199351
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1666199351
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1666199351
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1666199351
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1666199351
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1666199351
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1666199351
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1666199351
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1666199351
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1666199351
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1666199351
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1666199351
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1666199351
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1666199351
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1666199351
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1666199351
transform 1 0 47564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_513
timestamp 1666199351
transform 1 0 48300 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666199351
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666199351
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666199351
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666199351
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666199351
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666199351
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666199351
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666199351
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666199351
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666199351
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1666199351
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1666199351
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1666199351
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1666199351
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666199351
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666199351
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1666199351
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1666199351
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1666199351
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1666199351
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1666199351
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1666199351
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1666199351
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1666199351
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1666199351
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1666199351
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666199351
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1666199351
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1666199351
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1666199351
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1666199351
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1666199351
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1666199351
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1666199351
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1666199351
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1666199351
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1666199351
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1666199351
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1666199351
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1666199351
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1666199351
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1666199351
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1666199351
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1666199351
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1666199351
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1666199351
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1666199351
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1666199351
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1666199351
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1666199351
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1666199351
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1666199351
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1666199351
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1666199351
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_513
timestamp 1666199351
transform 1 0 48300 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666199351
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666199351
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1666199351
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1666199351
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1666199351
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1666199351
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666199351
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1666199351
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1666199351
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1666199351
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1666199351
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666199351
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666199351
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666199351
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1666199351
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1666199351
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1666199351
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666199351
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1666199351
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1666199351
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1666199351
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1666199351
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1666199351
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1666199351
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1666199351
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1666199351
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1666199351
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1666199351
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1666199351
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1666199351
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1666199351
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1666199351
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1666199351
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1666199351
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1666199351
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1666199351
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1666199351
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1666199351
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1666199351
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1666199351
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1666199351
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1666199351
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1666199351
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1666199351
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1666199351
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1666199351
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1666199351
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1666199351
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1666199351
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1666199351
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1666199351
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1666199351
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1666199351
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1666199351
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_505
timestamp 1666199351
transform 1 0 47564 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_513
timestamp 1666199351
transform 1 0 48300 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1666199351
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1666199351
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666199351
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1666199351
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1666199351
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1666199351
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666199351
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1666199351
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666199351
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1666199351
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1666199351
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1666199351
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1666199351
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1666199351
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666199351
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1666199351
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1666199351
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1666199351
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1666199351
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1666199351
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1666199351
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1666199351
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1666199351
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1666199351
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1666199351
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1666199351
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1666199351
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1666199351
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1666199351
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1666199351
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1666199351
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1666199351
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1666199351
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1666199351
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1666199351
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1666199351
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1666199351
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1666199351
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1666199351
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1666199351
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1666199351
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1666199351
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1666199351
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1666199351
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1666199351
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1666199351
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1666199351
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1666199351
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1666199351
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1666199351
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1666199351
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1666199351
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1666199351
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1666199351
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_513
timestamp 1666199351
transform 1 0 48300 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1666199351
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666199351
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1666199351
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1666199351
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1666199351
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1666199351
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1666199351
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1666199351
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1666199351
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1666199351
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1666199351
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666199351
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1666199351
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1666199351
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1666199351
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1666199351
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1666199351
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1666199351
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1666199351
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1666199351
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1666199351
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1666199351
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1666199351
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1666199351
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1666199351
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1666199351
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1666199351
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1666199351
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1666199351
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1666199351
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1666199351
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1666199351
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1666199351
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1666199351
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1666199351
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1666199351
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1666199351
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1666199351
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1666199351
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1666199351
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1666199351
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1666199351
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1666199351
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1666199351
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1666199351
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1666199351
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1666199351
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1666199351
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1666199351
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1666199351
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1666199351
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1666199351
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1666199351
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1666199351
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1666199351
transform 1 0 47564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_513
timestamp 1666199351
transform 1 0 48300 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1666199351
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1666199351
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1666199351
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1666199351
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1666199351
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1666199351
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1666199351
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1666199351
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666199351
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1666199351
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1666199351
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1666199351
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1666199351
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1666199351
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666199351
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1666199351
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1666199351
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1666199351
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1666199351
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1666199351
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1666199351
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1666199351
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1666199351
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1666199351
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1666199351
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1666199351
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1666199351
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1666199351
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1666199351
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1666199351
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1666199351
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1666199351
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1666199351
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1666199351
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1666199351
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1666199351
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1666199351
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1666199351
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1666199351
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1666199351
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1666199351
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1666199351
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1666199351
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1666199351
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1666199351
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1666199351
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1666199351
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1666199351
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1666199351
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1666199351
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1666199351
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1666199351
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1666199351
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1666199351
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_513
timestamp 1666199351
transform 1 0 48300 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1666199351
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1666199351
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1666199351
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1666199351
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1666199351
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1666199351
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1666199351
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1666199351
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1666199351
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1666199351
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1666199351
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666199351
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1666199351
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1666199351
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1666199351
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1666199351
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1666199351
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666199351
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1666199351
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1666199351
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1666199351
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1666199351
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1666199351
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1666199351
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1666199351
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1666199351
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1666199351
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1666199351
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1666199351
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1666199351
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1666199351
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1666199351
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1666199351
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1666199351
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1666199351
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1666199351
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1666199351
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1666199351
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1666199351
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1666199351
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1666199351
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1666199351
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1666199351
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1666199351
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1666199351
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1666199351
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1666199351
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1666199351
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1666199351
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1666199351
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1666199351
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1666199351
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1666199351
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1666199351
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1666199351
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1666199351
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1666199351
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1666199351
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1666199351
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1666199351
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1666199351
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1666199351
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1666199351
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1666199351
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1666199351
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1666199351
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1666199351
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1666199351
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1666199351
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1666199351
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1666199351
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1666199351
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1666199351
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1666199351
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1666199351
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1666199351
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1666199351
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1666199351
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1666199351
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1666199351
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1666199351
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1666199351
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1666199351
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1666199351
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1666199351
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1666199351
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1666199351
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1666199351
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1666199351
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1666199351
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1666199351
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1666199351
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1666199351
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1666199351
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1666199351
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1666199351
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1666199351
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1666199351
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1666199351
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1666199351
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1666199351
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1666199351
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1666199351
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1666199351
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1666199351
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1666199351
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1666199351
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1666199351
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1666199351
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1666199351
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1666199351
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1666199351
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1666199351
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1666199351
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1666199351
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1666199351
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1666199351
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1666199351
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1666199351
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1666199351
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1666199351
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1666199351
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666199351
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1666199351
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1666199351
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1666199351
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1666199351
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1666199351
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1666199351
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1666199351
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1666199351
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1666199351
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1666199351
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1666199351
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1666199351
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1666199351
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1666199351
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1666199351
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1666199351
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1666199351
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1666199351
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1666199351
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1666199351
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1666199351
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1666199351
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1666199351
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1666199351
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1666199351
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1666199351
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1666199351
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1666199351
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1666199351
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1666199351
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1666199351
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1666199351
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1666199351
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1666199351
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1666199351
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1666199351
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1666199351
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1666199351
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1666199351
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1666199351
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1666199351
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1666199351
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1666199351
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1666199351
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1666199351
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1666199351
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1666199351
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1666199351
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1666199351
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1666199351
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1666199351
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1666199351
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1666199351
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1666199351
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1666199351
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1666199351
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1666199351
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1666199351
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1666199351
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1666199351
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1666199351
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1666199351
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1666199351
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1666199351
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1666199351
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1666199351
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1666199351
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1666199351
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1666199351
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1666199351
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1666199351
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1666199351
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1666199351
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1666199351
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1666199351
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1666199351
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1666199351
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1666199351
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1666199351
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1666199351
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1666199351
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1666199351
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1666199351
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1666199351
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1666199351
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1666199351
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1666199351
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1666199351
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1666199351
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1666199351
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1666199351
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1666199351
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1666199351
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1666199351
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1666199351
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1666199351
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1666199351
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1666199351
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_513
timestamp 1666199351
transform 1 0 48300 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1666199351
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1666199351
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1666199351
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1666199351
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1666199351
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1666199351
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1666199351
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1666199351
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1666199351
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1666199351
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1666199351
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1666199351
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1666199351
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1666199351
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1666199351
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1666199351
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1666199351
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1666199351
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1666199351
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1666199351
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1666199351
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1666199351
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1666199351
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1666199351
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1666199351
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1666199351
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1666199351
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1666199351
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1666199351
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1666199351
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1666199351
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1666199351
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1666199351
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1666199351
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1666199351
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1666199351
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1666199351
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1666199351
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1666199351
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1666199351
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1666199351
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1666199351
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1666199351
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1666199351
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1666199351
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1666199351
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1666199351
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1666199351
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1666199351
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1666199351
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1666199351
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1666199351
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1666199351
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1666199351
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_505
timestamp 1666199351
transform 1 0 47564 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_513
timestamp 1666199351
transform 1 0 48300 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1666199351
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1666199351
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1666199351
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1666199351
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1666199351
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1666199351
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1666199351
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1666199351
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1666199351
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1666199351
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1666199351
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1666199351
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1666199351
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1666199351
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1666199351
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1666199351
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1666199351
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1666199351
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1666199351
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1666199351
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1666199351
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1666199351
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1666199351
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1666199351
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1666199351
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1666199351
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1666199351
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1666199351
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1666199351
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1666199351
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1666199351
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1666199351
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1666199351
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1666199351
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1666199351
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1666199351
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1666199351
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1666199351
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1666199351
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1666199351
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1666199351
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1666199351
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1666199351
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1666199351
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1666199351
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1666199351
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1666199351
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1666199351
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1666199351
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1666199351
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1666199351
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1666199351
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1666199351
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1666199351
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_513
timestamp 1666199351
transform 1 0 48300 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1666199351
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1666199351
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1666199351
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1666199351
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1666199351
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1666199351
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1666199351
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1666199351
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1666199351
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1666199351
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1666199351
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1666199351
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1666199351
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1666199351
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1666199351
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1666199351
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1666199351
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1666199351
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1666199351
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1666199351
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1666199351
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1666199351
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1666199351
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1666199351
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1666199351
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1666199351
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1666199351
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1666199351
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1666199351
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1666199351
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1666199351
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1666199351
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1666199351
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1666199351
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1666199351
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1666199351
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1666199351
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1666199351
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1666199351
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1666199351
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1666199351
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1666199351
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1666199351
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1666199351
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1666199351
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1666199351
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1666199351
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1666199351
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1666199351
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1666199351
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1666199351
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1666199351
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1666199351
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1666199351
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_505
timestamp 1666199351
transform 1 0 47564 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_513
timestamp 1666199351
transform 1 0 48300 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1666199351
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1666199351
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1666199351
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1666199351
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1666199351
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1666199351
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1666199351
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1666199351
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1666199351
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1666199351
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1666199351
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1666199351
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1666199351
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1666199351
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1666199351
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1666199351
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1666199351
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1666199351
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1666199351
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1666199351
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1666199351
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1666199351
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1666199351
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1666199351
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1666199351
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1666199351
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1666199351
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1666199351
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1666199351
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1666199351
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1666199351
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1666199351
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1666199351
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1666199351
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1666199351
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1666199351
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1666199351
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1666199351
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1666199351
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1666199351
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1666199351
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1666199351
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1666199351
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1666199351
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1666199351
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1666199351
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1666199351
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1666199351
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1666199351
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1666199351
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1666199351
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1666199351
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1666199351
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1666199351
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_513
timestamp 1666199351
transform 1 0 48300 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1666199351
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1666199351
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1666199351
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1666199351
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1666199351
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1666199351
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1666199351
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1666199351
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1666199351
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1666199351
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1666199351
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1666199351
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1666199351
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1666199351
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1666199351
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1666199351
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1666199351
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1666199351
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1666199351
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1666199351
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1666199351
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1666199351
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1666199351
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1666199351
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1666199351
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1666199351
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1666199351
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1666199351
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1666199351
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1666199351
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1666199351
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1666199351
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1666199351
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1666199351
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1666199351
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1666199351
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1666199351
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1666199351
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1666199351
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1666199351
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1666199351
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1666199351
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1666199351
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1666199351
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1666199351
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1666199351
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1666199351
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1666199351
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1666199351
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1666199351
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1666199351
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1666199351
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1666199351
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1666199351
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_505
timestamp 1666199351
transform 1 0 47564 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_513
timestamp 1666199351
transform 1 0 48300 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1666199351
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1666199351
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1666199351
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1666199351
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1666199351
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1666199351
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1666199351
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1666199351
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1666199351
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1666199351
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1666199351
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1666199351
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1666199351
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1666199351
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1666199351
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1666199351
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1666199351
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1666199351
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1666199351
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1666199351
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1666199351
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1666199351
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1666199351
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1666199351
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1666199351
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1666199351
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1666199351
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1666199351
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1666199351
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1666199351
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1666199351
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1666199351
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1666199351
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1666199351
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1666199351
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1666199351
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1666199351
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1666199351
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1666199351
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1666199351
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1666199351
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1666199351
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1666199351
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1666199351
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1666199351
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1666199351
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1666199351
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1666199351
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1666199351
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1666199351
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1666199351
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1666199351
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1666199351
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1666199351
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_513
timestamp 1666199351
transform 1 0 48300 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1666199351
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1666199351
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1666199351
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1666199351
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1666199351
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1666199351
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1666199351
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1666199351
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1666199351
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1666199351
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1666199351
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1666199351
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1666199351
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1666199351
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1666199351
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1666199351
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1666199351
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1666199351
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1666199351
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1666199351
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1666199351
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1666199351
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1666199351
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1666199351
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1666199351
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1666199351
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1666199351
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1666199351
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1666199351
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1666199351
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1666199351
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1666199351
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1666199351
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1666199351
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1666199351
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1666199351
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1666199351
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1666199351
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1666199351
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1666199351
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1666199351
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1666199351
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1666199351
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1666199351
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1666199351
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1666199351
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1666199351
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1666199351
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1666199351
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1666199351
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1666199351
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1666199351
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1666199351
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1666199351
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_505
timestamp 1666199351
transform 1 0 47564 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_513
timestamp 1666199351
transform 1 0 48300 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1666199351
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1666199351
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1666199351
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1666199351
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1666199351
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1666199351
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1666199351
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1666199351
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1666199351
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1666199351
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1666199351
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1666199351
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1666199351
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1666199351
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1666199351
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1666199351
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1666199351
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1666199351
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1666199351
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1666199351
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1666199351
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1666199351
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1666199351
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1666199351
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1666199351
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1666199351
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1666199351
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_253
timestamp 1666199351
transform 1 0 24380 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_261
timestamp 1666199351
transform 1 0 25116 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_264
timestamp 1666199351
transform 1 0 25392 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_276
timestamp 1666199351
transform 1 0 26496 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_288
timestamp 1666199351
transform 1 0 27600 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_300
timestamp 1666199351
transform 1 0 28704 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_309
timestamp 1666199351
transform 1 0 29532 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_313
timestamp 1666199351
transform 1 0 29900 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_325
timestamp 1666199351
transform 1 0 31004 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_337
timestamp 1666199351
transform 1 0 32108 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_349
timestamp 1666199351
transform 1 0 33212 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_361
timestamp 1666199351
transform 1 0 34316 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1666199351
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1666199351
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1666199351
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1666199351
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1666199351
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1666199351
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1666199351
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1666199351
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1666199351
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1666199351
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1666199351
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1666199351
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1666199351
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1666199351
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1666199351
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_513
timestamp 1666199351
transform 1 0 48300 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1666199351
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1666199351
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1666199351
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1666199351
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1666199351
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1666199351
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1666199351
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1666199351
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1666199351
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1666199351
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1666199351
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1666199351
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1666199351
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1666199351
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1666199351
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1666199351
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1666199351
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1666199351
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1666199351
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1666199351
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1666199351
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1666199351
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1666199351
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1666199351
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1666199351
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1666199351
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1666199351
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_263
timestamp 1666199351
transform 1 0 25300 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_269
timestamp 1666199351
transform 1 0 25852 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_275
timestamp 1666199351
transform 1 0 26404 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1666199351
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_281
timestamp 1666199351
transform 1 0 26956 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_285
timestamp 1666199351
transform 1 0 27324 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_291
timestamp 1666199351
transform 1 0 27876 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_297
timestamp 1666199351
transform 1 0 28428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_305
timestamp 1666199351
transform 1 0 29164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_308
timestamp 1666199351
transform 1 0 29440 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_314
timestamp 1666199351
transform 1 0 29992 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_324
timestamp 1666199351
transform 1 0 30912 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_337
timestamp 1666199351
transform 1 0 32108 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_341
timestamp 1666199351
transform 1 0 32476 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_353
timestamp 1666199351
transform 1 0 33580 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1666199351
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_375
timestamp 1666199351
transform 1 0 35604 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_381
timestamp 1666199351
transform 1 0 36156 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_389
timestamp 1666199351
transform 1 0 36892 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1666199351
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1666199351
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1666199351
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1666199351
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1666199351
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1666199351
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1666199351
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1666199351
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1666199351
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1666199351
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1666199351
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1666199351
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1666199351
transform 1 0 47564 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_513
timestamp 1666199351
transform 1 0 48300 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1666199351
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1666199351
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1666199351
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1666199351
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1666199351
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1666199351
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1666199351
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1666199351
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1666199351
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1666199351
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1666199351
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1666199351
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1666199351
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1666199351
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1666199351
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1666199351
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1666199351
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1666199351
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1666199351
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1666199351
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1666199351
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1666199351
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1666199351
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1666199351
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_233
timestamp 1666199351
transform 1 0 22540 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_239
timestamp 1666199351
transform 1 0 23092 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_247
timestamp 1666199351
transform 1 0 23828 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1666199351
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_253
timestamp 1666199351
transform 1 0 24380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_257
timestamp 1666199351
transform 1 0 24748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_263
timestamp 1666199351
transform 1 0 25300 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_269
timestamp 1666199351
transform 1 0 25852 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_275
timestamp 1666199351
transform 1 0 26404 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_285
timestamp 1666199351
transform 1 0 27324 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_291
timestamp 1666199351
transform 1 0 27876 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_299
timestamp 1666199351
transform 1 0 28612 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_74_305
timestamp 1666199351
transform 1 0 29164 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_309
timestamp 1666199351
transform 1 0 29532 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_313
timestamp 1666199351
transform 1 0 29900 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_319
timestamp 1666199351
transform 1 0 30452 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_325
timestamp 1666199351
transform 1 0 31004 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_331
timestamp 1666199351
transform 1 0 31556 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_337
timestamp 1666199351
transform 1 0 32108 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_343
timestamp 1666199351
transform 1 0 32660 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_346
timestamp 1666199351
transform 1 0 32936 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_352
timestamp 1666199351
transform 1 0 33488 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_358
timestamp 1666199351
transform 1 0 34040 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_365
timestamp 1666199351
transform 1 0 34684 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_369
timestamp 1666199351
transform 1 0 35052 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_375
timestamp 1666199351
transform 1 0 35604 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_381
timestamp 1666199351
transform 1 0 36156 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_387
timestamp 1666199351
transform 1 0 36708 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_399
timestamp 1666199351
transform 1 0 37812 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_411
timestamp 1666199351
transform 1 0 38916 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1666199351
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1666199351
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1666199351
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1666199351
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1666199351
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1666199351
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1666199351
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1666199351
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1666199351
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1666199351
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_513
timestamp 1666199351
transform 1 0 48300 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1666199351
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1666199351
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1666199351
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1666199351
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1666199351
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1666199351
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1666199351
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1666199351
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1666199351
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1666199351
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1666199351
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1666199351
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1666199351
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1666199351
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1666199351
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1666199351
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1666199351
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1666199351
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1666199351
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1666199351
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1666199351
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1666199351
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1666199351
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1666199351
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_225
timestamp 1666199351
transform 1 0 21804 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_233
timestamp 1666199351
transform 1 0 22540 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_239
timestamp 1666199351
transform 1 0 23092 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_246
timestamp 1666199351
transform 1 0 23736 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_255
timestamp 1666199351
transform 1 0 24564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_264
timestamp 1666199351
transform 1 0 25392 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1666199351
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1666199351
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_281
timestamp 1666199351
transform 1 0 26956 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_290
timestamp 1666199351
transform 1 0 27784 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_296
timestamp 1666199351
transform 1 0 28336 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_300
timestamp 1666199351
transform 1 0 28704 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_313
timestamp 1666199351
transform 1 0 29900 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_319
timestamp 1666199351
transform 1 0 30452 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_328
timestamp 1666199351
transform 1 0 31280 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_334
timestamp 1666199351
transform 1 0 31832 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_337
timestamp 1666199351
transform 1 0 32108 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_344
timestamp 1666199351
transform 1 0 32752 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_351
timestamp 1666199351
transform 1 0 33396 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_358
timestamp 1666199351
transform 1 0 34040 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_365
timestamp 1666199351
transform 1 0 34684 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_371
timestamp 1666199351
transform 1 0 35236 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_377
timestamp 1666199351
transform 1 0 35788 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_383
timestamp 1666199351
transform 1 0 36340 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_390
timestamp 1666199351
transform 1 0 36984 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_393
timestamp 1666199351
transform 1 0 37260 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_397
timestamp 1666199351
transform 1 0 37628 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_403
timestamp 1666199351
transform 1 0 38180 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_409
timestamp 1666199351
transform 1 0 38732 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_415
timestamp 1666199351
transform 1 0 39284 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_427
timestamp 1666199351
transform 1 0 40388 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_439
timestamp 1666199351
transform 1 0 41492 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1666199351
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1666199351
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1666199351
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1666199351
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1666199351
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1666199351
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1666199351
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_505
timestamp 1666199351
transform 1 0 47564 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_513
timestamp 1666199351
transform 1 0 48300 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1666199351
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1666199351
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1666199351
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1666199351
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1666199351
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1666199351
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1666199351
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1666199351
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1666199351
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1666199351
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1666199351
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1666199351
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1666199351
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1666199351
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1666199351
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1666199351
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1666199351
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1666199351
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1666199351
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1666199351
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1666199351
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1666199351
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_209
timestamp 1666199351
transform 1 0 20332 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_213
timestamp 1666199351
transform 1 0 20700 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_219
timestamp 1666199351
transform 1 0 21252 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_226
timestamp 1666199351
transform 1 0 21896 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_232
timestamp 1666199351
transform 1 0 22448 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_246
timestamp 1666199351
transform 1 0 23736 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_76_253
timestamp 1666199351
transform 1 0 24380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_268
timestamp 1666199351
transform 1 0 25760 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_275
timestamp 1666199351
transform 1 0 26404 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_292
timestamp 1666199351
transform 1 0 27968 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_299
timestamp 1666199351
transform 1 0 28612 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_306
timestamp 1666199351
transform 1 0 29256 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_309
timestamp 1666199351
transform 1 0 29532 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_314
timestamp 1666199351
transform 1 0 29992 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_322
timestamp 1666199351
transform 1 0 30728 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_326
timestamp 1666199351
transform 1 0 31096 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_335
timestamp 1666199351
transform 1 0 31924 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_344
timestamp 1666199351
transform 1 0 32752 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_353
timestamp 1666199351
transform 1 0 33580 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_362
timestamp 1666199351
transform 1 0 34408 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_365
timestamp 1666199351
transform 1 0 34684 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_369
timestamp 1666199351
transform 1 0 35052 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_380
timestamp 1666199351
transform 1 0 36064 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_391
timestamp 1666199351
transform 1 0 37076 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_402
timestamp 1666199351
transform 1 0 38088 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_408
timestamp 1666199351
transform 1 0 38640 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_414
timestamp 1666199351
transform 1 0 39192 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_76_421
timestamp 1666199351
transform 1 0 39836 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_425
timestamp 1666199351
transform 1 0 40204 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_437
timestamp 1666199351
transform 1 0 41308 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_449
timestamp 1666199351
transform 1 0 42412 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_461
timestamp 1666199351
transform 1 0 43516 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_473
timestamp 1666199351
transform 1 0 44620 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1666199351
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1666199351
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1666199351
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_513
timestamp 1666199351
transform 1 0 48300 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1666199351
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1666199351
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1666199351
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1666199351
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1666199351
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1666199351
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1666199351
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1666199351
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1666199351
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1666199351
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1666199351
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1666199351
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1666199351
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1666199351
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1666199351
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1666199351
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1666199351
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1666199351
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1666199351
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1666199351
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_193
timestamp 1666199351
transform 1 0 18860 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_197
timestamp 1666199351
transform 1 0 19228 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_77_206
timestamp 1666199351
transform 1 0 20056 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_215
timestamp 1666199351
transform 1 0 20884 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_222
timestamp 1666199351
transform 1 0 21528 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_225
timestamp 1666199351
transform 1 0 21804 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_229
timestamp 1666199351
transform 1 0 22172 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_233
timestamp 1666199351
transform 1 0 22540 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_242
timestamp 1666199351
transform 1 0 23368 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_253
timestamp 1666199351
transform 1 0 24380 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_259
timestamp 1666199351
transform 1 0 24932 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_270
timestamp 1666199351
transform 1 0 25944 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_77_277
timestamp 1666199351
transform 1 0 26588 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_281
timestamp 1666199351
transform 1 0 26956 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_290
timestamp 1666199351
transform 1 0 27784 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_298
timestamp 1666199351
transform 1 0 28520 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_312
timestamp 1666199351
transform 1 0 29808 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_316
timestamp 1666199351
transform 1 0 30176 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_330
timestamp 1666199351
transform 1 0 31464 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_337
timestamp 1666199351
transform 1 0 32108 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_341
timestamp 1666199351
transform 1 0 32476 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_355
timestamp 1666199351
transform 1 0 33764 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_364
timestamp 1666199351
transform 1 0 34592 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_372
timestamp 1666199351
transform 1 0 35328 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_386
timestamp 1666199351
transform 1 0 36616 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_393
timestamp 1666199351
transform 1 0 37260 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_403
timestamp 1666199351
transform 1 0 38180 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_414
timestamp 1666199351
transform 1 0 39192 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_420
timestamp 1666199351
transform 1 0 39744 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_426
timestamp 1666199351
transform 1 0 40296 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_432
timestamp 1666199351
transform 1 0 40848 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_438
timestamp 1666199351
transform 1 0 41400 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_446
timestamp 1666199351
transform 1 0 42136 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1666199351
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1666199351
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1666199351
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1666199351
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1666199351
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1666199351
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_505
timestamp 1666199351
transform 1 0 47564 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_513
timestamp 1666199351
transform 1 0 48300 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1666199351
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1666199351
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1666199351
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1666199351
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1666199351
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1666199351
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1666199351
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1666199351
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1666199351
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1666199351
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1666199351
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1666199351
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1666199351
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1666199351
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1666199351
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1666199351
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1666199351
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1666199351
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1666199351
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_189
timestamp 1666199351
transform 1 0 18492 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_194
timestamp 1666199351
transform 1 0 18952 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_197
timestamp 1666199351
transform 1 0 19228 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_206
timestamp 1666199351
transform 1 0 20056 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_213
timestamp 1666199351
transform 1 0 20700 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_222
timestamp 1666199351
transform 1 0 21528 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_230
timestamp 1666199351
transform 1 0 22264 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_238
timestamp 1666199351
transform 1 0 23000 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_250
timestamp 1666199351
transform 1 0 24104 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_253
timestamp 1666199351
transform 1 0 24380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_258
timestamp 1666199351
transform 1 0 24840 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_262
timestamp 1666199351
transform 1 0 25208 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_272
timestamp 1666199351
transform 1 0 26128 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_283
timestamp 1666199351
transform 1 0 27140 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_295
timestamp 1666199351
transform 1 0 28244 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_306
timestamp 1666199351
transform 1 0 29256 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_309
timestamp 1666199351
transform 1 0 29532 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_324
timestamp 1666199351
transform 1 0 30912 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_332
timestamp 1666199351
transform 1 0 31648 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_341
timestamp 1666199351
transform 1 0 32476 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_347
timestamp 1666199351
transform 1 0 33028 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_358
timestamp 1666199351
transform 1 0 34040 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_365
timestamp 1666199351
transform 1 0 34684 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_380
timestamp 1666199351
transform 1 0 36064 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_388
timestamp 1666199351
transform 1 0 36800 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_398
timestamp 1666199351
transform 1 0 37720 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_410
timestamp 1666199351
transform 1 0 38824 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_78_417
timestamp 1666199351
transform 1 0 39468 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_421
timestamp 1666199351
transform 1 0 39836 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_425
timestamp 1666199351
transform 1 0 40204 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_431
timestamp 1666199351
transform 1 0 40756 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_437
timestamp 1666199351
transform 1 0 41308 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_443
timestamp 1666199351
transform 1 0 41860 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_449
timestamp 1666199351
transform 1 0 42412 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_461
timestamp 1666199351
transform 1 0 43516 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_473
timestamp 1666199351
transform 1 0 44620 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1666199351
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1666199351
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1666199351
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_513
timestamp 1666199351
transform 1 0 48300 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1666199351
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1666199351
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1666199351
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1666199351
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1666199351
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1666199351
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1666199351
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1666199351
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1666199351
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1666199351
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1666199351
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1666199351
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1666199351
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1666199351
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1666199351
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1666199351
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1666199351
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1666199351
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_169
timestamp 1666199351
transform 1 0 16652 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_177
timestamp 1666199351
transform 1 0 17388 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_181
timestamp 1666199351
transform 1 0 17756 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_188
timestamp 1666199351
transform 1 0 18400 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_195
timestamp 1666199351
transform 1 0 19044 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_202
timestamp 1666199351
transform 1 0 19688 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_211
timestamp 1666199351
transform 1 0 20516 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_79_222
timestamp 1666199351
transform 1 0 21528 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_225
timestamp 1666199351
transform 1 0 21804 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_237
timestamp 1666199351
transform 1 0 22908 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_248
timestamp 1666199351
transform 1 0 23920 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_259
timestamp 1666199351
transform 1 0 24932 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_263
timestamp 1666199351
transform 1 0 25300 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_267
timestamp 1666199351
transform 1 0 25668 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1666199351
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_281
timestamp 1666199351
transform 1 0 26956 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_285
timestamp 1666199351
transform 1 0 27324 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_298
timestamp 1666199351
transform 1 0 28520 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_310
timestamp 1666199351
transform 1 0 29624 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_322
timestamp 1666199351
transform 1 0 30728 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_333
timestamp 1666199351
transform 1 0 31740 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_337
timestamp 1666199351
transform 1 0 32108 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_346
timestamp 1666199351
transform 1 0 32936 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_350
timestamp 1666199351
transform 1 0 33304 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_360
timestamp 1666199351
transform 1 0 34224 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_371
timestamp 1666199351
transform 1 0 35236 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_382
timestamp 1666199351
transform 1 0 36248 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_389
timestamp 1666199351
transform 1 0 36892 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_79_393
timestamp 1666199351
transform 1 0 37260 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_407
timestamp 1666199351
transform 1 0 38548 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_414
timestamp 1666199351
transform 1 0 39192 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_421
timestamp 1666199351
transform 1 0 39836 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_428
timestamp 1666199351
transform 1 0 40480 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_435
timestamp 1666199351
transform 1 0 41124 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1666199351
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1666199351
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_449
timestamp 1666199351
transform 1 0 42412 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_453
timestamp 1666199351
transform 1 0 42780 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_465
timestamp 1666199351
transform 1 0 43884 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_477
timestamp 1666199351
transform 1 0 44988 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_489
timestamp 1666199351
transform 1 0 46092 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_501
timestamp 1666199351
transform 1 0 47196 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_505
timestamp 1666199351
transform 1 0 47564 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_513
timestamp 1666199351
transform 1 0 48300 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1666199351
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1666199351
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1666199351
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1666199351
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1666199351
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1666199351
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1666199351
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1666199351
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1666199351
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1666199351
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1666199351
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1666199351
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1666199351
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1666199351
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1666199351
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1666199351
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1666199351
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_165
timestamp 1666199351
transform 1 0 16284 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_171
timestamp 1666199351
transform 1 0 16836 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_178
timestamp 1666199351
transform 1 0 17480 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_185
timestamp 1666199351
transform 1 0 18124 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_194
timestamp 1666199351
transform 1 0 18952 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_197
timestamp 1666199351
transform 1 0 19228 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_208
timestamp 1666199351
transform 1 0 20240 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_212
timestamp 1666199351
transform 1 0 20608 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_218
timestamp 1666199351
transform 1 0 21160 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_227
timestamp 1666199351
transform 1 0 21988 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_236
timestamp 1666199351
transform 1 0 22816 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_249
timestamp 1666199351
transform 1 0 24012 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_253
timestamp 1666199351
transform 1 0 24380 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_263
timestamp 1666199351
transform 1 0 25300 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_269
timestamp 1666199351
transform 1 0 25852 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_280
timestamp 1666199351
transform 1 0 26864 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_286
timestamp 1666199351
transform 1 0 27416 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_294
timestamp 1666199351
transform 1 0 28152 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_298
timestamp 1666199351
transform 1 0 28520 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_306
timestamp 1666199351
transform 1 0 29256 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_309
timestamp 1666199351
transform 1 0 29532 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_318
timestamp 1666199351
transform 1 0 30360 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_325
timestamp 1666199351
transform 1 0 31004 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_329
timestamp 1666199351
transform 1 0 31372 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_337
timestamp 1666199351
transform 1 0 32108 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_344
timestamp 1666199351
transform 1 0 32752 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_348
timestamp 1666199351
transform 1 0 33120 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_362
timestamp 1666199351
transform 1 0 34408 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_365
timestamp 1666199351
transform 1 0 34684 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_376
timestamp 1666199351
transform 1 0 35696 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_380
timestamp 1666199351
transform 1 0 36064 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_389
timestamp 1666199351
transform 1 0 36892 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_400
timestamp 1666199351
transform 1 0 37904 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_404
timestamp 1666199351
transform 1 0 38272 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_412
timestamp 1666199351
transform 1 0 39008 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_418
timestamp 1666199351
transform 1 0 39560 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_421
timestamp 1666199351
transform 1 0 39836 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_426
timestamp 1666199351
transform 1 0 40296 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_433
timestamp 1666199351
transform 1 0 40940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_440
timestamp 1666199351
transform 1 0 41584 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_447
timestamp 1666199351
transform 1 0 42228 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_454
timestamp 1666199351
transform 1 0 42872 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_460
timestamp 1666199351
transform 1 0 43424 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_472
timestamp 1666199351
transform 1 0 44528 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1666199351
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1666199351
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1666199351
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_513
timestamp 1666199351
transform 1 0 48300 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1666199351
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1666199351
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1666199351
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1666199351
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1666199351
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1666199351
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_57
timestamp 1666199351
transform 1 0 6348 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_64
timestamp 1666199351
transform 1 0 6992 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_76
timestamp 1666199351
transform 1 0 8096 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_88
timestamp 1666199351
transform 1 0 9200 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_100
timestamp 1666199351
transform 1 0 10304 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1666199351
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1666199351
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_137
timestamp 1666199351
transform 1 0 13708 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_148
timestamp 1666199351
transform 1 0 14720 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_160
timestamp 1666199351
transform 1 0 15824 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_166
timestamp 1666199351
transform 1 0 16376 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_169
timestamp 1666199351
transform 1 0 16652 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_173
timestamp 1666199351
transform 1 0 17020 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_177
timestamp 1666199351
transform 1 0 17388 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_184
timestamp 1666199351
transform 1 0 18032 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_191
timestamp 1666199351
transform 1 0 18676 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_198
timestamp 1666199351
transform 1 0 19320 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_207
timestamp 1666199351
transform 1 0 20148 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_81_222
timestamp 1666199351
transform 1 0 21528 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_225
timestamp 1666199351
transform 1 0 21804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_229
timestamp 1666199351
transform 1 0 22172 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_235
timestamp 1666199351
transform 1 0 22724 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_248
timestamp 1666199351
transform 1 0 23920 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_254
timestamp 1666199351
transform 1 0 24472 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_265
timestamp 1666199351
transform 1 0 25484 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_278
timestamp 1666199351
transform 1 0 26680 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_281
timestamp 1666199351
transform 1 0 26956 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_291
timestamp 1666199351
transform 1 0 27876 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_300
timestamp 1666199351
transform 1 0 28704 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_312
timestamp 1666199351
transform 1 0 29808 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_326
timestamp 1666199351
transform 1 0 31096 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_333
timestamp 1666199351
transform 1 0 31740 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_337
timestamp 1666199351
transform 1 0 32108 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_342
timestamp 1666199351
transform 1 0 32568 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_356
timestamp 1666199351
transform 1 0 33856 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_360
timestamp 1666199351
transform 1 0 34224 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_368
timestamp 1666199351
transform 1 0 34960 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_381
timestamp 1666199351
transform 1 0 36156 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_388
timestamp 1666199351
transform 1 0 36800 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_393
timestamp 1666199351
transform 1 0 37260 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_404
timestamp 1666199351
transform 1 0 38272 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_415
timestamp 1666199351
transform 1 0 39284 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_422
timestamp 1666199351
transform 1 0 39928 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_429
timestamp 1666199351
transform 1 0 40572 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_436
timestamp 1666199351
transform 1 0 41216 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_443
timestamp 1666199351
transform 1 0 41860 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1666199351
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_449
timestamp 1666199351
transform 1 0 42412 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_454
timestamp 1666199351
transform 1 0 42872 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_461
timestamp 1666199351
transform 1 0 43516 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_468
timestamp 1666199351
transform 1 0 44160 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_475
timestamp 1666199351
transform 1 0 44804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_487
timestamp 1666199351
transform 1 0 45908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_499
timestamp 1666199351
transform 1 0 47012 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1666199351
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_505
timestamp 1666199351
transform 1 0 47564 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_513
timestamp 1666199351
transform 1 0 48300 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1666199351
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1666199351
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1666199351
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_29
timestamp 1666199351
transform 1 0 3772 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_40
timestamp 1666199351
transform 1 0 4784 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_47
timestamp 1666199351
transform 1 0 5428 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_54
timestamp 1666199351
transform 1 0 6072 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_57
timestamp 1666199351
transform 1 0 6348 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_66
timestamp 1666199351
transform 1 0 7176 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_73
timestamp 1666199351
transform 1 0 7820 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_80
timestamp 1666199351
transform 1 0 8464 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_85
timestamp 1666199351
transform 1 0 8924 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_90
timestamp 1666199351
transform 1 0 9384 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_96
timestamp 1666199351
transform 1 0 9936 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_100
timestamp 1666199351
transform 1 0 10304 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_106
timestamp 1666199351
transform 1 0 10856 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_110
timestamp 1666199351
transform 1 0 11224 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_113
timestamp 1666199351
transform 1 0 11500 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_124
timestamp 1666199351
transform 1 0 12512 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_132
timestamp 1666199351
transform 1 0 13248 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_136
timestamp 1666199351
transform 1 0 13616 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_141
timestamp 1666199351
transform 1 0 14076 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_152
timestamp 1666199351
transform 1 0 15088 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_159
timestamp 1666199351
transform 1 0 15732 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_166
timestamp 1666199351
transform 1 0 16376 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_169
timestamp 1666199351
transform 1 0 16652 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_173
timestamp 1666199351
transform 1 0 17020 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_180
timestamp 1666199351
transform 1 0 17664 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_187
timestamp 1666199351
transform 1 0 18308 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1666199351
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_197
timestamp 1666199351
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_208
timestamp 1666199351
transform 1 0 20240 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_221
timestamp 1666199351
transform 1 0 21436 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_225
timestamp 1666199351
transform 1 0 21804 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_235
timestamp 1666199351
transform 1 0 22724 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_241
timestamp 1666199351
transform 1 0 23276 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1666199351
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1666199351
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_262
timestamp 1666199351
transform 1 0 25208 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_273
timestamp 1666199351
transform 1 0 26220 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_279
timestamp 1666199351
transform 1 0 26772 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_281
timestamp 1666199351
transform 1 0 26956 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_286
timestamp 1666199351
transform 1 0 27416 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_293
timestamp 1666199351
transform 1 0 28060 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_82_306
timestamp 1666199351
transform 1 0 29256 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1666199351
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_314
timestamp 1666199351
transform 1 0 29992 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_318
timestamp 1666199351
transform 1 0 30360 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_326
timestamp 1666199351
transform 1 0 31096 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_333
timestamp 1666199351
transform 1 0 31740 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_337
timestamp 1666199351
transform 1 0 32108 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_346
timestamp 1666199351
transform 1 0 32936 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1666199351
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1666199351
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_365
timestamp 1666199351
transform 1 0 34684 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_370
timestamp 1666199351
transform 1 0 35144 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_377
timestamp 1666199351
transform 1 0 35788 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_384
timestamp 1666199351
transform 1 0 36432 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_390
timestamp 1666199351
transform 1 0 36984 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_393
timestamp 1666199351
transform 1 0 37260 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_402
timestamp 1666199351
transform 1 0 38088 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_409
timestamp 1666199351
transform 1 0 38732 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_416
timestamp 1666199351
transform 1 0 39376 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_421
timestamp 1666199351
transform 1 0 39836 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_426
timestamp 1666199351
transform 1 0 40296 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_433
timestamp 1666199351
transform 1 0 40940 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_440
timestamp 1666199351
transform 1 0 41584 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_446
timestamp 1666199351
transform 1 0 42136 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1666199351
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_454
timestamp 1666199351
transform 1 0 42872 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_461
timestamp 1666199351
transform 1 0 43516 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_468
timestamp 1666199351
transform 1 0 44160 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_474
timestamp 1666199351
transform 1 0 44712 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1666199351
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_482
timestamp 1666199351
transform 1 0 45448 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_489
timestamp 1666199351
transform 1 0 46092 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_496
timestamp 1666199351
transform 1 0 46736 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_505
timestamp 1666199351
transform 1 0 47564 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_513
timestamp 1666199351
transform 1 0 48300 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666199351
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666199351
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666199351
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666199351
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666199351
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666199351
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666199351
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666199351
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666199351
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666199351
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666199351
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666199351
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666199351
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666199351
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666199351
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666199351
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666199351
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666199351
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666199351
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666199351
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666199351
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666199351
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666199351
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666199351
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666199351
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666199351
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666199351
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666199351
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666199351
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666199351
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666199351
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666199351
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666199351
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666199351
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666199351
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666199351
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666199351
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666199351
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666199351
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666199351
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666199351
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666199351
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666199351
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666199351
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666199351
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666199351
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666199351
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666199351
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666199351
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666199351
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666199351
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666199351
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666199351
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666199351
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666199351
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666199351
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666199351
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666199351
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666199351
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666199351
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666199351
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666199351
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666199351
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666199351
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666199351
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666199351
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666199351
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666199351
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666199351
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666199351
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666199351
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666199351
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666199351
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666199351
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666199351
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666199351
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666199351
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666199351
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666199351
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666199351
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666199351
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666199351
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666199351
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666199351
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666199351
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666199351
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666199351
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666199351
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666199351
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666199351
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666199351
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666199351
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666199351
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666199351
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666199351
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666199351
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666199351
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666199351
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666199351
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666199351
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666199351
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666199351
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666199351
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666199351
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666199351
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666199351
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666199351
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666199351
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666199351
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666199351
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666199351
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666199351
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666199351
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666199351
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666199351
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666199351
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666199351
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666199351
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666199351
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666199351
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666199351
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666199351
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666199351
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666199351
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666199351
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666199351
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666199351
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666199351
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666199351
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666199351
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666199351
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666199351
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666199351
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666199351
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666199351
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666199351
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666199351
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666199351
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666199351
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666199351
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666199351
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666199351
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666199351
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666199351
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666199351
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666199351
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666199351
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666199351
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666199351
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666199351
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666199351
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666199351
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666199351
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666199351
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666199351
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666199351
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666199351
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666199351
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666199351
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666199351
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666199351
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666199351
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666199351
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666199351
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666199351
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666199351
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666199351
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666199351
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666199351
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666199351
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666199351
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666199351
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666199351
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666199351
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666199351
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666199351
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666199351
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666199351
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666199351
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666199351
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666199351
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666199351
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666199351
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666199351
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666199351
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666199351
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666199351
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666199351
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666199351
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666199351
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666199351
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666199351
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666199351
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666199351
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666199351
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666199351
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666199351
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666199351
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666199351
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666199351
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666199351
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666199351
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666199351
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666199351
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666199351
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666199351
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666199351
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666199351
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666199351
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666199351
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666199351
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666199351
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666199351
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666199351
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666199351
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666199351
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666199351
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666199351
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666199351
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666199351
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666199351
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666199351
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666199351
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666199351
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666199351
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666199351
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666199351
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666199351
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666199351
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666199351
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666199351
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666199351
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666199351
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666199351
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666199351
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666199351
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666199351
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666199351
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666199351
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666199351
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666199351
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666199351
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666199351
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666199351
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666199351
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666199351
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666199351
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666199351
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666199351
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666199351
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666199351
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666199351
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666199351
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666199351
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666199351
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666199351
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666199351
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666199351
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666199351
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666199351
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666199351
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666199351
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666199351
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666199351
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666199351
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666199351
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666199351
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666199351
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666199351
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666199351
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666199351
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666199351
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666199351
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666199351
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666199351
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666199351
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666199351
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666199351
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666199351
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666199351
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666199351
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666199351
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666199351
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666199351
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666199351
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666199351
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666199351
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666199351
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666199351
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666199351
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666199351
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666199351
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666199351
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666199351
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666199351
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666199351
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666199351
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666199351
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666199351
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666199351
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666199351
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666199351
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666199351
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666199351
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666199351
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666199351
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666199351
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666199351
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666199351
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666199351
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666199351
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666199351
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666199351
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666199351
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666199351
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666199351
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666199351
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666199351
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666199351
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666199351
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666199351
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666199351
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666199351
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666199351
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666199351
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666199351
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666199351
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666199351
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666199351
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666199351
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666199351
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666199351
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666199351
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666199351
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666199351
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666199351
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666199351
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666199351
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666199351
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666199351
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666199351
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666199351
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666199351
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666199351
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666199351
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666199351
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666199351
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666199351
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666199351
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666199351
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666199351
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666199351
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666199351
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666199351
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666199351
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666199351
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666199351
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666199351
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666199351
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666199351
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666199351
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666199351
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666199351
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666199351
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666199351
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666199351
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666199351
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666199351
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666199351
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666199351
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666199351
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666199351
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666199351
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666199351
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666199351
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666199351
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666199351
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666199351
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666199351
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666199351
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666199351
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666199351
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666199351
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666199351
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666199351
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666199351
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666199351
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666199351
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666199351
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666199351
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666199351
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666199351
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666199351
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666199351
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666199351
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666199351
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666199351
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666199351
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666199351
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666199351
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666199351
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666199351
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666199351
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666199351
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666199351
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666199351
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666199351
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666199351
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666199351
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666199351
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666199351
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666199351
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666199351
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666199351
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666199351
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666199351
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666199351
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666199351
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666199351
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666199351
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666199351
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666199351
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666199351
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666199351
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666199351
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666199351
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666199351
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666199351
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666199351
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666199351
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666199351
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666199351
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666199351
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666199351
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666199351
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666199351
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666199351
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666199351
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666199351
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666199351
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666199351
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666199351
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666199351
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666199351
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666199351
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666199351
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666199351
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666199351
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666199351
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666199351
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666199351
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666199351
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666199351
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666199351
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666199351
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666199351
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666199351
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666199351
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666199351
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666199351
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666199351
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666199351
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666199351
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666199351
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666199351
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666199351
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666199351
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666199351
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666199351
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666199351
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666199351
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666199351
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666199351
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666199351
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666199351
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666199351
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666199351
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666199351
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666199351
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666199351
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666199351
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666199351
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666199351
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666199351
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666199351
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666199351
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666199351
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666199351
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666199351
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666199351
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666199351
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666199351
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666199351
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666199351
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666199351
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666199351
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666199351
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666199351
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666199351
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666199351
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666199351
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666199351
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666199351
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666199351
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666199351
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666199351
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666199351
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666199351
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666199351
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666199351
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666199351
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666199351
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666199351
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666199351
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666199351
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666199351
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666199351
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666199351
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666199351
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666199351
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666199351
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666199351
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666199351
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666199351
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666199351
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666199351
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666199351
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666199351
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666199351
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666199351
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666199351
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666199351
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666199351
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666199351
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666199351
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666199351
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666199351
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666199351
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666199351
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666199351
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666199351
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666199351
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666199351
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666199351
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666199351
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666199351
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666199351
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666199351
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666199351
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666199351
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666199351
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666199351
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666199351
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666199351
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666199351
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666199351
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666199351
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666199351
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666199351
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666199351
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666199351
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666199351
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666199351
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666199351
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666199351
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666199351
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666199351
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666199351
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666199351
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666199351
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666199351
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666199351
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666199351
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666199351
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666199351
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666199351
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666199351
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666199351
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666199351
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666199351
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666199351
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666199351
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666199351
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666199351
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666199351
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666199351
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666199351
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666199351
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666199351
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666199351
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666199351
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666199351
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666199351
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666199351
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666199351
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666199351
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666199351
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666199351
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666199351
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666199351
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666199351
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666199351
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666199351
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666199351
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666199351
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666199351
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666199351
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666199351
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666199351
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666199351
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666199351
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666199351
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666199351
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666199351
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666199351
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666199351
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666199351
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666199351
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666199351
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666199351
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666199351
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666199351
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666199351
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666199351
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666199351
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666199351
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666199351
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666199351
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666199351
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666199351
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666199351
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666199351
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666199351
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666199351
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666199351
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666199351
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666199351
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666199351
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666199351
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666199351
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666199351
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666199351
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666199351
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666199351
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666199351
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666199351
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666199351
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666199351
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666199351
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666199351
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666199351
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666199351
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666199351
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666199351
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666199351
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666199351
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666199351
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666199351
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666199351
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666199351
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666199351
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666199351
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666199351
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666199351
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666199351
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666199351
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666199351
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666199351
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666199351
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666199351
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666199351
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666199351
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666199351
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666199351
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666199351
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666199351
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666199351
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666199351
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666199351
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666199351
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666199351
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666199351
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666199351
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666199351
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666199351
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666199351
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666199351
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666199351
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666199351
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666199351
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666199351
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666199351
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666199351
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666199351
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666199351
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666199351
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666199351
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666199351
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666199351
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666199351
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666199351
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666199351
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666199351
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666199351
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666199351
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666199351
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666199351
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666199351
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666199351
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666199351
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666199351
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666199351
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666199351
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666199351
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666199351
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666199351
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666199351
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666199351
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666199351
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666199351
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666199351
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666199351
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666199351
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666199351
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666199351
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666199351
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666199351
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666199351
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666199351
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666199351
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666199351
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666199351
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666199351
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666199351
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666199351
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666199351
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666199351
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666199351
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666199351
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666199351
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666199351
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666199351
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666199351
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666199351
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666199351
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666199351
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666199351
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666199351
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666199351
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666199351
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666199351
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666199351
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666199351
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666199351
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666199351
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666199351
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666199351
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666199351
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666199351
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666199351
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666199351
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666199351
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666199351
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666199351
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666199351
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666199351
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666199351
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666199351
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666199351
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666199351
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666199351
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666199351
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666199351
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666199351
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666199351
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666199351
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666199351
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666199351
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666199351
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666199351
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666199351
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666199351
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666199351
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666199351
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666199351
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666199351
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666199351
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666199351
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666199351
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666199351
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666199351
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666199351
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666199351
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666199351
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666199351
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666199351
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666199351
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666199351
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666199351
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666199351
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666199351
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666199351
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666199351
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666199351
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666199351
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666199351
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666199351
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666199351
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666199351
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666199351
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666199351
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666199351
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666199351
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666199351
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666199351
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666199351
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666199351
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666199351
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666199351
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666199351
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666199351
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666199351
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666199351
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666199351
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666199351
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666199351
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666199351
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666199351
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666199351
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666199351
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666199351
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666199351
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666199351
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666199351
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666199351
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666199351
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666199351
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666199351
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666199351
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666199351
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666199351
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666199351
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666199351
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666199351
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666199351
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666199351
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666199351
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666199351
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666199351
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666199351
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666199351
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666199351
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666199351
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666199351
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666199351
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666199351
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666199351
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666199351
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666199351
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666199351
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666199351
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666199351
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666199351
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666199351
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666199351
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666199351
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666199351
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666199351
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666199351
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666199351
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666199351
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666199351
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666199351
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666199351
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666199351
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666199351
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666199351
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666199351
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666199351
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666199351
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666199351
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666199351
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666199351
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666199351
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666199351
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666199351
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666199351
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666199351
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666199351
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666199351
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666199351
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666199351
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666199351
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666199351
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666199351
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666199351
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666199351
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666199351
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666199351
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666199351
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666199351
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666199351
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666199351
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666199351
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666199351
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666199351
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666199351
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666199351
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666199351
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666199351
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666199351
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666199351
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666199351
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666199351
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666199351
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666199351
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666199351
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666199351
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666199351
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666199351
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666199351
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666199351
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666199351
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666199351
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666199351
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666199351
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666199351
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666199351
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666199351
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666199351
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _170_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 21252 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _171_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 21620 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _172_
timestamp 1666199351
transform -1 0 22264 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _173_
timestamp 1666199351
transform 1 0 29716 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1666199351
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1666199351
transform -1 0 29992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1666199351
transform -1 0 30636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1666199351
transform -1 0 30636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1666199351
transform -1 0 29992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _179_
timestamp 1666199351
transform -1 0 27048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1666199351
transform -1 0 27692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1666199351
transform -1 0 28244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1666199351
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1666199351
transform 1 0 28428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1666199351
transform -1 0 26680 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _185_
timestamp 1666199351
transform -1 0 25300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1666199351
transform 1 0 26588 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1666199351
transform 1 0 25668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1666199351
transform -1 0 26036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1666199351
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1666199351
transform -1 0 24104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _191_
timestamp 1666199351
transform -1 0 22356 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1666199351
transform 1 0 24380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _193_
timestamp 1666199351
transform 1 0 24564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _194_
timestamp 1666199351
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _195_
timestamp 1666199351
transform 1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1666199351
transform -1 0 20516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _197_
timestamp 1666199351
transform -1 0 22540 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp 1666199351
transform 1 0 22632 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1666199351
transform 1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1666199351
transform 1 0 20148 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1666199351
transform -1 0 19596 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1666199351
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _203_
timestamp 1666199351
transform -1 0 20884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1666199351
transform -1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 1666199351
transform 1 0 19596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _206_
timestamp 1666199351
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _207_
timestamp 1666199351
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _208_
timestamp 1666199351
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _209_
timestamp 1666199351
transform -1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _210_
timestamp 1666199351
transform -1 0 29256 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _211_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 29256 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _212_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 30728 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _213_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 30912 0 1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _214_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 22816 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _215_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 29716 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _216_
timestamp 1666199351
transform -1 0 29808 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _217_
timestamp 1666199351
transform -1 0 23368 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _218_
timestamp 1666199351
transform -1 0 32568 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _219_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 27692 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_2  _220_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 28888 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _221_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 29256 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_2  _222_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 26036 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _223_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 27508 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1666199351
transform 1 0 28336 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _225_
timestamp 1666199351
transform -1 0 27784 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _226_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 23644 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1666199351
transform 1 0 24564 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _228_
timestamp 1666199351
transform -1 0 24564 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1666199351
transform -1 0 23736 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _230_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 23368 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _231_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 28612 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _232_
timestamp 1666199351
transform 1 0 23276 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _233_
timestamp 1666199351
transform -1 0 25668 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _234_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 24288 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _235_
timestamp 1666199351
transform -1 0 21528 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _236_
timestamp 1666199351
transform -1 0 39836 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _237_
timestamp 1666199351
transform -1 0 39008 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _238_
timestamp 1666199351
transform 1 0 37536 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _239_
timestamp 1666199351
transform -1 0 34408 0 1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _240_
timestamp 1666199351
transform -1 0 32752 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _241_
timestamp 1666199351
transform 1 0 38548 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _242_
timestamp 1666199351
transform -1 0 36064 0 1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _243_
timestamp 1666199351
transform -1 0 33580 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _244_
timestamp 1666199351
transform -1 0 39192 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _245_
timestamp 1666199351
transform 1 0 36892 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_2  _246_
timestamp 1666199351
transform 1 0 38088 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_2  _247_
timestamp 1666199351
transform -1 0 38548 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _248_
timestamp 1666199351
transform 1 0 37444 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_2  _249_
timestamp 1666199351
transform -1 0 36248 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _250_
timestamp 1666199351
transform 1 0 37444 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1666199351
transform -1 0 36984 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _252_
timestamp 1666199351
transform 1 0 35420 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _253_
timestamp 1666199351
transform -1 0 31924 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1666199351
transform 1 0 36616 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _255_
timestamp 1666199351
transform -1 0 32752 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1666199351
transform 1 0 33120 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _257_
timestamp 1666199351
transform 1 0 31740 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _258_
timestamp 1666199351
transform -1 0 38088 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _259_
timestamp 1666199351
transform 1 0 31464 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _260_
timestamp 1666199351
transform -1 0 40480 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _261_
timestamp 1666199351
transform 1 0 32292 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _262_
timestamp 1666199351
transform -1 0 28704 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _263_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 29808 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _264_
timestamp 1666199351
transform -1 0 22908 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _265_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 21988 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1666199351
transform -1 0 27416 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _267_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 25852 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_2  _268_
timestamp 1666199351
transform 1 0 25576 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _269_
timestamp 1666199351
transform 1 0 24840 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1666199351
transform -1 0 41860 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _271_
timestamp 1666199351
transform 1 0 35328 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_2  _272_
timestamp 1666199351
transform 1 0 35052 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _273_
timestamp 1666199351
transform 1 0 34316 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _274_
timestamp 1666199351
transform -1 0 20700 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _275_
timestamp 1666199351
transform -1 0 18952 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1666199351
transform 1 0 18676 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _277_
timestamp 1666199351
transform 1 0 18952 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _278_
timestamp 1666199351
transform -1 0 21436 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1666199351
transform -1 0 18032 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _280_
timestamp 1666199351
transform 1 0 17112 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _281_
timestamp 1666199351
transform -1 0 20240 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_2  _282_
timestamp 1666199351
transform 1 0 27140 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _283_
timestamp 1666199351
transform -1 0 27968 0 1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_1  _284_
timestamp 1666199351
transform -1 0 31740 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _285_
timestamp 1666199351
transform 1 0 27508 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _286_
timestamp 1666199351
transform 1 0 27140 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _287_
timestamp 1666199351
transform 1 0 26220 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_2  _288_
timestamp 1666199351
transform -1 0 37076 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _289_
timestamp 1666199351
transform 1 0 35420 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_1  _290_
timestamp 1666199351
transform -1 0 41584 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _291_
timestamp 1666199351
transform 1 0 38640 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _292_
timestamp 1666199351
transform 1 0 36156 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _293_
timestamp 1666199351
transform 1 0 37260 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _294_
timestamp 1666199351
transform -1 0 20148 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1666199351
transform 1 0 19780 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _296_
timestamp 1666199351
transform -1 0 18400 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _297_
timestamp 1666199351
transform -1 0 20516 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1666199351
transform -1 0 19044 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _299_
timestamp 1666199351
transform 1 0 17848 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _300_
timestamp 1666199351
transform -1 0 20240 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _301_
timestamp 1666199351
transform -1 0 27140 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _302_
timestamp 1666199351
transform 1 0 25760 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _303_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 24564 0 1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _304_
timestamp 1666199351
transform 1 0 24932 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _305_
timestamp 1666199351
transform 1 0 25300 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _306_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 25300 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _307_
timestamp 1666199351
transform 1 0 34592 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _308_
timestamp 1666199351
transform 1 0 33948 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _309_
timestamp 1666199351
transform 1 0 32568 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _310_
timestamp 1666199351
transform -1 0 34592 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _311_
timestamp 1666199351
transform -1 0 34040 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _312_
timestamp 1666199351
transform 1 0 33396 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _313_
timestamp 1666199351
transform -1 0 21528 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1666199351
transform -1 0 20884 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _315_
timestamp 1666199351
transform -1 0 20056 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _316_
timestamp 1666199351
transform -1 0 21160 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1666199351
transform -1 0 19688 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _318_
timestamp 1666199351
transform 1 0 18400 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _319_
timestamp 1666199351
transform -1 0 21528 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _320_
timestamp 1666199351
transform -1 0 24380 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _321_
timestamp 1666199351
transform -1 0 23000 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1666199351
transform -1 0 22540 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _323_
timestamp 1666199351
transform -1 0 23736 0 1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _324_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 22724 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _325_
timestamp 1666199351
transform 1 0 24656 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _326_
timestamp 1666199351
transform 1 0 24564 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _327_
timestamp 1666199351
transform -1 0 21988 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _328_
timestamp 1666199351
transform 1 0 32292 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _329_
timestamp 1666199351
transform -1 0 31740 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1666199351
transform -1 0 31096 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _331_
timestamp 1666199351
transform -1 0 31464 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_2  _332_
timestamp 1666199351
transform 1 0 33304 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _333_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 32936 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_2  _334_
timestamp 1666199351
transform 1 0 30452 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _335_
timestamp 1666199351
transform 1 0 30176 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_2  _336_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 23092 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_2  _337_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 23184 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _338_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 40940 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _339_
timestamp 1666199351
transform -1 0 40296 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _340_
timestamp 1666199351
transform -1 0 39468 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _341_
timestamp 1666199351
transform -1 0 41584 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _342_
timestamp 1666199351
transform -1 0 43516 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _343_
timestamp 1666199351
transform -1 0 42872 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _344_
timestamp 1666199351
transform -1 0 42872 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _345_
timestamp 1666199351
transform -1 0 44160 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _346_
timestamp 1666199351
transform -1 0 44804 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _347_
timestamp 1666199351
transform -1 0 46092 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _348_
timestamp 1666199351
transform 1 0 5796 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _349_
timestamp 1666199351
transform 1 0 6900 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _350_
timestamp 1666199351
transform 1 0 8188 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _351_
timestamp 1666199351
transform -1 0 26404 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _352_
timestamp 1666199351
transform -1 0 28060 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _353_
timestamp 1666199351
transform -1 0 31740 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _354_
timestamp 1666199351
transform -1 0 32752 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _355_
timestamp 1666199351
transform -1 0 29992 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _356_
timestamp 1666199351
transform -1 0 36432 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _357_
timestamp 1666199351
transform -1 0 36800 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _358_
timestamp 1666199351
transform -1 0 39376 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _359_
timestamp 1666199351
transform -1 0 34684 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _360_
timestamp 1666199351
transform -1 0 39928 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _361_
timestamp 1666199351
transform -1 0 40572 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _362_
timestamp 1666199351
transform -1 0 41216 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _363_
timestamp 1666199351
transform -1 0 40940 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _364_
timestamp 1666199351
transform -1 0 42872 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _365_
timestamp 1666199351
transform -1 0 41124 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _366_
timestamp 1666199351
transform -1 0 42228 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _367_
timestamp 1666199351
transform -1 0 43516 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _368_
timestamp 1666199351
transform -1 0 44160 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _369_
timestamp 1666199351
transform -1 0 45448 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _370_
timestamp 1666199351
transform -1 0 46736 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _371_
timestamp 1666199351
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _372_
timestamp 1666199351
transform 1 0 12144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _373_
timestamp 1666199351
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _374_
timestamp 1666199351
transform 1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _375_
timestamp 1666199351
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _376_
timestamp 1666199351
transform 1 0 13432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _377_
timestamp 1666199351
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _378_
timestamp 1666199351
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _379_
timestamp 1666199351
transform 1 0 13524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _380_
timestamp 1666199351
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _381_
timestamp 1666199351
transform 1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _382_
timestamp 1666199351
transform 1 0 14168 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _383_
timestamp 1666199351
transform 1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _384_
timestamp 1666199351
transform 1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _385_
timestamp 1666199351
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _386_
timestamp 1666199351
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _387_
timestamp 1666199351
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _388_
timestamp 1666199351
transform 1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _389_
timestamp 1666199351
transform 1 0 17020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _390_
timestamp 1666199351
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _391_
timestamp 1666199351
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _392_
timestamp 1666199351
transform 1 0 17848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _393_
timestamp 1666199351
transform 1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _394_
timestamp 1666199351
transform 1 0 16744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _395_
timestamp 1666199351
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _396_
timestamp 1666199351
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _397_
timestamp 1666199351
transform 1 0 19228 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _398_
timestamp 1666199351
transform 1 0 18676 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _399_
timestamp 1666199351
transform 1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _400_
timestamp 1666199351
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _401_
timestamp 1666199351
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _402_
timestamp 1666199351
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _403_
timestamp 1666199351
transform -1 0 32568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _404_
timestamp 1666199351
transform -1 0 31280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _405_
timestamp 1666199351
transform -1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _406_
timestamp 1666199351
transform -1 0 32568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _407_
timestamp 1666199351
transform -1 0 31924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _408_
timestamp 1666199351
transform -1 0 33856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _409_
timestamp 1666199351
transform -1 0 33212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _410_
timestamp 1666199351
transform -1 0 32568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _411_
timestamp 1666199351
transform -1 0 33856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _412_
timestamp 1666199351
transform -1 0 33212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _413_
timestamp 1666199351
transform -1 0 34500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _414_
timestamp 1666199351
transform -1 0 33856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _415_
timestamp 1666199351
transform -1 0 35144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _416_
timestamp 1666199351
transform -1 0 35144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _417_
timestamp 1666199351
transform -1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _418_
timestamp 1666199351
transform -1 0 35788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _419_
timestamp 1666199351
transform -1 0 35144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _420_
timestamp 1666199351
transform -1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _421_
timestamp 1666199351
transform -1 0 35788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _422_
timestamp 1666199351
transform -1 0 36432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _423_
timestamp 1666199351
transform -1 0 37720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _424_
timestamp 1666199351
transform -1 0 36432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _425_
timestamp 1666199351
transform -1 0 37720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _426_
timestamp 1666199351
transform -1 0 37076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _427_
timestamp 1666199351
transform -1 0 38364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _428_
timestamp 1666199351
transform -1 0 37720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _429_
timestamp 1666199351
transform -1 0 38364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _430_
timestamp 1666199351
transform -1 0 39008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _431_
timestamp 1666199351
transform -1 0 38364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _432_
timestamp 1666199351
transform -1 0 39008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _433_
timestamp 1666199351
transform -1 0 39008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _434_
timestamp 1666199351
transform -1 0 40296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _435_
timestamp 1666199351
transform -1 0 39652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _436_
timestamp 1666199351
transform -1 0 40296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _437_
timestamp 1666199351
transform -1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _438_
timestamp 1666199351
transform -1 0 40296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _439_
timestamp 1666199351
transform -1 0 41584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _440_
timestamp 1666199351
transform -1 0 40940 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _441_
timestamp 1666199351
transform -1 0 40940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _442_
timestamp 1666199351
transform -1 0 41584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _443_
timestamp 1666199351
transform -1 0 41584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _444_
timestamp 1666199351
transform -1 0 42872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _445_
timestamp 1666199351
transform -1 0 42228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _446_
timestamp 1666199351
transform -1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _447_
timestamp 1666199351
transform -1 0 42872 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _448_
timestamp 1666199351
transform -1 0 44160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _449_
timestamp 1666199351
transform -1 0 43516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _450_
timestamp 1666199351
transform 1 0 42688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _451_
timestamp 1666199351
transform -1 0 43608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _452_
timestamp 1666199351
transform -1 0 44160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _453_
timestamp 1666199351
transform -1 0 45448 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _454_
timestamp 1666199351
transform -1 0 44804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _455_
timestamp 1666199351
transform -1 0 46092 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _456_
timestamp 1666199351
transform -1 0 45448 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _457_
timestamp 1666199351
transform -1 0 45448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _458_
timestamp 1666199351
transform -1 0 46736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _459_
timestamp 1666199351
transform -1 0 46092 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _460_
timestamp 1666199351
transform -1 0 46092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _461_
timestamp 1666199351
transform -1 0 46736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _462_
timestamp 1666199351
transform -1 0 48024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _463_
timestamp 1666199351
transform -1 0 46736 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _464_
timestamp 1666199351
transform -1 0 47380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _465_
timestamp 1666199351
transform -1 0 48024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _466_
timestamp 1666199351
transform -1 0 48024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _470_
timestamp 1666199351
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _471_
timestamp 1666199351
transform 1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _472_
timestamp 1666199351
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _473_
timestamp 1666199351
transform 1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _474_
timestamp 1666199351
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _475_
timestamp 1666199351
transform 1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _476_
timestamp 1666199351
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _477_
timestamp 1666199351
transform 1 0 4968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _478_
timestamp 1666199351
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _479_
timestamp 1666199351
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _480_
timestamp 1666199351
transform 1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _481_
timestamp 1666199351
transform 1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _482_
timestamp 1666199351
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _483_
timestamp 1666199351
transform 1 0 6624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _484_
timestamp 1666199351
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _485_
timestamp 1666199351
transform 1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _486_
timestamp 1666199351
transform 1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _487_
timestamp 1666199351
transform 1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _488_
timestamp 1666199351
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _489_
timestamp 1666199351
transform 1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _490_
timestamp 1666199351
transform 1 0 7728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _491_
timestamp 1666199351
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _492_
timestamp 1666199351
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _493_
timestamp 1666199351
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _494_
timestamp 1666199351
transform 1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _495_
timestamp 1666199351
transform 1 0 9936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _496_
timestamp 1666199351
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _497_
timestamp 1666199351
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _498_
timestamp 1666199351
transform 1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _499_
timestamp 1666199351
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _500_
timestamp 1666199351
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _501_
timestamp 1666199351
transform 1 0 11500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _502_
timestamp 1666199351
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _503_
timestamp 1666199351
transform 1 0 18400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _504_
timestamp 1666199351
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _505_
timestamp 1666199351
transform 1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _506_
timestamp 1666199351
transform -1 0 21528 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _507_
timestamp 1666199351
transform 1 0 19044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _508_
timestamp 1666199351
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _509_
timestamp 1666199351
transform 1 0 18676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _510_
timestamp 1666199351
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _511_
timestamp 1666199351
transform 1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _512_
timestamp 1666199351
transform -1 0 23184 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _513_
timestamp 1666199351
transform 1 0 22540 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _514_
timestamp 1666199351
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _515_
timestamp 1666199351
transform 1 0 20608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _516_
timestamp 1666199351
transform 1 0 23184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _517_
timestamp 1666199351
transform 1 0 23276 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _518_
timestamp 1666199351
transform 1 0 23920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _519_
timestamp 1666199351
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _520_
timestamp 1666199351
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _521_
timestamp 1666199351
transform 1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _522_
timestamp 1666199351
transform 1 0 25024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _523_
timestamp 1666199351
transform -1 0 26220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _524_
timestamp 1666199351
transform -1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _525_
timestamp 1666199351
transform -1 0 29992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _526_
timestamp 1666199351
transform 1 0 26404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _527_
timestamp 1666199351
transform -1 0 28704 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _528_
timestamp 1666199351
transform -1 0 27600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _529_
timestamp 1666199351
transform -1 0 31004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _530_
timestamp 1666199351
transform -1 0 30636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _531_
timestamp 1666199351
transform -1 0 29348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _532_
timestamp 1666199351
transform -1 0 30636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _533_
timestamp 1666199351
transform -1 0 31280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _534_
timestamp 1666199351
transform 1 0 28428 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _535_
timestamp 1666199351
transform 1 0 4508 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _536_
timestamp 1666199351
transform 1 0 5152 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _537_
timestamp 1666199351
transform 1 0 6716 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _538_
timestamp 1666199351
transform 1 0 7544 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _539_
timestamp 1666199351
transform -1 0 9384 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _540_
timestamp 1666199351
transform 1 0 10028 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _541_
timestamp 1666199351
transform 1 0 10948 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _542_
timestamp 1666199351
transform 1 0 12236 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _543_
timestamp 1666199351
transform 1 0 13340 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _544_
timestamp 1666199351
transform 1 0 14444 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _545_
timestamp 1666199351
transform 1 0 14812 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _546_
timestamp 1666199351
transform 1 0 15456 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _547_
timestamp 1666199351
transform 1 0 16100 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _548_
timestamp 1666199351
transform 1 0 16100 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _549_
timestamp 1666199351
transform 1 0 17204 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _550_
timestamp 1666199351
transform 1 0 17388 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _551_
timestamp 1666199351
transform 1 0 18032 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _552_
timestamp 1666199351
transform 1 0 19044 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _553_
timestamp 1666199351
transform 1 0 18676 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _554_
timestamp 1666199351
transform -1 0 26588 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _555_
timestamp 1666199351
transform -1 0 29992 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _556_
timestamp 1666199351
transform -1 0 31004 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _557_
timestamp 1666199351
transform -1 0 35144 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _558_
timestamp 1666199351
transform -1 0 35788 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _559_
timestamp 1666199351
transform 1 0 31004 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _560_
timestamp 1666199351
transform -1 0 38732 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _561_
timestamp 1666199351
transform -1 0 34040 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _562_
timestamp 1666199351
transform -1 0 40296 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _563_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 20332 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _564_
timestamp 1666199351
transform 1 0 20608 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _565_
timestamp 1666199351
transform 1 0 20792 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _566_
timestamp 1666199351
transform 1 0 21252 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _567_
timestamp 1666199351
transform 1 0 21988 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _568_
timestamp 1666199351
transform 1 0 21528 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _569_
timestamp 1666199351
transform 1 0 22540 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _570_
timestamp 1666199351
transform 1 0 22632 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _571_
timestamp 1666199351
transform 1 0 22724 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _572_
timestamp 1666199351
transform 1 0 22908 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _573_
timestamp 1666199351
transform 1 0 23184 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _574_
timestamp 1666199351
transform 1 0 24564 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _575_
timestamp 1666199351
transform 1 0 23920 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _576_
timestamp 1666199351
transform 1 0 24104 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _577_
timestamp 1666199351
transform 1 0 24564 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _578_
timestamp 1666199351
transform 1 0 24564 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _579_
timestamp 1666199351
transform 1 0 25116 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _580_
timestamp 1666199351
transform 1 0 25208 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _581_
timestamp 1666199351
transform 1 0 25300 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _582_
timestamp 1666199351
transform 1 0 25668 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _583_
timestamp 1666199351
transform 1 0 25852 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _584_
timestamp 1666199351
transform -1 0 27968 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _585_
timestamp 1666199351
transform -1 0 27508 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _586_
timestamp 1666199351
transform 1 0 27140 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _587_
timestamp 1666199351
transform -1 0 28060 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _588_
timestamp 1666199351
transform 1 0 27324 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _589_
timestamp 1666199351
transform -1 0 28704 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _590_
timestamp 1666199351
transform -1 0 29164 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _591_
timestamp 1666199351
transform -1 0 29256 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _592_
timestamp 1666199351
transform -1 0 29348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _593_
timestamp 1666199351
transform -1 0 30360 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _594_
timestamp 1666199351
transform 1 0 29072 0 -1 43520
box -38 -48 866 592
<< labels >>
flabel metal2 s 3974 49200 4030 50000 0 FreeSans 224 90 0 0 io_active
port 0 nsew signal input
flabel metal2 s 4342 49200 4398 50000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 15382 49200 15438 50000 0 FreeSans 224 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s 16486 49200 16542 50000 0 FreeSans 224 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal2 s 17590 49200 17646 50000 0 FreeSans 224 90 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 18694 49200 18750 50000 0 FreeSans 224 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 19798 49200 19854 50000 0 FreeSans 224 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal2 s 20902 49200 20958 50000 0 FreeSans 224 90 0 0 io_in[15]
port 7 nsew signal input
flabel metal2 s 22006 49200 22062 50000 0 FreeSans 224 90 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 23110 49200 23166 50000 0 FreeSans 224 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 24214 49200 24270 50000 0 FreeSans 224 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 25318 49200 25374 50000 0 FreeSans 224 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal2 s 5446 49200 5502 50000 0 FreeSans 224 90 0 0 io_in[1]
port 12 nsew signal input
flabel metal2 s 26422 49200 26478 50000 0 FreeSans 224 90 0 0 io_in[20]
port 13 nsew signal input
flabel metal2 s 27526 49200 27582 50000 0 FreeSans 224 90 0 0 io_in[21]
port 14 nsew signal input
flabel metal2 s 28630 49200 28686 50000 0 FreeSans 224 90 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 29734 49200 29790 50000 0 FreeSans 224 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 30838 49200 30894 50000 0 FreeSans 224 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 31942 49200 31998 50000 0 FreeSans 224 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 33046 49200 33102 50000 0 FreeSans 224 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal2 s 34150 49200 34206 50000 0 FreeSans 224 90 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 35254 49200 35310 50000 0 FreeSans 224 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 36358 49200 36414 50000 0 FreeSans 224 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 6550 49200 6606 50000 0 FreeSans 224 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal2 s 37462 49200 37518 50000 0 FreeSans 224 90 0 0 io_in[30]
port 24 nsew signal input
flabel metal2 s 38566 49200 38622 50000 0 FreeSans 224 90 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 39670 49200 39726 50000 0 FreeSans 224 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal2 s 40774 49200 40830 50000 0 FreeSans 224 90 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 41878 49200 41934 50000 0 FreeSans 224 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 42982 49200 43038 50000 0 FreeSans 224 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal2 s 44086 49200 44142 50000 0 FreeSans 224 90 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 45190 49200 45246 50000 0 FreeSans 224 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 7654 49200 7710 50000 0 FreeSans 224 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal2 s 8758 49200 8814 50000 0 FreeSans 224 90 0 0 io_in[4]
port 33 nsew signal input
flabel metal2 s 9862 49200 9918 50000 0 FreeSans 224 90 0 0 io_in[5]
port 34 nsew signal input
flabel metal2 s 10966 49200 11022 50000 0 FreeSans 224 90 0 0 io_in[6]
port 35 nsew signal input
flabel metal2 s 12070 49200 12126 50000 0 FreeSans 224 90 0 0 io_in[7]
port 36 nsew signal input
flabel metal2 s 13174 49200 13230 50000 0 FreeSans 224 90 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 14278 49200 14334 50000 0 FreeSans 224 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 4710 49200 4766 50000 0 FreeSans 224 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal2 s 15750 49200 15806 50000 0 FreeSans 224 90 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal2 s 16854 49200 16910 50000 0 FreeSans 224 90 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal2 s 17958 49200 18014 50000 0 FreeSans 224 90 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal2 s 19062 49200 19118 50000 0 FreeSans 224 90 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal2 s 20166 49200 20222 50000 0 FreeSans 224 90 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 21270 49200 21326 50000 0 FreeSans 224 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal2 s 22374 49200 22430 50000 0 FreeSans 224 90 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 23478 49200 23534 50000 0 FreeSans 224 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 24582 49200 24638 50000 0 FreeSans 224 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 25686 49200 25742 50000 0 FreeSans 224 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal2 s 5814 49200 5870 50000 0 FreeSans 224 90 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal2 s 26790 49200 26846 50000 0 FreeSans 224 90 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal2 s 27894 49200 27950 50000 0 FreeSans 224 90 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 28998 49200 29054 50000 0 FreeSans 224 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 30102 49200 30158 50000 0 FreeSans 224 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 31206 49200 31262 50000 0 FreeSans 224 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal2 s 32310 49200 32366 50000 0 FreeSans 224 90 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal2 s 33414 49200 33470 50000 0 FreeSans 224 90 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 34518 49200 34574 50000 0 FreeSans 224 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal2 s 35622 49200 35678 50000 0 FreeSans 224 90 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal2 s 36726 49200 36782 50000 0 FreeSans 224 90 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 6918 49200 6974 50000 0 FreeSans 224 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal2 s 37830 49200 37886 50000 0 FreeSans 224 90 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal2 s 38934 49200 38990 50000 0 FreeSans 224 90 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal2 s 40038 49200 40094 50000 0 FreeSans 224 90 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal2 s 41142 49200 41198 50000 0 FreeSans 224 90 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal2 s 42246 49200 42302 50000 0 FreeSans 224 90 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal2 s 43350 49200 43406 50000 0 FreeSans 224 90 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal2 s 44454 49200 44510 50000 0 FreeSans 224 90 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal2 s 45558 49200 45614 50000 0 FreeSans 224 90 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 8022 49200 8078 50000 0 FreeSans 224 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal2 s 9126 49200 9182 50000 0 FreeSans 224 90 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal2 s 10230 49200 10286 50000 0 FreeSans 224 90 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal2 s 11334 49200 11390 50000 0 FreeSans 224 90 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 12438 49200 12494 50000 0 FreeSans 224 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 13542 49200 13598 50000 0 FreeSans 224 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 14646 49200 14702 50000 0 FreeSans 224 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal2 s 5078 49200 5134 50000 0 FreeSans 224 90 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal2 s 16118 49200 16174 50000 0 FreeSans 224 90 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal2 s 17222 49200 17278 50000 0 FreeSans 224 90 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal2 s 18326 49200 18382 50000 0 FreeSans 224 90 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal2 s 19430 49200 19486 50000 0 FreeSans 224 90 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal2 s 20534 49200 20590 50000 0 FreeSans 224 90 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal2 s 21638 49200 21694 50000 0 FreeSans 224 90 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal2 s 22742 49200 22798 50000 0 FreeSans 224 90 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 23846 49200 23902 50000 0 FreeSans 224 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal2 s 24950 49200 25006 50000 0 FreeSans 224 90 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal2 s 26054 49200 26110 50000 0 FreeSans 224 90 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 6182 49200 6238 50000 0 FreeSans 224 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 27158 49200 27214 50000 0 FreeSans 224 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal2 s 28262 49200 28318 50000 0 FreeSans 224 90 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 29366 49200 29422 50000 0 FreeSans 224 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal2 s 30470 49200 30526 50000 0 FreeSans 224 90 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 31574 49200 31630 50000 0 FreeSans 224 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 32678 49200 32734 50000 0 FreeSans 224 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal2 s 33782 49200 33838 50000 0 FreeSans 224 90 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 34886 49200 34942 50000 0 FreeSans 224 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 35990 49200 36046 50000 0 FreeSans 224 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal2 s 37094 49200 37150 50000 0 FreeSans 224 90 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 7286 49200 7342 50000 0 FreeSans 224 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal2 s 38198 49200 38254 50000 0 FreeSans 224 90 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal2 s 39302 49200 39358 50000 0 FreeSans 224 90 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal2 s 40406 49200 40462 50000 0 FreeSans 224 90 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal2 s 41510 49200 41566 50000 0 FreeSans 224 90 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal2 s 42614 49200 42670 50000 0 FreeSans 224 90 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal2 s 43718 49200 43774 50000 0 FreeSans 224 90 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 44822 49200 44878 50000 0 FreeSans 224 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal2 s 45926 49200 45982 50000 0 FreeSans 224 90 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal2 s 8390 49200 8446 50000 0 FreeSans 224 90 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal2 s 9494 49200 9550 50000 0 FreeSans 224 90 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 10598 49200 10654 50000 0 FreeSans 224 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 11702 49200 11758 50000 0 FreeSans 224 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal2 s 12806 49200 12862 50000 0 FreeSans 224 90 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 13910 49200 13966 50000 0 FreeSans 224 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal2 s 15014 49200 15070 50000 0 FreeSans 224 90 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 115 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 116 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 117 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 118 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 119 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 120 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 121 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 122 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 123 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 124 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 125 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 126 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 127 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 128 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 129 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 130 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 131 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 132 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 133 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 134 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 135 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 136 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 137 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 138 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 139 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 140 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 141 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 142 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 143 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 144 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 145 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 146 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 147 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 148 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 149 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 150 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 151 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 152 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 153 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 154 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 155 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 156 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 157 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 158 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 159 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 160 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 161 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 162 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 163 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 164 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 165 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 166 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 167 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 168 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 169 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 170 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 171 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 172 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 173 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 174 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 175 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 176 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 177 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 178 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 179 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 180 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 181 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 182 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 183 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 184 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 185 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 186 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 187 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 188 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 189 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 190 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 191 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 192 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 193 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 194 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 195 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 196 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 197 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 198 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 199 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 200 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 201 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 202 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 203 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 204 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 205 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 206 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 207 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 208 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 209 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 210 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 211 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 212 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 213 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 214 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 215 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 216 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 217 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 218 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 219 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 220 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 221 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 222 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 223 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 224 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 225 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 226 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 227 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 228 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 229 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 230 nsew signal input
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 231 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 232 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 233 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 234 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 235 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 236 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 237 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 238 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 239 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 240 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 241 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 242 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 243 nsew signal tristate
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 244 nsew signal tristate
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 245 nsew signal tristate
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 246 nsew signal tristate
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 247 nsew signal tristate
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 248 nsew signal tristate
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 249 nsew signal tristate
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 250 nsew signal tristate
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 251 nsew signal tristate
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 252 nsew signal tristate
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 253 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 254 nsew signal tristate
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 255 nsew signal tristate
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 256 nsew signal tristate
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 257 nsew signal tristate
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 258 nsew signal tristate
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 259 nsew signal tristate
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 260 nsew signal tristate
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 261 nsew signal tristate
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 262 nsew signal tristate
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 263 nsew signal tristate
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 264 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 265 nsew signal tristate
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 266 nsew signal tristate
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 267 nsew signal tristate
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 268 nsew signal tristate
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 269 nsew signal tristate
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 270 nsew signal tristate
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 271 nsew signal tristate
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 272 nsew signal tristate
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 273 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 274 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 275 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 276 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 277 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 278 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 279 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 280 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 281 nsew signal tristate
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 282 nsew signal tristate
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 283 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 284 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 285 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 286 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 287 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 288 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 289 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 290 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 291 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 292 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 293 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 294 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 295 nsew signal tristate
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 296 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 297 nsew signal tristate
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 298 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 299 nsew signal tristate
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 300 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 301 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 302 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 303 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 304 nsew signal tristate
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 305 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 306 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 307 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 308 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 309 nsew signal tristate
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 310 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 311 nsew signal tristate
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 312 nsew signal tristate
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 313 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 314 nsew signal tristate
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 315 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 316 nsew signal tristate
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 317 nsew signal tristate
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 318 nsew signal tristate
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 319 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 320 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 321 nsew signal tristate
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 322 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 323 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 324 nsew signal tristate
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 325 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 326 nsew signal tristate
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 327 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 328 nsew signal tristate
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 329 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 330 nsew signal tristate
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 331 nsew signal tristate
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 332 nsew signal tristate
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 333 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 334 nsew signal tristate
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 335 nsew signal tristate
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 336 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 337 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 338 nsew signal tristate
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 339 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 340 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 341 nsew signal tristate
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 342 nsew signal tristate
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 343 nsew signal tristate
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 344 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 345 nsew signal tristate
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 346 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 347 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 348 nsew signal tristate
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 349 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 350 nsew signal tristate
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 351 nsew signal tristate
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 352 nsew signal tristate
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 353 nsew signal tristate
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 354 nsew signal tristate
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 355 nsew signal tristate
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 356 nsew signal tristate
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 357 nsew signal tristate
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 358 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 359 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 360 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 361 nsew signal tristate
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 362 nsew signal tristate
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 363 nsew signal tristate
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 364 nsew signal tristate
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 365 nsew signal tristate
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 366 nsew signal tristate
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 367 nsew signal tristate
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 368 nsew signal tristate
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 369 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 370 nsew signal tristate
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 371 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 372 nsew signal input
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 373 nsew signal input
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 374 nsew signal input
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 375 nsew signal input
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 376 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 377 nsew signal input
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 378 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 379 nsew signal input
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 380 nsew signal input
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 381 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 382 nsew signal input
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 383 nsew signal input
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 384 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 385 nsew signal input
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 386 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 387 nsew signal input
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 388 nsew signal input
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 389 nsew signal input
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 390 nsew signal input
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 391 nsew signal input
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 392 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 393 nsew signal input
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 394 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 395 nsew signal input
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 396 nsew signal input
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 397 nsew signal input
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 398 nsew signal input
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 399 nsew signal input
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 400 nsew signal input
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 401 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 402 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 403 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 404 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 405 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 406 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 407 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 408 nsew signal input
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 409 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 410 nsew signal input
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 411 nsew signal input
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 412 nsew signal input
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 413 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 414 nsew signal input
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 415 nsew signal input
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 416 nsew signal input
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 417 nsew signal input
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 418 nsew signal input
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 419 nsew signal input
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 420 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 421 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 422 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 423 nsew signal input
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 424 nsew signal input
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 425 nsew signal input
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 426 nsew signal input
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 427 nsew signal input
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 428 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 429 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 430 nsew signal input
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 431 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 432 nsew signal input
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 433 nsew signal input
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 434 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 435 nsew signal input
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 436 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 437 nsew signal input
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 438 nsew signal input
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 439 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 440 nsew signal input
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 441 nsew signal input
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 442 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 443 nsew signal input
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 444 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 445 nsew signal input
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 446 nsew signal input
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 447 nsew signal input
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 448 nsew signal input
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 449 nsew signal input
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 450 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 451 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 452 nsew signal input
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 453 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 454 nsew signal input
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 455 nsew signal input
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 456 nsew signal input
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 457 nsew signal input
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 458 nsew signal input
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 459 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 460 nsew signal input
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 461 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 462 nsew signal input
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 463 nsew signal input
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 464 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 465 nsew signal input
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 466 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 467 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 468 nsew signal input
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 469 nsew signal input
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 470 nsew signal input
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 471 nsew signal input
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 472 nsew signal input
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 473 nsew signal input
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 474 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 475 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 476 nsew signal input
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 477 nsew signal input
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 478 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 479 nsew signal input
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 480 nsew signal input
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 481 nsew signal input
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 482 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 483 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 484 nsew signal input
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 485 nsew signal input
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 486 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 487 nsew signal input
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 488 nsew signal input
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 489 nsew signal input
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 490 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 491 nsew signal input
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 492 nsew signal input
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 493 nsew signal input
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 494 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 495 nsew signal input
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 496 nsew signal input
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 497 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 498 nsew signal input
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 34928 2128 35248 47376 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 19568 2128 19888 47376 0 FreeSans 1920 90 0 0 vssd1
port 500 nsew ground bidirectional
flabel metal2 s 2410 0 2466 800 0 FreeSans 224 90 0 0 wb_clk_i
port 501 nsew signal input
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 wb_rst_i
port 502 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 503 nsew signal tristate
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 504 nsew signal input
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 505 nsew signal input
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 506 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 507 nsew signal input
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 508 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 509 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 510 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 511 nsew signal input
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 512 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 513 nsew signal input
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 514 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 515 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 516 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 517 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 518 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 519 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 520 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 521 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 522 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 523 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 524 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 525 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 526 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 527 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 528 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 529 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 530 nsew signal input
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 531 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 532 nsew signal input
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 533 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 534 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 535 nsew signal input
flabel metal2 s 2686 0 2742 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 536 nsew signal input
flabel metal2 s 3054 0 3110 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 537 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 538 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 539 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 540 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 541 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 542 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 543 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 544 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 545 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 546 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 547 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 548 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 549 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 550 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 551 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 552 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 553 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 554 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 555 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 556 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 557 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 558 nsew signal input
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 559 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 560 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 561 nsew signal input
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 562 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 563 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 564 nsew signal input
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 565 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 566 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 567 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 568 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 569 nsew signal tristate
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 570 nsew signal tristate
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 571 nsew signal tristate
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 572 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 573 nsew signal tristate
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 574 nsew signal tristate
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 575 nsew signal tristate
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 576 nsew signal tristate
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 577 nsew signal tristate
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 578 nsew signal tristate
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 579 nsew signal tristate
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 580 nsew signal tristate
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 581 nsew signal tristate
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 582 nsew signal tristate
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 583 nsew signal tristate
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 584 nsew signal tristate
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 585 nsew signal tristate
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 586 nsew signal tristate
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 587 nsew signal tristate
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 588 nsew signal tristate
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 589 nsew signal tristate
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 590 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 591 nsew signal tristate
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 592 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 593 nsew signal tristate
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 594 nsew signal tristate
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 595 nsew signal tristate
flabel metal2 s 4894 0 4950 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 596 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 597 nsew signal tristate
flabel metal2 s 5446 0 5502 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 598 nsew signal tristate
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 599 nsew signal tristate
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 600 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 601 nsew signal input
flabel metal2 s 3606 0 3662 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 602 nsew signal input
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 603 nsew signal input
flabel metal2 s 4342 0 4398 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 604 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 605 nsew signal input
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 wbs_we_i
port 606 nsew signal input
rlabel metal1 24978 47328 24978 47328 0 vccd1
rlabel metal1 24978 46784 24978 46784 0 vssd1
rlabel metal2 18722 3264 18722 3264 0 _000_
rlabel metal1 28106 45968 28106 45968 0 _001_
rlabel metal1 28704 46002 28704 46002 0 _002_
rlabel metal2 30590 45764 30590 45764 0 _003_
rlabel metal1 29762 44982 29762 44982 0 _004_
rlabel metal2 22402 45390 22402 45390 0 _005_
rlabel metal2 29670 45084 29670 45084 0 _006_
rlabel metal1 25675 43758 25675 43758 0 _007_
rlabel viali 24150 44369 24150 44369 0 _008_
rlabel metal1 29118 45560 29118 45560 0 _009_
rlabel metal2 27830 45050 27830 45050 0 _010_
rlabel metal2 28658 45050 28658 45050 0 _011_
rlabel metal2 27278 44608 27278 44608 0 _012_
rlabel metal1 26864 44438 26864 44438 0 _013_
rlabel metal1 27968 43690 27968 43690 0 _014_
rlabel metal1 25484 44302 25484 44302 0 _015_
rlabel metal1 23966 44812 23966 44812 0 _016_
rlabel metal1 23690 44302 23690 44302 0 _017_
rlabel metal1 24081 45458 24081 45458 0 _018_
rlabel metal1 26884 45526 26884 45526 0 _019_
rlabel metal1 22586 45492 22586 45492 0 _020_
rlabel metal2 23690 46716 23690 46716 0 _021_
rlabel metal1 22402 45356 22402 45356 0 _022_
rlabel metal2 21390 46274 21390 46274 0 _023_
rlabel metal1 39330 45254 39330 45254 0 _024_
rlabel metal1 38272 46138 38272 46138 0 _025_
rlabel metal2 37674 46104 37674 46104 0 _026_
rlabel metal2 32706 44574 32706 44574 0 _027_
rlabel metal2 32154 44370 32154 44370 0 _028_
rlabel metal2 38686 44608 38686 44608 0 _029_
rlabel metal2 33074 44540 33074 44540 0 _030_
rlabel metal1 32154 44880 32154 44880 0 _031_
rlabel metal2 37214 45084 37214 45084 0 _032_
rlabel metal2 37674 44574 37674 44574 0 _033_
rlabel metal1 38318 45050 38318 45050 0 _034_
rlabel metal1 37306 43758 37306 43758 0 _035_
rlabel metal1 35880 44302 35880 44302 0 _036_
rlabel metal2 36846 43690 36846 43690 0 _037_
rlabel metal2 34546 44166 34546 44166 0 _038_
rlabel metal2 32338 44897 32338 44897 0 _039_
rlabel metal1 32844 44846 32844 44846 0 _040_
rlabel metal2 31510 46444 31510 46444 0 _041_
rlabel metal1 32706 46988 32706 46988 0 _042_
rlabel metal2 29486 46308 29486 46308 0 _043_
rlabel metal1 40250 45356 40250 45356 0 _044_
rlabel metal2 29302 46818 29302 46818 0 _045_
rlabel metal2 28290 46886 28290 46886 0 _046_
rlabel metal2 26634 46750 26634 46750 0 _047_
rlabel metal1 25944 46682 25944 46682 0 _048_
rlabel metal1 25576 46614 25576 46614 0 _049_
rlabel metal1 21298 47056 21298 47056 0 _050_
rlabel metal2 41722 46189 41722 46189 0 _051_
rlabel metal2 35374 46172 35374 46172 0 _052_
rlabel metal1 35006 46138 35006 46138 0 _053_
rlabel metal1 20010 46886 20010 46886 0 _054_
rlabel metal1 20838 45968 20838 45968 0 _055_
rlabel metal2 18998 44540 18998 44540 0 _056_
rlabel metal1 17526 46546 17526 46546 0 _057_
rlabel metal2 27646 43588 27646 43588 0 _058_
rlabel metal1 26772 43826 26772 43826 0 _059_
rlabel metal1 27462 46580 27462 46580 0 _060_
rlabel metal1 27738 46138 27738 46138 0 _061_
rlabel metal1 26910 46002 26910 46002 0 _062_
rlabel metal1 20746 45458 20746 45458 0 _063_
rlabel metal2 36570 44166 36570 44166 0 _064_
rlabel metal1 37168 44506 37168 44506 0 _065_
rlabel metal2 41262 47260 41262 47260 0 _066_
rlabel metal2 38502 46393 38502 46393 0 _067_
rlabel metal1 37306 45934 37306 45934 0 _068_
rlabel metal1 17802 45526 17802 45526 0 _069_
rlabel metal1 19136 44506 19136 44506 0 _070_
rlabel metal1 18676 45526 18676 45526 0 _071_
rlabel metal1 26496 44914 26496 44914 0 _072_
rlabel metal1 26128 43350 26128 43350 0 _073_
rlabel metal2 25714 43520 25714 43520 0 _074_
rlabel metal1 25484 43282 25484 43282 0 _075_
rlabel metal2 25530 44642 25530 44642 0 _076_
rlabel metal1 21160 45934 21160 45934 0 _077_
rlabel metal1 34408 45458 34408 45458 0 _078_
rlabel metal1 34224 43962 34224 43962 0 _079_
rlabel metal1 34040 44438 34040 44438 0 _080_
rlabel metal1 34086 44370 34086 44370 0 _081_
rlabel metal2 33626 45220 33626 45220 0 _082_
rlabel metal2 21482 45730 21482 45730 0 _083_
rlabel metal1 20378 44506 20378 44506 0 _084_
rlabel metal1 19274 45254 19274 45254 0 _085_
rlabel metal1 23644 43758 23644 43758 0 _086_
rlabel metal2 22402 43962 22402 43962 0 _087_
rlabel metal1 22540 46546 22540 46546 0 _088_
rlabel metal1 23092 46002 23092 46002 0 _089_
rlabel via1 23321 46546 23321 46546 0 _090_
rlabel metal1 21758 45968 21758 45968 0 _091_
rlabel metal1 23276 45934 23276 45934 0 _092_
rlabel metal2 32430 44812 32430 44812 0 _093_
rlabel metal2 30958 44132 30958 44132 0 _094_
rlabel metal2 31050 46138 31050 46138 0 _095_
rlabel metal1 33120 46546 33120 46546 0 _096_
rlabel metal1 30498 46580 30498 46580 0 _097_
rlabel metal2 23690 46087 23690 46087 0 _098_
rlabel metal1 22494 5236 22494 5236 0 _099_
rlabel metal1 24380 4590 24380 4590 0 _100_
rlabel metal1 31004 2414 31004 2414 0 _101_
rlabel via1 27922 4590 27922 4590 0 _102_
rlabel metal2 25714 5134 25714 5134 0 _103_
rlabel metal2 24426 5984 24426 5984 0 _104_
rlabel metal2 22310 5678 22310 5678 0 _105_
rlabel metal1 20378 4182 20378 4182 0 _106_
rlabel metal1 19826 3094 19826 3094 0 _107_
rlabel metal1 20562 4522 20562 4522 0 _108_
rlabel metal1 21114 5610 21114 5610 0 _109_
rlabel metal1 20286 3366 20286 3366 0 _110_
rlabel metal2 18170 3434 18170 3434 0 _111_
rlabel metal1 20516 2550 20516 2550 0 _112_
rlabel metal1 22448 2346 22448 2346 0 _113_
rlabel metal1 22954 4488 22954 4488 0 _114_
rlabel metal1 23138 5304 23138 5304 0 _115_
rlabel metal2 23414 5848 23414 5848 0 _116_
rlabel metal1 24794 3400 24794 3400 0 _117_
rlabel metal2 24150 3230 24150 3230 0 _118_
rlabel metal1 24150 3706 24150 3706 0 _119_
rlabel metal2 24794 6120 24794 6120 0 _120_
rlabel metal2 24518 5848 24518 5848 0 _121_
rlabel metal1 24426 2482 24426 2482 0 _122_
rlabel metal1 25438 2312 25438 2312 0 _123_
rlabel metal1 25714 3706 25714 3706 0 _124_
rlabel metal2 25806 5032 25806 5032 0 _125_
rlabel metal2 26726 6120 26726 6120 0 _126_
rlabel metal1 27140 2550 27140 2550 0 _127_
rlabel metal1 28474 2618 28474 2618 0 _128_
rlabel metal1 27324 2618 27324 2618 0 _129_
rlabel metal2 27830 5678 27830 5678 0 _130_
rlabel metal2 27554 5202 27554 5202 0 _131_
rlabel metal1 28474 3400 28474 3400 0 _132_
rlabel metal1 30406 2618 30406 2618 0 _133_
rlabel metal1 29762 4522 29762 4522 0 _134_
rlabel metal1 29486 4182 29486 4182 0 _135_
rlabel metal1 30820 3094 30820 3094 0 _136_
rlabel metal2 22770 44982 22770 44982 0 _137_
rlabel metal1 19550 4046 19550 4046 0 _138_
rlabel metal1 19688 2958 19688 2958 0 _139_
rlabel metal2 20930 5372 20930 5372 0 _140_
rlabel metal2 21390 5916 21390 5916 0 _141_
rlabel metal1 22126 4012 22126 4012 0 _142_
rlabel metal1 19090 2550 19090 2550 0 _143_
rlabel metal1 22678 2924 22678 2924 0 _144_
rlabel metal1 20838 2482 20838 2482 0 _145_
rlabel metal1 20332 3910 20332 3910 0 _146_
rlabel metal2 23046 6018 23046 6018 0 _147_
rlabel metal1 23046 5746 23046 5746 0 _148_
rlabel metal1 23966 3570 23966 3570 0 _149_
rlabel metal1 21482 2618 21482 2618 0 _150_
rlabel metal2 23414 3876 23414 3876 0 _151_
rlabel metal2 24702 5916 24702 5916 0 _152_
rlabel metal1 24426 6222 24426 6222 0 _153_
rlabel metal1 23368 2618 23368 2618 0 _154_
rlabel metal1 25346 2516 25346 2516 0 _155_
rlabel metal1 24104 3978 24104 3978 0 _156_
rlabel metal1 25530 5134 25530 5134 0 _157_
rlabel metal2 25990 6052 25990 6052 0 _158_
rlabel metal2 27830 2788 27830 2788 0 _159_
rlabel metal1 28980 2550 28980 2550 0 _160_
rlabel metal2 26634 3536 26634 3536 0 _161_
rlabel metal1 28198 5134 28198 5134 0 _162_
rlabel metal2 27462 5916 27462 5916 0 _163_
rlabel metal2 30774 3230 30774 3230 0 _164_
rlabel metal1 29532 3094 29532 3094 0 _165_
rlabel metal2 29118 4828 29118 4828 0 _166_
rlabel metal1 29808 4046 29808 4046 0 _167_
rlabel metal2 31050 2788 31050 2788 0 _168_
rlabel metal1 28934 43214 28934 43214 0 _169_
rlabel metal2 28382 44336 28382 44336 0 _595_
rlabel metal2 24610 45900 24610 45900 0 _596_
rlabel metal1 23920 43282 23920 43282 0 _597_
rlabel metal1 37260 43282 37260 43282 0 _598_
rlabel metal1 32936 43962 32936 43962 0 _599_
rlabel metal1 33120 43282 33120 43282 0 _600_
rlabel metal2 18722 45356 18722 45356 0 _601_
rlabel metal2 17986 46750 17986 46750 0 _602_
rlabel metal1 19964 44370 19964 44370 0 _603_
rlabel metal1 19550 45390 19550 45390 0 _604_
rlabel metal2 20838 44574 20838 44574 0 _605_
rlabel metal1 19642 45492 19642 45492 0 _606_
rlabel metal2 22494 44574 22494 44574 0 _607_
rlabel metal2 31050 44506 31050 44506 0 _608_
rlabel metal1 21160 44370 21160 44370 0 active
rlabel metal2 24334 47957 24334 47957 0 io_in[18]
rlabel metal1 27646 45934 27646 45934 0 io_in[19]
rlabel metal1 26128 46138 26128 46138 0 io_in[20]
rlabel metal2 16974 47430 16974 47430 0 io_in[21]
rlabel metal2 28658 47984 28658 47984 0 io_in[22]
rlabel via1 29193 45458 29193 45458 0 io_in[23]
rlabel metal1 30590 45458 30590 45458 0 io_in[24]
rlabel metal2 31970 47066 31970 47066 0 io_in[25]
rlabel metal1 34546 46580 34546 46580 0 io_in[26]
rlabel metal1 38916 46478 38916 46478 0 io_in[27]
rlabel metal1 35328 45526 35328 45526 0 io_in[28]
rlabel metal2 41998 47294 41998 47294 0 io_in[29]
rlabel metal1 37720 45390 37720 45390 0 io_in[30]
rlabel metal1 38455 45458 38455 45458 0 io_in[31]
rlabel viali 37858 46548 37858 46548 0 io_in[32]
rlabel metal1 40158 45934 40158 45934 0 io_in[33]
rlabel metal2 41906 48222 41906 48222 0 io_in[34]
rlabel metal2 43010 47593 43010 47593 0 io_in[35]
rlabel metal1 44344 47226 44344 47226 0 io_in[36]
rlabel metal1 42550 45050 42550 45050 0 io_in[37]
rlabel metal2 4738 48256 4738 48256 0 io_oeb[0]
rlabel metal1 15410 47226 15410 47226 0 io_oeb[10]
rlabel metal1 16284 47158 16284 47158 0 io_oeb[11]
rlabel metal1 17204 46478 17204 46478 0 io_oeb[12]
rlabel metal1 17710 47226 17710 47226 0 io_oeb[13]
rlabel metal2 20049 49300 20049 49300 0 io_oeb[14]
rlabel metal2 17618 47328 17618 47328 0 io_oeb[15]
rlabel metal1 20194 47124 20194 47124 0 io_oeb[16]
rlabel metal1 19435 46478 19435 46478 0 io_oeb[17]
rlabel metal2 18906 47396 18906 47396 0 io_oeb[18]
rlabel metal1 26312 44370 26312 44370 0 io_oeb[19]
rlabel metal1 5612 47226 5612 47226 0 io_oeb[1]
rlabel metal1 28290 47226 28290 47226 0 io_oeb[20]
rlabel metal1 29348 46138 29348 46138 0 io_oeb[21]
rlabel metal1 34822 47022 34822 47022 0 io_oeb[22]
rlabel metal2 34546 46886 34546 46886 0 io_oeb[23]
rlabel metal2 31234 46284 31234 46284 0 io_oeb[24]
rlabel metal1 38502 46988 38502 46988 0 io_oeb[25]
rlabel metal1 33626 43282 33626 43282 0 io_oeb[26]
rlabel metal1 40112 47022 40112 47022 0 io_oeb[27]
rlabel metal2 40710 46937 40710 46937 0 io_oeb[28]
rlabel metal1 40020 46002 40020 46002 0 io_oeb[29]
rlabel metal2 6946 47916 6946 47916 0 io_oeb[2]
rlabel metal2 39238 45322 39238 45322 0 io_oeb[30]
rlabel metal1 40158 46138 40158 46138 0 io_oeb[31]
rlabel metal2 43286 46852 43286 46852 0 io_oeb[32]
rlabel metal2 41170 47848 41170 47848 0 io_oeb[33]
rlabel metal1 42458 46138 42458 46138 0 io_oeb[34]
rlabel metal1 43654 47226 43654 47226 0 io_oeb[35]
rlabel metal2 44574 47923 44574 47923 0 io_oeb[36]
rlabel metal2 45862 48263 45862 48263 0 io_oeb[37]
rlabel metal2 7774 48263 7774 48263 0 io_oeb[3]
rlabel metal2 9154 48256 9154 48256 0 io_oeb[4]
rlabel metal2 10258 48256 10258 48256 0 io_oeb[5]
rlabel metal2 11178 48263 11178 48263 0 io_oeb[6]
rlabel metal2 12466 48256 12466 48256 0 io_oeb[7]
rlabel metal2 13570 48256 13570 48256 0 io_oeb[8]
rlabel metal2 14674 47916 14674 47916 0 io_oeb[9]
rlabel metal2 5106 48426 5106 48426 0 io_out[0]
rlabel metal1 18676 47022 18676 47022 0 io_out[10]
rlabel metal1 17710 45594 17710 45594 0 io_out[11]
rlabel metal2 18354 47950 18354 47950 0 io_out[12]
rlabel metal2 23966 46852 23966 46852 0 io_out[13]
rlabel metal2 20417 49300 20417 49300 0 io_out[14]
rlabel metal2 19734 45968 19734 45968 0 io_out[15]
rlabel metal2 22823 49300 22823 49300 0 io_out[16]
rlabel metal2 23874 47950 23874 47950 0 io_out[17]
rlabel metal1 25576 43962 25576 43962 0 io_out[18]
rlabel metal1 27830 46988 27830 46988 0 io_out[19]
rlabel metal2 6026 48263 6026 48263 0 io_out[1]
rlabel metal1 31188 47022 31188 47022 0 io_out[20]
rlabel metal1 32522 45866 32522 45866 0 io_out[21]
rlabel metal1 29578 43962 29578 43962 0 io_out[22]
rlabel metal2 30498 48222 30498 48222 0 io_out[23]
rlabel metal2 36570 46886 36570 46886 0 io_out[24]
rlabel metal1 35926 47226 35926 47226 0 io_out[25]
rlabel metal1 34178 43282 34178 43282 0 io_out[26]
rlabel metal1 38732 46342 38732 46342 0 io_out[27]
rlabel metal1 39698 46478 39698 46478 0 io_out[28]
rlabel metal1 40986 46580 40986 46580 0 io_out[29]
rlabel metal2 7130 48263 7130 48263 0 io_out[2]
rlabel metal1 39468 46070 39468 46070 0 io_out[30]
rlabel metal2 39330 48256 39330 48256 0 io_out[31]
rlabel metal1 40664 45322 40664 45322 0 io_out[32]
rlabel metal1 41768 46138 41768 46138 0 io_out[33]
rlabel metal1 42964 46546 42964 46546 0 io_out[34]
rlabel metal2 43930 47923 43930 47923 0 io_out[35]
rlabel metal1 45034 47226 45034 47226 0 io_out[36]
rlabel metal1 46230 47226 46230 47226 0 io_out[37]
rlabel metal2 8418 48256 8418 48256 0 io_out[3]
rlabel metal2 9522 47729 9522 47729 0 io_out[4]
rlabel metal2 9706 45465 9706 45465 0 io_out[5]
rlabel metal2 11730 48358 11730 48358 0 io_out[6]
rlabel metal2 12834 47678 12834 47678 0 io_out[7]
rlabel metal2 13938 47814 13938 47814 0 io_out[8]
rlabel metal2 15042 47848 15042 47848 0 io_out[9]
rlabel metal2 12282 1588 12282 1588 0 la_data_out[0]
rlabel metal2 39882 1588 39882 1588 0 la_data_out[100]
rlabel metal2 40158 1792 40158 1792 0 la_data_out[101]
rlabel metal2 40434 2132 40434 2132 0 la_data_out[102]
rlabel metal2 40710 1860 40710 1860 0 la_data_out[103]
rlabel metal2 40986 2132 40986 2132 0 la_data_out[104]
rlabel metal2 41262 1622 41262 1622 0 la_data_out[105]
rlabel metal2 41538 2132 41538 2132 0 la_data_out[106]
rlabel metal2 41814 1588 41814 1588 0 la_data_out[107]
rlabel metal2 42090 1792 42090 1792 0 la_data_out[108]
rlabel metal2 42366 1656 42366 1656 0 la_data_out[109]
rlabel metal2 15042 2336 15042 2336 0 la_data_out[10]
rlabel metal2 42642 1860 42642 1860 0 la_data_out[110]
rlabel metal2 42918 2132 42918 2132 0 la_data_out[111]
rlabel metal2 43194 2132 43194 2132 0 la_data_out[112]
rlabel metal2 43470 1792 43470 1792 0 la_data_out[113]
rlabel metal2 43746 1622 43746 1622 0 la_data_out[114]
rlabel metal2 44022 1792 44022 1792 0 la_data_out[115]
rlabel metal2 44298 1554 44298 1554 0 la_data_out[116]
rlabel metal2 44574 1860 44574 1860 0 la_data_out[117]
rlabel metal2 44850 2132 44850 2132 0 la_data_out[118]
rlabel metal2 45126 1656 45126 1656 0 la_data_out[119]
rlabel metal1 14858 2958 14858 2958 0 la_data_out[11]
rlabel metal2 45402 1792 45402 1792 0 la_data_out[120]
rlabel metal2 45678 2132 45678 2132 0 la_data_out[121]
rlabel metal2 45954 1792 45954 1792 0 la_data_out[122]
rlabel metal2 46230 1588 46230 1588 0 la_data_out[123]
rlabel metal2 46506 2132 46506 2132 0 la_data_out[124]
rlabel metal2 46782 2132 46782 2132 0 la_data_out[125]
rlabel metal2 47058 1792 47058 1792 0 la_data_out[126]
rlabel metal2 47334 2132 47334 2132 0 la_data_out[127]
rlabel metal2 15594 1588 15594 1588 0 la_data_out[12]
rlabel metal1 15456 3570 15456 3570 0 la_data_out[13]
rlabel metal2 16146 2336 16146 2336 0 la_data_out[14]
rlabel metal1 16054 3502 16054 3502 0 la_data_out[15]
rlabel metal1 15870 2890 15870 2890 0 la_data_out[16]
rlabel metal1 16652 3638 16652 3638 0 la_data_out[17]
rlabel metal2 17250 2336 17250 2336 0 la_data_out[18]
rlabel metal1 16606 2958 16606 2958 0 la_data_out[19]
rlabel metal1 12466 3502 12466 3502 0 la_data_out[1]
rlabel metal2 17802 1622 17802 1622 0 la_data_out[20]
rlabel metal2 18078 2676 18078 2676 0 la_data_out[21]
rlabel metal1 17940 2890 17940 2890 0 la_data_out[22]
rlabel metal2 18630 1299 18630 1299 0 la_data_out[23]
rlabel metal1 18446 3910 18446 3910 0 la_data_out[24]
rlabel metal2 19182 1690 19182 1690 0 la_data_out[25]
rlabel metal2 19458 2880 19458 2880 0 la_data_out[26]
rlabel metal2 19734 1367 19734 1367 0 la_data_out[27]
rlabel metal2 20010 1316 20010 1316 0 la_data_out[28]
rlabel metal1 18952 3570 18952 3570 0 la_data_out[29]
rlabel metal2 12834 1622 12834 1622 0 la_data_out[2]
rlabel metal1 19090 2822 19090 2822 0 la_data_out[30]
rlabel metal2 20838 1520 20838 1520 0 la_data_out[31]
rlabel metal2 21114 2404 21114 2404 0 la_data_out[32]
rlabel metal2 21390 1860 21390 1860 0 la_data_out[33]
rlabel metal1 21620 4522 21620 4522 0 la_data_out[34]
rlabel metal2 21942 3288 21942 3288 0 la_data_out[35]
rlabel metal2 22218 2404 22218 2404 0 la_data_out[36]
rlabel metal2 22494 2098 22494 2098 0 la_data_out[37]
rlabel metal2 22770 1860 22770 1860 0 la_data_out[38]
rlabel metal2 23046 1622 23046 1622 0 la_data_out[39]
rlabel metal1 13064 3502 13064 3502 0 la_data_out[3]
rlabel metal2 23322 2710 23322 2710 0 la_data_out[40]
rlabel metal2 23598 2914 23598 2914 0 la_data_out[41]
rlabel metal2 23874 3288 23874 3288 0 la_data_out[42]
rlabel metal2 24150 1231 24150 1231 0 la_data_out[43]
rlabel metal2 24426 1860 24426 1860 0 la_data_out[44]
rlabel metal2 24702 2370 24702 2370 0 la_data_out[45]
rlabel metal2 24978 3254 24978 3254 0 la_data_out[46]
rlabel metal2 25254 3458 25254 3458 0 la_data_out[47]
rlabel metal2 25530 1860 25530 1860 0 la_data_out[48]
rlabel metal2 25806 1622 25806 1622 0 la_data_out[49]
rlabel metal1 12926 2890 12926 2890 0 la_data_out[4]
rlabel metal2 26082 2404 26082 2404 0 la_data_out[50]
rlabel metal2 26358 2914 26358 2914 0 la_data_out[51]
rlabel metal2 26634 1843 26634 1843 0 la_data_out[52]
rlabel metal2 26910 1860 26910 1860 0 la_data_out[53]
rlabel metal2 27186 2166 27186 2166 0 la_data_out[54]
rlabel metal2 27462 2404 27462 2404 0 la_data_out[55]
rlabel metal2 27738 1571 27738 1571 0 la_data_out[56]
rlabel metal2 28014 3288 28014 3288 0 la_data_out[57]
rlabel metal2 28290 2166 28290 2166 0 la_data_out[58]
rlabel metal2 28566 1860 28566 1860 0 la_data_out[59]
rlabel metal2 13662 2132 13662 2132 0 la_data_out[5]
rlabel metal2 28842 2710 28842 2710 0 la_data_out[60]
rlabel metal2 29118 2404 29118 2404 0 la_data_out[61]
rlabel metal2 29394 1860 29394 1860 0 la_data_out[62]
rlabel metal2 29670 3831 29670 3831 0 la_data_out[63]
rlabel metal2 29946 1656 29946 1656 0 la_data_out[64]
rlabel metal2 30222 2166 30222 2166 0 la_data_out[65]
rlabel metal2 30498 1554 30498 1554 0 la_data_out[66]
rlabel metal2 30774 1792 30774 1792 0 la_data_out[67]
rlabel metal2 31050 1299 31050 1299 0 la_data_out[68]
rlabel metal2 31326 1622 31326 1622 0 la_data_out[69]
rlabel metal1 13524 2822 13524 2822 0 la_data_out[6]
rlabel metal2 31602 1826 31602 1826 0 la_data_out[70]
rlabel metal2 31878 2132 31878 2132 0 la_data_out[71]
rlabel metal2 32154 1860 32154 1860 0 la_data_out[72]
rlabel metal2 32430 2132 32430 2132 0 la_data_out[73]
rlabel metal2 32706 1894 32706 1894 0 la_data_out[74]
rlabel metal2 32982 2200 32982 2200 0 la_data_out[75]
rlabel metal2 33258 1656 33258 1656 0 la_data_out[76]
rlabel metal2 33534 1826 33534 1826 0 la_data_out[77]
rlabel metal2 33810 1588 33810 1588 0 la_data_out[78]
rlabel metal2 34086 1860 34086 1860 0 la_data_out[79]
rlabel metal2 14214 1656 14214 1656 0 la_data_out[7]
rlabel metal2 34362 2132 34362 2132 0 la_data_out[80]
rlabel metal2 34638 1622 34638 1622 0 la_data_out[81]
rlabel metal2 34914 1299 34914 1299 0 la_data_out[82]
rlabel metal2 35190 1095 35190 1095 0 la_data_out[83]
rlabel metal2 35466 1656 35466 1656 0 la_data_out[84]
rlabel metal2 35742 2132 35742 2132 0 la_data_out[85]
rlabel metal2 36018 1792 36018 1792 0 la_data_out[86]
rlabel metal2 36294 2132 36294 2132 0 la_data_out[87]
rlabel metal2 36570 1588 36570 1588 0 la_data_out[88]
rlabel metal2 36846 2200 36846 2200 0 la_data_out[89]
rlabel metal1 14122 2890 14122 2890 0 la_data_out[8]
rlabel metal2 37122 1860 37122 1860 0 la_data_out[90]
rlabel metal2 37398 1622 37398 1622 0 la_data_out[91]
rlabel metal2 37674 2132 37674 2132 0 la_data_out[92]
rlabel metal2 37950 1826 37950 1826 0 la_data_out[93]
rlabel metal2 38226 2132 38226 2132 0 la_data_out[94]
rlabel metal2 38502 1656 38502 1656 0 la_data_out[95]
rlabel metal2 38778 1860 38778 1860 0 la_data_out[96]
rlabel metal2 39054 1792 39054 1792 0 la_data_out[97]
rlabel metal2 39330 1622 39330 1622 0 la_data_out[98]
rlabel metal2 39606 2132 39606 2132 0 la_data_out[99]
rlabel metal2 14766 1622 14766 1622 0 la_data_out[9]
rlabel metal2 2622 1588 2622 1588 0 wbs_ack_o
rlabel metal2 3174 1792 3174 1792 0 wbs_dat_o[0]
rlabel metal2 6302 1826 6302 1826 0 wbs_dat_o[10]
rlabel metal2 6578 1792 6578 1792 0 wbs_dat_o[11]
rlabel metal2 6854 2132 6854 2132 0 wbs_dat_o[12]
rlabel metal2 7130 1656 7130 1656 0 wbs_dat_o[13]
rlabel metal1 6463 2414 6463 2414 0 wbs_dat_o[14]
rlabel metal2 7682 2132 7682 2132 0 wbs_dat_o[15]
rlabel metal2 7958 1860 7958 1860 0 wbs_dat_o[16]
rlabel metal2 8234 1622 8234 1622 0 wbs_dat_o[17]
rlabel metal2 8510 2132 8510 2132 0 wbs_dat_o[18]
rlabel metal2 8786 1826 8786 1826 0 wbs_dat_o[19]
rlabel metal2 3542 1622 3542 1622 0 wbs_dat_o[1]
rlabel metal2 9062 1792 9062 1792 0 wbs_dat_o[20]
rlabel metal2 9338 2132 9338 2132 0 wbs_dat_o[21]
rlabel metal2 9614 1656 9614 1656 0 wbs_dat_o[22]
rlabel metal2 9890 1860 9890 1860 0 wbs_dat_o[23]
rlabel metal2 10166 2132 10166 2132 0 wbs_dat_o[24]
rlabel metal2 10442 1622 10442 1622 0 wbs_dat_o[25]
rlabel metal2 10718 1792 10718 1792 0 wbs_dat_o[26]
rlabel metal2 10994 2132 10994 2132 0 wbs_dat_o[27]
rlabel metal2 11270 1826 11270 1826 0 wbs_dat_o[28]
rlabel metal2 11546 1656 11546 1656 0 wbs_dat_o[29]
rlabel metal2 3910 1792 3910 1792 0 wbs_dat_o[2]
rlabel metal2 11822 2132 11822 2132 0 wbs_dat_o[30]
rlabel metal2 12098 1792 12098 1792 0 wbs_dat_o[31]
rlabel metal2 4278 1656 4278 1656 0 wbs_dat_o[3]
rlabel metal2 4646 1588 4646 1588 0 wbs_dat_o[4]
rlabel metal2 4922 1826 4922 1826 0 wbs_dat_o[5]
rlabel metal2 5198 2132 5198 2132 0 wbs_dat_o[6]
rlabel metal2 5474 1860 5474 1860 0 wbs_dat_o[7]
rlabel metal2 5750 1588 5750 1588 0 wbs_dat_o[8]
rlabel metal2 6026 2132 6026 2132 0 wbs_dat_o[9]
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
