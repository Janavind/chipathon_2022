magic
tech sky130B
magscale 1 2
timestamp 1666199351
use sky130_fd_pr__dfl1sd2__example_55959141808515  sky130_fd_pr__dfl1sd2__example_55959141808515_0
timestamp 1666199351
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808515  sky130_fd_pr__dfl1sd2__example_55959141808515_1
timestamp 1666199351
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808515  sky130_fd_pr__dfl1sd2__example_55959141808515_2
timestamp 1666199351
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808340  sky130_fd_pr__dfl1sd__example_55959141808340_0
timestamp 1666199351
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808340  sky130_fd_pr__dfl1sd__example_55959141808340_1
timestamp 1666199351
transform 1 0 568 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 28908838
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 28906240
<< end >>
