magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 643 203
rect 29 -17 63 21
<< scnmos >>
rect 84 47 114 177
rect 169 47 199 177
rect 255 47 285 177
rect 327 47 357 177
rect 423 47 453 177
rect 507 47 537 177
<< scpmoshvt >>
rect 83 297 113 497
rect 169 297 199 497
rect 255 297 285 497
rect 339 297 369 497
rect 423 297 453 497
rect 507 297 537 497
<< ndiff >>
rect 27 157 84 177
rect 27 123 39 157
rect 73 123 84 157
rect 27 89 84 123
rect 27 55 39 89
rect 73 55 84 89
rect 27 47 84 55
rect 114 47 169 177
rect 199 157 255 177
rect 199 123 210 157
rect 244 123 255 157
rect 199 89 255 123
rect 199 55 210 89
rect 244 55 255 89
rect 199 47 255 55
rect 285 47 327 177
rect 357 89 423 177
rect 357 55 368 89
rect 402 55 423 89
rect 357 47 423 55
rect 453 169 507 177
rect 453 135 463 169
rect 497 135 507 169
rect 453 101 507 135
rect 453 67 463 101
rect 497 67 507 101
rect 453 47 507 67
rect 537 165 617 177
rect 537 131 575 165
rect 609 131 617 165
rect 537 93 617 131
rect 537 59 575 93
rect 609 59 617 93
rect 537 47 617 59
<< pdiff >>
rect 27 477 83 497
rect 27 443 38 477
rect 72 443 83 477
rect 27 409 83 443
rect 27 375 38 409
rect 72 375 83 409
rect 27 297 83 375
rect 113 489 169 497
rect 113 455 124 489
rect 158 455 169 489
rect 113 297 169 455
rect 199 477 255 497
rect 199 443 210 477
rect 244 443 255 477
rect 199 405 255 443
rect 199 371 210 405
rect 244 371 255 405
rect 199 297 255 371
rect 285 489 339 497
rect 285 455 295 489
rect 329 455 339 489
rect 285 297 339 455
rect 369 489 423 497
rect 369 455 379 489
rect 413 455 423 489
rect 369 421 423 455
rect 369 387 379 421
rect 413 387 423 421
rect 369 297 423 387
rect 453 407 507 497
rect 453 373 463 407
rect 497 373 507 407
rect 453 339 507 373
rect 453 305 463 339
rect 497 305 507 339
rect 453 297 507 305
rect 537 477 609 497
rect 537 443 567 477
rect 601 443 609 477
rect 537 409 609 443
rect 537 375 567 409
rect 601 375 609 409
rect 537 297 609 375
<< ndiffc >>
rect 39 123 73 157
rect 39 55 73 89
rect 210 123 244 157
rect 210 55 244 89
rect 368 55 402 89
rect 463 135 497 169
rect 463 67 497 101
rect 575 131 609 165
rect 575 59 609 93
<< pdiffc >>
rect 38 443 72 477
rect 38 375 72 409
rect 124 455 158 489
rect 210 443 244 477
rect 210 371 244 405
rect 295 455 329 489
rect 379 455 413 489
rect 379 387 413 421
rect 463 373 497 407
rect 463 305 497 339
rect 567 443 601 477
rect 567 375 601 409
<< poly >>
rect 83 497 113 523
rect 169 497 199 523
rect 255 497 285 523
rect 339 497 369 523
rect 423 497 453 523
rect 507 497 537 523
rect 83 261 113 297
rect 169 265 199 297
rect 255 265 285 297
rect 339 265 369 297
rect 47 259 113 261
rect 47 249 114 259
rect 47 215 63 249
rect 97 215 114 249
rect 47 203 114 215
rect 84 177 114 203
rect 163 249 285 265
rect 163 215 173 249
rect 207 215 241 249
rect 275 215 285 249
rect 163 199 285 215
rect 169 177 199 199
rect 255 177 285 199
rect 327 249 381 265
rect 327 215 337 249
rect 371 215 381 249
rect 327 199 381 215
rect 423 261 453 297
rect 507 261 537 297
rect 423 249 623 261
rect 423 215 573 249
rect 607 215 623 249
rect 423 203 623 215
rect 327 177 357 199
rect 423 177 453 203
rect 507 177 537 203
rect 84 21 114 47
rect 169 21 199 47
rect 255 21 285 47
rect 327 21 357 47
rect 423 21 453 47
rect 507 21 537 47
<< polycont >>
rect 63 215 97 249
rect 173 215 207 249
rect 241 215 275 249
rect 337 215 371 249
rect 573 215 607 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 22 477 74 493
rect 22 443 38 477
rect 72 443 74 477
rect 108 489 174 527
rect 108 455 124 489
rect 158 455 174 489
rect 210 477 244 493
rect 22 421 74 443
rect 210 421 244 443
rect 295 489 329 527
rect 295 439 329 455
rect 363 489 618 493
rect 363 455 379 489
rect 413 477 618 489
rect 413 457 567 477
rect 413 455 429 457
rect 22 409 244 421
rect 22 375 38 409
rect 72 405 244 409
rect 363 421 429 455
rect 557 443 567 457
rect 601 443 618 477
rect 363 405 379 421
rect 72 375 210 405
rect 22 371 210 375
rect 244 387 379 405
rect 413 387 429 421
rect 244 371 429 387
rect 463 407 523 423
rect 497 373 523 407
rect 463 339 523 373
rect 557 409 618 443
rect 557 375 567 409
rect 601 375 618 409
rect 557 359 618 375
rect 29 299 386 335
rect 29 249 129 299
rect 29 215 63 249
rect 97 215 129 249
rect 29 207 129 215
rect 163 249 285 265
rect 163 215 173 249
rect 207 215 241 249
rect 275 215 285 249
rect 321 249 386 299
rect 497 305 523 339
rect 321 215 337 249
rect 371 215 387 249
rect 163 199 285 215
rect 20 157 79 173
rect 463 169 523 305
rect 560 249 615 325
rect 560 215 573 249
rect 607 215 615 249
rect 560 199 615 215
rect 20 123 39 157
rect 73 123 79 157
rect 20 89 79 123
rect 20 55 39 89
rect 73 55 79 89
rect 20 17 79 55
rect 191 123 210 157
rect 244 135 463 157
rect 497 135 523 169
rect 244 123 523 135
rect 191 89 260 123
rect 459 101 523 123
rect 191 55 210 89
rect 244 55 260 89
rect 191 51 260 55
rect 352 55 368 89
rect 402 55 418 89
rect 352 17 418 55
rect 459 67 463 101
rect 497 67 523 101
rect 459 51 523 67
rect 559 131 575 165
rect 609 131 625 165
rect 559 93 625 131
rect 559 59 575 93
rect 609 59 625 93
rect 559 17 625 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 581 221 615 255 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 581 289 615 323 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 340 180 0 0 A2
port 2 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 340 180 0 0 A1
port 1 nsew signal input
flabel locali s 489 85 523 119 0 FreeSans 340 180 0 0 Y
port 8 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a21oi_2
rlabel metal1 s 0 -48 644 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 4037950
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4032086
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
