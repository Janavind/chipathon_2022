magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 2000 203
rect 29 -17 63 21
<< scnmos >>
rect 82 47 112 177
rect 166 47 196 177
rect 250 47 280 177
rect 334 47 364 177
rect 418 47 448 177
rect 502 47 532 177
rect 586 47 616 177
rect 670 47 700 177
rect 858 47 888 177
rect 942 47 972 177
rect 1026 47 1056 177
rect 1110 47 1140 177
rect 1194 47 1224 177
rect 1278 47 1308 177
rect 1362 47 1392 177
rect 1446 47 1476 177
rect 1636 47 1666 177
rect 1720 47 1750 177
rect 1804 47 1834 177
rect 1888 47 1918 177
<< scpmoshvt >>
rect 82 297 112 497
rect 166 297 196 497
rect 250 297 280 497
rect 334 297 364 497
rect 418 297 448 497
rect 502 297 532 497
rect 586 297 616 497
rect 670 297 700 497
rect 858 297 888 497
rect 942 297 972 497
rect 1026 297 1056 497
rect 1110 297 1140 497
rect 1194 297 1224 497
rect 1278 297 1308 497
rect 1362 297 1392 497
rect 1446 297 1476 497
rect 1636 297 1666 497
rect 1720 297 1750 497
rect 1804 297 1834 497
rect 1888 297 1918 497
<< ndiff >>
rect 27 95 82 177
rect 27 61 38 95
rect 72 61 82 95
rect 27 47 82 61
rect 112 163 166 177
rect 112 129 122 163
rect 156 129 166 163
rect 112 95 166 129
rect 112 61 122 95
rect 156 61 166 95
rect 112 47 166 61
rect 196 95 250 177
rect 196 61 206 95
rect 240 61 250 95
rect 196 47 250 61
rect 280 163 334 177
rect 280 129 290 163
rect 324 129 334 163
rect 280 95 334 129
rect 280 61 290 95
rect 324 61 334 95
rect 280 47 334 61
rect 364 95 418 177
rect 364 61 374 95
rect 408 61 418 95
rect 364 47 418 61
rect 448 163 502 177
rect 448 129 458 163
rect 492 129 502 163
rect 448 95 502 129
rect 448 61 458 95
rect 492 61 502 95
rect 448 47 502 61
rect 532 95 586 177
rect 532 61 542 95
rect 576 61 586 95
rect 532 47 586 61
rect 616 163 670 177
rect 616 129 626 163
rect 660 129 670 163
rect 616 95 670 129
rect 616 61 626 95
rect 660 61 670 95
rect 616 47 670 61
rect 700 163 752 177
rect 700 129 710 163
rect 744 129 752 163
rect 700 95 752 129
rect 700 61 710 95
rect 744 61 752 95
rect 700 47 752 61
rect 806 95 858 177
rect 806 61 814 95
rect 848 61 858 95
rect 806 47 858 61
rect 888 163 942 177
rect 888 129 898 163
rect 932 129 942 163
rect 888 47 942 129
rect 972 95 1026 177
rect 972 61 982 95
rect 1016 61 1026 95
rect 972 47 1026 61
rect 1056 163 1110 177
rect 1056 129 1066 163
rect 1100 129 1110 163
rect 1056 47 1110 129
rect 1140 163 1194 177
rect 1140 129 1150 163
rect 1184 129 1194 163
rect 1140 95 1194 129
rect 1140 61 1150 95
rect 1184 61 1194 95
rect 1140 47 1194 61
rect 1224 95 1278 177
rect 1224 61 1234 95
rect 1268 61 1278 95
rect 1224 47 1278 61
rect 1308 163 1362 177
rect 1308 129 1318 163
rect 1352 129 1362 163
rect 1308 95 1362 129
rect 1308 61 1318 95
rect 1352 61 1362 95
rect 1308 47 1362 61
rect 1392 95 1446 177
rect 1392 61 1402 95
rect 1436 61 1446 95
rect 1392 47 1446 61
rect 1476 163 1528 177
rect 1476 129 1486 163
rect 1520 129 1528 163
rect 1476 95 1528 129
rect 1476 61 1486 95
rect 1520 61 1528 95
rect 1476 47 1528 61
rect 1584 95 1636 177
rect 1584 61 1592 95
rect 1626 61 1636 95
rect 1584 47 1636 61
rect 1666 163 1720 177
rect 1666 129 1676 163
rect 1710 129 1720 163
rect 1666 95 1720 129
rect 1666 61 1676 95
rect 1710 61 1720 95
rect 1666 47 1720 61
rect 1750 95 1804 177
rect 1750 61 1760 95
rect 1794 61 1804 95
rect 1750 47 1804 61
rect 1834 163 1888 177
rect 1834 129 1844 163
rect 1878 129 1888 163
rect 1834 95 1888 129
rect 1834 61 1844 95
rect 1878 61 1888 95
rect 1834 47 1888 61
rect 1918 95 1974 177
rect 1918 61 1928 95
rect 1962 61 1974 95
rect 1918 47 1974 61
<< pdiff >>
rect 27 477 82 497
rect 27 443 38 477
rect 72 443 82 477
rect 27 409 82 443
rect 27 375 38 409
rect 72 375 82 409
rect 27 297 82 375
rect 112 485 166 497
rect 112 451 122 485
rect 156 451 166 485
rect 112 297 166 451
rect 196 477 250 497
rect 196 443 206 477
rect 240 443 250 477
rect 196 409 250 443
rect 196 375 206 409
rect 240 375 250 409
rect 196 297 250 375
rect 280 485 334 497
rect 280 451 290 485
rect 324 451 334 485
rect 280 297 334 451
rect 364 477 418 497
rect 364 443 374 477
rect 408 443 418 477
rect 364 409 418 443
rect 364 375 374 409
rect 408 375 418 409
rect 364 297 418 375
rect 448 409 502 497
rect 448 375 458 409
rect 492 375 502 409
rect 448 297 502 375
rect 532 477 586 497
rect 532 443 542 477
rect 576 443 586 477
rect 532 297 586 443
rect 616 409 670 497
rect 616 375 626 409
rect 660 375 670 409
rect 616 297 670 375
rect 700 477 752 497
rect 700 443 710 477
rect 744 443 752 477
rect 700 409 752 443
rect 700 375 710 409
rect 744 375 752 409
rect 700 297 752 375
rect 806 477 858 497
rect 806 443 814 477
rect 848 443 858 477
rect 806 409 858 443
rect 806 375 814 409
rect 848 375 858 409
rect 806 297 858 375
rect 888 485 942 497
rect 888 451 898 485
rect 932 451 942 485
rect 888 297 942 451
rect 972 477 1026 497
rect 972 443 982 477
rect 1016 443 1026 477
rect 972 409 1026 443
rect 972 375 982 409
rect 1016 375 1026 409
rect 972 297 1026 375
rect 1056 485 1110 497
rect 1056 451 1066 485
rect 1100 451 1110 485
rect 1056 297 1110 451
rect 1140 477 1194 497
rect 1140 443 1150 477
rect 1184 443 1194 477
rect 1140 409 1194 443
rect 1140 375 1150 409
rect 1184 375 1194 409
rect 1140 297 1194 375
rect 1224 485 1278 497
rect 1224 451 1234 485
rect 1268 451 1278 485
rect 1224 297 1278 451
rect 1308 477 1362 497
rect 1308 443 1318 477
rect 1352 443 1362 477
rect 1308 409 1362 443
rect 1308 375 1318 409
rect 1352 375 1362 409
rect 1308 341 1362 375
rect 1308 307 1318 341
rect 1352 307 1362 341
rect 1308 297 1362 307
rect 1392 485 1446 497
rect 1392 451 1402 485
rect 1436 451 1446 485
rect 1392 297 1446 451
rect 1476 477 1528 497
rect 1476 443 1486 477
rect 1520 443 1528 477
rect 1476 409 1528 443
rect 1476 375 1486 409
rect 1520 375 1528 409
rect 1476 361 1528 375
rect 1582 409 1636 497
rect 1582 375 1592 409
rect 1626 375 1636 409
rect 1476 297 1526 361
rect 1582 346 1636 375
rect 1580 339 1636 346
rect 1580 305 1592 339
rect 1626 305 1636 339
rect 1580 297 1636 305
rect 1666 485 1720 497
rect 1666 451 1676 485
rect 1710 451 1720 485
rect 1666 417 1720 451
rect 1666 383 1676 417
rect 1710 383 1720 417
rect 1666 297 1720 383
rect 1750 409 1804 497
rect 1750 375 1760 409
rect 1794 375 1804 409
rect 1750 341 1804 375
rect 1750 307 1760 341
rect 1794 307 1804 341
rect 1750 297 1804 307
rect 1834 477 1888 497
rect 1834 443 1844 477
rect 1878 443 1888 477
rect 1834 409 1888 443
rect 1834 375 1844 409
rect 1878 375 1888 409
rect 1834 297 1888 375
rect 1918 477 1974 497
rect 1918 443 1928 477
rect 1962 443 1974 477
rect 1918 409 1974 443
rect 1918 375 1928 409
rect 1962 375 1974 409
rect 1918 341 1974 375
rect 1918 307 1928 341
rect 1962 307 1974 341
rect 1918 297 1974 307
<< ndiffc >>
rect 38 61 72 95
rect 122 129 156 163
rect 122 61 156 95
rect 206 61 240 95
rect 290 129 324 163
rect 290 61 324 95
rect 374 61 408 95
rect 458 129 492 163
rect 458 61 492 95
rect 542 61 576 95
rect 626 129 660 163
rect 626 61 660 95
rect 710 129 744 163
rect 710 61 744 95
rect 814 61 848 95
rect 898 129 932 163
rect 982 61 1016 95
rect 1066 129 1100 163
rect 1150 129 1184 163
rect 1150 61 1184 95
rect 1234 61 1268 95
rect 1318 129 1352 163
rect 1318 61 1352 95
rect 1402 61 1436 95
rect 1486 129 1520 163
rect 1486 61 1520 95
rect 1592 61 1626 95
rect 1676 129 1710 163
rect 1676 61 1710 95
rect 1760 61 1794 95
rect 1844 129 1878 163
rect 1844 61 1878 95
rect 1928 61 1962 95
<< pdiffc >>
rect 38 443 72 477
rect 38 375 72 409
rect 122 451 156 485
rect 206 443 240 477
rect 206 375 240 409
rect 290 451 324 485
rect 374 443 408 477
rect 374 375 408 409
rect 458 375 492 409
rect 542 443 576 477
rect 626 375 660 409
rect 710 443 744 477
rect 710 375 744 409
rect 814 443 848 477
rect 814 375 848 409
rect 898 451 932 485
rect 982 443 1016 477
rect 982 375 1016 409
rect 1066 451 1100 485
rect 1150 443 1184 477
rect 1150 375 1184 409
rect 1234 451 1268 485
rect 1318 443 1352 477
rect 1318 375 1352 409
rect 1318 307 1352 341
rect 1402 451 1436 485
rect 1486 443 1520 477
rect 1486 375 1520 409
rect 1592 375 1626 409
rect 1592 305 1626 339
rect 1676 451 1710 485
rect 1676 383 1710 417
rect 1760 375 1794 409
rect 1760 307 1794 341
rect 1844 443 1878 477
rect 1844 375 1878 409
rect 1928 443 1962 477
rect 1928 375 1962 409
rect 1928 307 1962 341
<< poly >>
rect 82 497 112 523
rect 166 497 196 523
rect 250 497 280 523
rect 334 497 364 523
rect 418 497 448 523
rect 502 497 532 523
rect 586 497 616 523
rect 670 497 700 523
rect 858 497 888 523
rect 942 497 972 523
rect 1026 497 1056 523
rect 1110 497 1140 523
rect 1194 497 1224 523
rect 1278 497 1308 523
rect 1362 497 1392 523
rect 1446 497 1476 523
rect 1636 497 1666 523
rect 1720 497 1750 523
rect 1804 497 1834 523
rect 1888 497 1918 523
rect 82 265 112 297
rect 166 265 196 297
rect 250 265 280 297
rect 334 265 364 297
rect 82 249 364 265
rect 82 215 102 249
rect 136 215 170 249
rect 204 215 238 249
rect 272 215 306 249
rect 340 215 364 249
rect 82 199 364 215
rect 82 177 112 199
rect 166 177 196 199
rect 250 177 280 199
rect 334 177 364 199
rect 418 265 448 297
rect 502 265 532 297
rect 586 265 616 297
rect 670 265 700 297
rect 858 265 888 297
rect 942 265 972 297
rect 1026 265 1056 297
rect 1110 265 1140 297
rect 418 249 1140 265
rect 418 215 610 249
rect 644 215 678 249
rect 712 215 746 249
rect 780 215 814 249
rect 848 215 882 249
rect 916 215 950 249
rect 984 215 1140 249
rect 418 199 1140 215
rect 418 177 448 199
rect 502 177 532 199
rect 586 177 616 199
rect 670 177 700 199
rect 858 177 888 199
rect 942 177 972 199
rect 1026 177 1056 199
rect 1110 177 1140 199
rect 1194 265 1224 297
rect 1278 265 1308 297
rect 1362 265 1392 297
rect 1446 265 1476 297
rect 1194 249 1476 265
rect 1194 215 1217 249
rect 1251 215 1285 249
rect 1319 215 1353 249
rect 1387 215 1421 249
rect 1455 215 1476 249
rect 1194 199 1476 215
rect 1194 177 1224 199
rect 1278 177 1308 199
rect 1362 177 1392 199
rect 1446 177 1476 199
rect 1636 265 1666 297
rect 1720 265 1750 297
rect 1804 265 1834 297
rect 1888 265 1918 297
rect 1636 249 1918 265
rect 1636 215 1724 249
rect 1758 215 1792 249
rect 1826 215 1860 249
rect 1894 215 1918 249
rect 1636 199 1918 215
rect 1636 177 1666 199
rect 1720 177 1750 199
rect 1804 177 1834 199
rect 1888 177 1918 199
rect 82 21 112 47
rect 166 21 196 47
rect 250 21 280 47
rect 334 21 364 47
rect 418 21 448 47
rect 502 21 532 47
rect 586 21 616 47
rect 670 21 700 47
rect 858 21 888 47
rect 942 21 972 47
rect 1026 21 1056 47
rect 1110 21 1140 47
rect 1194 21 1224 47
rect 1278 21 1308 47
rect 1362 21 1392 47
rect 1446 21 1476 47
rect 1636 21 1666 47
rect 1720 21 1750 47
rect 1804 21 1834 47
rect 1888 21 1918 47
<< polycont >>
rect 102 215 136 249
rect 170 215 204 249
rect 238 215 272 249
rect 306 215 340 249
rect 610 215 644 249
rect 678 215 712 249
rect 746 215 780 249
rect 814 215 848 249
rect 882 215 916 249
rect 950 215 984 249
rect 1217 215 1251 249
rect 1285 215 1319 249
rect 1353 215 1387 249
rect 1421 215 1455 249
rect 1724 215 1758 249
rect 1792 215 1826 249
rect 1860 215 1894 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 17 477 80 493
rect 17 443 38 477
rect 72 443 80 477
rect 17 409 80 443
rect 114 485 164 527
rect 114 451 122 485
rect 156 451 164 485
rect 114 435 164 451
rect 198 477 248 493
rect 198 443 206 477
rect 240 443 248 477
rect 17 375 38 409
rect 72 401 80 409
rect 198 409 248 443
rect 282 485 332 527
rect 282 451 290 485
rect 324 451 332 485
rect 282 435 332 451
rect 366 477 752 493
rect 366 443 374 477
rect 408 459 542 477
rect 408 443 416 459
rect 198 401 206 409
rect 72 375 206 401
rect 240 401 248 409
rect 366 409 416 443
rect 534 443 542 459
rect 576 459 710 477
rect 576 443 584 459
rect 534 425 584 443
rect 702 443 710 459
rect 744 443 752 477
rect 366 401 374 409
rect 240 375 374 401
rect 408 375 416 409
rect 17 357 416 375
rect 450 409 500 425
rect 450 375 458 409
rect 492 391 500 409
rect 618 409 668 425
rect 618 391 626 409
rect 492 375 626 391
rect 660 375 668 409
rect 450 357 668 375
rect 702 409 752 443
rect 702 375 710 409
rect 744 375 752 409
rect 702 359 752 375
rect 806 477 856 493
rect 806 443 814 477
rect 848 443 856 477
rect 806 409 856 443
rect 890 485 940 527
rect 890 451 898 485
rect 932 451 940 485
rect 890 435 940 451
rect 974 477 1024 493
rect 974 443 982 477
rect 1016 443 1024 477
rect 806 375 814 409
rect 848 401 856 409
rect 974 409 1024 443
rect 1058 485 1108 527
rect 1058 451 1066 485
rect 1100 451 1108 485
rect 1058 435 1108 451
rect 1142 477 1192 493
rect 1142 443 1150 477
rect 1184 443 1192 477
rect 974 401 982 409
rect 848 375 982 401
rect 1016 401 1024 409
rect 1142 409 1192 443
rect 1226 485 1276 527
rect 1226 451 1234 485
rect 1268 451 1276 485
rect 1226 435 1276 451
rect 1310 477 1360 493
rect 1310 443 1318 477
rect 1352 443 1360 477
rect 1142 401 1150 409
rect 1016 375 1150 401
rect 1184 401 1192 409
rect 1310 409 1360 443
rect 1394 485 1444 527
rect 1394 451 1402 485
rect 1436 451 1444 485
rect 1394 435 1444 451
rect 1478 485 1886 493
rect 1478 477 1676 485
rect 1478 443 1486 477
rect 1520 459 1676 477
rect 1520 443 1528 459
rect 1310 401 1318 409
rect 1184 375 1318 401
rect 1352 401 1360 409
rect 1478 409 1528 443
rect 1668 451 1676 459
rect 1710 477 1886 485
rect 1710 459 1844 477
rect 1710 451 1718 459
rect 1478 401 1486 409
rect 1352 375 1486 401
rect 1520 375 1528 409
rect 806 357 1528 375
rect 1576 409 1634 425
rect 1576 375 1592 409
rect 1626 375 1634 409
rect 450 323 484 357
rect 1310 341 1360 357
rect 17 289 397 323
rect 431 289 484 323
rect 526 289 1233 323
rect 1310 307 1318 341
rect 1352 307 1360 341
rect 1576 339 1634 375
rect 1668 417 1718 451
rect 1836 443 1844 459
rect 1878 443 1886 477
rect 1668 383 1676 417
rect 1710 383 1718 417
rect 1668 367 1718 383
rect 1752 409 1802 425
rect 1752 375 1760 409
rect 1794 375 1802 409
rect 1310 291 1360 307
rect 1452 289 1501 323
rect 1535 289 1542 323
rect 1576 305 1592 339
rect 1626 333 1634 339
rect 1752 341 1802 375
rect 1836 409 1886 443
rect 1836 375 1844 409
rect 1878 375 1886 409
rect 1836 359 1886 375
rect 1920 477 2007 493
rect 1920 443 1928 477
rect 1962 443 2007 477
rect 1920 409 2007 443
rect 1920 375 1928 409
rect 1962 375 2007 409
rect 1752 333 1760 341
rect 1626 307 1760 333
rect 1794 325 1802 341
rect 1920 341 2007 375
rect 1920 325 1928 341
rect 1794 307 1928 325
rect 1962 307 2007 341
rect 1626 305 2007 307
rect 1576 289 2007 305
rect 17 181 51 289
rect 526 255 560 289
rect 1199 255 1233 289
rect 1508 255 1542 289
rect 85 249 560 255
rect 85 215 102 249
rect 136 215 170 249
rect 204 215 238 249
rect 272 215 306 249
rect 340 215 560 249
rect 594 249 1148 255
rect 594 215 610 249
rect 644 215 678 249
rect 712 215 746 249
rect 780 215 814 249
rect 848 215 882 249
rect 916 215 950 249
rect 984 221 1148 249
rect 1199 249 1474 255
rect 984 215 1000 221
rect 1199 215 1217 249
rect 1251 215 1285 249
rect 1319 215 1353 249
rect 1387 215 1421 249
rect 1455 215 1474 249
rect 1508 249 1913 255
rect 1508 221 1724 249
rect 1708 215 1724 221
rect 1758 215 1792 249
rect 1826 215 1860 249
rect 1894 215 1913 249
rect 1030 181 1041 187
rect 17 163 676 181
rect 17 147 122 163
rect 106 129 122 147
rect 156 145 290 163
rect 156 129 172 145
rect 17 95 72 113
rect 17 61 38 95
rect 17 17 72 61
rect 106 95 172 129
rect 274 129 290 145
rect 324 145 458 163
rect 324 129 340 145
rect 106 61 122 95
rect 156 61 172 95
rect 106 51 172 61
rect 206 95 240 111
rect 206 17 240 61
rect 274 95 340 129
rect 442 129 458 145
rect 492 145 626 163
rect 492 129 508 145
rect 274 61 290 95
rect 324 61 340 95
rect 274 51 340 61
rect 374 95 408 111
rect 374 17 408 61
rect 442 95 508 129
rect 610 129 626 145
rect 660 129 676 163
rect 442 61 458 95
rect 492 61 508 95
rect 442 51 508 61
rect 542 95 576 111
rect 542 17 576 61
rect 610 95 676 129
rect 610 61 626 95
rect 660 61 676 95
rect 610 51 676 61
rect 710 163 764 179
rect 744 129 764 163
rect 833 163 1041 181
rect 1075 163 1116 187
rect 833 129 898 163
rect 932 153 1041 163
rect 932 129 1066 153
rect 1100 129 1116 163
rect 1150 163 1536 181
rect 1184 145 1318 163
rect 1184 129 1200 145
rect 710 95 764 129
rect 1150 95 1200 129
rect 1302 129 1318 145
rect 1352 145 1486 163
rect 1352 129 1368 145
rect 744 61 764 95
rect 710 17 764 61
rect 798 61 814 95
rect 848 61 982 95
rect 1016 61 1150 95
rect 1184 61 1200 95
rect 798 51 1200 61
rect 1234 95 1268 111
rect 1234 17 1268 61
rect 1302 95 1368 129
rect 1470 129 1486 145
rect 1520 129 1536 163
rect 1570 153 1593 187
rect 1627 181 1661 187
rect 1947 181 2007 289
rect 1627 163 2007 181
rect 1627 153 1676 163
rect 1570 145 1676 153
rect 1302 61 1318 95
rect 1352 61 1368 95
rect 1302 51 1368 61
rect 1402 95 1436 111
rect 1402 17 1436 61
rect 1470 95 1536 129
rect 1660 129 1676 145
rect 1710 147 1844 163
rect 1710 129 1726 147
rect 1470 61 1486 95
rect 1520 61 1536 95
rect 1470 51 1536 61
rect 1592 95 1626 111
rect 1592 17 1626 61
rect 1660 95 1726 129
rect 1828 129 1844 147
rect 1878 147 2007 163
rect 1878 129 1894 147
rect 1660 61 1676 95
rect 1710 61 1726 95
rect 1660 51 1726 61
rect 1760 95 1794 111
rect 1760 17 1794 61
rect 1828 95 1894 129
rect 1828 61 1844 95
rect 1878 61 1894 95
rect 1828 51 1894 61
rect 1928 95 1962 111
rect 1928 17 1962 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 397 289 431 323
rect 1501 289 1535 323
rect 1041 163 1075 187
rect 1041 153 1066 163
rect 1066 153 1075 163
rect 1593 153 1627 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 385 323 443 329
rect 385 289 397 323
rect 431 320 443 323
rect 1489 323 1547 329
rect 1489 320 1501 323
rect 431 292 1501 320
rect 431 289 443 292
rect 385 283 443 289
rect 1489 289 1501 292
rect 1535 289 1547 323
rect 1489 283 1547 289
rect 1029 187 1087 193
rect 1029 153 1041 187
rect 1075 184 1087 187
rect 1581 187 1639 193
rect 1581 184 1593 187
rect 1075 156 1593 184
rect 1075 153 1087 156
rect 1029 147 1087 153
rect 1581 153 1593 156
rect 1627 153 1639 187
rect 1581 147 1639 153
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel locali s 1961 357 1995 391 0 FreeSans 400 0 0 0 X
port 7 nsew signal output
flabel locali s 765 221 799 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 xor2_4
rlabel locali s 1947 181 2007 289 1 X
port 7 nsew signal output
rlabel locali s 1920 325 2007 493 1 X
port 7 nsew signal output
rlabel locali s 1828 51 1894 147 1 X
port 7 nsew signal output
rlabel locali s 1752 333 1802 425 1 X
port 7 nsew signal output
rlabel locali s 1660 51 1726 145 1 X
port 7 nsew signal output
rlabel locali s 1576 333 1634 425 1 X
port 7 nsew signal output
rlabel locali s 1576 325 1802 333 1 X
port 7 nsew signal output
rlabel locali s 1576 289 2007 325 1 X
port 7 nsew signal output
rlabel locali s 1570 181 1661 187 1 X
port 7 nsew signal output
rlabel locali s 1570 147 2007 181 1 X
port 7 nsew signal output
rlabel locali s 1570 145 1726 147 1 X
port 7 nsew signal output
rlabel metal1 s 1581 184 1639 193 1 X
port 7 nsew signal output
rlabel metal1 s 1581 147 1639 156 1 X
port 7 nsew signal output
rlabel metal1 s 1029 184 1087 193 1 X
port 7 nsew signal output
rlabel metal1 s 1029 156 1639 184 1 X
port 7 nsew signal output
rlabel metal1 s 1029 147 1087 156 1 X
port 7 nsew signal output
rlabel metal1 s 0 -48 2024 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2024 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_END 661364
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 646958
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 10.120 0.000 
<< end >>
