magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1165 203
rect 29 -17 63 21
<< locali >>
rect 1005 325 1055 425
rect 141 289 376 323
rect 141 255 175 289
rect 342 255 376 289
rect 109 215 175 255
rect 342 215 646 255
rect 1005 283 1179 325
rect 1097 181 1179 283
rect 725 145 1179 181
rect 725 129 791 145
rect 997 129 1063 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 24 427 80 493
rect 114 427 164 527
rect 198 459 416 493
rect 198 427 248 459
rect 366 427 416 459
rect 29 425 63 427
rect 213 425 247 427
rect 457 425 520 493
rect 554 427 604 527
rect 282 391 332 425
rect 478 391 520 425
rect 638 391 688 493
rect 722 427 783 527
rect 817 459 1139 493
rect 817 391 971 459
rect 24 357 444 391
rect 478 357 971 391
rect 24 181 58 357
rect 410 323 444 357
rect 1089 359 1139 459
rect 410 289 957 323
rect 209 221 213 255
rect 247 221 308 255
rect 209 215 308 221
rect 684 221 765 255
rect 799 221 818 255
rect 684 215 818 221
rect 923 249 957 289
rect 923 215 1055 249
rect 24 145 340 181
rect 38 17 72 111
rect 106 51 172 145
rect 206 17 240 111
rect 274 51 340 145
rect 462 145 680 181
rect 374 17 408 111
rect 462 51 528 145
rect 562 17 596 111
rect 630 95 680 145
rect 630 51 876 95
rect 929 17 963 111
rect 1097 17 1131 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 213 221 247 255
rect 765 221 799 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 201 255 259 261
rect 201 221 213 255
rect 247 252 259 255
rect 753 255 811 261
rect 753 252 765 255
rect 247 224 765 252
rect 247 221 259 224
rect 201 215 259 221
rect 753 221 765 224
rect 799 221 811 255
rect 753 215 811 221
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< obsm1 >>
rect 17 456 75 465
rect 201 456 259 465
rect 17 428 259 456
rect 17 419 75 428
rect 201 419 259 428
<< labels >>
rlabel locali s 342 215 646 255 6 A
port 1 nsew signal input
rlabel locali s 342 255 376 289 6 A
port 1 nsew signal input
rlabel locali s 109 215 175 255 6 A
port 1 nsew signal input
rlabel locali s 141 255 175 289 6 A
port 1 nsew signal input
rlabel locali s 141 289 376 323 6 A
port 1 nsew signal input
rlabel metal1 s 753 215 811 224 6 B
port 2 nsew signal input
rlabel metal1 s 201 215 259 224 6 B
port 2 nsew signal input
rlabel metal1 s 201 224 811 252 6 B
port 2 nsew signal input
rlabel metal1 s 753 252 811 261 6 B
port 2 nsew signal input
rlabel metal1 s 201 252 259 261 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 1196 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 1165 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 997 129 1063 145 6 X
port 7 nsew signal output
rlabel locali s 725 129 791 145 6 X
port 7 nsew signal output
rlabel locali s 725 145 1179 181 6 X
port 7 nsew signal output
rlabel locali s 1097 181 1179 283 6 X
port 7 nsew signal output
rlabel locali s 1005 283 1179 325 6 X
port 7 nsew signal output
rlabel locali s 1005 325 1055 425 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1196 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 646902
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 637824
<< end >>
