magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< locali >>
rect 2459 1416 2912 1450
rect 1488 1372 1504 1406
rect 1538 1372 1554 1406
rect 1504 1298 1538 1314
rect 1504 1248 1538 1264
rect 1504 1106 1538 1122
rect 1504 1056 1538 1072
rect 1488 964 1504 998
rect 1538 964 1554 998
rect 2459 920 2912 954
rect 921 705 1095 739
rect 1129 705 1145 739
rect 921 626 955 705
rect 2459 626 2912 660
rect 380 610 414 626
rect 1488 582 1504 616
rect 1538 582 1554 616
rect 380 560 414 576
rect 1504 508 1538 524
rect 1504 458 1538 474
rect 921 310 1015 344
rect 1049 310 1065 344
rect 1504 316 1538 332
rect 380 214 414 230
rect 380 164 414 180
rect 921 130 955 310
rect 1504 266 1538 282
rect 1488 174 1504 208
rect 1538 174 1554 208
rect 2459 130 2912 164
<< viali >>
rect 1504 1372 1538 1406
rect 1504 1264 1538 1298
rect 1504 1072 1538 1106
rect 1504 964 1538 998
rect 1095 705 1129 739
rect 380 576 414 610
rect 1504 582 1538 616
rect 1504 474 1538 508
rect 1015 310 1049 344
rect 380 180 414 214
rect 1504 282 1538 316
rect 1504 174 1538 208
<< metal1 >>
rect 80 1307 108 1500
rect 160 1415 188 1500
rect 142 1363 148 1415
rect 200 1363 206 1415
rect 62 1255 68 1307
rect 120 1255 126 1307
rect 80 229 108 1255
rect 160 625 188 1363
rect 1018 1121 1046 1500
rect 1006 1115 1058 1121
rect 1006 1057 1058 1063
rect 148 619 200 625
rect 142 567 148 619
rect 200 567 206 619
rect 365 567 371 619
rect 423 567 429 619
rect 148 561 200 567
rect 68 223 120 229
rect 62 171 68 223
rect 120 171 126 223
rect 68 165 120 171
rect 80 80 108 165
rect 160 80 188 561
rect 504 421 532 790
rect 776 421 804 790
rect 486 369 492 421
rect 544 369 550 421
rect 758 369 764 421
rect 816 369 822 421
rect 365 171 371 223
rect 423 171 429 223
rect 504 80 532 369
rect 776 80 804 369
rect 1018 356 1046 1057
rect 1098 751 1126 1500
rect 1178 1313 1206 1500
rect 1258 1421 1286 1500
rect 1246 1415 1298 1421
rect 1240 1363 1246 1415
rect 1298 1363 1304 1415
rect 1489 1363 1495 1415
rect 1547 1363 1553 1415
rect 1246 1357 1298 1363
rect 1166 1307 1218 1313
rect 1160 1255 1166 1307
rect 1218 1255 1224 1307
rect 1166 1249 1218 1255
rect 1089 739 1135 751
rect 1089 705 1095 739
rect 1129 705 1135 739
rect 1089 693 1135 705
rect 1098 631 1126 693
rect 1086 625 1138 631
rect 1086 567 1138 573
rect 1009 344 1055 356
rect 1009 331 1015 344
rect 1006 325 1015 331
rect 1049 331 1055 344
rect 1049 325 1058 331
rect 1006 267 1058 273
rect 1018 80 1046 267
rect 1098 223 1126 567
rect 1178 523 1206 1249
rect 1258 1013 1286 1357
rect 1489 1255 1495 1307
rect 1547 1255 1553 1307
rect 1664 1218 1712 1610
rect 2088 1218 2138 1612
rect 1656 1166 1662 1218
rect 1714 1166 1720 1218
rect 2081 1166 2087 1218
rect 2139 1166 2145 1218
rect 2478 1211 2506 1580
rect 2750 1211 2778 1580
rect 1489 1063 1495 1115
rect 1547 1063 1553 1115
rect 1246 1007 1298 1013
rect 1489 955 1495 1007
rect 1547 955 1553 1007
rect 1246 949 1298 955
rect 1166 517 1218 523
rect 1166 459 1218 465
rect 1086 217 1138 223
rect 1086 159 1138 165
rect 1098 80 1126 159
rect 1178 80 1206 459
rect 1258 80 1286 949
rect 1489 573 1495 625
rect 1547 573 1553 625
rect 1489 465 1495 517
rect 1547 465 1553 517
rect 1664 428 1712 1166
rect 2088 428 2138 1166
rect 2460 1159 2466 1211
rect 2518 1159 2524 1211
rect 2732 1159 2738 1211
rect 2790 1159 2796 1211
rect 1656 376 1662 428
rect 1714 376 1720 428
rect 2081 376 2087 428
rect 2139 376 2145 428
rect 2478 421 2506 1159
rect 2750 421 2778 1159
rect 1489 273 1495 325
rect 1547 273 1553 325
rect 1489 165 1495 217
rect 1547 165 1553 217
rect 1664 80 1712 376
rect 2088 80 2138 376
rect 2460 369 2466 421
rect 2518 369 2524 421
rect 2732 369 2738 421
rect 2790 369 2796 421
rect 2478 80 2506 369
rect 2750 80 2778 369
<< via1 >>
rect 148 1363 200 1415
rect 68 1255 120 1307
rect 1006 1063 1058 1115
rect 148 567 200 619
rect 371 610 423 619
rect 371 576 380 610
rect 380 576 414 610
rect 414 576 423 610
rect 371 567 423 576
rect 68 171 120 223
rect 492 369 544 421
rect 764 369 816 421
rect 371 214 423 223
rect 371 180 380 214
rect 380 180 414 214
rect 414 180 423 214
rect 371 171 423 180
rect 1246 1363 1298 1415
rect 1495 1406 1547 1415
rect 1495 1372 1504 1406
rect 1504 1372 1538 1406
rect 1538 1372 1547 1406
rect 1495 1363 1547 1372
rect 1166 1255 1218 1307
rect 1086 573 1138 625
rect 1006 310 1015 325
rect 1015 310 1049 325
rect 1049 310 1058 325
rect 1006 273 1058 310
rect 1495 1298 1547 1307
rect 1495 1264 1504 1298
rect 1504 1264 1538 1298
rect 1538 1264 1547 1298
rect 1495 1255 1547 1264
rect 1662 1166 1714 1218
rect 2087 1166 2139 1218
rect 1495 1106 1547 1115
rect 1495 1072 1504 1106
rect 1504 1072 1538 1106
rect 1538 1072 1547 1106
rect 1495 1063 1547 1072
rect 1246 955 1298 1007
rect 1495 998 1547 1007
rect 1495 964 1504 998
rect 1504 964 1538 998
rect 1538 964 1547 998
rect 1495 955 1547 964
rect 1166 465 1218 517
rect 1086 165 1138 217
rect 1495 616 1547 625
rect 1495 582 1504 616
rect 1504 582 1538 616
rect 1538 582 1547 616
rect 1495 573 1547 582
rect 1495 508 1547 517
rect 1495 474 1504 508
rect 1504 474 1538 508
rect 1538 474 1547 508
rect 1495 465 1547 474
rect 2466 1159 2518 1211
rect 2738 1159 2790 1211
rect 1662 376 1714 428
rect 2087 376 2139 428
rect 1495 316 1547 325
rect 1495 282 1504 316
rect 1504 282 1538 316
rect 1538 282 1547 316
rect 1495 273 1547 282
rect 1495 208 1547 217
rect 1495 174 1504 208
rect 1504 174 1538 208
rect 1538 174 1547 208
rect 1495 165 1547 174
rect 2466 369 2518 421
rect 2738 369 2790 421
<< metal2 >>
rect 148 1415 200 1421
rect 1246 1415 1298 1421
rect 1240 1403 1246 1415
rect 200 1375 1246 1403
rect 1240 1363 1246 1375
rect 1298 1403 1304 1415
rect 1489 1403 1495 1415
rect 1298 1375 1495 1403
rect 1298 1363 1304 1375
rect 1489 1363 1495 1375
rect 1547 1363 1553 1415
rect 148 1357 200 1363
rect 1246 1357 1298 1363
rect 68 1307 120 1313
rect 1166 1307 1218 1313
rect 1495 1307 1547 1313
rect 1160 1295 1166 1307
rect 120 1267 1166 1295
rect 1160 1255 1166 1267
rect 1218 1295 1224 1307
rect 1218 1267 1495 1295
rect 1218 1255 1224 1267
rect 68 1249 120 1255
rect 1166 1249 1218 1255
rect 1495 1249 1547 1255
rect 1660 1220 1716 1229
rect 1660 1155 1716 1164
rect 2085 1220 2141 1229
rect 2085 1155 2141 1164
rect 2464 1213 2520 1222
rect 2464 1148 2520 1157
rect 2736 1213 2792 1222
rect 2736 1148 2792 1157
rect 1495 1115 1547 1121
rect 1000 1063 1006 1115
rect 1058 1103 1064 1115
rect 1058 1075 1495 1103
rect 1058 1063 1064 1075
rect 1495 1057 1547 1063
rect 1240 955 1246 1007
rect 1298 995 1304 1007
rect 1489 995 1495 1007
rect 1298 967 1495 995
rect 1298 955 1304 967
rect 1489 955 1495 967
rect 1547 955 1553 1007
rect 148 619 200 625
rect 371 619 423 625
rect 200 579 371 607
rect 148 561 200 567
rect 1080 573 1086 625
rect 1138 613 1144 625
rect 1489 613 1495 625
rect 1138 585 1495 613
rect 1138 573 1144 585
rect 1489 573 1495 585
rect 1547 573 1553 625
rect 371 561 423 567
rect 1495 517 1547 523
rect 1160 465 1166 517
rect 1218 505 1224 517
rect 1218 477 1495 505
rect 1218 465 1224 477
rect 1495 459 1547 465
rect 490 423 546 432
rect 490 358 546 367
rect 762 423 818 432
rect 762 358 818 367
rect 1660 430 1716 439
rect 1660 365 1716 374
rect 2085 430 2141 439
rect 2085 365 2141 374
rect 2464 423 2520 432
rect 2464 358 2520 367
rect 2736 423 2792 432
rect 2736 358 2792 367
rect 1495 325 1547 331
rect 1000 273 1006 325
rect 1058 313 1064 325
rect 1058 285 1495 313
rect 1058 273 1064 285
rect 1495 267 1547 273
rect 68 223 120 229
rect 371 223 423 229
rect 120 183 371 211
rect 68 165 120 171
rect 371 165 423 171
rect 1080 165 1086 217
rect 1138 205 1144 217
rect 1489 205 1495 217
rect 1138 177 1495 205
rect 1138 165 1144 177
rect 1489 165 1495 177
rect 1547 165 1553 217
<< via2 >>
rect 1660 1218 1716 1220
rect 1660 1166 1662 1218
rect 1662 1166 1714 1218
rect 1714 1166 1716 1218
rect 1660 1164 1716 1166
rect 2085 1218 2141 1220
rect 2085 1166 2087 1218
rect 2087 1166 2139 1218
rect 2139 1166 2141 1218
rect 2085 1164 2141 1166
rect 2464 1211 2520 1213
rect 2464 1159 2466 1211
rect 2466 1159 2518 1211
rect 2518 1159 2520 1211
rect 2464 1157 2520 1159
rect 2736 1211 2792 1213
rect 2736 1159 2738 1211
rect 2738 1159 2790 1211
rect 2790 1159 2792 1211
rect 2736 1157 2792 1159
rect 490 421 546 423
rect 490 369 492 421
rect 492 369 544 421
rect 544 369 546 421
rect 490 367 546 369
rect 762 421 818 423
rect 762 369 764 421
rect 764 369 816 421
rect 816 369 818 421
rect 762 367 818 369
rect 1660 428 1716 430
rect 1660 376 1662 428
rect 1662 376 1714 428
rect 1714 376 1716 428
rect 1660 374 1716 376
rect 2085 428 2141 430
rect 2085 376 2087 428
rect 2087 376 2139 428
rect 2139 376 2141 428
rect 2085 374 2141 376
rect 2464 421 2520 423
rect 2464 369 2466 421
rect 2466 369 2518 421
rect 2518 369 2520 421
rect 2464 367 2520 369
rect 2736 421 2792 423
rect 2736 369 2738 421
rect 2738 369 2790 421
rect 2790 369 2792 421
rect 2736 367 2792 369
<< metal3 >>
rect 1639 1220 1737 1241
rect 1639 1164 1660 1220
rect 1716 1164 1737 1220
rect 1639 1143 1737 1164
rect 2064 1220 2162 1241
rect 2064 1164 2085 1220
rect 2141 1164 2162 1220
rect 2064 1143 2162 1164
rect 2443 1213 2541 1234
rect 2443 1157 2464 1213
rect 2520 1157 2541 1213
rect 2443 1136 2541 1157
rect 2715 1213 2813 1234
rect 2715 1157 2736 1213
rect 2792 1157 2813 1213
rect 2715 1136 2813 1157
rect 469 423 567 444
rect 469 367 490 423
rect 546 367 567 423
rect 469 346 567 367
rect 741 423 839 444
rect 741 367 762 423
rect 818 367 839 423
rect 741 346 839 367
rect 1639 430 1737 451
rect 1639 374 1660 430
rect 1716 374 1737 430
rect 1639 353 1737 374
rect 2064 430 2162 451
rect 2064 374 2085 430
rect 2141 374 2162 430
rect 2064 353 2162 374
rect 2443 423 2541 444
rect 2443 367 2464 423
rect 2520 367 2541 423
rect 2443 346 2541 367
rect 2715 423 2813 444
rect 2715 367 2736 423
rect 2792 367 2813 423
rect 2715 346 2813 367
use and2_dec  and2_dec_0
timestamp 1666199351
transform 1 0 1418 0 -1 1580
box 70 -56 1512 490
use and2_dec  and2_dec_1
timestamp 1666199351
transform 1 0 1418 0 1 790
box 70 -56 1512 490
use and2_dec  and2_dec_2
timestamp 1666199351
transform 1 0 1418 0 -1 790
box 70 -56 1512 490
use and2_dec  and2_dec_3
timestamp 1666199351
transform 1 0 1418 0 1 0
box 70 -56 1512 490
use contact_7  contact_7_0
timestamp 1666199351
transform 1 0 1492 0 1 1248
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1666199351
transform 1 0 1492 0 1 1056
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1666199351
transform 1 0 1492 0 1 458
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1666199351
transform 1 0 1492 0 1 266
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1666199351
transform 1 0 368 0 1 560
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1666199351
transform 1 0 368 0 1 164
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1666199351
transform 1 0 1656 0 1 1160
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1666199351
transform 1 0 1656 0 1 1160
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1666199351
transform 1 0 2460 0 1 1153
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1666199351
transform 1 0 2460 0 1 1153
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1666199351
transform 1 0 1656 0 1 370
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1666199351
transform 1 0 1656 0 1 370
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1666199351
transform 1 0 2460 0 1 363
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1666199351
transform 1 0 2460 0 1 363
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1666199351
transform 1 0 486 0 1 363
box 0 0 1 1
use contact_8  contact_8_9
timestamp 1666199351
transform 1 0 486 0 1 363
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1666199351
transform 1 0 2081 0 1 1160
box 0 0 1 1
use contact_8  contact_8_11
timestamp 1666199351
transform 1 0 2081 0 1 1160
box 0 0 1 1
use contact_8  contact_8_12
timestamp 1666199351
transform 1 0 2732 0 1 1153
box 0 0 1 1
use contact_8  contact_8_13
timestamp 1666199351
transform 1 0 2732 0 1 1153
box 0 0 1 1
use contact_8  contact_8_14
timestamp 1666199351
transform 1 0 2081 0 1 370
box 0 0 1 1
use contact_8  contact_8_15
timestamp 1666199351
transform 1 0 2081 0 1 370
box 0 0 1 1
use contact_8  contact_8_16
timestamp 1666199351
transform 1 0 2732 0 1 363
box 0 0 1 1
use contact_8  contact_8_17
timestamp 1666199351
transform 1 0 2732 0 1 363
box 0 0 1 1
use contact_8  contact_8_18
timestamp 1666199351
transform 1 0 758 0 1 363
box 0 0 1 1
use contact_8  contact_8_19
timestamp 1666199351
transform 1 0 758 0 1 363
box 0 0 1 1
use contact_8  contact_8_20
timestamp 1666199351
transform 1 0 1489 0 1 1249
box 0 0 1 1
use contact_8  contact_8_21
timestamp 1666199351
transform 1 0 1489 0 1 1057
box 0 0 1 1
use contact_8  contact_8_22
timestamp 1666199351
transform 1 0 1489 0 1 459
box 0 0 1 1
use contact_8  contact_8_23
timestamp 1666199351
transform 1 0 1489 0 1 267
box 0 0 1 1
use contact_8  contact_8_24
timestamp 1666199351
transform 1 0 1240 0 1 1357
box 0 0 1 1
use contact_8  contact_8_25
timestamp 1666199351
transform 1 0 142 0 1 1357
box 0 0 1 1
use contact_8  contact_8_26
timestamp 1666199351
transform 1 0 1160 0 1 1249
box 0 0 1 1
use contact_8  contact_8_27
timestamp 1666199351
transform 1 0 62 0 1 1249
box 0 0 1 1
use contact_8  contact_8_28
timestamp 1666199351
transform 1 0 142 0 1 561
box 0 0 1 1
use contact_8  contact_8_29
timestamp 1666199351
transform 1 0 365 0 1 561
box 0 0 1 1
use contact_8  contact_8_30
timestamp 1666199351
transform 1 0 62 0 1 165
box 0 0 1 1
use contact_8  contact_8_31
timestamp 1666199351
transform 1 0 365 0 1 165
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1666199351
transform 1 0 1655 0 1 1155
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1666199351
transform 1 0 1655 0 1 1155
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1666199351
transform 1 0 2459 0 1 1148
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1666199351
transform 1 0 2459 0 1 1148
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1666199351
transform 1 0 1655 0 1 365
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1666199351
transform 1 0 1655 0 1 365
box 0 0 1 1
use contact_9  contact_9_6
timestamp 1666199351
transform 1 0 2459 0 1 358
box 0 0 1 1
use contact_9  contact_9_7
timestamp 1666199351
transform 1 0 2459 0 1 358
box 0 0 1 1
use contact_9  contact_9_8
timestamp 1666199351
transform 1 0 485 0 1 358
box 0 0 1 1
use contact_9  contact_9_9
timestamp 1666199351
transform 1 0 485 0 1 358
box 0 0 1 1
use contact_9  contact_9_10
timestamp 1666199351
transform 1 0 2080 0 1 1155
box 0 0 1 1
use contact_9  contact_9_11
timestamp 1666199351
transform 1 0 2080 0 1 1155
box 0 0 1 1
use contact_9  contact_9_12
timestamp 1666199351
transform 1 0 2731 0 1 1148
box 0 0 1 1
use contact_9  contact_9_13
timestamp 1666199351
transform 1 0 2731 0 1 1148
box 0 0 1 1
use contact_9  contact_9_14
timestamp 1666199351
transform 1 0 2080 0 1 365
box 0 0 1 1
use contact_9  contact_9_15
timestamp 1666199351
transform 1 0 2080 0 1 365
box 0 0 1 1
use contact_9  contact_9_16
timestamp 1666199351
transform 1 0 2731 0 1 358
box 0 0 1 1
use contact_9  contact_9_17
timestamp 1666199351
transform 1 0 2731 0 1 358
box 0 0 1 1
use contact_9  contact_9_18
timestamp 1666199351
transform 1 0 757 0 1 358
box 0 0 1 1
use contact_9  contact_9_19
timestamp 1666199351
transform 1 0 757 0 1 358
box 0 0 1 1
use contact_26  contact_26_0
timestamp 1666199351
transform 1 0 1079 0 1 693
box 0 0 1 1
use contact_26  contact_26_1
timestamp 1666199351
transform 1 0 999 0 1 298
box 0 0 1 1
use contact_27  contact_27_0
timestamp 1666199351
transform 1 0 1240 0 1 1357
box 0 0 1 1
use contact_27  contact_27_1
timestamp 1666199351
transform 1 0 1160 0 1 1249
box 0 0 1 1
use contact_27  contact_27_2
timestamp 1666199351
transform 1 0 1240 0 1 949
box 0 0 1 1
use contact_27  contact_27_3
timestamp 1666199351
transform 1 0 1000 0 1 1057
box 0 0 1 1
use contact_27  contact_27_4
timestamp 1666199351
transform 1 0 1080 0 1 567
box 0 0 1 1
use contact_27  contact_27_5
timestamp 1666199351
transform 1 0 1160 0 1 459
box 0 0 1 1
use contact_27  contact_27_6
timestamp 1666199351
transform 1 0 1080 0 1 159
box 0 0 1 1
use contact_27  contact_27_7
timestamp 1666199351
transform 1 0 1000 0 1 267
box 0 0 1 1
use contact_28  contact_28_0
timestamp 1666199351
transform 1 0 1488 0 1 1366
box 0 0 1 1
use contact_28  contact_28_1
timestamp 1666199351
transform 1 0 1488 0 1 958
box 0 0 1 1
use contact_28  contact_28_2
timestamp 1666199351
transform 1 0 1488 0 1 576
box 0 0 1 1
use contact_28  contact_28_3
timestamp 1666199351
transform 1 0 1488 0 1 168
box 0 0 1 1
use contact_29  contact_29_0
timestamp 1666199351
transform 1 0 1489 0 1 1363
box 0 0 1 1
use contact_29  contact_29_1
timestamp 1666199351
transform 1 0 1489 0 1 955
box 0 0 1 1
use contact_29  contact_29_2
timestamp 1666199351
transform 1 0 1489 0 1 573
box 0 0 1 1
use contact_29  contact_29_3
timestamp 1666199351
transform 1 0 1489 0 1 165
box 0 0 1 1
use pinv_dec  pinv_dec_0
timestamp 1666199351
transform 1 0 320 0 -1 790
box 44 0 636 490
use pinv_dec  pinv_dec_1
timestamp 1666199351
transform 1 0 320 0 1 0
box 44 0 636 490
<< labels >>
rlabel locali s 2685 643 2685 643 4 out_1
port 4 nsew
rlabel locali s 2685 147 2685 147 4 out_0
port 3 nsew
rlabel locali s 2685 937 2685 937 4 out_2
port 5 nsew
rlabel locali s 2685 1433 2685 1433 4 out_3
port 6 nsew
rlabel metal1 s 94 197 94 197 4 in_0
port 1 nsew
rlabel metal1 s 174 593 174 593 4 in_1
port 2 nsew
rlabel metal3 s 790 395 790 395 4 vdd
port 7 nsew
rlabel metal3 s 2113 402 2113 402 4 vdd
port 7 nsew
rlabel metal3 s 2113 1192 2113 1192 4 vdd
port 7 nsew
rlabel metal3 s 2764 1185 2764 1185 4 vdd
port 7 nsew
rlabel metal3 s 2764 395 2764 395 4 vdd
port 7 nsew
rlabel metal3 s 2492 395 2492 395 4 gnd
port 8 nsew
rlabel metal3 s 2492 1185 2492 1185 4 gnd
port 8 nsew
rlabel metal3 s 1688 402 1688 402 4 gnd
port 8 nsew
rlabel metal3 s 1688 1192 1688 1192 4 gnd
port 8 nsew
rlabel metal3 s 518 395 518 395 4 gnd
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 2912 1580
string GDS_END 112658
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 103804
<< end >>
