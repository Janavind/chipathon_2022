magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< metal4 >>
rect 0 39427 254 39451
rect 14746 39427 15000 39451
rect 0 39416 15000 39427
rect 0 39180 241 39416
rect 477 39180 568 39416
rect 804 39180 895 39416
rect 1131 39180 1222 39416
rect 1458 39180 1549 39416
rect 1785 39180 1876 39416
rect 2112 39180 2203 39416
rect 2439 39180 2530 39416
rect 2766 39180 2857 39416
rect 3093 39180 3184 39416
rect 3420 39180 3511 39416
rect 3747 39180 3838 39416
rect 4074 39180 4165 39416
rect 4401 39180 4492 39416
rect 4728 39180 4819 39416
rect 5055 39180 5146 39416
rect 5382 39180 5473 39416
rect 5709 39180 5800 39416
rect 6036 39180 6127 39416
rect 6363 39180 6454 39416
rect 6690 39180 6781 39416
rect 7017 39180 7108 39416
rect 7344 39180 7435 39416
rect 7671 39180 7762 39416
rect 7998 39180 8089 39416
rect 8325 39180 8415 39416
rect 8651 39180 8741 39416
rect 8977 39180 9067 39416
rect 9303 39180 9393 39416
rect 9629 39180 9719 39416
rect 9955 39180 10045 39416
rect 10281 39180 10371 39416
rect 10607 39180 10697 39416
rect 10933 39180 11023 39416
rect 11259 39180 11349 39416
rect 11585 39180 11675 39416
rect 11911 39180 12001 39416
rect 12237 39180 12327 39416
rect 12563 39180 12653 39416
rect 12889 39180 12979 39416
rect 13215 39180 13305 39416
rect 13541 39180 13631 39416
rect 13867 39180 13957 39416
rect 14193 39180 14283 39416
rect 14519 39180 14609 39416
rect 14845 39180 15000 39416
rect 0 39092 15000 39180
rect 0 38856 241 39092
rect 477 38856 568 39092
rect 804 38856 895 39092
rect 1131 38856 1222 39092
rect 1458 38856 1549 39092
rect 1785 38856 1876 39092
rect 2112 38856 2203 39092
rect 2439 38856 2530 39092
rect 2766 38856 2857 39092
rect 3093 38856 3184 39092
rect 3420 38856 3511 39092
rect 3747 38856 3838 39092
rect 4074 38856 4165 39092
rect 4401 38856 4492 39092
rect 4728 38856 4819 39092
rect 5055 38856 5146 39092
rect 5382 38856 5473 39092
rect 5709 38856 5800 39092
rect 6036 38856 6127 39092
rect 6363 38856 6454 39092
rect 6690 38856 6781 39092
rect 7017 38856 7108 39092
rect 7344 38856 7435 39092
rect 7671 38856 7762 39092
rect 7998 38856 8089 39092
rect 8325 38856 8415 39092
rect 8651 38856 8741 39092
rect 8977 38856 9067 39092
rect 9303 38856 9393 39092
rect 9629 38856 9719 39092
rect 9955 38856 10045 39092
rect 10281 38856 10371 39092
rect 10607 38856 10697 39092
rect 10933 38856 11023 39092
rect 11259 38856 11349 39092
rect 11585 38856 11675 39092
rect 11911 38856 12001 39092
rect 12237 38856 12327 39092
rect 12563 38856 12653 39092
rect 12889 38856 12979 39092
rect 13215 38856 13305 39092
rect 13541 38856 13631 39092
rect 13867 38856 13957 39092
rect 14193 38856 14283 39092
rect 14519 38856 14609 39092
rect 14845 38856 15000 39092
rect 0 38768 15000 38856
rect 0 38532 241 38768
rect 477 38532 568 38768
rect 804 38532 895 38768
rect 1131 38532 1222 38768
rect 1458 38532 1549 38768
rect 1785 38532 1876 38768
rect 2112 38532 2203 38768
rect 2439 38532 2530 38768
rect 2766 38532 2857 38768
rect 3093 38532 3184 38768
rect 3420 38532 3511 38768
rect 3747 38532 3838 38768
rect 4074 38532 4165 38768
rect 4401 38532 4492 38768
rect 4728 38532 4819 38768
rect 5055 38532 5146 38768
rect 5382 38532 5473 38768
rect 5709 38532 5800 38768
rect 6036 38532 6127 38768
rect 6363 38532 6454 38768
rect 6690 38532 6781 38768
rect 7017 38532 7108 38768
rect 7344 38532 7435 38768
rect 7671 38532 7762 38768
rect 7998 38532 8089 38768
rect 8325 38532 8415 38768
rect 8651 38532 8741 38768
rect 8977 38532 9067 38768
rect 9303 38532 9393 38768
rect 9629 38532 9719 38768
rect 9955 38532 10045 38768
rect 10281 38532 10371 38768
rect 10607 38532 10697 38768
rect 10933 38532 11023 38768
rect 11259 38532 11349 38768
rect 11585 38532 11675 38768
rect 11911 38532 12001 38768
rect 12237 38532 12327 38768
rect 12563 38532 12653 38768
rect 12889 38532 12979 38768
rect 13215 38532 13305 38768
rect 13541 38532 13631 38768
rect 13867 38532 13957 38768
rect 14193 38532 14283 38768
rect 14519 38532 14609 38768
rect 14845 38532 15000 38768
rect 0 38444 15000 38532
rect 0 38208 241 38444
rect 477 38208 568 38444
rect 804 38208 895 38444
rect 1131 38208 1222 38444
rect 1458 38208 1549 38444
rect 1785 38208 1876 38444
rect 2112 38208 2203 38444
rect 2439 38208 2530 38444
rect 2766 38208 2857 38444
rect 3093 38208 3184 38444
rect 3420 38208 3511 38444
rect 3747 38208 3838 38444
rect 4074 38208 4165 38444
rect 4401 38208 4492 38444
rect 4728 38208 4819 38444
rect 5055 38208 5146 38444
rect 5382 38208 5473 38444
rect 5709 38208 5800 38444
rect 6036 38208 6127 38444
rect 6363 38208 6454 38444
rect 6690 38208 6781 38444
rect 7017 38208 7108 38444
rect 7344 38208 7435 38444
rect 7671 38208 7762 38444
rect 7998 38208 8089 38444
rect 8325 38208 8415 38444
rect 8651 38208 8741 38444
rect 8977 38208 9067 38444
rect 9303 38208 9393 38444
rect 9629 38208 9719 38444
rect 9955 38208 10045 38444
rect 10281 38208 10371 38444
rect 10607 38208 10697 38444
rect 10933 38208 11023 38444
rect 11259 38208 11349 38444
rect 11585 38208 11675 38444
rect 11911 38208 12001 38444
rect 12237 38208 12327 38444
rect 12563 38208 12653 38444
rect 12889 38208 12979 38444
rect 13215 38208 13305 38444
rect 13541 38208 13631 38444
rect 13867 38208 13957 38444
rect 14193 38208 14283 38444
rect 14519 38208 14609 38444
rect 14845 38208 15000 38444
rect 0 38120 15000 38208
rect 0 37884 241 38120
rect 477 37884 568 38120
rect 804 37884 895 38120
rect 1131 37884 1222 38120
rect 1458 37884 1549 38120
rect 1785 37884 1876 38120
rect 2112 37884 2203 38120
rect 2439 37884 2530 38120
rect 2766 37884 2857 38120
rect 3093 37884 3184 38120
rect 3420 37884 3511 38120
rect 3747 37884 3838 38120
rect 4074 37884 4165 38120
rect 4401 37884 4492 38120
rect 4728 37884 4819 38120
rect 5055 37884 5146 38120
rect 5382 37884 5473 38120
rect 5709 37884 5800 38120
rect 6036 37884 6127 38120
rect 6363 37884 6454 38120
rect 6690 37884 6781 38120
rect 7017 37884 7108 38120
rect 7344 37884 7435 38120
rect 7671 37884 7762 38120
rect 7998 37884 8089 38120
rect 8325 37884 8415 38120
rect 8651 37884 8741 38120
rect 8977 37884 9067 38120
rect 9303 37884 9393 38120
rect 9629 37884 9719 38120
rect 9955 37884 10045 38120
rect 10281 37884 10371 38120
rect 10607 37884 10697 38120
rect 10933 37884 11023 38120
rect 11259 37884 11349 38120
rect 11585 37884 11675 38120
rect 11911 37884 12001 38120
rect 12237 37884 12327 38120
rect 12563 37884 12653 38120
rect 12889 37884 12979 38120
rect 13215 37884 13305 38120
rect 13541 37884 13631 38120
rect 13867 37884 13957 38120
rect 14193 37884 14283 38120
rect 14519 37884 14609 38120
rect 14845 37884 15000 38120
rect 0 37796 15000 37884
rect 0 37560 241 37796
rect 477 37560 568 37796
rect 804 37560 895 37796
rect 1131 37560 1222 37796
rect 1458 37560 1549 37796
rect 1785 37560 1876 37796
rect 2112 37560 2203 37796
rect 2439 37560 2530 37796
rect 2766 37560 2857 37796
rect 3093 37560 3184 37796
rect 3420 37560 3511 37796
rect 3747 37560 3838 37796
rect 4074 37560 4165 37796
rect 4401 37560 4492 37796
rect 4728 37560 4819 37796
rect 5055 37560 5146 37796
rect 5382 37560 5473 37796
rect 5709 37560 5800 37796
rect 6036 37560 6127 37796
rect 6363 37560 6454 37796
rect 6690 37560 6781 37796
rect 7017 37560 7108 37796
rect 7344 37560 7435 37796
rect 7671 37560 7762 37796
rect 7998 37560 8089 37796
rect 8325 37560 8415 37796
rect 8651 37560 8741 37796
rect 8977 37560 9067 37796
rect 9303 37560 9393 37796
rect 9629 37560 9719 37796
rect 9955 37560 10045 37796
rect 10281 37560 10371 37796
rect 10607 37560 10697 37796
rect 10933 37560 11023 37796
rect 11259 37560 11349 37796
rect 11585 37560 11675 37796
rect 11911 37560 12001 37796
rect 12237 37560 12327 37796
rect 12563 37560 12653 37796
rect 12889 37560 12979 37796
rect 13215 37560 13305 37796
rect 13541 37560 13631 37796
rect 13867 37560 13957 37796
rect 14193 37560 14283 37796
rect 14519 37560 14609 37796
rect 14845 37560 15000 37796
rect 0 37472 15000 37560
rect 0 37236 241 37472
rect 477 37236 568 37472
rect 804 37236 895 37472
rect 1131 37236 1222 37472
rect 1458 37236 1549 37472
rect 1785 37236 1876 37472
rect 2112 37236 2203 37472
rect 2439 37236 2530 37472
rect 2766 37236 2857 37472
rect 3093 37236 3184 37472
rect 3420 37236 3511 37472
rect 3747 37236 3838 37472
rect 4074 37236 4165 37472
rect 4401 37236 4492 37472
rect 4728 37236 4819 37472
rect 5055 37236 5146 37472
rect 5382 37236 5473 37472
rect 5709 37236 5800 37472
rect 6036 37236 6127 37472
rect 6363 37236 6454 37472
rect 6690 37236 6781 37472
rect 7017 37236 7108 37472
rect 7344 37236 7435 37472
rect 7671 37236 7762 37472
rect 7998 37236 8089 37472
rect 8325 37236 8415 37472
rect 8651 37236 8741 37472
rect 8977 37236 9067 37472
rect 9303 37236 9393 37472
rect 9629 37236 9719 37472
rect 9955 37236 10045 37472
rect 10281 37236 10371 37472
rect 10607 37236 10697 37472
rect 10933 37236 11023 37472
rect 11259 37236 11349 37472
rect 11585 37236 11675 37472
rect 11911 37236 12001 37472
rect 12237 37236 12327 37472
rect 12563 37236 12653 37472
rect 12889 37236 12979 37472
rect 13215 37236 13305 37472
rect 13541 37236 13631 37472
rect 13867 37236 13957 37472
rect 14193 37236 14283 37472
rect 14519 37236 14609 37472
rect 14845 37236 15000 37472
rect 0 37148 15000 37236
rect 0 36912 241 37148
rect 477 36912 568 37148
rect 804 36912 895 37148
rect 1131 36912 1222 37148
rect 1458 36912 1549 37148
rect 1785 36912 1876 37148
rect 2112 36912 2203 37148
rect 2439 36912 2530 37148
rect 2766 36912 2857 37148
rect 3093 36912 3184 37148
rect 3420 36912 3511 37148
rect 3747 36912 3838 37148
rect 4074 36912 4165 37148
rect 4401 36912 4492 37148
rect 4728 36912 4819 37148
rect 5055 36912 5146 37148
rect 5382 36912 5473 37148
rect 5709 36912 5800 37148
rect 6036 36912 6127 37148
rect 6363 36912 6454 37148
rect 6690 36912 6781 37148
rect 7017 36912 7108 37148
rect 7344 36912 7435 37148
rect 7671 36912 7762 37148
rect 7998 36912 8089 37148
rect 8325 36912 8415 37148
rect 8651 36912 8741 37148
rect 8977 36912 9067 37148
rect 9303 36912 9393 37148
rect 9629 36912 9719 37148
rect 9955 36912 10045 37148
rect 10281 36912 10371 37148
rect 10607 36912 10697 37148
rect 10933 36912 11023 37148
rect 11259 36912 11349 37148
rect 11585 36912 11675 37148
rect 11911 36912 12001 37148
rect 12237 36912 12327 37148
rect 12563 36912 12653 37148
rect 12889 36912 12979 37148
rect 13215 36912 13305 37148
rect 13541 36912 13631 37148
rect 13867 36912 13957 37148
rect 14193 36912 14283 37148
rect 14519 36912 14609 37148
rect 14845 36912 15000 37148
rect 0 36824 15000 36912
rect 0 36588 241 36824
rect 477 36588 568 36824
rect 804 36588 895 36824
rect 1131 36588 1222 36824
rect 1458 36588 1549 36824
rect 1785 36588 1876 36824
rect 2112 36588 2203 36824
rect 2439 36588 2530 36824
rect 2766 36588 2857 36824
rect 3093 36588 3184 36824
rect 3420 36588 3511 36824
rect 3747 36588 3838 36824
rect 4074 36588 4165 36824
rect 4401 36588 4492 36824
rect 4728 36588 4819 36824
rect 5055 36588 5146 36824
rect 5382 36588 5473 36824
rect 5709 36588 5800 36824
rect 6036 36588 6127 36824
rect 6363 36588 6454 36824
rect 6690 36588 6781 36824
rect 7017 36588 7108 36824
rect 7344 36588 7435 36824
rect 7671 36588 7762 36824
rect 7998 36588 8089 36824
rect 8325 36588 8415 36824
rect 8651 36588 8741 36824
rect 8977 36588 9067 36824
rect 9303 36588 9393 36824
rect 9629 36588 9719 36824
rect 9955 36588 10045 36824
rect 10281 36588 10371 36824
rect 10607 36588 10697 36824
rect 10933 36588 11023 36824
rect 11259 36588 11349 36824
rect 11585 36588 11675 36824
rect 11911 36588 12001 36824
rect 12237 36588 12327 36824
rect 12563 36588 12653 36824
rect 12889 36588 12979 36824
rect 13215 36588 13305 36824
rect 13541 36588 13631 36824
rect 13867 36588 13957 36824
rect 14193 36588 14283 36824
rect 14519 36588 14609 36824
rect 14845 36588 15000 36824
rect 0 36500 15000 36588
rect 0 36264 241 36500
rect 477 36264 568 36500
rect 804 36264 895 36500
rect 1131 36264 1222 36500
rect 1458 36264 1549 36500
rect 1785 36264 1876 36500
rect 2112 36264 2203 36500
rect 2439 36264 2530 36500
rect 2766 36264 2857 36500
rect 3093 36264 3184 36500
rect 3420 36264 3511 36500
rect 3747 36264 3838 36500
rect 4074 36264 4165 36500
rect 4401 36264 4492 36500
rect 4728 36264 4819 36500
rect 5055 36264 5146 36500
rect 5382 36264 5473 36500
rect 5709 36264 5800 36500
rect 6036 36264 6127 36500
rect 6363 36264 6454 36500
rect 6690 36264 6781 36500
rect 7017 36264 7108 36500
rect 7344 36264 7435 36500
rect 7671 36264 7762 36500
rect 7998 36264 8089 36500
rect 8325 36264 8415 36500
rect 8651 36264 8741 36500
rect 8977 36264 9067 36500
rect 9303 36264 9393 36500
rect 9629 36264 9719 36500
rect 9955 36264 10045 36500
rect 10281 36264 10371 36500
rect 10607 36264 10697 36500
rect 10933 36264 11023 36500
rect 11259 36264 11349 36500
rect 11585 36264 11675 36500
rect 11911 36264 12001 36500
rect 12237 36264 12327 36500
rect 12563 36264 12653 36500
rect 12889 36264 12979 36500
rect 13215 36264 13305 36500
rect 13541 36264 13631 36500
rect 13867 36264 13957 36500
rect 14193 36264 14283 36500
rect 14519 36264 14609 36500
rect 14845 36264 15000 36500
rect 0 36176 15000 36264
rect 0 35940 241 36176
rect 477 35940 568 36176
rect 804 35940 895 36176
rect 1131 35940 1222 36176
rect 1458 35940 1549 36176
rect 1785 35940 1876 36176
rect 2112 35940 2203 36176
rect 2439 35940 2530 36176
rect 2766 35940 2857 36176
rect 3093 35940 3184 36176
rect 3420 35940 3511 36176
rect 3747 35940 3838 36176
rect 4074 35940 4165 36176
rect 4401 35940 4492 36176
rect 4728 35940 4819 36176
rect 5055 35940 5146 36176
rect 5382 35940 5473 36176
rect 5709 35940 5800 36176
rect 6036 35940 6127 36176
rect 6363 35940 6454 36176
rect 6690 35940 6781 36176
rect 7017 35940 7108 36176
rect 7344 35940 7435 36176
rect 7671 35940 7762 36176
rect 7998 35940 8089 36176
rect 8325 35940 8415 36176
rect 8651 35940 8741 36176
rect 8977 35940 9067 36176
rect 9303 35940 9393 36176
rect 9629 35940 9719 36176
rect 9955 35940 10045 36176
rect 10281 35940 10371 36176
rect 10607 35940 10697 36176
rect 10933 35940 11023 36176
rect 11259 35940 11349 36176
rect 11585 35940 11675 36176
rect 11911 35940 12001 36176
rect 12237 35940 12327 36176
rect 12563 35940 12653 36176
rect 12889 35940 12979 36176
rect 13215 35940 13305 36176
rect 13541 35940 13631 36176
rect 13867 35940 13957 36176
rect 14193 35940 14283 36176
rect 14519 35940 14609 36176
rect 14845 35940 15000 36176
rect 0 35852 15000 35940
rect 0 35616 241 35852
rect 477 35616 568 35852
rect 804 35616 895 35852
rect 1131 35616 1222 35852
rect 1458 35616 1549 35852
rect 1785 35616 1876 35852
rect 2112 35616 2203 35852
rect 2439 35616 2530 35852
rect 2766 35616 2857 35852
rect 3093 35616 3184 35852
rect 3420 35616 3511 35852
rect 3747 35616 3838 35852
rect 4074 35616 4165 35852
rect 4401 35616 4492 35852
rect 4728 35616 4819 35852
rect 5055 35616 5146 35852
rect 5382 35616 5473 35852
rect 5709 35616 5800 35852
rect 6036 35616 6127 35852
rect 6363 35616 6454 35852
rect 6690 35616 6781 35852
rect 7017 35616 7108 35852
rect 7344 35616 7435 35852
rect 7671 35616 7762 35852
rect 7998 35616 8089 35852
rect 8325 35616 8415 35852
rect 8651 35616 8741 35852
rect 8977 35616 9067 35852
rect 9303 35616 9393 35852
rect 9629 35616 9719 35852
rect 9955 35616 10045 35852
rect 10281 35616 10371 35852
rect 10607 35616 10697 35852
rect 10933 35616 11023 35852
rect 11259 35616 11349 35852
rect 11585 35616 11675 35852
rect 11911 35616 12001 35852
rect 12237 35616 12327 35852
rect 12563 35616 12653 35852
rect 12889 35616 12979 35852
rect 13215 35616 13305 35852
rect 13541 35616 13631 35852
rect 13867 35616 13957 35852
rect 14193 35616 14283 35852
rect 14519 35616 14609 35852
rect 14845 35616 15000 35852
rect 0 35528 15000 35616
rect 0 35292 241 35528
rect 477 35292 568 35528
rect 804 35292 895 35528
rect 1131 35292 1222 35528
rect 1458 35292 1549 35528
rect 1785 35292 1876 35528
rect 2112 35292 2203 35528
rect 2439 35292 2530 35528
rect 2766 35292 2857 35528
rect 3093 35292 3184 35528
rect 3420 35292 3511 35528
rect 3747 35292 3838 35528
rect 4074 35292 4165 35528
rect 4401 35292 4492 35528
rect 4728 35292 4819 35528
rect 5055 35292 5146 35528
rect 5382 35292 5473 35528
rect 5709 35292 5800 35528
rect 6036 35292 6127 35528
rect 6363 35292 6454 35528
rect 6690 35292 6781 35528
rect 7017 35292 7108 35528
rect 7344 35292 7435 35528
rect 7671 35292 7762 35528
rect 7998 35292 8089 35528
rect 8325 35292 8415 35528
rect 8651 35292 8741 35528
rect 8977 35292 9067 35528
rect 9303 35292 9393 35528
rect 9629 35292 9719 35528
rect 9955 35292 10045 35528
rect 10281 35292 10371 35528
rect 10607 35292 10697 35528
rect 10933 35292 11023 35528
rect 11259 35292 11349 35528
rect 11585 35292 11675 35528
rect 11911 35292 12001 35528
rect 12237 35292 12327 35528
rect 12563 35292 12653 35528
rect 12889 35292 12979 35528
rect 13215 35292 13305 35528
rect 13541 35292 13631 35528
rect 13867 35292 13957 35528
rect 14193 35292 14283 35528
rect 14519 35292 14609 35528
rect 14845 35292 15000 35528
rect 0 35204 15000 35292
rect 0 34968 241 35204
rect 477 34968 568 35204
rect 804 34968 895 35204
rect 1131 34968 1222 35204
rect 1458 34968 1549 35204
rect 1785 34968 1876 35204
rect 2112 34968 2203 35204
rect 2439 34968 2530 35204
rect 2766 34968 2857 35204
rect 3093 34968 3184 35204
rect 3420 34968 3511 35204
rect 3747 34968 3838 35204
rect 4074 34968 4165 35204
rect 4401 34968 4492 35204
rect 4728 34968 4819 35204
rect 5055 34968 5146 35204
rect 5382 34968 5473 35204
rect 5709 34968 5800 35204
rect 6036 34968 6127 35204
rect 6363 34968 6454 35204
rect 6690 34968 6781 35204
rect 7017 34968 7108 35204
rect 7344 34968 7435 35204
rect 7671 34968 7762 35204
rect 7998 34968 8089 35204
rect 8325 34968 8415 35204
rect 8651 34968 8741 35204
rect 8977 34968 9067 35204
rect 9303 34968 9393 35204
rect 9629 34968 9719 35204
rect 9955 34968 10045 35204
rect 10281 34968 10371 35204
rect 10607 34968 10697 35204
rect 10933 34968 11023 35204
rect 11259 34968 11349 35204
rect 11585 34968 11675 35204
rect 11911 34968 12001 35204
rect 12237 34968 12327 35204
rect 12563 34968 12653 35204
rect 12889 34968 12979 35204
rect 13215 34968 13305 35204
rect 13541 34968 13631 35204
rect 13867 34968 13957 35204
rect 14193 34968 14283 35204
rect 14519 34968 14609 35204
rect 14845 34968 15000 35204
rect 0 34880 15000 34968
rect 0 34644 241 34880
rect 477 34644 568 34880
rect 804 34644 895 34880
rect 1131 34644 1222 34880
rect 1458 34644 1549 34880
rect 1785 34644 1876 34880
rect 2112 34644 2203 34880
rect 2439 34644 2530 34880
rect 2766 34644 2857 34880
rect 3093 34644 3184 34880
rect 3420 34644 3511 34880
rect 3747 34644 3838 34880
rect 4074 34644 4165 34880
rect 4401 34644 4492 34880
rect 4728 34644 4819 34880
rect 5055 34644 5146 34880
rect 5382 34644 5473 34880
rect 5709 34644 5800 34880
rect 6036 34644 6127 34880
rect 6363 34644 6454 34880
rect 6690 34644 6781 34880
rect 7017 34644 7108 34880
rect 7344 34644 7435 34880
rect 7671 34644 7762 34880
rect 7998 34644 8089 34880
rect 8325 34644 8415 34880
rect 8651 34644 8741 34880
rect 8977 34644 9067 34880
rect 9303 34644 9393 34880
rect 9629 34644 9719 34880
rect 9955 34644 10045 34880
rect 10281 34644 10371 34880
rect 10607 34644 10697 34880
rect 10933 34644 11023 34880
rect 11259 34644 11349 34880
rect 11585 34644 11675 34880
rect 11911 34644 12001 34880
rect 12237 34644 12327 34880
rect 12563 34644 12653 34880
rect 12889 34644 12979 34880
rect 13215 34644 13305 34880
rect 13541 34644 13631 34880
rect 13867 34644 13957 34880
rect 14193 34644 14283 34880
rect 14519 34644 14609 34880
rect 14845 34644 15000 34880
rect 0 34633 15000 34644
rect 0 34608 254 34633
rect 14746 34608 15000 34633
rect 0 18424 254 18451
rect 14746 18424 15000 18451
rect 0 18423 15000 18424
rect 0 18187 143 18423
rect 379 18187 465 18423
rect 701 18187 787 18423
rect 1023 18187 1109 18423
rect 1345 18187 1431 18423
rect 1667 18187 1753 18423
rect 1989 18187 2075 18423
rect 2311 18187 2397 18423
rect 2633 18187 2719 18423
rect 2955 18187 3041 18423
rect 3277 18187 3363 18423
rect 3599 18187 3685 18423
rect 3921 18187 4007 18423
rect 4243 18187 4329 18423
rect 4565 18187 4651 18423
rect 4887 18187 4973 18423
rect 5209 18187 5295 18423
rect 5531 18187 5617 18423
rect 5853 18187 5938 18423
rect 6174 18187 6259 18423
rect 6495 18187 6580 18423
rect 6816 18187 6901 18423
rect 7137 18187 7222 18423
rect 7458 18187 7543 18423
rect 7779 18187 7864 18423
rect 8100 18187 8185 18423
rect 8421 18187 8506 18423
rect 8742 18187 8827 18423
rect 9063 18187 9148 18423
rect 9384 18187 9469 18423
rect 9705 18187 9790 18423
rect 10026 18187 10111 18423
rect 10347 18187 10432 18423
rect 10668 18187 10753 18423
rect 10989 18187 11074 18423
rect 11310 18187 11395 18423
rect 11631 18187 11716 18423
rect 11952 18187 12037 18423
rect 12273 18187 12358 18423
rect 12594 18187 12679 18423
rect 12915 18187 13000 18423
rect 13236 18187 13321 18423
rect 13557 18187 13642 18423
rect 13878 18187 13963 18423
rect 14199 18187 14284 18423
rect 14520 18187 14605 18423
rect 14841 18187 15000 18423
rect 0 18087 15000 18187
rect 0 17851 143 18087
rect 379 17851 465 18087
rect 701 17851 787 18087
rect 1023 17851 1109 18087
rect 1345 17851 1431 18087
rect 1667 17851 1753 18087
rect 1989 17851 2075 18087
rect 2311 17851 2397 18087
rect 2633 17851 2719 18087
rect 2955 17851 3041 18087
rect 3277 17851 3363 18087
rect 3599 17851 3685 18087
rect 3921 17851 4007 18087
rect 4243 17851 4329 18087
rect 4565 17851 4651 18087
rect 4887 17851 4973 18087
rect 5209 17851 5295 18087
rect 5531 17851 5617 18087
rect 5853 17851 5938 18087
rect 6174 17851 6259 18087
rect 6495 17851 6580 18087
rect 6816 17851 6901 18087
rect 7137 17851 7222 18087
rect 7458 17851 7543 18087
rect 7779 17851 7864 18087
rect 8100 17851 8185 18087
rect 8421 17851 8506 18087
rect 8742 17851 8827 18087
rect 9063 17851 9148 18087
rect 9384 17851 9469 18087
rect 9705 17851 9790 18087
rect 10026 17851 10111 18087
rect 10347 17851 10432 18087
rect 10668 17851 10753 18087
rect 10989 17851 11074 18087
rect 11310 17851 11395 18087
rect 11631 17851 11716 18087
rect 11952 17851 12037 18087
rect 12273 17851 12358 18087
rect 12594 17851 12679 18087
rect 12915 17851 13000 18087
rect 13236 17851 13321 18087
rect 13557 17851 13642 18087
rect 13878 17851 13963 18087
rect 14199 17851 14284 18087
rect 14520 17851 14605 18087
rect 14841 17851 15000 18087
rect 0 17751 15000 17851
rect 0 17515 143 17751
rect 379 17515 465 17751
rect 701 17515 787 17751
rect 1023 17515 1109 17751
rect 1345 17515 1431 17751
rect 1667 17515 1753 17751
rect 1989 17515 2075 17751
rect 2311 17515 2397 17751
rect 2633 17515 2719 17751
rect 2955 17515 3041 17751
rect 3277 17515 3363 17751
rect 3599 17515 3685 17751
rect 3921 17515 4007 17751
rect 4243 17515 4329 17751
rect 4565 17515 4651 17751
rect 4887 17515 4973 17751
rect 5209 17515 5295 17751
rect 5531 17515 5617 17751
rect 5853 17515 5938 17751
rect 6174 17515 6259 17751
rect 6495 17515 6580 17751
rect 6816 17515 6901 17751
rect 7137 17515 7222 17751
rect 7458 17515 7543 17751
rect 7779 17515 7864 17751
rect 8100 17515 8185 17751
rect 8421 17515 8506 17751
rect 8742 17515 8827 17751
rect 9063 17515 9148 17751
rect 9384 17515 9469 17751
rect 9705 17515 9790 17751
rect 10026 17515 10111 17751
rect 10347 17515 10432 17751
rect 10668 17515 10753 17751
rect 10989 17515 11074 17751
rect 11310 17515 11395 17751
rect 11631 17515 11716 17751
rect 11952 17515 12037 17751
rect 12273 17515 12358 17751
rect 12594 17515 12679 17751
rect 12915 17515 13000 17751
rect 13236 17515 13321 17751
rect 13557 17515 13642 17751
rect 13878 17515 13963 17751
rect 14199 17515 14284 17751
rect 14520 17515 14605 17751
rect 14841 17515 15000 17751
rect 0 17415 15000 17515
rect 0 17179 143 17415
rect 379 17179 465 17415
rect 701 17179 787 17415
rect 1023 17179 1109 17415
rect 1345 17179 1431 17415
rect 1667 17179 1753 17415
rect 1989 17179 2075 17415
rect 2311 17179 2397 17415
rect 2633 17179 2719 17415
rect 2955 17179 3041 17415
rect 3277 17179 3363 17415
rect 3599 17179 3685 17415
rect 3921 17179 4007 17415
rect 4243 17179 4329 17415
rect 4565 17179 4651 17415
rect 4887 17179 4973 17415
rect 5209 17179 5295 17415
rect 5531 17179 5617 17415
rect 5853 17179 5938 17415
rect 6174 17179 6259 17415
rect 6495 17179 6580 17415
rect 6816 17179 6901 17415
rect 7137 17179 7222 17415
rect 7458 17179 7543 17415
rect 7779 17179 7864 17415
rect 8100 17179 8185 17415
rect 8421 17179 8506 17415
rect 8742 17179 8827 17415
rect 9063 17179 9148 17415
rect 9384 17179 9469 17415
rect 9705 17179 9790 17415
rect 10026 17179 10111 17415
rect 10347 17179 10432 17415
rect 10668 17179 10753 17415
rect 10989 17179 11074 17415
rect 11310 17179 11395 17415
rect 11631 17179 11716 17415
rect 11952 17179 12037 17415
rect 12273 17179 12358 17415
rect 12594 17179 12679 17415
rect 12915 17179 13000 17415
rect 13236 17179 13321 17415
rect 13557 17179 13642 17415
rect 13878 17179 13963 17415
rect 14199 17179 14284 17415
rect 14520 17179 14605 17415
rect 14841 17179 15000 17415
rect 0 17079 15000 17179
rect 0 16843 143 17079
rect 379 16843 465 17079
rect 701 16843 787 17079
rect 1023 16843 1109 17079
rect 1345 16843 1431 17079
rect 1667 16843 1753 17079
rect 1989 16843 2075 17079
rect 2311 16843 2397 17079
rect 2633 16843 2719 17079
rect 2955 16843 3041 17079
rect 3277 16843 3363 17079
rect 3599 16843 3685 17079
rect 3921 16843 4007 17079
rect 4243 16843 4329 17079
rect 4565 16843 4651 17079
rect 4887 16843 4973 17079
rect 5209 16843 5295 17079
rect 5531 16843 5617 17079
rect 5853 16843 5938 17079
rect 6174 16843 6259 17079
rect 6495 16843 6580 17079
rect 6816 16843 6901 17079
rect 7137 16843 7222 17079
rect 7458 16843 7543 17079
rect 7779 16843 7864 17079
rect 8100 16843 8185 17079
rect 8421 16843 8506 17079
rect 8742 16843 8827 17079
rect 9063 16843 9148 17079
rect 9384 16843 9469 17079
rect 9705 16843 9790 17079
rect 10026 16843 10111 17079
rect 10347 16843 10432 17079
rect 10668 16843 10753 17079
rect 10989 16843 11074 17079
rect 11310 16843 11395 17079
rect 11631 16843 11716 17079
rect 11952 16843 12037 17079
rect 12273 16843 12358 17079
rect 12594 16843 12679 17079
rect 12915 16843 13000 17079
rect 13236 16843 13321 17079
rect 13557 16843 13642 17079
rect 13878 16843 13963 17079
rect 14199 16843 14284 17079
rect 14520 16843 14605 17079
rect 14841 16843 15000 17079
rect 0 16743 15000 16843
rect 0 16507 143 16743
rect 379 16507 465 16743
rect 701 16507 787 16743
rect 1023 16507 1109 16743
rect 1345 16507 1431 16743
rect 1667 16507 1753 16743
rect 1989 16507 2075 16743
rect 2311 16507 2397 16743
rect 2633 16507 2719 16743
rect 2955 16507 3041 16743
rect 3277 16507 3363 16743
rect 3599 16507 3685 16743
rect 3921 16507 4007 16743
rect 4243 16507 4329 16743
rect 4565 16507 4651 16743
rect 4887 16507 4973 16743
rect 5209 16507 5295 16743
rect 5531 16507 5617 16743
rect 5853 16507 5938 16743
rect 6174 16507 6259 16743
rect 6495 16507 6580 16743
rect 6816 16507 6901 16743
rect 7137 16507 7222 16743
rect 7458 16507 7543 16743
rect 7779 16507 7864 16743
rect 8100 16507 8185 16743
rect 8421 16507 8506 16743
rect 8742 16507 8827 16743
rect 9063 16507 9148 16743
rect 9384 16507 9469 16743
rect 9705 16507 9790 16743
rect 10026 16507 10111 16743
rect 10347 16507 10432 16743
rect 10668 16507 10753 16743
rect 10989 16507 11074 16743
rect 11310 16507 11395 16743
rect 11631 16507 11716 16743
rect 11952 16507 12037 16743
rect 12273 16507 12358 16743
rect 12594 16507 12679 16743
rect 12915 16507 13000 16743
rect 13236 16507 13321 16743
rect 13557 16507 13642 16743
rect 13878 16507 13963 16743
rect 14199 16507 14284 16743
rect 14520 16507 14605 16743
rect 14841 16507 15000 16743
rect 0 16407 15000 16507
rect 0 16171 143 16407
rect 379 16171 465 16407
rect 701 16171 787 16407
rect 1023 16171 1109 16407
rect 1345 16171 1431 16407
rect 1667 16171 1753 16407
rect 1989 16171 2075 16407
rect 2311 16171 2397 16407
rect 2633 16171 2719 16407
rect 2955 16171 3041 16407
rect 3277 16171 3363 16407
rect 3599 16171 3685 16407
rect 3921 16171 4007 16407
rect 4243 16171 4329 16407
rect 4565 16171 4651 16407
rect 4887 16171 4973 16407
rect 5209 16171 5295 16407
rect 5531 16171 5617 16407
rect 5853 16171 5938 16407
rect 6174 16171 6259 16407
rect 6495 16171 6580 16407
rect 6816 16171 6901 16407
rect 7137 16171 7222 16407
rect 7458 16171 7543 16407
rect 7779 16171 7864 16407
rect 8100 16171 8185 16407
rect 8421 16171 8506 16407
rect 8742 16171 8827 16407
rect 9063 16171 9148 16407
rect 9384 16171 9469 16407
rect 9705 16171 9790 16407
rect 10026 16171 10111 16407
rect 10347 16171 10432 16407
rect 10668 16171 10753 16407
rect 10989 16171 11074 16407
rect 11310 16171 11395 16407
rect 11631 16171 11716 16407
rect 11952 16171 12037 16407
rect 12273 16171 12358 16407
rect 12594 16171 12679 16407
rect 12915 16171 13000 16407
rect 13236 16171 13321 16407
rect 13557 16171 13642 16407
rect 13878 16171 13963 16407
rect 14199 16171 14284 16407
rect 14520 16171 14605 16407
rect 14841 16171 15000 16407
rect 0 16071 15000 16171
rect 0 15835 143 16071
rect 379 15835 465 16071
rect 701 15835 787 16071
rect 1023 15835 1109 16071
rect 1345 15835 1431 16071
rect 1667 15835 1753 16071
rect 1989 15835 2075 16071
rect 2311 15835 2397 16071
rect 2633 15835 2719 16071
rect 2955 15835 3041 16071
rect 3277 15835 3363 16071
rect 3599 15835 3685 16071
rect 3921 15835 4007 16071
rect 4243 15835 4329 16071
rect 4565 15835 4651 16071
rect 4887 15835 4973 16071
rect 5209 15835 5295 16071
rect 5531 15835 5617 16071
rect 5853 15835 5938 16071
rect 6174 15835 6259 16071
rect 6495 15835 6580 16071
rect 6816 15835 6901 16071
rect 7137 15835 7222 16071
rect 7458 15835 7543 16071
rect 7779 15835 7864 16071
rect 8100 15835 8185 16071
rect 8421 15835 8506 16071
rect 8742 15835 8827 16071
rect 9063 15835 9148 16071
rect 9384 15835 9469 16071
rect 9705 15835 9790 16071
rect 10026 15835 10111 16071
rect 10347 15835 10432 16071
rect 10668 15835 10753 16071
rect 10989 15835 11074 16071
rect 11310 15835 11395 16071
rect 11631 15835 11716 16071
rect 11952 15835 12037 16071
rect 12273 15835 12358 16071
rect 12594 15835 12679 16071
rect 12915 15835 13000 16071
rect 13236 15835 13321 16071
rect 13557 15835 13642 16071
rect 13878 15835 13963 16071
rect 14199 15835 14284 16071
rect 14520 15835 14605 16071
rect 14841 15835 15000 16071
rect 0 15735 15000 15835
rect 0 15499 143 15735
rect 379 15499 465 15735
rect 701 15499 787 15735
rect 1023 15499 1109 15735
rect 1345 15499 1431 15735
rect 1667 15499 1753 15735
rect 1989 15499 2075 15735
rect 2311 15499 2397 15735
rect 2633 15499 2719 15735
rect 2955 15499 3041 15735
rect 3277 15499 3363 15735
rect 3599 15499 3685 15735
rect 3921 15499 4007 15735
rect 4243 15499 4329 15735
rect 4565 15499 4651 15735
rect 4887 15499 4973 15735
rect 5209 15499 5295 15735
rect 5531 15499 5617 15735
rect 5853 15499 5938 15735
rect 6174 15499 6259 15735
rect 6495 15499 6580 15735
rect 6816 15499 6901 15735
rect 7137 15499 7222 15735
rect 7458 15499 7543 15735
rect 7779 15499 7864 15735
rect 8100 15499 8185 15735
rect 8421 15499 8506 15735
rect 8742 15499 8827 15735
rect 9063 15499 9148 15735
rect 9384 15499 9469 15735
rect 9705 15499 9790 15735
rect 10026 15499 10111 15735
rect 10347 15499 10432 15735
rect 10668 15499 10753 15735
rect 10989 15499 11074 15735
rect 11310 15499 11395 15735
rect 11631 15499 11716 15735
rect 11952 15499 12037 15735
rect 12273 15499 12358 15735
rect 12594 15499 12679 15735
rect 12915 15499 13000 15735
rect 13236 15499 13321 15735
rect 13557 15499 13642 15735
rect 13878 15499 13963 15735
rect 14199 15499 14284 15735
rect 14520 15499 14605 15735
rect 14841 15499 15000 15735
rect 0 15399 15000 15499
rect 0 15163 143 15399
rect 379 15163 465 15399
rect 701 15163 787 15399
rect 1023 15163 1109 15399
rect 1345 15163 1431 15399
rect 1667 15163 1753 15399
rect 1989 15163 2075 15399
rect 2311 15163 2397 15399
rect 2633 15163 2719 15399
rect 2955 15163 3041 15399
rect 3277 15163 3363 15399
rect 3599 15163 3685 15399
rect 3921 15163 4007 15399
rect 4243 15163 4329 15399
rect 4565 15163 4651 15399
rect 4887 15163 4973 15399
rect 5209 15163 5295 15399
rect 5531 15163 5617 15399
rect 5853 15163 5938 15399
rect 6174 15163 6259 15399
rect 6495 15163 6580 15399
rect 6816 15163 6901 15399
rect 7137 15163 7222 15399
rect 7458 15163 7543 15399
rect 7779 15163 7864 15399
rect 8100 15163 8185 15399
rect 8421 15163 8506 15399
rect 8742 15163 8827 15399
rect 9063 15163 9148 15399
rect 9384 15163 9469 15399
rect 9705 15163 9790 15399
rect 10026 15163 10111 15399
rect 10347 15163 10432 15399
rect 10668 15163 10753 15399
rect 10989 15163 11074 15399
rect 11310 15163 11395 15399
rect 11631 15163 11716 15399
rect 11952 15163 12037 15399
rect 12273 15163 12358 15399
rect 12594 15163 12679 15399
rect 12915 15163 13000 15399
rect 13236 15163 13321 15399
rect 13557 15163 13642 15399
rect 13878 15163 13963 15399
rect 14199 15163 14284 15399
rect 14520 15163 14605 15399
rect 14841 15163 15000 15399
rect 0 15063 15000 15163
rect 0 14827 143 15063
rect 379 14827 465 15063
rect 701 14827 787 15063
rect 1023 14827 1109 15063
rect 1345 14827 1431 15063
rect 1667 14827 1753 15063
rect 1989 14827 2075 15063
rect 2311 14827 2397 15063
rect 2633 14827 2719 15063
rect 2955 14827 3041 15063
rect 3277 14827 3363 15063
rect 3599 14827 3685 15063
rect 3921 14827 4007 15063
rect 4243 14827 4329 15063
rect 4565 14827 4651 15063
rect 4887 14827 4973 15063
rect 5209 14827 5295 15063
rect 5531 14827 5617 15063
rect 5853 14827 5938 15063
rect 6174 14827 6259 15063
rect 6495 14827 6580 15063
rect 6816 14827 6901 15063
rect 7137 14827 7222 15063
rect 7458 14827 7543 15063
rect 7779 14827 7864 15063
rect 8100 14827 8185 15063
rect 8421 14827 8506 15063
rect 8742 14827 8827 15063
rect 9063 14827 9148 15063
rect 9384 14827 9469 15063
rect 9705 14827 9790 15063
rect 10026 14827 10111 15063
rect 10347 14827 10432 15063
rect 10668 14827 10753 15063
rect 10989 14827 11074 15063
rect 11310 14827 11395 15063
rect 11631 14827 11716 15063
rect 11952 14827 12037 15063
rect 12273 14827 12358 15063
rect 12594 14827 12679 15063
rect 12915 14827 13000 15063
rect 13236 14827 13321 15063
rect 13557 14827 13642 15063
rect 13878 14827 13963 15063
rect 14199 14827 14284 15063
rect 14520 14827 14605 15063
rect 14841 14827 15000 15063
rect 0 14727 15000 14827
rect 0 14491 143 14727
rect 379 14491 465 14727
rect 701 14491 787 14727
rect 1023 14491 1109 14727
rect 1345 14491 1431 14727
rect 1667 14491 1753 14727
rect 1989 14491 2075 14727
rect 2311 14491 2397 14727
rect 2633 14491 2719 14727
rect 2955 14491 3041 14727
rect 3277 14491 3363 14727
rect 3599 14491 3685 14727
rect 3921 14491 4007 14727
rect 4243 14491 4329 14727
rect 4565 14491 4651 14727
rect 4887 14491 4973 14727
rect 5209 14491 5295 14727
rect 5531 14491 5617 14727
rect 5853 14491 5938 14727
rect 6174 14491 6259 14727
rect 6495 14491 6580 14727
rect 6816 14491 6901 14727
rect 7137 14491 7222 14727
rect 7458 14491 7543 14727
rect 7779 14491 7864 14727
rect 8100 14491 8185 14727
rect 8421 14491 8506 14727
rect 8742 14491 8827 14727
rect 9063 14491 9148 14727
rect 9384 14491 9469 14727
rect 9705 14491 9790 14727
rect 10026 14491 10111 14727
rect 10347 14491 10432 14727
rect 10668 14491 10753 14727
rect 10989 14491 11074 14727
rect 11310 14491 11395 14727
rect 11631 14491 11716 14727
rect 11952 14491 12037 14727
rect 12273 14491 12358 14727
rect 12594 14491 12679 14727
rect 12915 14491 13000 14727
rect 13236 14491 13321 14727
rect 13557 14491 13642 14727
rect 13878 14491 13963 14727
rect 14199 14491 14284 14727
rect 14520 14491 14605 14727
rect 14841 14491 15000 14727
rect 0 14391 15000 14491
rect 0 14155 143 14391
rect 379 14155 465 14391
rect 701 14155 787 14391
rect 1023 14155 1109 14391
rect 1345 14155 1431 14391
rect 1667 14155 1753 14391
rect 1989 14155 2075 14391
rect 2311 14155 2397 14391
rect 2633 14155 2719 14391
rect 2955 14155 3041 14391
rect 3277 14155 3363 14391
rect 3599 14155 3685 14391
rect 3921 14155 4007 14391
rect 4243 14155 4329 14391
rect 4565 14155 4651 14391
rect 4887 14155 4973 14391
rect 5209 14155 5295 14391
rect 5531 14155 5617 14391
rect 5853 14155 5938 14391
rect 6174 14155 6259 14391
rect 6495 14155 6580 14391
rect 6816 14155 6901 14391
rect 7137 14155 7222 14391
rect 7458 14155 7543 14391
rect 7779 14155 7864 14391
rect 8100 14155 8185 14391
rect 8421 14155 8506 14391
rect 8742 14155 8827 14391
rect 9063 14155 9148 14391
rect 9384 14155 9469 14391
rect 9705 14155 9790 14391
rect 10026 14155 10111 14391
rect 10347 14155 10432 14391
rect 10668 14155 10753 14391
rect 10989 14155 11074 14391
rect 11310 14155 11395 14391
rect 11631 14155 11716 14391
rect 11952 14155 12037 14391
rect 12273 14155 12358 14391
rect 12594 14155 12679 14391
rect 12915 14155 13000 14391
rect 13236 14155 13321 14391
rect 13557 14155 13642 14391
rect 13878 14155 13963 14391
rect 14199 14155 14284 14391
rect 14520 14155 14605 14391
rect 14841 14155 15000 14391
rect 0 14055 15000 14155
rect 0 13819 143 14055
rect 379 13819 465 14055
rect 701 13819 787 14055
rect 1023 13819 1109 14055
rect 1345 13819 1431 14055
rect 1667 13819 1753 14055
rect 1989 13819 2075 14055
rect 2311 13819 2397 14055
rect 2633 13819 2719 14055
rect 2955 13819 3041 14055
rect 3277 13819 3363 14055
rect 3599 13819 3685 14055
rect 3921 13819 4007 14055
rect 4243 13819 4329 14055
rect 4565 13819 4651 14055
rect 4887 13819 4973 14055
rect 5209 13819 5295 14055
rect 5531 13819 5617 14055
rect 5853 13819 5938 14055
rect 6174 13819 6259 14055
rect 6495 13819 6580 14055
rect 6816 13819 6901 14055
rect 7137 13819 7222 14055
rect 7458 13819 7543 14055
rect 7779 13819 7864 14055
rect 8100 13819 8185 14055
rect 8421 13819 8506 14055
rect 8742 13819 8827 14055
rect 9063 13819 9148 14055
rect 9384 13819 9469 14055
rect 9705 13819 9790 14055
rect 10026 13819 10111 14055
rect 10347 13819 10432 14055
rect 10668 13819 10753 14055
rect 10989 13819 11074 14055
rect 11310 13819 11395 14055
rect 11631 13819 11716 14055
rect 11952 13819 12037 14055
rect 12273 13819 12358 14055
rect 12594 13819 12679 14055
rect 12915 13819 13000 14055
rect 13236 13819 13321 14055
rect 13557 13819 13642 14055
rect 13878 13819 13963 14055
rect 14199 13819 14284 14055
rect 14520 13819 14605 14055
rect 14841 13819 15000 14055
rect 0 13719 15000 13819
rect 0 13483 143 13719
rect 379 13483 465 13719
rect 701 13483 787 13719
rect 1023 13483 1109 13719
rect 1345 13483 1431 13719
rect 1667 13483 1753 13719
rect 1989 13483 2075 13719
rect 2311 13483 2397 13719
rect 2633 13483 2719 13719
rect 2955 13483 3041 13719
rect 3277 13483 3363 13719
rect 3599 13483 3685 13719
rect 3921 13483 4007 13719
rect 4243 13483 4329 13719
rect 4565 13483 4651 13719
rect 4887 13483 4973 13719
rect 5209 13483 5295 13719
rect 5531 13483 5617 13719
rect 5853 13483 5938 13719
rect 6174 13483 6259 13719
rect 6495 13483 6580 13719
rect 6816 13483 6901 13719
rect 7137 13483 7222 13719
rect 7458 13483 7543 13719
rect 7779 13483 7864 13719
rect 8100 13483 8185 13719
rect 8421 13483 8506 13719
rect 8742 13483 8827 13719
rect 9063 13483 9148 13719
rect 9384 13483 9469 13719
rect 9705 13483 9790 13719
rect 10026 13483 10111 13719
rect 10347 13483 10432 13719
rect 10668 13483 10753 13719
rect 10989 13483 11074 13719
rect 11310 13483 11395 13719
rect 11631 13483 11716 13719
rect 11952 13483 12037 13719
rect 12273 13483 12358 13719
rect 12594 13483 12679 13719
rect 12915 13483 13000 13719
rect 13236 13483 13321 13719
rect 13557 13483 13642 13719
rect 13878 13483 13963 13719
rect 14199 13483 14284 13719
rect 14520 13483 14605 13719
rect 14841 13483 15000 13719
rect 0 13482 15000 13483
rect 0 13458 254 13482
rect 14746 13458 15000 13482
rect 0 13114 254 13158
rect 14746 13114 15000 13158
rect 0 12878 143 13114
rect 379 12878 465 13114
rect 701 12878 787 13114
rect 1023 12878 1109 13114
rect 1345 12878 1431 13114
rect 1667 12878 1753 13114
rect 1989 12878 2075 13114
rect 2311 12878 2397 13114
rect 2633 12878 2719 13114
rect 2955 12878 3041 13114
rect 3277 12878 3363 13114
rect 3599 12878 3685 13114
rect 3921 12878 4007 13114
rect 4243 12878 4329 13114
rect 4565 12878 4651 13114
rect 4887 12878 4973 13114
rect 5209 12878 5294 13114
rect 5530 12878 5615 13114
rect 5851 12878 5936 13114
rect 6172 12878 6257 13114
rect 6493 12878 6578 13114
rect 6814 12878 6899 13114
rect 7135 12878 7220 13114
rect 7456 12878 7541 13114
rect 7777 12878 7862 13114
rect 8098 12878 8183 13114
rect 8419 12878 8504 13114
rect 8740 12878 8825 13114
rect 9061 12878 9146 13114
rect 9382 12878 9467 13114
rect 9703 12878 9788 13114
rect 10024 12878 10109 13114
rect 10345 12878 10430 13114
rect 10666 12878 10751 13114
rect 10987 12878 11072 13114
rect 11308 12878 11393 13114
rect 11629 12878 11714 13114
rect 11950 12878 12035 13114
rect 12271 12878 12356 13114
rect 12592 12878 12677 13114
rect 12913 12878 12998 13114
rect 13234 12878 13319 13114
rect 13555 12878 13640 13114
rect 13876 12878 13961 13114
rect 14197 12878 14282 13114
rect 14518 12878 14603 13114
rect 14839 12878 15000 13114
rect 0 12548 15000 12878
rect 0 12312 143 12548
rect 379 12312 465 12548
rect 701 12312 787 12548
rect 1023 12312 1109 12548
rect 1345 12312 1431 12548
rect 1667 12312 1753 12548
rect 1989 12312 2075 12548
rect 2311 12312 2397 12548
rect 2633 12312 2719 12548
rect 2955 12312 3041 12548
rect 3277 12312 3363 12548
rect 3599 12312 3685 12548
rect 3921 12312 4007 12548
rect 4243 12312 4329 12548
rect 4565 12312 4651 12548
rect 4887 12312 4973 12548
rect 5209 12312 5294 12548
rect 5530 12312 5615 12548
rect 5851 12312 5936 12548
rect 6172 12312 6257 12548
rect 6493 12312 6578 12548
rect 6814 12312 6899 12548
rect 7135 12312 7220 12548
rect 7456 12312 7541 12548
rect 7777 12312 7862 12548
rect 8098 12312 8183 12548
rect 8419 12312 8504 12548
rect 8740 12312 8825 12548
rect 9061 12312 9146 12548
rect 9382 12312 9467 12548
rect 9703 12312 9788 12548
rect 10024 12312 10109 12548
rect 10345 12312 10430 12548
rect 10666 12312 10751 12548
rect 10987 12312 11072 12548
rect 11308 12312 11393 12548
rect 11629 12312 11714 12548
rect 11950 12312 12035 12548
rect 12271 12312 12356 12548
rect 12592 12312 12677 12548
rect 12913 12312 12998 12548
rect 13234 12312 13319 12548
rect 13555 12312 13640 12548
rect 13876 12312 13961 12548
rect 14197 12312 14282 12548
rect 14518 12312 14603 12548
rect 14839 12312 15000 12548
rect 0 12268 254 12312
rect 14746 12268 15000 12312
rect 0 11944 254 11988
rect 14746 11944 15000 11988
rect 0 11708 143 11944
rect 379 11708 465 11944
rect 701 11708 787 11944
rect 1023 11708 1109 11944
rect 1345 11708 1431 11944
rect 1667 11708 1753 11944
rect 1989 11708 2075 11944
rect 2311 11708 2397 11944
rect 2633 11708 2719 11944
rect 2955 11708 3041 11944
rect 3277 11708 3363 11944
rect 3599 11708 3685 11944
rect 3921 11708 4007 11944
rect 4243 11708 4329 11944
rect 4565 11708 4651 11944
rect 4887 11708 4973 11944
rect 5209 11708 5294 11944
rect 5530 11708 5615 11944
rect 5851 11708 5936 11944
rect 6172 11708 6257 11944
rect 6493 11708 6578 11944
rect 6814 11708 6899 11944
rect 7135 11708 7220 11944
rect 7456 11708 7541 11944
rect 7777 11708 7862 11944
rect 8098 11708 8183 11944
rect 8419 11708 8504 11944
rect 8740 11708 8825 11944
rect 9061 11708 9146 11944
rect 9382 11708 9467 11944
rect 9703 11708 9788 11944
rect 10024 11708 10109 11944
rect 10345 11708 10430 11944
rect 10666 11708 10751 11944
rect 10987 11708 11072 11944
rect 11308 11708 11393 11944
rect 11629 11708 11714 11944
rect 11950 11708 12035 11944
rect 12271 11708 12356 11944
rect 12592 11708 12677 11944
rect 12913 11708 12998 11944
rect 13234 11708 13319 11944
rect 13555 11708 13640 11944
rect 13876 11708 13961 11944
rect 14197 11708 14282 11944
rect 14518 11708 14603 11944
rect 14839 11708 15000 11944
rect 0 11378 15000 11708
rect 0 11142 143 11378
rect 379 11142 465 11378
rect 701 11142 787 11378
rect 1023 11142 1109 11378
rect 1345 11142 1431 11378
rect 1667 11142 1753 11378
rect 1989 11142 2075 11378
rect 2311 11142 2397 11378
rect 2633 11142 2719 11378
rect 2955 11142 3041 11378
rect 3277 11142 3363 11378
rect 3599 11142 3685 11378
rect 3921 11142 4007 11378
rect 4243 11142 4329 11378
rect 4565 11142 4651 11378
rect 4887 11142 4973 11378
rect 5209 11142 5294 11378
rect 5530 11142 5615 11378
rect 5851 11142 5936 11378
rect 6172 11142 6257 11378
rect 6493 11142 6578 11378
rect 6814 11142 6899 11378
rect 7135 11142 7220 11378
rect 7456 11142 7541 11378
rect 7777 11142 7862 11378
rect 8098 11142 8183 11378
rect 8419 11142 8504 11378
rect 8740 11142 8825 11378
rect 9061 11142 9146 11378
rect 9382 11142 9467 11378
rect 9703 11142 9788 11378
rect 10024 11142 10109 11378
rect 10345 11142 10430 11378
rect 10666 11142 10751 11378
rect 10987 11142 11072 11378
rect 11308 11142 11393 11378
rect 11629 11142 11714 11378
rect 11950 11142 12035 11378
rect 12271 11142 12356 11378
rect 12592 11142 12677 11378
rect 12913 11142 12998 11378
rect 13234 11142 13319 11378
rect 13555 11142 13640 11378
rect 13876 11142 13961 11378
rect 14197 11142 14282 11378
rect 14518 11142 14603 11378
rect 14839 11142 15000 11378
rect 0 11098 254 11142
rect 14746 11098 15000 11142
rect 0 10732 254 10798
rect 14746 10732 15000 10798
rect 0 10076 254 10672
rect 14746 10076 15000 10672
rect 0 9780 254 10016
rect 14746 9780 15000 10016
rect 0 9124 254 9720
rect 14746 9124 15000 9720
rect 0 8998 254 9064
rect 14746 8998 15000 9064
rect 0 8654 254 8698
rect 14746 8654 15000 8698
rect 0 8418 143 8654
rect 379 8418 465 8654
rect 701 8418 787 8654
rect 1023 8418 1109 8654
rect 1345 8418 1431 8654
rect 1667 8418 1753 8654
rect 1989 8418 2075 8654
rect 2311 8418 2397 8654
rect 2633 8418 2719 8654
rect 2955 8418 3041 8654
rect 3277 8418 3363 8654
rect 3599 8418 3685 8654
rect 3921 8418 4007 8654
rect 4243 8418 4329 8654
rect 4565 8418 4651 8654
rect 4887 8418 4973 8654
rect 5209 8418 5295 8654
rect 5531 8418 5617 8654
rect 5853 8418 5938 8654
rect 6174 8418 6259 8654
rect 6495 8418 6580 8654
rect 6816 8418 6901 8654
rect 7137 8418 7222 8654
rect 7458 8418 7543 8654
rect 7779 8418 7864 8654
rect 8100 8418 8185 8654
rect 8421 8418 8506 8654
rect 8742 8418 8827 8654
rect 9063 8418 9148 8654
rect 9384 8418 9469 8654
rect 9705 8418 9790 8654
rect 10026 8418 10111 8654
rect 10347 8418 10432 8654
rect 10668 8418 10753 8654
rect 10989 8418 11074 8654
rect 11310 8418 11395 8654
rect 11631 8418 11716 8654
rect 11952 8418 12037 8654
rect 12273 8418 12358 8654
rect 12594 8418 12679 8654
rect 12915 8418 13000 8654
rect 13236 8418 13321 8654
rect 13557 8418 13642 8654
rect 13878 8418 13963 8654
rect 14199 8418 14284 8654
rect 14520 8418 14605 8654
rect 14841 8418 15000 8654
rect 0 8048 15000 8418
rect 0 7812 143 8048
rect 379 7812 465 8048
rect 701 7812 787 8048
rect 1023 7812 1109 8048
rect 1345 7812 1431 8048
rect 1667 7812 1753 8048
rect 1989 7812 2075 8048
rect 2311 7812 2397 8048
rect 2633 7812 2719 8048
rect 2955 7812 3041 8048
rect 3277 7812 3363 8048
rect 3599 7812 3685 8048
rect 3921 7812 4007 8048
rect 4243 7812 4329 8048
rect 4565 7812 4651 8048
rect 4887 7812 4973 8048
rect 5209 7812 5295 8048
rect 5531 7812 5617 8048
rect 5853 7812 5938 8048
rect 6174 7812 6259 8048
rect 6495 7812 6580 8048
rect 6816 7812 6901 8048
rect 7137 7812 7222 8048
rect 7458 7812 7543 8048
rect 7779 7812 7864 8048
rect 8100 7812 8185 8048
rect 8421 7812 8506 8048
rect 8742 7812 8827 8048
rect 9063 7812 9148 8048
rect 9384 7812 9469 8048
rect 9705 7812 9790 8048
rect 10026 7812 10111 8048
rect 10347 7812 10432 8048
rect 10668 7812 10753 8048
rect 10989 7812 11074 8048
rect 11310 7812 11395 8048
rect 11631 7812 11716 8048
rect 11952 7812 12037 8048
rect 12273 7812 12358 8048
rect 12594 7812 12679 8048
rect 12915 7812 13000 8048
rect 13236 7812 13321 8048
rect 13557 7812 13642 8048
rect 13878 7812 13963 8048
rect 14199 7812 14284 8048
rect 14520 7812 14605 8048
rect 14841 7812 15000 8048
rect 0 7768 254 7812
rect 14746 7768 15000 7812
rect 0 7444 254 7488
rect 14746 7444 15000 7488
rect 0 7208 143 7444
rect 379 7208 465 7444
rect 701 7208 787 7444
rect 1023 7208 1109 7444
rect 1345 7208 1431 7444
rect 1667 7208 1753 7444
rect 1989 7208 2075 7444
rect 2311 7208 2397 7444
rect 2633 7208 2719 7444
rect 2955 7208 3041 7444
rect 3277 7208 3363 7444
rect 3599 7208 3685 7444
rect 3921 7208 4007 7444
rect 4243 7208 4329 7444
rect 4565 7208 4651 7444
rect 4887 7208 4973 7444
rect 5209 7208 5295 7444
rect 5531 7208 5617 7444
rect 5853 7208 5938 7444
rect 6174 7208 6259 7444
rect 6495 7208 6580 7444
rect 6816 7208 6901 7444
rect 7137 7208 7222 7444
rect 7458 7208 7543 7444
rect 7779 7208 7864 7444
rect 8100 7208 8185 7444
rect 8421 7208 8506 7444
rect 8742 7208 8827 7444
rect 9063 7208 9148 7444
rect 9384 7208 9469 7444
rect 9705 7208 9790 7444
rect 10026 7208 10111 7444
rect 10347 7208 10432 7444
rect 10668 7208 10753 7444
rect 10989 7208 11074 7444
rect 11310 7208 11395 7444
rect 11631 7208 11716 7444
rect 11952 7208 12037 7444
rect 12273 7208 12358 7444
rect 12594 7208 12679 7444
rect 12915 7208 13000 7444
rect 13236 7208 13321 7444
rect 13557 7208 13642 7444
rect 13878 7208 13963 7444
rect 14199 7208 14284 7444
rect 14520 7208 14605 7444
rect 14841 7208 15000 7444
rect 0 7078 15000 7208
rect 0 6842 143 7078
rect 379 6842 465 7078
rect 701 6842 787 7078
rect 1023 6842 1109 7078
rect 1345 6842 1431 7078
rect 1667 6842 1753 7078
rect 1989 6842 2075 7078
rect 2311 6842 2397 7078
rect 2633 6842 2719 7078
rect 2955 6842 3041 7078
rect 3277 6842 3363 7078
rect 3599 6842 3685 7078
rect 3921 6842 4007 7078
rect 4243 6842 4329 7078
rect 4565 6842 4651 7078
rect 4887 6842 4973 7078
rect 5209 6842 5295 7078
rect 5531 6842 5617 7078
rect 5853 6842 5938 7078
rect 6174 6842 6259 7078
rect 6495 6842 6580 7078
rect 6816 6842 6901 7078
rect 7137 6842 7222 7078
rect 7458 6842 7543 7078
rect 7779 6842 7864 7078
rect 8100 6842 8185 7078
rect 8421 6842 8506 7078
rect 8742 6842 8827 7078
rect 9063 6842 9148 7078
rect 9384 6842 9469 7078
rect 9705 6842 9790 7078
rect 10026 6842 10111 7078
rect 10347 6842 10432 7078
rect 10668 6842 10753 7078
rect 10989 6842 11074 7078
rect 11310 6842 11395 7078
rect 11631 6842 11716 7078
rect 11952 6842 12037 7078
rect 12273 6842 12358 7078
rect 12594 6842 12679 7078
rect 12915 6842 13000 7078
rect 13236 6842 13321 7078
rect 13557 6842 13642 7078
rect 13878 6842 13963 7078
rect 14199 6842 14284 7078
rect 14520 6842 14605 7078
rect 14841 6842 15000 7078
rect 0 6798 254 6842
rect 14746 6798 15000 6842
rect 0 6474 254 6518
rect 14746 6474 15000 6518
rect 0 6238 143 6474
rect 379 6238 465 6474
rect 701 6238 787 6474
rect 1023 6238 1109 6474
rect 1345 6238 1431 6474
rect 1667 6238 1753 6474
rect 1989 6238 2075 6474
rect 2311 6238 2397 6474
rect 2633 6238 2719 6474
rect 2955 6238 3041 6474
rect 3277 6238 3363 6474
rect 3599 6238 3685 6474
rect 3921 6238 4007 6474
rect 4243 6238 4329 6474
rect 4565 6238 4651 6474
rect 4887 6238 4973 6474
rect 5209 6238 5295 6474
rect 5531 6238 5617 6474
rect 5853 6238 5938 6474
rect 6174 6238 6259 6474
rect 6495 6238 6580 6474
rect 6816 6238 6901 6474
rect 7137 6238 7222 6474
rect 7458 6238 7543 6474
rect 7779 6238 7864 6474
rect 8100 6238 8185 6474
rect 8421 6238 8506 6474
rect 8742 6238 8827 6474
rect 9063 6238 9148 6474
rect 9384 6238 9469 6474
rect 9705 6238 9790 6474
rect 10026 6238 10111 6474
rect 10347 6238 10432 6474
rect 10668 6238 10753 6474
rect 10989 6238 11074 6474
rect 11310 6238 11395 6474
rect 11631 6238 11716 6474
rect 11952 6238 12037 6474
rect 12273 6238 12358 6474
rect 12594 6238 12679 6474
rect 12915 6238 13000 6474
rect 13236 6238 13321 6474
rect 13557 6238 13642 6474
rect 13878 6238 13963 6474
rect 14199 6238 14284 6474
rect 14520 6238 14605 6474
rect 14841 6238 15000 6474
rect 0 6108 15000 6238
rect 0 5872 143 6108
rect 379 5872 465 6108
rect 701 5872 787 6108
rect 1023 5872 1109 6108
rect 1345 5872 1431 6108
rect 1667 5872 1753 6108
rect 1989 5872 2075 6108
rect 2311 5872 2397 6108
rect 2633 5872 2719 6108
rect 2955 5872 3041 6108
rect 3277 5872 3363 6108
rect 3599 5872 3685 6108
rect 3921 5872 4007 6108
rect 4243 5872 4329 6108
rect 4565 5872 4651 6108
rect 4887 5872 4973 6108
rect 5209 5872 5295 6108
rect 5531 5872 5617 6108
rect 5853 5872 5938 6108
rect 6174 5872 6259 6108
rect 6495 5872 6580 6108
rect 6816 5872 6901 6108
rect 7137 5872 7222 6108
rect 7458 5872 7543 6108
rect 7779 5872 7864 6108
rect 8100 5872 8185 6108
rect 8421 5872 8506 6108
rect 8742 5872 8827 6108
rect 9063 5872 9148 6108
rect 9384 5872 9469 6108
rect 9705 5872 9790 6108
rect 10026 5872 10111 6108
rect 10347 5872 10432 6108
rect 10668 5872 10753 6108
rect 10989 5872 11074 6108
rect 11310 5872 11395 6108
rect 11631 5872 11716 6108
rect 11952 5872 12037 6108
rect 12273 5872 12358 6108
rect 12594 5872 12679 6108
rect 12915 5872 13000 6108
rect 13236 5872 13321 6108
rect 13557 5872 13642 6108
rect 13878 5872 13963 6108
rect 14199 5872 14284 6108
rect 14520 5872 14605 6108
rect 14841 5872 15000 6108
rect 0 5828 254 5872
rect 14746 5828 15000 5872
rect 0 5504 254 5548
rect 14746 5504 15000 5548
rect 0 5268 143 5504
rect 379 5268 465 5504
rect 701 5268 787 5504
rect 1023 5268 1109 5504
rect 1345 5268 1431 5504
rect 1667 5268 1753 5504
rect 1989 5268 2075 5504
rect 2311 5268 2397 5504
rect 2633 5268 2719 5504
rect 2955 5268 3041 5504
rect 3277 5268 3363 5504
rect 3599 5268 3685 5504
rect 3921 5268 4007 5504
rect 4243 5268 4329 5504
rect 4565 5268 4651 5504
rect 4887 5268 4973 5504
rect 5209 5268 5295 5504
rect 5531 5268 5617 5504
rect 5853 5268 5938 5504
rect 6174 5268 6259 5504
rect 6495 5268 6580 5504
rect 6816 5268 6901 5504
rect 7137 5268 7222 5504
rect 7458 5268 7543 5504
rect 7779 5268 7864 5504
rect 8100 5268 8185 5504
rect 8421 5268 8506 5504
rect 8742 5268 8827 5504
rect 9063 5268 9148 5504
rect 9384 5268 9469 5504
rect 9705 5268 9790 5504
rect 10026 5268 10111 5504
rect 10347 5268 10432 5504
rect 10668 5268 10753 5504
rect 10989 5268 11074 5504
rect 11310 5268 11395 5504
rect 11631 5268 11716 5504
rect 11952 5268 12037 5504
rect 12273 5268 12358 5504
rect 12594 5268 12679 5504
rect 12915 5268 13000 5504
rect 13236 5268 13321 5504
rect 13557 5268 13642 5504
rect 13878 5268 13963 5504
rect 14199 5268 14284 5504
rect 14520 5268 14605 5504
rect 14841 5268 15000 5504
rect 0 4898 15000 5268
rect 0 4662 143 4898
rect 379 4662 465 4898
rect 701 4662 787 4898
rect 1023 4662 1109 4898
rect 1345 4662 1431 4898
rect 1667 4662 1753 4898
rect 1989 4662 2075 4898
rect 2311 4662 2397 4898
rect 2633 4662 2719 4898
rect 2955 4662 3041 4898
rect 3277 4662 3363 4898
rect 3599 4662 3685 4898
rect 3921 4662 4007 4898
rect 4243 4662 4329 4898
rect 4565 4662 4651 4898
rect 4887 4662 4973 4898
rect 5209 4662 5295 4898
rect 5531 4662 5617 4898
rect 5853 4662 5938 4898
rect 6174 4662 6259 4898
rect 6495 4662 6580 4898
rect 6816 4662 6901 4898
rect 7137 4662 7222 4898
rect 7458 4662 7543 4898
rect 7779 4662 7864 4898
rect 8100 4662 8185 4898
rect 8421 4662 8506 4898
rect 8742 4662 8827 4898
rect 9063 4662 9148 4898
rect 9384 4662 9469 4898
rect 9705 4662 9790 4898
rect 10026 4662 10111 4898
rect 10347 4662 10432 4898
rect 10668 4662 10753 4898
rect 10989 4662 11074 4898
rect 11310 4662 11395 4898
rect 11631 4662 11716 4898
rect 11952 4662 12037 4898
rect 12273 4662 12358 4898
rect 12594 4662 12679 4898
rect 12915 4662 13000 4898
rect 13236 4662 13321 4898
rect 13557 4662 13642 4898
rect 13878 4662 13963 4898
rect 14199 4662 14284 4898
rect 14520 4662 14605 4898
rect 14841 4662 15000 4898
rect 0 4618 254 4662
rect 14746 4618 15000 4662
rect 0 4294 254 4338
rect 14746 4294 15000 4338
rect 0 4058 143 4294
rect 379 4058 465 4294
rect 701 4058 787 4294
rect 1023 4058 1109 4294
rect 1345 4058 1431 4294
rect 1667 4058 1753 4294
rect 1989 4058 2075 4294
rect 2311 4058 2397 4294
rect 2633 4058 2719 4294
rect 2955 4058 3041 4294
rect 3277 4058 3363 4294
rect 3599 4058 3685 4294
rect 3921 4058 4007 4294
rect 4243 4058 4329 4294
rect 4565 4058 4651 4294
rect 4887 4058 4973 4294
rect 5209 4058 5295 4294
rect 5531 4058 5617 4294
rect 5853 4058 5938 4294
rect 6174 4058 6259 4294
rect 6495 4058 6580 4294
rect 6816 4058 6901 4294
rect 7137 4058 7222 4294
rect 7458 4058 7543 4294
rect 7779 4058 7864 4294
rect 8100 4058 8185 4294
rect 8421 4058 8506 4294
rect 8742 4058 8827 4294
rect 9063 4058 9148 4294
rect 9384 4058 9469 4294
rect 9705 4058 9790 4294
rect 10026 4058 10111 4294
rect 10347 4058 10432 4294
rect 10668 4058 10753 4294
rect 10989 4058 11074 4294
rect 11310 4058 11395 4294
rect 11631 4058 11716 4294
rect 11952 4058 12037 4294
rect 12273 4058 12358 4294
rect 12594 4058 12679 4294
rect 12915 4058 13000 4294
rect 13236 4058 13321 4294
rect 13557 4058 13642 4294
rect 13878 4058 13963 4294
rect 14199 4058 14284 4294
rect 14520 4058 14605 4294
rect 14841 4058 15000 4294
rect 0 3688 15000 4058
rect 0 3452 143 3688
rect 379 3452 465 3688
rect 701 3452 787 3688
rect 1023 3452 1109 3688
rect 1345 3452 1431 3688
rect 1667 3452 1753 3688
rect 1989 3452 2075 3688
rect 2311 3452 2397 3688
rect 2633 3452 2719 3688
rect 2955 3452 3041 3688
rect 3277 3452 3363 3688
rect 3599 3452 3685 3688
rect 3921 3452 4007 3688
rect 4243 3452 4329 3688
rect 4565 3452 4651 3688
rect 4887 3452 4973 3688
rect 5209 3452 5295 3688
rect 5531 3452 5617 3688
rect 5853 3452 5938 3688
rect 6174 3452 6259 3688
rect 6495 3452 6580 3688
rect 6816 3452 6901 3688
rect 7137 3452 7222 3688
rect 7458 3452 7543 3688
rect 7779 3452 7864 3688
rect 8100 3452 8185 3688
rect 8421 3452 8506 3688
rect 8742 3452 8827 3688
rect 9063 3452 9148 3688
rect 9384 3452 9469 3688
rect 9705 3452 9790 3688
rect 10026 3452 10111 3688
rect 10347 3452 10432 3688
rect 10668 3452 10753 3688
rect 10989 3452 11074 3688
rect 11310 3452 11395 3688
rect 11631 3452 11716 3688
rect 11952 3452 12037 3688
rect 12273 3452 12358 3688
rect 12594 3452 12679 3688
rect 12915 3452 13000 3688
rect 13236 3452 13321 3688
rect 13557 3452 13642 3688
rect 13878 3452 13963 3688
rect 14199 3452 14284 3688
rect 14520 3452 14605 3688
rect 14841 3452 15000 3688
rect 0 3408 254 3452
rect 14746 3408 15000 3452
rect 0 3084 193 3128
rect 14807 3084 15000 3128
rect 0 2848 143 3084
rect 379 2848 465 3084
rect 701 2848 787 3084
rect 1023 2848 1109 3084
rect 1345 2848 1431 3084
rect 1667 2848 1753 3084
rect 1989 2848 2075 3084
rect 2311 2848 2397 3084
rect 2633 2848 2719 3084
rect 2955 2848 3041 3084
rect 3277 2848 3363 3084
rect 3599 2848 3685 3084
rect 3921 2848 4007 3084
rect 4243 2848 4329 3084
rect 4565 2848 4651 3084
rect 4887 2848 4973 3084
rect 5209 2848 5295 3084
rect 5531 2848 5617 3084
rect 5853 2848 5938 3084
rect 6174 2848 6259 3084
rect 6495 2848 6580 3084
rect 6816 2848 6901 3084
rect 7137 2848 7222 3084
rect 7458 2848 7543 3084
rect 7779 2848 7864 3084
rect 8100 2848 8185 3084
rect 8421 2848 8506 3084
rect 8742 2848 8827 3084
rect 9063 2848 9148 3084
rect 9384 2848 9469 3084
rect 9705 2848 9790 3084
rect 10026 2848 10111 3084
rect 10347 2848 10432 3084
rect 10668 2848 10753 3084
rect 10989 2848 11074 3084
rect 11310 2848 11395 3084
rect 11631 2848 11716 3084
rect 11952 2848 12037 3084
rect 12273 2848 12358 3084
rect 12594 2848 12679 3084
rect 12915 2848 13000 3084
rect 13236 2848 13321 3084
rect 13557 2848 13642 3084
rect 13878 2848 13963 3084
rect 14199 2848 14284 3084
rect 14520 2848 14605 3084
rect 14841 2848 15000 3084
rect 0 2718 15000 2848
rect 0 2482 143 2718
rect 379 2482 465 2718
rect 701 2482 787 2718
rect 1023 2482 1109 2718
rect 1345 2482 1431 2718
rect 1667 2482 1753 2718
rect 1989 2482 2075 2718
rect 2311 2482 2397 2718
rect 2633 2482 2719 2718
rect 2955 2482 3041 2718
rect 3277 2482 3363 2718
rect 3599 2482 3685 2718
rect 3921 2482 4007 2718
rect 4243 2482 4329 2718
rect 4565 2482 4651 2718
rect 4887 2482 4973 2718
rect 5209 2482 5295 2718
rect 5531 2482 5617 2718
rect 5853 2482 5938 2718
rect 6174 2482 6259 2718
rect 6495 2482 6580 2718
rect 6816 2482 6901 2718
rect 7137 2482 7222 2718
rect 7458 2482 7543 2718
rect 7779 2482 7864 2718
rect 8100 2482 8185 2718
rect 8421 2482 8506 2718
rect 8742 2482 8827 2718
rect 9063 2482 9148 2718
rect 9384 2482 9469 2718
rect 9705 2482 9790 2718
rect 10026 2482 10111 2718
rect 10347 2482 10432 2718
rect 10668 2482 10753 2718
rect 10989 2482 11074 2718
rect 11310 2482 11395 2718
rect 11631 2482 11716 2718
rect 11952 2482 12037 2718
rect 12273 2482 12358 2718
rect 12594 2482 12679 2718
rect 12915 2482 13000 2718
rect 13236 2482 13321 2718
rect 13557 2482 13642 2718
rect 13878 2482 13963 2718
rect 14199 2482 14284 2718
rect 14520 2482 14605 2718
rect 14841 2482 15000 2718
rect 0 2438 193 2482
rect 14807 2438 15000 2482
rect 0 2114 254 2158
rect 14746 2114 15000 2158
rect 0 1878 143 2114
rect 379 1878 465 2114
rect 701 1878 787 2114
rect 1023 1878 1109 2114
rect 1345 1878 1431 2114
rect 1667 1878 1753 2114
rect 1989 1878 2075 2114
rect 2311 1878 2397 2114
rect 2633 1878 2719 2114
rect 2955 1878 3041 2114
rect 3277 1878 3363 2114
rect 3599 1878 3685 2114
rect 3921 1878 4007 2114
rect 4243 1878 4329 2114
rect 4565 1878 4651 2114
rect 4887 1878 4973 2114
rect 5209 1878 5295 2114
rect 5531 1878 5617 2114
rect 5853 1878 5938 2114
rect 6174 1878 6259 2114
rect 6495 1878 6580 2114
rect 6816 1878 6901 2114
rect 7137 1878 7222 2114
rect 7458 1878 7543 2114
rect 7779 1878 7864 2114
rect 8100 1878 8185 2114
rect 8421 1878 8506 2114
rect 8742 1878 8827 2114
rect 9063 1878 9148 2114
rect 9384 1878 9469 2114
rect 9705 1878 9790 2114
rect 10026 1878 10111 2114
rect 10347 1878 10432 2114
rect 10668 1878 10753 2114
rect 10989 1878 11074 2114
rect 11310 1878 11395 2114
rect 11631 1878 11716 2114
rect 11952 1878 12037 2114
rect 12273 1878 12358 2114
rect 12594 1878 12679 2114
rect 12915 1878 13000 2114
rect 13236 1878 13321 2114
rect 13557 1878 13642 2114
rect 13878 1878 13963 2114
rect 14199 1878 14284 2114
rect 14520 1878 14605 2114
rect 14841 1878 15000 2114
rect 0 1508 15000 1878
rect 0 1272 143 1508
rect 379 1272 465 1508
rect 701 1272 787 1508
rect 1023 1272 1109 1508
rect 1345 1272 1431 1508
rect 1667 1272 1753 1508
rect 1989 1272 2075 1508
rect 2311 1272 2397 1508
rect 2633 1272 2719 1508
rect 2955 1272 3041 1508
rect 3277 1272 3363 1508
rect 3599 1272 3685 1508
rect 3921 1272 4007 1508
rect 4243 1272 4329 1508
rect 4565 1272 4651 1508
rect 4887 1272 4973 1508
rect 5209 1272 5295 1508
rect 5531 1272 5617 1508
rect 5853 1272 5938 1508
rect 6174 1272 6259 1508
rect 6495 1272 6580 1508
rect 6816 1272 6901 1508
rect 7137 1272 7222 1508
rect 7458 1272 7543 1508
rect 7779 1272 7864 1508
rect 8100 1272 8185 1508
rect 8421 1272 8506 1508
rect 8742 1272 8827 1508
rect 9063 1272 9148 1508
rect 9384 1272 9469 1508
rect 9705 1272 9790 1508
rect 10026 1272 10111 1508
rect 10347 1272 10432 1508
rect 10668 1272 10753 1508
rect 10989 1272 11074 1508
rect 11310 1272 11395 1508
rect 11631 1272 11716 1508
rect 11952 1272 12037 1508
rect 12273 1272 12358 1508
rect 12594 1272 12679 1508
rect 12915 1272 13000 1508
rect 13236 1272 13321 1508
rect 13557 1272 13642 1508
rect 13878 1272 13963 1508
rect 14199 1272 14284 1508
rect 14520 1272 14605 1508
rect 14841 1272 15000 1508
rect 0 1228 254 1272
rect 14746 1228 15000 1272
rect 0 904 254 948
rect 14746 904 15000 948
rect 0 903 15000 904
rect 0 667 143 903
rect 379 667 465 903
rect 701 667 787 903
rect 1023 667 1109 903
rect 1345 667 1431 903
rect 1667 667 1753 903
rect 1989 667 2075 903
rect 2311 667 2397 903
rect 2633 667 2719 903
rect 2955 667 3041 903
rect 3277 667 3363 903
rect 3599 667 3685 903
rect 3921 667 4007 903
rect 4243 667 4329 903
rect 4565 667 4651 903
rect 4887 667 4973 903
rect 5209 667 5295 903
rect 5531 667 5617 903
rect 5853 667 5938 903
rect 6174 667 6259 903
rect 6495 667 6580 903
rect 6816 667 6901 903
rect 7137 667 7222 903
rect 7458 667 7543 903
rect 7779 667 7864 903
rect 8100 667 8185 903
rect 8421 667 8506 903
rect 8742 667 8827 903
rect 9063 667 9148 903
rect 9384 667 9469 903
rect 9705 667 9790 903
rect 10026 667 10111 903
rect 10347 667 10432 903
rect 10668 667 10753 903
rect 10989 667 11074 903
rect 11310 667 11395 903
rect 11631 667 11716 903
rect 11952 667 12037 903
rect 12273 667 12358 903
rect 12594 667 12679 903
rect 12915 667 13000 903
rect 13236 667 13321 903
rect 13557 667 13642 903
rect 13878 667 13963 903
rect 14199 667 14284 903
rect 14520 667 14605 903
rect 14841 667 15000 903
rect 0 521 15000 667
rect 0 285 143 521
rect 379 285 465 521
rect 701 285 787 521
rect 1023 285 1109 521
rect 1345 285 1431 521
rect 1667 285 1753 521
rect 1989 285 2075 521
rect 2311 285 2397 521
rect 2633 285 2719 521
rect 2955 285 3041 521
rect 3277 285 3363 521
rect 3599 285 3685 521
rect 3921 285 4007 521
rect 4243 285 4329 521
rect 4565 285 4651 521
rect 4887 285 4973 521
rect 5209 285 5295 521
rect 5531 285 5617 521
rect 5853 285 5938 521
rect 6174 285 6259 521
rect 6495 285 6580 521
rect 6816 285 6901 521
rect 7137 285 7222 521
rect 7458 285 7543 521
rect 7779 285 7864 521
rect 8100 285 8185 521
rect 8421 285 8506 521
rect 8742 285 8827 521
rect 9063 285 9148 521
rect 9384 285 9469 521
rect 9705 285 9790 521
rect 10026 285 10111 521
rect 10347 285 10432 521
rect 10668 285 10753 521
rect 10989 285 11074 521
rect 11310 285 11395 521
rect 11631 285 11716 521
rect 11952 285 12037 521
rect 12273 285 12358 521
rect 12594 285 12679 521
rect 12915 285 13000 521
rect 13236 285 13321 521
rect 13557 285 13642 521
rect 13878 285 13963 521
rect 14199 285 14284 521
rect 14520 285 14605 521
rect 14841 285 15000 521
rect 0 139 15000 285
rect 0 -97 143 139
rect 379 -97 465 139
rect 701 -97 787 139
rect 1023 -97 1109 139
rect 1345 -97 1431 139
rect 1667 -97 1753 139
rect 1989 -97 2075 139
rect 2311 -97 2397 139
rect 2633 -97 2719 139
rect 2955 -97 3041 139
rect 3277 -97 3363 139
rect 3599 -97 3685 139
rect 3921 -97 4007 139
rect 4243 -97 4329 139
rect 4565 -97 4651 139
rect 4887 -97 4973 139
rect 5209 -97 5295 139
rect 5531 -97 5617 139
rect 5853 -97 5938 139
rect 6174 -97 6259 139
rect 6495 -97 6580 139
rect 6816 -97 6901 139
rect 7137 -97 7222 139
rect 7458 -97 7543 139
rect 7779 -97 7864 139
rect 8100 -97 8185 139
rect 8421 -97 8506 139
rect 8742 -97 8827 139
rect 9063 -97 9148 139
rect 9384 -97 9469 139
rect 9705 -97 9790 139
rect 10026 -97 10111 139
rect 10347 -97 10432 139
rect 10668 -97 10753 139
rect 10989 -97 11074 139
rect 11310 -97 11395 139
rect 11631 -97 11716 139
rect 11952 -97 12037 139
rect 12273 -97 12358 139
rect 12594 -97 12679 139
rect 12915 -97 13000 139
rect 13236 -97 13321 139
rect 13557 -97 13642 139
rect 13878 -97 13963 139
rect 14199 -97 14284 139
rect 14520 -97 14605 139
rect 14841 -97 15000 139
rect 0 -98 15000 -97
rect 0 -142 254 -98
rect 14746 -142 15000 -98
<< via4 >>
rect 241 39180 477 39416
rect 568 39180 804 39416
rect 895 39180 1131 39416
rect 1222 39180 1458 39416
rect 1549 39180 1785 39416
rect 1876 39180 2112 39416
rect 2203 39180 2439 39416
rect 2530 39180 2766 39416
rect 2857 39180 3093 39416
rect 3184 39180 3420 39416
rect 3511 39180 3747 39416
rect 3838 39180 4074 39416
rect 4165 39180 4401 39416
rect 4492 39180 4728 39416
rect 4819 39180 5055 39416
rect 5146 39180 5382 39416
rect 5473 39180 5709 39416
rect 5800 39180 6036 39416
rect 6127 39180 6363 39416
rect 6454 39180 6690 39416
rect 6781 39180 7017 39416
rect 7108 39180 7344 39416
rect 7435 39180 7671 39416
rect 7762 39180 7998 39416
rect 8089 39180 8325 39416
rect 8415 39180 8651 39416
rect 8741 39180 8977 39416
rect 9067 39180 9303 39416
rect 9393 39180 9629 39416
rect 9719 39180 9955 39416
rect 10045 39180 10281 39416
rect 10371 39180 10607 39416
rect 10697 39180 10933 39416
rect 11023 39180 11259 39416
rect 11349 39180 11585 39416
rect 11675 39180 11911 39416
rect 12001 39180 12237 39416
rect 12327 39180 12563 39416
rect 12653 39180 12889 39416
rect 12979 39180 13215 39416
rect 13305 39180 13541 39416
rect 13631 39180 13867 39416
rect 13957 39180 14193 39416
rect 14283 39180 14519 39416
rect 14609 39180 14845 39416
rect 241 38856 477 39092
rect 568 38856 804 39092
rect 895 38856 1131 39092
rect 1222 38856 1458 39092
rect 1549 38856 1785 39092
rect 1876 38856 2112 39092
rect 2203 38856 2439 39092
rect 2530 38856 2766 39092
rect 2857 38856 3093 39092
rect 3184 38856 3420 39092
rect 3511 38856 3747 39092
rect 3838 38856 4074 39092
rect 4165 38856 4401 39092
rect 4492 38856 4728 39092
rect 4819 38856 5055 39092
rect 5146 38856 5382 39092
rect 5473 38856 5709 39092
rect 5800 38856 6036 39092
rect 6127 38856 6363 39092
rect 6454 38856 6690 39092
rect 6781 38856 7017 39092
rect 7108 38856 7344 39092
rect 7435 38856 7671 39092
rect 7762 38856 7998 39092
rect 8089 38856 8325 39092
rect 8415 38856 8651 39092
rect 8741 38856 8977 39092
rect 9067 38856 9303 39092
rect 9393 38856 9629 39092
rect 9719 38856 9955 39092
rect 10045 38856 10281 39092
rect 10371 38856 10607 39092
rect 10697 38856 10933 39092
rect 11023 38856 11259 39092
rect 11349 38856 11585 39092
rect 11675 38856 11911 39092
rect 12001 38856 12237 39092
rect 12327 38856 12563 39092
rect 12653 38856 12889 39092
rect 12979 38856 13215 39092
rect 13305 38856 13541 39092
rect 13631 38856 13867 39092
rect 13957 38856 14193 39092
rect 14283 38856 14519 39092
rect 14609 38856 14845 39092
rect 241 38532 477 38768
rect 568 38532 804 38768
rect 895 38532 1131 38768
rect 1222 38532 1458 38768
rect 1549 38532 1785 38768
rect 1876 38532 2112 38768
rect 2203 38532 2439 38768
rect 2530 38532 2766 38768
rect 2857 38532 3093 38768
rect 3184 38532 3420 38768
rect 3511 38532 3747 38768
rect 3838 38532 4074 38768
rect 4165 38532 4401 38768
rect 4492 38532 4728 38768
rect 4819 38532 5055 38768
rect 5146 38532 5382 38768
rect 5473 38532 5709 38768
rect 5800 38532 6036 38768
rect 6127 38532 6363 38768
rect 6454 38532 6690 38768
rect 6781 38532 7017 38768
rect 7108 38532 7344 38768
rect 7435 38532 7671 38768
rect 7762 38532 7998 38768
rect 8089 38532 8325 38768
rect 8415 38532 8651 38768
rect 8741 38532 8977 38768
rect 9067 38532 9303 38768
rect 9393 38532 9629 38768
rect 9719 38532 9955 38768
rect 10045 38532 10281 38768
rect 10371 38532 10607 38768
rect 10697 38532 10933 38768
rect 11023 38532 11259 38768
rect 11349 38532 11585 38768
rect 11675 38532 11911 38768
rect 12001 38532 12237 38768
rect 12327 38532 12563 38768
rect 12653 38532 12889 38768
rect 12979 38532 13215 38768
rect 13305 38532 13541 38768
rect 13631 38532 13867 38768
rect 13957 38532 14193 38768
rect 14283 38532 14519 38768
rect 14609 38532 14845 38768
rect 241 38208 477 38444
rect 568 38208 804 38444
rect 895 38208 1131 38444
rect 1222 38208 1458 38444
rect 1549 38208 1785 38444
rect 1876 38208 2112 38444
rect 2203 38208 2439 38444
rect 2530 38208 2766 38444
rect 2857 38208 3093 38444
rect 3184 38208 3420 38444
rect 3511 38208 3747 38444
rect 3838 38208 4074 38444
rect 4165 38208 4401 38444
rect 4492 38208 4728 38444
rect 4819 38208 5055 38444
rect 5146 38208 5382 38444
rect 5473 38208 5709 38444
rect 5800 38208 6036 38444
rect 6127 38208 6363 38444
rect 6454 38208 6690 38444
rect 6781 38208 7017 38444
rect 7108 38208 7344 38444
rect 7435 38208 7671 38444
rect 7762 38208 7998 38444
rect 8089 38208 8325 38444
rect 8415 38208 8651 38444
rect 8741 38208 8977 38444
rect 9067 38208 9303 38444
rect 9393 38208 9629 38444
rect 9719 38208 9955 38444
rect 10045 38208 10281 38444
rect 10371 38208 10607 38444
rect 10697 38208 10933 38444
rect 11023 38208 11259 38444
rect 11349 38208 11585 38444
rect 11675 38208 11911 38444
rect 12001 38208 12237 38444
rect 12327 38208 12563 38444
rect 12653 38208 12889 38444
rect 12979 38208 13215 38444
rect 13305 38208 13541 38444
rect 13631 38208 13867 38444
rect 13957 38208 14193 38444
rect 14283 38208 14519 38444
rect 14609 38208 14845 38444
rect 241 37884 477 38120
rect 568 37884 804 38120
rect 895 37884 1131 38120
rect 1222 37884 1458 38120
rect 1549 37884 1785 38120
rect 1876 37884 2112 38120
rect 2203 37884 2439 38120
rect 2530 37884 2766 38120
rect 2857 37884 3093 38120
rect 3184 37884 3420 38120
rect 3511 37884 3747 38120
rect 3838 37884 4074 38120
rect 4165 37884 4401 38120
rect 4492 37884 4728 38120
rect 4819 37884 5055 38120
rect 5146 37884 5382 38120
rect 5473 37884 5709 38120
rect 5800 37884 6036 38120
rect 6127 37884 6363 38120
rect 6454 37884 6690 38120
rect 6781 37884 7017 38120
rect 7108 37884 7344 38120
rect 7435 37884 7671 38120
rect 7762 37884 7998 38120
rect 8089 37884 8325 38120
rect 8415 37884 8651 38120
rect 8741 37884 8977 38120
rect 9067 37884 9303 38120
rect 9393 37884 9629 38120
rect 9719 37884 9955 38120
rect 10045 37884 10281 38120
rect 10371 37884 10607 38120
rect 10697 37884 10933 38120
rect 11023 37884 11259 38120
rect 11349 37884 11585 38120
rect 11675 37884 11911 38120
rect 12001 37884 12237 38120
rect 12327 37884 12563 38120
rect 12653 37884 12889 38120
rect 12979 37884 13215 38120
rect 13305 37884 13541 38120
rect 13631 37884 13867 38120
rect 13957 37884 14193 38120
rect 14283 37884 14519 38120
rect 14609 37884 14845 38120
rect 241 37560 477 37796
rect 568 37560 804 37796
rect 895 37560 1131 37796
rect 1222 37560 1458 37796
rect 1549 37560 1785 37796
rect 1876 37560 2112 37796
rect 2203 37560 2439 37796
rect 2530 37560 2766 37796
rect 2857 37560 3093 37796
rect 3184 37560 3420 37796
rect 3511 37560 3747 37796
rect 3838 37560 4074 37796
rect 4165 37560 4401 37796
rect 4492 37560 4728 37796
rect 4819 37560 5055 37796
rect 5146 37560 5382 37796
rect 5473 37560 5709 37796
rect 5800 37560 6036 37796
rect 6127 37560 6363 37796
rect 6454 37560 6690 37796
rect 6781 37560 7017 37796
rect 7108 37560 7344 37796
rect 7435 37560 7671 37796
rect 7762 37560 7998 37796
rect 8089 37560 8325 37796
rect 8415 37560 8651 37796
rect 8741 37560 8977 37796
rect 9067 37560 9303 37796
rect 9393 37560 9629 37796
rect 9719 37560 9955 37796
rect 10045 37560 10281 37796
rect 10371 37560 10607 37796
rect 10697 37560 10933 37796
rect 11023 37560 11259 37796
rect 11349 37560 11585 37796
rect 11675 37560 11911 37796
rect 12001 37560 12237 37796
rect 12327 37560 12563 37796
rect 12653 37560 12889 37796
rect 12979 37560 13215 37796
rect 13305 37560 13541 37796
rect 13631 37560 13867 37796
rect 13957 37560 14193 37796
rect 14283 37560 14519 37796
rect 14609 37560 14845 37796
rect 241 37236 477 37472
rect 568 37236 804 37472
rect 895 37236 1131 37472
rect 1222 37236 1458 37472
rect 1549 37236 1785 37472
rect 1876 37236 2112 37472
rect 2203 37236 2439 37472
rect 2530 37236 2766 37472
rect 2857 37236 3093 37472
rect 3184 37236 3420 37472
rect 3511 37236 3747 37472
rect 3838 37236 4074 37472
rect 4165 37236 4401 37472
rect 4492 37236 4728 37472
rect 4819 37236 5055 37472
rect 5146 37236 5382 37472
rect 5473 37236 5709 37472
rect 5800 37236 6036 37472
rect 6127 37236 6363 37472
rect 6454 37236 6690 37472
rect 6781 37236 7017 37472
rect 7108 37236 7344 37472
rect 7435 37236 7671 37472
rect 7762 37236 7998 37472
rect 8089 37236 8325 37472
rect 8415 37236 8651 37472
rect 8741 37236 8977 37472
rect 9067 37236 9303 37472
rect 9393 37236 9629 37472
rect 9719 37236 9955 37472
rect 10045 37236 10281 37472
rect 10371 37236 10607 37472
rect 10697 37236 10933 37472
rect 11023 37236 11259 37472
rect 11349 37236 11585 37472
rect 11675 37236 11911 37472
rect 12001 37236 12237 37472
rect 12327 37236 12563 37472
rect 12653 37236 12889 37472
rect 12979 37236 13215 37472
rect 13305 37236 13541 37472
rect 13631 37236 13867 37472
rect 13957 37236 14193 37472
rect 14283 37236 14519 37472
rect 14609 37236 14845 37472
rect 241 36912 477 37148
rect 568 36912 804 37148
rect 895 36912 1131 37148
rect 1222 36912 1458 37148
rect 1549 36912 1785 37148
rect 1876 36912 2112 37148
rect 2203 36912 2439 37148
rect 2530 36912 2766 37148
rect 2857 36912 3093 37148
rect 3184 36912 3420 37148
rect 3511 36912 3747 37148
rect 3838 36912 4074 37148
rect 4165 36912 4401 37148
rect 4492 36912 4728 37148
rect 4819 36912 5055 37148
rect 5146 36912 5382 37148
rect 5473 36912 5709 37148
rect 5800 36912 6036 37148
rect 6127 36912 6363 37148
rect 6454 36912 6690 37148
rect 6781 36912 7017 37148
rect 7108 36912 7344 37148
rect 7435 36912 7671 37148
rect 7762 36912 7998 37148
rect 8089 36912 8325 37148
rect 8415 36912 8651 37148
rect 8741 36912 8977 37148
rect 9067 36912 9303 37148
rect 9393 36912 9629 37148
rect 9719 36912 9955 37148
rect 10045 36912 10281 37148
rect 10371 36912 10607 37148
rect 10697 36912 10933 37148
rect 11023 36912 11259 37148
rect 11349 36912 11585 37148
rect 11675 36912 11911 37148
rect 12001 36912 12237 37148
rect 12327 36912 12563 37148
rect 12653 36912 12889 37148
rect 12979 36912 13215 37148
rect 13305 36912 13541 37148
rect 13631 36912 13867 37148
rect 13957 36912 14193 37148
rect 14283 36912 14519 37148
rect 14609 36912 14845 37148
rect 241 36588 477 36824
rect 568 36588 804 36824
rect 895 36588 1131 36824
rect 1222 36588 1458 36824
rect 1549 36588 1785 36824
rect 1876 36588 2112 36824
rect 2203 36588 2439 36824
rect 2530 36588 2766 36824
rect 2857 36588 3093 36824
rect 3184 36588 3420 36824
rect 3511 36588 3747 36824
rect 3838 36588 4074 36824
rect 4165 36588 4401 36824
rect 4492 36588 4728 36824
rect 4819 36588 5055 36824
rect 5146 36588 5382 36824
rect 5473 36588 5709 36824
rect 5800 36588 6036 36824
rect 6127 36588 6363 36824
rect 6454 36588 6690 36824
rect 6781 36588 7017 36824
rect 7108 36588 7344 36824
rect 7435 36588 7671 36824
rect 7762 36588 7998 36824
rect 8089 36588 8325 36824
rect 8415 36588 8651 36824
rect 8741 36588 8977 36824
rect 9067 36588 9303 36824
rect 9393 36588 9629 36824
rect 9719 36588 9955 36824
rect 10045 36588 10281 36824
rect 10371 36588 10607 36824
rect 10697 36588 10933 36824
rect 11023 36588 11259 36824
rect 11349 36588 11585 36824
rect 11675 36588 11911 36824
rect 12001 36588 12237 36824
rect 12327 36588 12563 36824
rect 12653 36588 12889 36824
rect 12979 36588 13215 36824
rect 13305 36588 13541 36824
rect 13631 36588 13867 36824
rect 13957 36588 14193 36824
rect 14283 36588 14519 36824
rect 14609 36588 14845 36824
rect 241 36264 477 36500
rect 568 36264 804 36500
rect 895 36264 1131 36500
rect 1222 36264 1458 36500
rect 1549 36264 1785 36500
rect 1876 36264 2112 36500
rect 2203 36264 2439 36500
rect 2530 36264 2766 36500
rect 2857 36264 3093 36500
rect 3184 36264 3420 36500
rect 3511 36264 3747 36500
rect 3838 36264 4074 36500
rect 4165 36264 4401 36500
rect 4492 36264 4728 36500
rect 4819 36264 5055 36500
rect 5146 36264 5382 36500
rect 5473 36264 5709 36500
rect 5800 36264 6036 36500
rect 6127 36264 6363 36500
rect 6454 36264 6690 36500
rect 6781 36264 7017 36500
rect 7108 36264 7344 36500
rect 7435 36264 7671 36500
rect 7762 36264 7998 36500
rect 8089 36264 8325 36500
rect 8415 36264 8651 36500
rect 8741 36264 8977 36500
rect 9067 36264 9303 36500
rect 9393 36264 9629 36500
rect 9719 36264 9955 36500
rect 10045 36264 10281 36500
rect 10371 36264 10607 36500
rect 10697 36264 10933 36500
rect 11023 36264 11259 36500
rect 11349 36264 11585 36500
rect 11675 36264 11911 36500
rect 12001 36264 12237 36500
rect 12327 36264 12563 36500
rect 12653 36264 12889 36500
rect 12979 36264 13215 36500
rect 13305 36264 13541 36500
rect 13631 36264 13867 36500
rect 13957 36264 14193 36500
rect 14283 36264 14519 36500
rect 14609 36264 14845 36500
rect 241 35940 477 36176
rect 568 35940 804 36176
rect 895 35940 1131 36176
rect 1222 35940 1458 36176
rect 1549 35940 1785 36176
rect 1876 35940 2112 36176
rect 2203 35940 2439 36176
rect 2530 35940 2766 36176
rect 2857 35940 3093 36176
rect 3184 35940 3420 36176
rect 3511 35940 3747 36176
rect 3838 35940 4074 36176
rect 4165 35940 4401 36176
rect 4492 35940 4728 36176
rect 4819 35940 5055 36176
rect 5146 35940 5382 36176
rect 5473 35940 5709 36176
rect 5800 35940 6036 36176
rect 6127 35940 6363 36176
rect 6454 35940 6690 36176
rect 6781 35940 7017 36176
rect 7108 35940 7344 36176
rect 7435 35940 7671 36176
rect 7762 35940 7998 36176
rect 8089 35940 8325 36176
rect 8415 35940 8651 36176
rect 8741 35940 8977 36176
rect 9067 35940 9303 36176
rect 9393 35940 9629 36176
rect 9719 35940 9955 36176
rect 10045 35940 10281 36176
rect 10371 35940 10607 36176
rect 10697 35940 10933 36176
rect 11023 35940 11259 36176
rect 11349 35940 11585 36176
rect 11675 35940 11911 36176
rect 12001 35940 12237 36176
rect 12327 35940 12563 36176
rect 12653 35940 12889 36176
rect 12979 35940 13215 36176
rect 13305 35940 13541 36176
rect 13631 35940 13867 36176
rect 13957 35940 14193 36176
rect 14283 35940 14519 36176
rect 14609 35940 14845 36176
rect 241 35616 477 35852
rect 568 35616 804 35852
rect 895 35616 1131 35852
rect 1222 35616 1458 35852
rect 1549 35616 1785 35852
rect 1876 35616 2112 35852
rect 2203 35616 2439 35852
rect 2530 35616 2766 35852
rect 2857 35616 3093 35852
rect 3184 35616 3420 35852
rect 3511 35616 3747 35852
rect 3838 35616 4074 35852
rect 4165 35616 4401 35852
rect 4492 35616 4728 35852
rect 4819 35616 5055 35852
rect 5146 35616 5382 35852
rect 5473 35616 5709 35852
rect 5800 35616 6036 35852
rect 6127 35616 6363 35852
rect 6454 35616 6690 35852
rect 6781 35616 7017 35852
rect 7108 35616 7344 35852
rect 7435 35616 7671 35852
rect 7762 35616 7998 35852
rect 8089 35616 8325 35852
rect 8415 35616 8651 35852
rect 8741 35616 8977 35852
rect 9067 35616 9303 35852
rect 9393 35616 9629 35852
rect 9719 35616 9955 35852
rect 10045 35616 10281 35852
rect 10371 35616 10607 35852
rect 10697 35616 10933 35852
rect 11023 35616 11259 35852
rect 11349 35616 11585 35852
rect 11675 35616 11911 35852
rect 12001 35616 12237 35852
rect 12327 35616 12563 35852
rect 12653 35616 12889 35852
rect 12979 35616 13215 35852
rect 13305 35616 13541 35852
rect 13631 35616 13867 35852
rect 13957 35616 14193 35852
rect 14283 35616 14519 35852
rect 14609 35616 14845 35852
rect 241 35292 477 35528
rect 568 35292 804 35528
rect 895 35292 1131 35528
rect 1222 35292 1458 35528
rect 1549 35292 1785 35528
rect 1876 35292 2112 35528
rect 2203 35292 2439 35528
rect 2530 35292 2766 35528
rect 2857 35292 3093 35528
rect 3184 35292 3420 35528
rect 3511 35292 3747 35528
rect 3838 35292 4074 35528
rect 4165 35292 4401 35528
rect 4492 35292 4728 35528
rect 4819 35292 5055 35528
rect 5146 35292 5382 35528
rect 5473 35292 5709 35528
rect 5800 35292 6036 35528
rect 6127 35292 6363 35528
rect 6454 35292 6690 35528
rect 6781 35292 7017 35528
rect 7108 35292 7344 35528
rect 7435 35292 7671 35528
rect 7762 35292 7998 35528
rect 8089 35292 8325 35528
rect 8415 35292 8651 35528
rect 8741 35292 8977 35528
rect 9067 35292 9303 35528
rect 9393 35292 9629 35528
rect 9719 35292 9955 35528
rect 10045 35292 10281 35528
rect 10371 35292 10607 35528
rect 10697 35292 10933 35528
rect 11023 35292 11259 35528
rect 11349 35292 11585 35528
rect 11675 35292 11911 35528
rect 12001 35292 12237 35528
rect 12327 35292 12563 35528
rect 12653 35292 12889 35528
rect 12979 35292 13215 35528
rect 13305 35292 13541 35528
rect 13631 35292 13867 35528
rect 13957 35292 14193 35528
rect 14283 35292 14519 35528
rect 14609 35292 14845 35528
rect 241 34968 477 35204
rect 568 34968 804 35204
rect 895 34968 1131 35204
rect 1222 34968 1458 35204
rect 1549 34968 1785 35204
rect 1876 34968 2112 35204
rect 2203 34968 2439 35204
rect 2530 34968 2766 35204
rect 2857 34968 3093 35204
rect 3184 34968 3420 35204
rect 3511 34968 3747 35204
rect 3838 34968 4074 35204
rect 4165 34968 4401 35204
rect 4492 34968 4728 35204
rect 4819 34968 5055 35204
rect 5146 34968 5382 35204
rect 5473 34968 5709 35204
rect 5800 34968 6036 35204
rect 6127 34968 6363 35204
rect 6454 34968 6690 35204
rect 6781 34968 7017 35204
rect 7108 34968 7344 35204
rect 7435 34968 7671 35204
rect 7762 34968 7998 35204
rect 8089 34968 8325 35204
rect 8415 34968 8651 35204
rect 8741 34968 8977 35204
rect 9067 34968 9303 35204
rect 9393 34968 9629 35204
rect 9719 34968 9955 35204
rect 10045 34968 10281 35204
rect 10371 34968 10607 35204
rect 10697 34968 10933 35204
rect 11023 34968 11259 35204
rect 11349 34968 11585 35204
rect 11675 34968 11911 35204
rect 12001 34968 12237 35204
rect 12327 34968 12563 35204
rect 12653 34968 12889 35204
rect 12979 34968 13215 35204
rect 13305 34968 13541 35204
rect 13631 34968 13867 35204
rect 13957 34968 14193 35204
rect 14283 34968 14519 35204
rect 14609 34968 14845 35204
rect 241 34644 477 34880
rect 568 34644 804 34880
rect 895 34644 1131 34880
rect 1222 34644 1458 34880
rect 1549 34644 1785 34880
rect 1876 34644 2112 34880
rect 2203 34644 2439 34880
rect 2530 34644 2766 34880
rect 2857 34644 3093 34880
rect 3184 34644 3420 34880
rect 3511 34644 3747 34880
rect 3838 34644 4074 34880
rect 4165 34644 4401 34880
rect 4492 34644 4728 34880
rect 4819 34644 5055 34880
rect 5146 34644 5382 34880
rect 5473 34644 5709 34880
rect 5800 34644 6036 34880
rect 6127 34644 6363 34880
rect 6454 34644 6690 34880
rect 6781 34644 7017 34880
rect 7108 34644 7344 34880
rect 7435 34644 7671 34880
rect 7762 34644 7998 34880
rect 8089 34644 8325 34880
rect 8415 34644 8651 34880
rect 8741 34644 8977 34880
rect 9067 34644 9303 34880
rect 9393 34644 9629 34880
rect 9719 34644 9955 34880
rect 10045 34644 10281 34880
rect 10371 34644 10607 34880
rect 10697 34644 10933 34880
rect 11023 34644 11259 34880
rect 11349 34644 11585 34880
rect 11675 34644 11911 34880
rect 12001 34644 12237 34880
rect 12327 34644 12563 34880
rect 12653 34644 12889 34880
rect 12979 34644 13215 34880
rect 13305 34644 13541 34880
rect 13631 34644 13867 34880
rect 13957 34644 14193 34880
rect 14283 34644 14519 34880
rect 14609 34644 14845 34880
rect 143 18187 379 18423
rect 465 18187 701 18423
rect 787 18187 1023 18423
rect 1109 18187 1345 18423
rect 1431 18187 1667 18423
rect 1753 18187 1989 18423
rect 2075 18187 2311 18423
rect 2397 18187 2633 18423
rect 2719 18187 2955 18423
rect 3041 18187 3277 18423
rect 3363 18187 3599 18423
rect 3685 18187 3921 18423
rect 4007 18187 4243 18423
rect 4329 18187 4565 18423
rect 4651 18187 4887 18423
rect 4973 18187 5209 18423
rect 5295 18187 5531 18423
rect 5617 18187 5853 18423
rect 5938 18187 6174 18423
rect 6259 18187 6495 18423
rect 6580 18187 6816 18423
rect 6901 18187 7137 18423
rect 7222 18187 7458 18423
rect 7543 18187 7779 18423
rect 7864 18187 8100 18423
rect 8185 18187 8421 18423
rect 8506 18187 8742 18423
rect 8827 18187 9063 18423
rect 9148 18187 9384 18423
rect 9469 18187 9705 18423
rect 9790 18187 10026 18423
rect 10111 18187 10347 18423
rect 10432 18187 10668 18423
rect 10753 18187 10989 18423
rect 11074 18187 11310 18423
rect 11395 18187 11631 18423
rect 11716 18187 11952 18423
rect 12037 18187 12273 18423
rect 12358 18187 12594 18423
rect 12679 18187 12915 18423
rect 13000 18187 13236 18423
rect 13321 18187 13557 18423
rect 13642 18187 13878 18423
rect 13963 18187 14199 18423
rect 14284 18187 14520 18423
rect 14605 18187 14841 18423
rect 143 17851 379 18087
rect 465 17851 701 18087
rect 787 17851 1023 18087
rect 1109 17851 1345 18087
rect 1431 17851 1667 18087
rect 1753 17851 1989 18087
rect 2075 17851 2311 18087
rect 2397 17851 2633 18087
rect 2719 17851 2955 18087
rect 3041 17851 3277 18087
rect 3363 17851 3599 18087
rect 3685 17851 3921 18087
rect 4007 17851 4243 18087
rect 4329 17851 4565 18087
rect 4651 17851 4887 18087
rect 4973 17851 5209 18087
rect 5295 17851 5531 18087
rect 5617 17851 5853 18087
rect 5938 17851 6174 18087
rect 6259 17851 6495 18087
rect 6580 17851 6816 18087
rect 6901 17851 7137 18087
rect 7222 17851 7458 18087
rect 7543 17851 7779 18087
rect 7864 17851 8100 18087
rect 8185 17851 8421 18087
rect 8506 17851 8742 18087
rect 8827 17851 9063 18087
rect 9148 17851 9384 18087
rect 9469 17851 9705 18087
rect 9790 17851 10026 18087
rect 10111 17851 10347 18087
rect 10432 17851 10668 18087
rect 10753 17851 10989 18087
rect 11074 17851 11310 18087
rect 11395 17851 11631 18087
rect 11716 17851 11952 18087
rect 12037 17851 12273 18087
rect 12358 17851 12594 18087
rect 12679 17851 12915 18087
rect 13000 17851 13236 18087
rect 13321 17851 13557 18087
rect 13642 17851 13878 18087
rect 13963 17851 14199 18087
rect 14284 17851 14520 18087
rect 14605 17851 14841 18087
rect 143 17515 379 17751
rect 465 17515 701 17751
rect 787 17515 1023 17751
rect 1109 17515 1345 17751
rect 1431 17515 1667 17751
rect 1753 17515 1989 17751
rect 2075 17515 2311 17751
rect 2397 17515 2633 17751
rect 2719 17515 2955 17751
rect 3041 17515 3277 17751
rect 3363 17515 3599 17751
rect 3685 17515 3921 17751
rect 4007 17515 4243 17751
rect 4329 17515 4565 17751
rect 4651 17515 4887 17751
rect 4973 17515 5209 17751
rect 5295 17515 5531 17751
rect 5617 17515 5853 17751
rect 5938 17515 6174 17751
rect 6259 17515 6495 17751
rect 6580 17515 6816 17751
rect 6901 17515 7137 17751
rect 7222 17515 7458 17751
rect 7543 17515 7779 17751
rect 7864 17515 8100 17751
rect 8185 17515 8421 17751
rect 8506 17515 8742 17751
rect 8827 17515 9063 17751
rect 9148 17515 9384 17751
rect 9469 17515 9705 17751
rect 9790 17515 10026 17751
rect 10111 17515 10347 17751
rect 10432 17515 10668 17751
rect 10753 17515 10989 17751
rect 11074 17515 11310 17751
rect 11395 17515 11631 17751
rect 11716 17515 11952 17751
rect 12037 17515 12273 17751
rect 12358 17515 12594 17751
rect 12679 17515 12915 17751
rect 13000 17515 13236 17751
rect 13321 17515 13557 17751
rect 13642 17515 13878 17751
rect 13963 17515 14199 17751
rect 14284 17515 14520 17751
rect 14605 17515 14841 17751
rect 143 17179 379 17415
rect 465 17179 701 17415
rect 787 17179 1023 17415
rect 1109 17179 1345 17415
rect 1431 17179 1667 17415
rect 1753 17179 1989 17415
rect 2075 17179 2311 17415
rect 2397 17179 2633 17415
rect 2719 17179 2955 17415
rect 3041 17179 3277 17415
rect 3363 17179 3599 17415
rect 3685 17179 3921 17415
rect 4007 17179 4243 17415
rect 4329 17179 4565 17415
rect 4651 17179 4887 17415
rect 4973 17179 5209 17415
rect 5295 17179 5531 17415
rect 5617 17179 5853 17415
rect 5938 17179 6174 17415
rect 6259 17179 6495 17415
rect 6580 17179 6816 17415
rect 6901 17179 7137 17415
rect 7222 17179 7458 17415
rect 7543 17179 7779 17415
rect 7864 17179 8100 17415
rect 8185 17179 8421 17415
rect 8506 17179 8742 17415
rect 8827 17179 9063 17415
rect 9148 17179 9384 17415
rect 9469 17179 9705 17415
rect 9790 17179 10026 17415
rect 10111 17179 10347 17415
rect 10432 17179 10668 17415
rect 10753 17179 10989 17415
rect 11074 17179 11310 17415
rect 11395 17179 11631 17415
rect 11716 17179 11952 17415
rect 12037 17179 12273 17415
rect 12358 17179 12594 17415
rect 12679 17179 12915 17415
rect 13000 17179 13236 17415
rect 13321 17179 13557 17415
rect 13642 17179 13878 17415
rect 13963 17179 14199 17415
rect 14284 17179 14520 17415
rect 14605 17179 14841 17415
rect 143 16843 379 17079
rect 465 16843 701 17079
rect 787 16843 1023 17079
rect 1109 16843 1345 17079
rect 1431 16843 1667 17079
rect 1753 16843 1989 17079
rect 2075 16843 2311 17079
rect 2397 16843 2633 17079
rect 2719 16843 2955 17079
rect 3041 16843 3277 17079
rect 3363 16843 3599 17079
rect 3685 16843 3921 17079
rect 4007 16843 4243 17079
rect 4329 16843 4565 17079
rect 4651 16843 4887 17079
rect 4973 16843 5209 17079
rect 5295 16843 5531 17079
rect 5617 16843 5853 17079
rect 5938 16843 6174 17079
rect 6259 16843 6495 17079
rect 6580 16843 6816 17079
rect 6901 16843 7137 17079
rect 7222 16843 7458 17079
rect 7543 16843 7779 17079
rect 7864 16843 8100 17079
rect 8185 16843 8421 17079
rect 8506 16843 8742 17079
rect 8827 16843 9063 17079
rect 9148 16843 9384 17079
rect 9469 16843 9705 17079
rect 9790 16843 10026 17079
rect 10111 16843 10347 17079
rect 10432 16843 10668 17079
rect 10753 16843 10989 17079
rect 11074 16843 11310 17079
rect 11395 16843 11631 17079
rect 11716 16843 11952 17079
rect 12037 16843 12273 17079
rect 12358 16843 12594 17079
rect 12679 16843 12915 17079
rect 13000 16843 13236 17079
rect 13321 16843 13557 17079
rect 13642 16843 13878 17079
rect 13963 16843 14199 17079
rect 14284 16843 14520 17079
rect 14605 16843 14841 17079
rect 143 16507 379 16743
rect 465 16507 701 16743
rect 787 16507 1023 16743
rect 1109 16507 1345 16743
rect 1431 16507 1667 16743
rect 1753 16507 1989 16743
rect 2075 16507 2311 16743
rect 2397 16507 2633 16743
rect 2719 16507 2955 16743
rect 3041 16507 3277 16743
rect 3363 16507 3599 16743
rect 3685 16507 3921 16743
rect 4007 16507 4243 16743
rect 4329 16507 4565 16743
rect 4651 16507 4887 16743
rect 4973 16507 5209 16743
rect 5295 16507 5531 16743
rect 5617 16507 5853 16743
rect 5938 16507 6174 16743
rect 6259 16507 6495 16743
rect 6580 16507 6816 16743
rect 6901 16507 7137 16743
rect 7222 16507 7458 16743
rect 7543 16507 7779 16743
rect 7864 16507 8100 16743
rect 8185 16507 8421 16743
rect 8506 16507 8742 16743
rect 8827 16507 9063 16743
rect 9148 16507 9384 16743
rect 9469 16507 9705 16743
rect 9790 16507 10026 16743
rect 10111 16507 10347 16743
rect 10432 16507 10668 16743
rect 10753 16507 10989 16743
rect 11074 16507 11310 16743
rect 11395 16507 11631 16743
rect 11716 16507 11952 16743
rect 12037 16507 12273 16743
rect 12358 16507 12594 16743
rect 12679 16507 12915 16743
rect 13000 16507 13236 16743
rect 13321 16507 13557 16743
rect 13642 16507 13878 16743
rect 13963 16507 14199 16743
rect 14284 16507 14520 16743
rect 14605 16507 14841 16743
rect 143 16171 379 16407
rect 465 16171 701 16407
rect 787 16171 1023 16407
rect 1109 16171 1345 16407
rect 1431 16171 1667 16407
rect 1753 16171 1989 16407
rect 2075 16171 2311 16407
rect 2397 16171 2633 16407
rect 2719 16171 2955 16407
rect 3041 16171 3277 16407
rect 3363 16171 3599 16407
rect 3685 16171 3921 16407
rect 4007 16171 4243 16407
rect 4329 16171 4565 16407
rect 4651 16171 4887 16407
rect 4973 16171 5209 16407
rect 5295 16171 5531 16407
rect 5617 16171 5853 16407
rect 5938 16171 6174 16407
rect 6259 16171 6495 16407
rect 6580 16171 6816 16407
rect 6901 16171 7137 16407
rect 7222 16171 7458 16407
rect 7543 16171 7779 16407
rect 7864 16171 8100 16407
rect 8185 16171 8421 16407
rect 8506 16171 8742 16407
rect 8827 16171 9063 16407
rect 9148 16171 9384 16407
rect 9469 16171 9705 16407
rect 9790 16171 10026 16407
rect 10111 16171 10347 16407
rect 10432 16171 10668 16407
rect 10753 16171 10989 16407
rect 11074 16171 11310 16407
rect 11395 16171 11631 16407
rect 11716 16171 11952 16407
rect 12037 16171 12273 16407
rect 12358 16171 12594 16407
rect 12679 16171 12915 16407
rect 13000 16171 13236 16407
rect 13321 16171 13557 16407
rect 13642 16171 13878 16407
rect 13963 16171 14199 16407
rect 14284 16171 14520 16407
rect 14605 16171 14841 16407
rect 143 15835 379 16071
rect 465 15835 701 16071
rect 787 15835 1023 16071
rect 1109 15835 1345 16071
rect 1431 15835 1667 16071
rect 1753 15835 1989 16071
rect 2075 15835 2311 16071
rect 2397 15835 2633 16071
rect 2719 15835 2955 16071
rect 3041 15835 3277 16071
rect 3363 15835 3599 16071
rect 3685 15835 3921 16071
rect 4007 15835 4243 16071
rect 4329 15835 4565 16071
rect 4651 15835 4887 16071
rect 4973 15835 5209 16071
rect 5295 15835 5531 16071
rect 5617 15835 5853 16071
rect 5938 15835 6174 16071
rect 6259 15835 6495 16071
rect 6580 15835 6816 16071
rect 6901 15835 7137 16071
rect 7222 15835 7458 16071
rect 7543 15835 7779 16071
rect 7864 15835 8100 16071
rect 8185 15835 8421 16071
rect 8506 15835 8742 16071
rect 8827 15835 9063 16071
rect 9148 15835 9384 16071
rect 9469 15835 9705 16071
rect 9790 15835 10026 16071
rect 10111 15835 10347 16071
rect 10432 15835 10668 16071
rect 10753 15835 10989 16071
rect 11074 15835 11310 16071
rect 11395 15835 11631 16071
rect 11716 15835 11952 16071
rect 12037 15835 12273 16071
rect 12358 15835 12594 16071
rect 12679 15835 12915 16071
rect 13000 15835 13236 16071
rect 13321 15835 13557 16071
rect 13642 15835 13878 16071
rect 13963 15835 14199 16071
rect 14284 15835 14520 16071
rect 14605 15835 14841 16071
rect 143 15499 379 15735
rect 465 15499 701 15735
rect 787 15499 1023 15735
rect 1109 15499 1345 15735
rect 1431 15499 1667 15735
rect 1753 15499 1989 15735
rect 2075 15499 2311 15735
rect 2397 15499 2633 15735
rect 2719 15499 2955 15735
rect 3041 15499 3277 15735
rect 3363 15499 3599 15735
rect 3685 15499 3921 15735
rect 4007 15499 4243 15735
rect 4329 15499 4565 15735
rect 4651 15499 4887 15735
rect 4973 15499 5209 15735
rect 5295 15499 5531 15735
rect 5617 15499 5853 15735
rect 5938 15499 6174 15735
rect 6259 15499 6495 15735
rect 6580 15499 6816 15735
rect 6901 15499 7137 15735
rect 7222 15499 7458 15735
rect 7543 15499 7779 15735
rect 7864 15499 8100 15735
rect 8185 15499 8421 15735
rect 8506 15499 8742 15735
rect 8827 15499 9063 15735
rect 9148 15499 9384 15735
rect 9469 15499 9705 15735
rect 9790 15499 10026 15735
rect 10111 15499 10347 15735
rect 10432 15499 10668 15735
rect 10753 15499 10989 15735
rect 11074 15499 11310 15735
rect 11395 15499 11631 15735
rect 11716 15499 11952 15735
rect 12037 15499 12273 15735
rect 12358 15499 12594 15735
rect 12679 15499 12915 15735
rect 13000 15499 13236 15735
rect 13321 15499 13557 15735
rect 13642 15499 13878 15735
rect 13963 15499 14199 15735
rect 14284 15499 14520 15735
rect 14605 15499 14841 15735
rect 143 15163 379 15399
rect 465 15163 701 15399
rect 787 15163 1023 15399
rect 1109 15163 1345 15399
rect 1431 15163 1667 15399
rect 1753 15163 1989 15399
rect 2075 15163 2311 15399
rect 2397 15163 2633 15399
rect 2719 15163 2955 15399
rect 3041 15163 3277 15399
rect 3363 15163 3599 15399
rect 3685 15163 3921 15399
rect 4007 15163 4243 15399
rect 4329 15163 4565 15399
rect 4651 15163 4887 15399
rect 4973 15163 5209 15399
rect 5295 15163 5531 15399
rect 5617 15163 5853 15399
rect 5938 15163 6174 15399
rect 6259 15163 6495 15399
rect 6580 15163 6816 15399
rect 6901 15163 7137 15399
rect 7222 15163 7458 15399
rect 7543 15163 7779 15399
rect 7864 15163 8100 15399
rect 8185 15163 8421 15399
rect 8506 15163 8742 15399
rect 8827 15163 9063 15399
rect 9148 15163 9384 15399
rect 9469 15163 9705 15399
rect 9790 15163 10026 15399
rect 10111 15163 10347 15399
rect 10432 15163 10668 15399
rect 10753 15163 10989 15399
rect 11074 15163 11310 15399
rect 11395 15163 11631 15399
rect 11716 15163 11952 15399
rect 12037 15163 12273 15399
rect 12358 15163 12594 15399
rect 12679 15163 12915 15399
rect 13000 15163 13236 15399
rect 13321 15163 13557 15399
rect 13642 15163 13878 15399
rect 13963 15163 14199 15399
rect 14284 15163 14520 15399
rect 14605 15163 14841 15399
rect 143 14827 379 15063
rect 465 14827 701 15063
rect 787 14827 1023 15063
rect 1109 14827 1345 15063
rect 1431 14827 1667 15063
rect 1753 14827 1989 15063
rect 2075 14827 2311 15063
rect 2397 14827 2633 15063
rect 2719 14827 2955 15063
rect 3041 14827 3277 15063
rect 3363 14827 3599 15063
rect 3685 14827 3921 15063
rect 4007 14827 4243 15063
rect 4329 14827 4565 15063
rect 4651 14827 4887 15063
rect 4973 14827 5209 15063
rect 5295 14827 5531 15063
rect 5617 14827 5853 15063
rect 5938 14827 6174 15063
rect 6259 14827 6495 15063
rect 6580 14827 6816 15063
rect 6901 14827 7137 15063
rect 7222 14827 7458 15063
rect 7543 14827 7779 15063
rect 7864 14827 8100 15063
rect 8185 14827 8421 15063
rect 8506 14827 8742 15063
rect 8827 14827 9063 15063
rect 9148 14827 9384 15063
rect 9469 14827 9705 15063
rect 9790 14827 10026 15063
rect 10111 14827 10347 15063
rect 10432 14827 10668 15063
rect 10753 14827 10989 15063
rect 11074 14827 11310 15063
rect 11395 14827 11631 15063
rect 11716 14827 11952 15063
rect 12037 14827 12273 15063
rect 12358 14827 12594 15063
rect 12679 14827 12915 15063
rect 13000 14827 13236 15063
rect 13321 14827 13557 15063
rect 13642 14827 13878 15063
rect 13963 14827 14199 15063
rect 14284 14827 14520 15063
rect 14605 14827 14841 15063
rect 143 14491 379 14727
rect 465 14491 701 14727
rect 787 14491 1023 14727
rect 1109 14491 1345 14727
rect 1431 14491 1667 14727
rect 1753 14491 1989 14727
rect 2075 14491 2311 14727
rect 2397 14491 2633 14727
rect 2719 14491 2955 14727
rect 3041 14491 3277 14727
rect 3363 14491 3599 14727
rect 3685 14491 3921 14727
rect 4007 14491 4243 14727
rect 4329 14491 4565 14727
rect 4651 14491 4887 14727
rect 4973 14491 5209 14727
rect 5295 14491 5531 14727
rect 5617 14491 5853 14727
rect 5938 14491 6174 14727
rect 6259 14491 6495 14727
rect 6580 14491 6816 14727
rect 6901 14491 7137 14727
rect 7222 14491 7458 14727
rect 7543 14491 7779 14727
rect 7864 14491 8100 14727
rect 8185 14491 8421 14727
rect 8506 14491 8742 14727
rect 8827 14491 9063 14727
rect 9148 14491 9384 14727
rect 9469 14491 9705 14727
rect 9790 14491 10026 14727
rect 10111 14491 10347 14727
rect 10432 14491 10668 14727
rect 10753 14491 10989 14727
rect 11074 14491 11310 14727
rect 11395 14491 11631 14727
rect 11716 14491 11952 14727
rect 12037 14491 12273 14727
rect 12358 14491 12594 14727
rect 12679 14491 12915 14727
rect 13000 14491 13236 14727
rect 13321 14491 13557 14727
rect 13642 14491 13878 14727
rect 13963 14491 14199 14727
rect 14284 14491 14520 14727
rect 14605 14491 14841 14727
rect 143 14155 379 14391
rect 465 14155 701 14391
rect 787 14155 1023 14391
rect 1109 14155 1345 14391
rect 1431 14155 1667 14391
rect 1753 14155 1989 14391
rect 2075 14155 2311 14391
rect 2397 14155 2633 14391
rect 2719 14155 2955 14391
rect 3041 14155 3277 14391
rect 3363 14155 3599 14391
rect 3685 14155 3921 14391
rect 4007 14155 4243 14391
rect 4329 14155 4565 14391
rect 4651 14155 4887 14391
rect 4973 14155 5209 14391
rect 5295 14155 5531 14391
rect 5617 14155 5853 14391
rect 5938 14155 6174 14391
rect 6259 14155 6495 14391
rect 6580 14155 6816 14391
rect 6901 14155 7137 14391
rect 7222 14155 7458 14391
rect 7543 14155 7779 14391
rect 7864 14155 8100 14391
rect 8185 14155 8421 14391
rect 8506 14155 8742 14391
rect 8827 14155 9063 14391
rect 9148 14155 9384 14391
rect 9469 14155 9705 14391
rect 9790 14155 10026 14391
rect 10111 14155 10347 14391
rect 10432 14155 10668 14391
rect 10753 14155 10989 14391
rect 11074 14155 11310 14391
rect 11395 14155 11631 14391
rect 11716 14155 11952 14391
rect 12037 14155 12273 14391
rect 12358 14155 12594 14391
rect 12679 14155 12915 14391
rect 13000 14155 13236 14391
rect 13321 14155 13557 14391
rect 13642 14155 13878 14391
rect 13963 14155 14199 14391
rect 14284 14155 14520 14391
rect 14605 14155 14841 14391
rect 143 13819 379 14055
rect 465 13819 701 14055
rect 787 13819 1023 14055
rect 1109 13819 1345 14055
rect 1431 13819 1667 14055
rect 1753 13819 1989 14055
rect 2075 13819 2311 14055
rect 2397 13819 2633 14055
rect 2719 13819 2955 14055
rect 3041 13819 3277 14055
rect 3363 13819 3599 14055
rect 3685 13819 3921 14055
rect 4007 13819 4243 14055
rect 4329 13819 4565 14055
rect 4651 13819 4887 14055
rect 4973 13819 5209 14055
rect 5295 13819 5531 14055
rect 5617 13819 5853 14055
rect 5938 13819 6174 14055
rect 6259 13819 6495 14055
rect 6580 13819 6816 14055
rect 6901 13819 7137 14055
rect 7222 13819 7458 14055
rect 7543 13819 7779 14055
rect 7864 13819 8100 14055
rect 8185 13819 8421 14055
rect 8506 13819 8742 14055
rect 8827 13819 9063 14055
rect 9148 13819 9384 14055
rect 9469 13819 9705 14055
rect 9790 13819 10026 14055
rect 10111 13819 10347 14055
rect 10432 13819 10668 14055
rect 10753 13819 10989 14055
rect 11074 13819 11310 14055
rect 11395 13819 11631 14055
rect 11716 13819 11952 14055
rect 12037 13819 12273 14055
rect 12358 13819 12594 14055
rect 12679 13819 12915 14055
rect 13000 13819 13236 14055
rect 13321 13819 13557 14055
rect 13642 13819 13878 14055
rect 13963 13819 14199 14055
rect 14284 13819 14520 14055
rect 14605 13819 14841 14055
rect 143 13483 379 13719
rect 465 13483 701 13719
rect 787 13483 1023 13719
rect 1109 13483 1345 13719
rect 1431 13483 1667 13719
rect 1753 13483 1989 13719
rect 2075 13483 2311 13719
rect 2397 13483 2633 13719
rect 2719 13483 2955 13719
rect 3041 13483 3277 13719
rect 3363 13483 3599 13719
rect 3685 13483 3921 13719
rect 4007 13483 4243 13719
rect 4329 13483 4565 13719
rect 4651 13483 4887 13719
rect 4973 13483 5209 13719
rect 5295 13483 5531 13719
rect 5617 13483 5853 13719
rect 5938 13483 6174 13719
rect 6259 13483 6495 13719
rect 6580 13483 6816 13719
rect 6901 13483 7137 13719
rect 7222 13483 7458 13719
rect 7543 13483 7779 13719
rect 7864 13483 8100 13719
rect 8185 13483 8421 13719
rect 8506 13483 8742 13719
rect 8827 13483 9063 13719
rect 9148 13483 9384 13719
rect 9469 13483 9705 13719
rect 9790 13483 10026 13719
rect 10111 13483 10347 13719
rect 10432 13483 10668 13719
rect 10753 13483 10989 13719
rect 11074 13483 11310 13719
rect 11395 13483 11631 13719
rect 11716 13483 11952 13719
rect 12037 13483 12273 13719
rect 12358 13483 12594 13719
rect 12679 13483 12915 13719
rect 13000 13483 13236 13719
rect 13321 13483 13557 13719
rect 13642 13483 13878 13719
rect 13963 13483 14199 13719
rect 14284 13483 14520 13719
rect 14605 13483 14841 13719
rect 143 12878 379 13114
rect 465 12878 701 13114
rect 787 12878 1023 13114
rect 1109 12878 1345 13114
rect 1431 12878 1667 13114
rect 1753 12878 1989 13114
rect 2075 12878 2311 13114
rect 2397 12878 2633 13114
rect 2719 12878 2955 13114
rect 3041 12878 3277 13114
rect 3363 12878 3599 13114
rect 3685 12878 3921 13114
rect 4007 12878 4243 13114
rect 4329 12878 4565 13114
rect 4651 12878 4887 13114
rect 4973 12878 5209 13114
rect 5294 12878 5530 13114
rect 5615 12878 5851 13114
rect 5936 12878 6172 13114
rect 6257 12878 6493 13114
rect 6578 12878 6814 13114
rect 6899 12878 7135 13114
rect 7220 12878 7456 13114
rect 7541 12878 7777 13114
rect 7862 12878 8098 13114
rect 8183 12878 8419 13114
rect 8504 12878 8740 13114
rect 8825 12878 9061 13114
rect 9146 12878 9382 13114
rect 9467 12878 9703 13114
rect 9788 12878 10024 13114
rect 10109 12878 10345 13114
rect 10430 12878 10666 13114
rect 10751 12878 10987 13114
rect 11072 12878 11308 13114
rect 11393 12878 11629 13114
rect 11714 12878 11950 13114
rect 12035 12878 12271 13114
rect 12356 12878 12592 13114
rect 12677 12878 12913 13114
rect 12998 12878 13234 13114
rect 13319 12878 13555 13114
rect 13640 12878 13876 13114
rect 13961 12878 14197 13114
rect 14282 12878 14518 13114
rect 14603 12878 14839 13114
rect 143 12312 379 12548
rect 465 12312 701 12548
rect 787 12312 1023 12548
rect 1109 12312 1345 12548
rect 1431 12312 1667 12548
rect 1753 12312 1989 12548
rect 2075 12312 2311 12548
rect 2397 12312 2633 12548
rect 2719 12312 2955 12548
rect 3041 12312 3277 12548
rect 3363 12312 3599 12548
rect 3685 12312 3921 12548
rect 4007 12312 4243 12548
rect 4329 12312 4565 12548
rect 4651 12312 4887 12548
rect 4973 12312 5209 12548
rect 5294 12312 5530 12548
rect 5615 12312 5851 12548
rect 5936 12312 6172 12548
rect 6257 12312 6493 12548
rect 6578 12312 6814 12548
rect 6899 12312 7135 12548
rect 7220 12312 7456 12548
rect 7541 12312 7777 12548
rect 7862 12312 8098 12548
rect 8183 12312 8419 12548
rect 8504 12312 8740 12548
rect 8825 12312 9061 12548
rect 9146 12312 9382 12548
rect 9467 12312 9703 12548
rect 9788 12312 10024 12548
rect 10109 12312 10345 12548
rect 10430 12312 10666 12548
rect 10751 12312 10987 12548
rect 11072 12312 11308 12548
rect 11393 12312 11629 12548
rect 11714 12312 11950 12548
rect 12035 12312 12271 12548
rect 12356 12312 12592 12548
rect 12677 12312 12913 12548
rect 12998 12312 13234 12548
rect 13319 12312 13555 12548
rect 13640 12312 13876 12548
rect 13961 12312 14197 12548
rect 14282 12312 14518 12548
rect 14603 12312 14839 12548
rect 143 11708 379 11944
rect 465 11708 701 11944
rect 787 11708 1023 11944
rect 1109 11708 1345 11944
rect 1431 11708 1667 11944
rect 1753 11708 1989 11944
rect 2075 11708 2311 11944
rect 2397 11708 2633 11944
rect 2719 11708 2955 11944
rect 3041 11708 3277 11944
rect 3363 11708 3599 11944
rect 3685 11708 3921 11944
rect 4007 11708 4243 11944
rect 4329 11708 4565 11944
rect 4651 11708 4887 11944
rect 4973 11708 5209 11944
rect 5294 11708 5530 11944
rect 5615 11708 5851 11944
rect 5936 11708 6172 11944
rect 6257 11708 6493 11944
rect 6578 11708 6814 11944
rect 6899 11708 7135 11944
rect 7220 11708 7456 11944
rect 7541 11708 7777 11944
rect 7862 11708 8098 11944
rect 8183 11708 8419 11944
rect 8504 11708 8740 11944
rect 8825 11708 9061 11944
rect 9146 11708 9382 11944
rect 9467 11708 9703 11944
rect 9788 11708 10024 11944
rect 10109 11708 10345 11944
rect 10430 11708 10666 11944
rect 10751 11708 10987 11944
rect 11072 11708 11308 11944
rect 11393 11708 11629 11944
rect 11714 11708 11950 11944
rect 12035 11708 12271 11944
rect 12356 11708 12592 11944
rect 12677 11708 12913 11944
rect 12998 11708 13234 11944
rect 13319 11708 13555 11944
rect 13640 11708 13876 11944
rect 13961 11708 14197 11944
rect 14282 11708 14518 11944
rect 14603 11708 14839 11944
rect 143 11142 379 11378
rect 465 11142 701 11378
rect 787 11142 1023 11378
rect 1109 11142 1345 11378
rect 1431 11142 1667 11378
rect 1753 11142 1989 11378
rect 2075 11142 2311 11378
rect 2397 11142 2633 11378
rect 2719 11142 2955 11378
rect 3041 11142 3277 11378
rect 3363 11142 3599 11378
rect 3685 11142 3921 11378
rect 4007 11142 4243 11378
rect 4329 11142 4565 11378
rect 4651 11142 4887 11378
rect 4973 11142 5209 11378
rect 5294 11142 5530 11378
rect 5615 11142 5851 11378
rect 5936 11142 6172 11378
rect 6257 11142 6493 11378
rect 6578 11142 6814 11378
rect 6899 11142 7135 11378
rect 7220 11142 7456 11378
rect 7541 11142 7777 11378
rect 7862 11142 8098 11378
rect 8183 11142 8419 11378
rect 8504 11142 8740 11378
rect 8825 11142 9061 11378
rect 9146 11142 9382 11378
rect 9467 11142 9703 11378
rect 9788 11142 10024 11378
rect 10109 11142 10345 11378
rect 10430 11142 10666 11378
rect 10751 11142 10987 11378
rect 11072 11142 11308 11378
rect 11393 11142 11629 11378
rect 11714 11142 11950 11378
rect 12035 11142 12271 11378
rect 12356 11142 12592 11378
rect 12677 11142 12913 11378
rect 12998 11142 13234 11378
rect 13319 11142 13555 11378
rect 13640 11142 13876 11378
rect 13961 11142 14197 11378
rect 14282 11142 14518 11378
rect 14603 11142 14839 11378
rect 143 8418 379 8654
rect 465 8418 701 8654
rect 787 8418 1023 8654
rect 1109 8418 1345 8654
rect 1431 8418 1667 8654
rect 1753 8418 1989 8654
rect 2075 8418 2311 8654
rect 2397 8418 2633 8654
rect 2719 8418 2955 8654
rect 3041 8418 3277 8654
rect 3363 8418 3599 8654
rect 3685 8418 3921 8654
rect 4007 8418 4243 8654
rect 4329 8418 4565 8654
rect 4651 8418 4887 8654
rect 4973 8418 5209 8654
rect 5295 8418 5531 8654
rect 5617 8418 5853 8654
rect 5938 8418 6174 8654
rect 6259 8418 6495 8654
rect 6580 8418 6816 8654
rect 6901 8418 7137 8654
rect 7222 8418 7458 8654
rect 7543 8418 7779 8654
rect 7864 8418 8100 8654
rect 8185 8418 8421 8654
rect 8506 8418 8742 8654
rect 8827 8418 9063 8654
rect 9148 8418 9384 8654
rect 9469 8418 9705 8654
rect 9790 8418 10026 8654
rect 10111 8418 10347 8654
rect 10432 8418 10668 8654
rect 10753 8418 10989 8654
rect 11074 8418 11310 8654
rect 11395 8418 11631 8654
rect 11716 8418 11952 8654
rect 12037 8418 12273 8654
rect 12358 8418 12594 8654
rect 12679 8418 12915 8654
rect 13000 8418 13236 8654
rect 13321 8418 13557 8654
rect 13642 8418 13878 8654
rect 13963 8418 14199 8654
rect 14284 8418 14520 8654
rect 14605 8418 14841 8654
rect 143 7812 379 8048
rect 465 7812 701 8048
rect 787 7812 1023 8048
rect 1109 7812 1345 8048
rect 1431 7812 1667 8048
rect 1753 7812 1989 8048
rect 2075 7812 2311 8048
rect 2397 7812 2633 8048
rect 2719 7812 2955 8048
rect 3041 7812 3277 8048
rect 3363 7812 3599 8048
rect 3685 7812 3921 8048
rect 4007 7812 4243 8048
rect 4329 7812 4565 8048
rect 4651 7812 4887 8048
rect 4973 7812 5209 8048
rect 5295 7812 5531 8048
rect 5617 7812 5853 8048
rect 5938 7812 6174 8048
rect 6259 7812 6495 8048
rect 6580 7812 6816 8048
rect 6901 7812 7137 8048
rect 7222 7812 7458 8048
rect 7543 7812 7779 8048
rect 7864 7812 8100 8048
rect 8185 7812 8421 8048
rect 8506 7812 8742 8048
rect 8827 7812 9063 8048
rect 9148 7812 9384 8048
rect 9469 7812 9705 8048
rect 9790 7812 10026 8048
rect 10111 7812 10347 8048
rect 10432 7812 10668 8048
rect 10753 7812 10989 8048
rect 11074 7812 11310 8048
rect 11395 7812 11631 8048
rect 11716 7812 11952 8048
rect 12037 7812 12273 8048
rect 12358 7812 12594 8048
rect 12679 7812 12915 8048
rect 13000 7812 13236 8048
rect 13321 7812 13557 8048
rect 13642 7812 13878 8048
rect 13963 7812 14199 8048
rect 14284 7812 14520 8048
rect 14605 7812 14841 8048
rect 143 7208 379 7444
rect 465 7208 701 7444
rect 787 7208 1023 7444
rect 1109 7208 1345 7444
rect 1431 7208 1667 7444
rect 1753 7208 1989 7444
rect 2075 7208 2311 7444
rect 2397 7208 2633 7444
rect 2719 7208 2955 7444
rect 3041 7208 3277 7444
rect 3363 7208 3599 7444
rect 3685 7208 3921 7444
rect 4007 7208 4243 7444
rect 4329 7208 4565 7444
rect 4651 7208 4887 7444
rect 4973 7208 5209 7444
rect 5295 7208 5531 7444
rect 5617 7208 5853 7444
rect 5938 7208 6174 7444
rect 6259 7208 6495 7444
rect 6580 7208 6816 7444
rect 6901 7208 7137 7444
rect 7222 7208 7458 7444
rect 7543 7208 7779 7444
rect 7864 7208 8100 7444
rect 8185 7208 8421 7444
rect 8506 7208 8742 7444
rect 8827 7208 9063 7444
rect 9148 7208 9384 7444
rect 9469 7208 9705 7444
rect 9790 7208 10026 7444
rect 10111 7208 10347 7444
rect 10432 7208 10668 7444
rect 10753 7208 10989 7444
rect 11074 7208 11310 7444
rect 11395 7208 11631 7444
rect 11716 7208 11952 7444
rect 12037 7208 12273 7444
rect 12358 7208 12594 7444
rect 12679 7208 12915 7444
rect 13000 7208 13236 7444
rect 13321 7208 13557 7444
rect 13642 7208 13878 7444
rect 13963 7208 14199 7444
rect 14284 7208 14520 7444
rect 14605 7208 14841 7444
rect 143 6842 379 7078
rect 465 6842 701 7078
rect 787 6842 1023 7078
rect 1109 6842 1345 7078
rect 1431 6842 1667 7078
rect 1753 6842 1989 7078
rect 2075 6842 2311 7078
rect 2397 6842 2633 7078
rect 2719 6842 2955 7078
rect 3041 6842 3277 7078
rect 3363 6842 3599 7078
rect 3685 6842 3921 7078
rect 4007 6842 4243 7078
rect 4329 6842 4565 7078
rect 4651 6842 4887 7078
rect 4973 6842 5209 7078
rect 5295 6842 5531 7078
rect 5617 6842 5853 7078
rect 5938 6842 6174 7078
rect 6259 6842 6495 7078
rect 6580 6842 6816 7078
rect 6901 6842 7137 7078
rect 7222 6842 7458 7078
rect 7543 6842 7779 7078
rect 7864 6842 8100 7078
rect 8185 6842 8421 7078
rect 8506 6842 8742 7078
rect 8827 6842 9063 7078
rect 9148 6842 9384 7078
rect 9469 6842 9705 7078
rect 9790 6842 10026 7078
rect 10111 6842 10347 7078
rect 10432 6842 10668 7078
rect 10753 6842 10989 7078
rect 11074 6842 11310 7078
rect 11395 6842 11631 7078
rect 11716 6842 11952 7078
rect 12037 6842 12273 7078
rect 12358 6842 12594 7078
rect 12679 6842 12915 7078
rect 13000 6842 13236 7078
rect 13321 6842 13557 7078
rect 13642 6842 13878 7078
rect 13963 6842 14199 7078
rect 14284 6842 14520 7078
rect 14605 6842 14841 7078
rect 143 6238 379 6474
rect 465 6238 701 6474
rect 787 6238 1023 6474
rect 1109 6238 1345 6474
rect 1431 6238 1667 6474
rect 1753 6238 1989 6474
rect 2075 6238 2311 6474
rect 2397 6238 2633 6474
rect 2719 6238 2955 6474
rect 3041 6238 3277 6474
rect 3363 6238 3599 6474
rect 3685 6238 3921 6474
rect 4007 6238 4243 6474
rect 4329 6238 4565 6474
rect 4651 6238 4887 6474
rect 4973 6238 5209 6474
rect 5295 6238 5531 6474
rect 5617 6238 5853 6474
rect 5938 6238 6174 6474
rect 6259 6238 6495 6474
rect 6580 6238 6816 6474
rect 6901 6238 7137 6474
rect 7222 6238 7458 6474
rect 7543 6238 7779 6474
rect 7864 6238 8100 6474
rect 8185 6238 8421 6474
rect 8506 6238 8742 6474
rect 8827 6238 9063 6474
rect 9148 6238 9384 6474
rect 9469 6238 9705 6474
rect 9790 6238 10026 6474
rect 10111 6238 10347 6474
rect 10432 6238 10668 6474
rect 10753 6238 10989 6474
rect 11074 6238 11310 6474
rect 11395 6238 11631 6474
rect 11716 6238 11952 6474
rect 12037 6238 12273 6474
rect 12358 6238 12594 6474
rect 12679 6238 12915 6474
rect 13000 6238 13236 6474
rect 13321 6238 13557 6474
rect 13642 6238 13878 6474
rect 13963 6238 14199 6474
rect 14284 6238 14520 6474
rect 14605 6238 14841 6474
rect 143 5872 379 6108
rect 465 5872 701 6108
rect 787 5872 1023 6108
rect 1109 5872 1345 6108
rect 1431 5872 1667 6108
rect 1753 5872 1989 6108
rect 2075 5872 2311 6108
rect 2397 5872 2633 6108
rect 2719 5872 2955 6108
rect 3041 5872 3277 6108
rect 3363 5872 3599 6108
rect 3685 5872 3921 6108
rect 4007 5872 4243 6108
rect 4329 5872 4565 6108
rect 4651 5872 4887 6108
rect 4973 5872 5209 6108
rect 5295 5872 5531 6108
rect 5617 5872 5853 6108
rect 5938 5872 6174 6108
rect 6259 5872 6495 6108
rect 6580 5872 6816 6108
rect 6901 5872 7137 6108
rect 7222 5872 7458 6108
rect 7543 5872 7779 6108
rect 7864 5872 8100 6108
rect 8185 5872 8421 6108
rect 8506 5872 8742 6108
rect 8827 5872 9063 6108
rect 9148 5872 9384 6108
rect 9469 5872 9705 6108
rect 9790 5872 10026 6108
rect 10111 5872 10347 6108
rect 10432 5872 10668 6108
rect 10753 5872 10989 6108
rect 11074 5872 11310 6108
rect 11395 5872 11631 6108
rect 11716 5872 11952 6108
rect 12037 5872 12273 6108
rect 12358 5872 12594 6108
rect 12679 5872 12915 6108
rect 13000 5872 13236 6108
rect 13321 5872 13557 6108
rect 13642 5872 13878 6108
rect 13963 5872 14199 6108
rect 14284 5872 14520 6108
rect 14605 5872 14841 6108
rect 143 5268 379 5504
rect 465 5268 701 5504
rect 787 5268 1023 5504
rect 1109 5268 1345 5504
rect 1431 5268 1667 5504
rect 1753 5268 1989 5504
rect 2075 5268 2311 5504
rect 2397 5268 2633 5504
rect 2719 5268 2955 5504
rect 3041 5268 3277 5504
rect 3363 5268 3599 5504
rect 3685 5268 3921 5504
rect 4007 5268 4243 5504
rect 4329 5268 4565 5504
rect 4651 5268 4887 5504
rect 4973 5268 5209 5504
rect 5295 5268 5531 5504
rect 5617 5268 5853 5504
rect 5938 5268 6174 5504
rect 6259 5268 6495 5504
rect 6580 5268 6816 5504
rect 6901 5268 7137 5504
rect 7222 5268 7458 5504
rect 7543 5268 7779 5504
rect 7864 5268 8100 5504
rect 8185 5268 8421 5504
rect 8506 5268 8742 5504
rect 8827 5268 9063 5504
rect 9148 5268 9384 5504
rect 9469 5268 9705 5504
rect 9790 5268 10026 5504
rect 10111 5268 10347 5504
rect 10432 5268 10668 5504
rect 10753 5268 10989 5504
rect 11074 5268 11310 5504
rect 11395 5268 11631 5504
rect 11716 5268 11952 5504
rect 12037 5268 12273 5504
rect 12358 5268 12594 5504
rect 12679 5268 12915 5504
rect 13000 5268 13236 5504
rect 13321 5268 13557 5504
rect 13642 5268 13878 5504
rect 13963 5268 14199 5504
rect 14284 5268 14520 5504
rect 14605 5268 14841 5504
rect 143 4662 379 4898
rect 465 4662 701 4898
rect 787 4662 1023 4898
rect 1109 4662 1345 4898
rect 1431 4662 1667 4898
rect 1753 4662 1989 4898
rect 2075 4662 2311 4898
rect 2397 4662 2633 4898
rect 2719 4662 2955 4898
rect 3041 4662 3277 4898
rect 3363 4662 3599 4898
rect 3685 4662 3921 4898
rect 4007 4662 4243 4898
rect 4329 4662 4565 4898
rect 4651 4662 4887 4898
rect 4973 4662 5209 4898
rect 5295 4662 5531 4898
rect 5617 4662 5853 4898
rect 5938 4662 6174 4898
rect 6259 4662 6495 4898
rect 6580 4662 6816 4898
rect 6901 4662 7137 4898
rect 7222 4662 7458 4898
rect 7543 4662 7779 4898
rect 7864 4662 8100 4898
rect 8185 4662 8421 4898
rect 8506 4662 8742 4898
rect 8827 4662 9063 4898
rect 9148 4662 9384 4898
rect 9469 4662 9705 4898
rect 9790 4662 10026 4898
rect 10111 4662 10347 4898
rect 10432 4662 10668 4898
rect 10753 4662 10989 4898
rect 11074 4662 11310 4898
rect 11395 4662 11631 4898
rect 11716 4662 11952 4898
rect 12037 4662 12273 4898
rect 12358 4662 12594 4898
rect 12679 4662 12915 4898
rect 13000 4662 13236 4898
rect 13321 4662 13557 4898
rect 13642 4662 13878 4898
rect 13963 4662 14199 4898
rect 14284 4662 14520 4898
rect 14605 4662 14841 4898
rect 143 4058 379 4294
rect 465 4058 701 4294
rect 787 4058 1023 4294
rect 1109 4058 1345 4294
rect 1431 4058 1667 4294
rect 1753 4058 1989 4294
rect 2075 4058 2311 4294
rect 2397 4058 2633 4294
rect 2719 4058 2955 4294
rect 3041 4058 3277 4294
rect 3363 4058 3599 4294
rect 3685 4058 3921 4294
rect 4007 4058 4243 4294
rect 4329 4058 4565 4294
rect 4651 4058 4887 4294
rect 4973 4058 5209 4294
rect 5295 4058 5531 4294
rect 5617 4058 5853 4294
rect 5938 4058 6174 4294
rect 6259 4058 6495 4294
rect 6580 4058 6816 4294
rect 6901 4058 7137 4294
rect 7222 4058 7458 4294
rect 7543 4058 7779 4294
rect 7864 4058 8100 4294
rect 8185 4058 8421 4294
rect 8506 4058 8742 4294
rect 8827 4058 9063 4294
rect 9148 4058 9384 4294
rect 9469 4058 9705 4294
rect 9790 4058 10026 4294
rect 10111 4058 10347 4294
rect 10432 4058 10668 4294
rect 10753 4058 10989 4294
rect 11074 4058 11310 4294
rect 11395 4058 11631 4294
rect 11716 4058 11952 4294
rect 12037 4058 12273 4294
rect 12358 4058 12594 4294
rect 12679 4058 12915 4294
rect 13000 4058 13236 4294
rect 13321 4058 13557 4294
rect 13642 4058 13878 4294
rect 13963 4058 14199 4294
rect 14284 4058 14520 4294
rect 14605 4058 14841 4294
rect 143 3452 379 3688
rect 465 3452 701 3688
rect 787 3452 1023 3688
rect 1109 3452 1345 3688
rect 1431 3452 1667 3688
rect 1753 3452 1989 3688
rect 2075 3452 2311 3688
rect 2397 3452 2633 3688
rect 2719 3452 2955 3688
rect 3041 3452 3277 3688
rect 3363 3452 3599 3688
rect 3685 3452 3921 3688
rect 4007 3452 4243 3688
rect 4329 3452 4565 3688
rect 4651 3452 4887 3688
rect 4973 3452 5209 3688
rect 5295 3452 5531 3688
rect 5617 3452 5853 3688
rect 5938 3452 6174 3688
rect 6259 3452 6495 3688
rect 6580 3452 6816 3688
rect 6901 3452 7137 3688
rect 7222 3452 7458 3688
rect 7543 3452 7779 3688
rect 7864 3452 8100 3688
rect 8185 3452 8421 3688
rect 8506 3452 8742 3688
rect 8827 3452 9063 3688
rect 9148 3452 9384 3688
rect 9469 3452 9705 3688
rect 9790 3452 10026 3688
rect 10111 3452 10347 3688
rect 10432 3452 10668 3688
rect 10753 3452 10989 3688
rect 11074 3452 11310 3688
rect 11395 3452 11631 3688
rect 11716 3452 11952 3688
rect 12037 3452 12273 3688
rect 12358 3452 12594 3688
rect 12679 3452 12915 3688
rect 13000 3452 13236 3688
rect 13321 3452 13557 3688
rect 13642 3452 13878 3688
rect 13963 3452 14199 3688
rect 14284 3452 14520 3688
rect 14605 3452 14841 3688
rect 143 2848 379 3084
rect 465 2848 701 3084
rect 787 2848 1023 3084
rect 1109 2848 1345 3084
rect 1431 2848 1667 3084
rect 1753 2848 1989 3084
rect 2075 2848 2311 3084
rect 2397 2848 2633 3084
rect 2719 2848 2955 3084
rect 3041 2848 3277 3084
rect 3363 2848 3599 3084
rect 3685 2848 3921 3084
rect 4007 2848 4243 3084
rect 4329 2848 4565 3084
rect 4651 2848 4887 3084
rect 4973 2848 5209 3084
rect 5295 2848 5531 3084
rect 5617 2848 5853 3084
rect 5938 2848 6174 3084
rect 6259 2848 6495 3084
rect 6580 2848 6816 3084
rect 6901 2848 7137 3084
rect 7222 2848 7458 3084
rect 7543 2848 7779 3084
rect 7864 2848 8100 3084
rect 8185 2848 8421 3084
rect 8506 2848 8742 3084
rect 8827 2848 9063 3084
rect 9148 2848 9384 3084
rect 9469 2848 9705 3084
rect 9790 2848 10026 3084
rect 10111 2848 10347 3084
rect 10432 2848 10668 3084
rect 10753 2848 10989 3084
rect 11074 2848 11310 3084
rect 11395 2848 11631 3084
rect 11716 2848 11952 3084
rect 12037 2848 12273 3084
rect 12358 2848 12594 3084
rect 12679 2848 12915 3084
rect 13000 2848 13236 3084
rect 13321 2848 13557 3084
rect 13642 2848 13878 3084
rect 13963 2848 14199 3084
rect 14284 2848 14520 3084
rect 14605 2848 14841 3084
rect 143 2482 379 2718
rect 465 2482 701 2718
rect 787 2482 1023 2718
rect 1109 2482 1345 2718
rect 1431 2482 1667 2718
rect 1753 2482 1989 2718
rect 2075 2482 2311 2718
rect 2397 2482 2633 2718
rect 2719 2482 2955 2718
rect 3041 2482 3277 2718
rect 3363 2482 3599 2718
rect 3685 2482 3921 2718
rect 4007 2482 4243 2718
rect 4329 2482 4565 2718
rect 4651 2482 4887 2718
rect 4973 2482 5209 2718
rect 5295 2482 5531 2718
rect 5617 2482 5853 2718
rect 5938 2482 6174 2718
rect 6259 2482 6495 2718
rect 6580 2482 6816 2718
rect 6901 2482 7137 2718
rect 7222 2482 7458 2718
rect 7543 2482 7779 2718
rect 7864 2482 8100 2718
rect 8185 2482 8421 2718
rect 8506 2482 8742 2718
rect 8827 2482 9063 2718
rect 9148 2482 9384 2718
rect 9469 2482 9705 2718
rect 9790 2482 10026 2718
rect 10111 2482 10347 2718
rect 10432 2482 10668 2718
rect 10753 2482 10989 2718
rect 11074 2482 11310 2718
rect 11395 2482 11631 2718
rect 11716 2482 11952 2718
rect 12037 2482 12273 2718
rect 12358 2482 12594 2718
rect 12679 2482 12915 2718
rect 13000 2482 13236 2718
rect 13321 2482 13557 2718
rect 13642 2482 13878 2718
rect 13963 2482 14199 2718
rect 14284 2482 14520 2718
rect 14605 2482 14841 2718
rect 143 1878 379 2114
rect 465 1878 701 2114
rect 787 1878 1023 2114
rect 1109 1878 1345 2114
rect 1431 1878 1667 2114
rect 1753 1878 1989 2114
rect 2075 1878 2311 2114
rect 2397 1878 2633 2114
rect 2719 1878 2955 2114
rect 3041 1878 3277 2114
rect 3363 1878 3599 2114
rect 3685 1878 3921 2114
rect 4007 1878 4243 2114
rect 4329 1878 4565 2114
rect 4651 1878 4887 2114
rect 4973 1878 5209 2114
rect 5295 1878 5531 2114
rect 5617 1878 5853 2114
rect 5938 1878 6174 2114
rect 6259 1878 6495 2114
rect 6580 1878 6816 2114
rect 6901 1878 7137 2114
rect 7222 1878 7458 2114
rect 7543 1878 7779 2114
rect 7864 1878 8100 2114
rect 8185 1878 8421 2114
rect 8506 1878 8742 2114
rect 8827 1878 9063 2114
rect 9148 1878 9384 2114
rect 9469 1878 9705 2114
rect 9790 1878 10026 2114
rect 10111 1878 10347 2114
rect 10432 1878 10668 2114
rect 10753 1878 10989 2114
rect 11074 1878 11310 2114
rect 11395 1878 11631 2114
rect 11716 1878 11952 2114
rect 12037 1878 12273 2114
rect 12358 1878 12594 2114
rect 12679 1878 12915 2114
rect 13000 1878 13236 2114
rect 13321 1878 13557 2114
rect 13642 1878 13878 2114
rect 13963 1878 14199 2114
rect 14284 1878 14520 2114
rect 14605 1878 14841 2114
rect 143 1272 379 1508
rect 465 1272 701 1508
rect 787 1272 1023 1508
rect 1109 1272 1345 1508
rect 1431 1272 1667 1508
rect 1753 1272 1989 1508
rect 2075 1272 2311 1508
rect 2397 1272 2633 1508
rect 2719 1272 2955 1508
rect 3041 1272 3277 1508
rect 3363 1272 3599 1508
rect 3685 1272 3921 1508
rect 4007 1272 4243 1508
rect 4329 1272 4565 1508
rect 4651 1272 4887 1508
rect 4973 1272 5209 1508
rect 5295 1272 5531 1508
rect 5617 1272 5853 1508
rect 5938 1272 6174 1508
rect 6259 1272 6495 1508
rect 6580 1272 6816 1508
rect 6901 1272 7137 1508
rect 7222 1272 7458 1508
rect 7543 1272 7779 1508
rect 7864 1272 8100 1508
rect 8185 1272 8421 1508
rect 8506 1272 8742 1508
rect 8827 1272 9063 1508
rect 9148 1272 9384 1508
rect 9469 1272 9705 1508
rect 9790 1272 10026 1508
rect 10111 1272 10347 1508
rect 10432 1272 10668 1508
rect 10753 1272 10989 1508
rect 11074 1272 11310 1508
rect 11395 1272 11631 1508
rect 11716 1272 11952 1508
rect 12037 1272 12273 1508
rect 12358 1272 12594 1508
rect 12679 1272 12915 1508
rect 13000 1272 13236 1508
rect 13321 1272 13557 1508
rect 13642 1272 13878 1508
rect 13963 1272 14199 1508
rect 14284 1272 14520 1508
rect 14605 1272 14841 1508
rect 143 667 379 903
rect 465 667 701 903
rect 787 667 1023 903
rect 1109 667 1345 903
rect 1431 667 1667 903
rect 1753 667 1989 903
rect 2075 667 2311 903
rect 2397 667 2633 903
rect 2719 667 2955 903
rect 3041 667 3277 903
rect 3363 667 3599 903
rect 3685 667 3921 903
rect 4007 667 4243 903
rect 4329 667 4565 903
rect 4651 667 4887 903
rect 4973 667 5209 903
rect 5295 667 5531 903
rect 5617 667 5853 903
rect 5938 667 6174 903
rect 6259 667 6495 903
rect 6580 667 6816 903
rect 6901 667 7137 903
rect 7222 667 7458 903
rect 7543 667 7779 903
rect 7864 667 8100 903
rect 8185 667 8421 903
rect 8506 667 8742 903
rect 8827 667 9063 903
rect 9148 667 9384 903
rect 9469 667 9705 903
rect 9790 667 10026 903
rect 10111 667 10347 903
rect 10432 667 10668 903
rect 10753 667 10989 903
rect 11074 667 11310 903
rect 11395 667 11631 903
rect 11716 667 11952 903
rect 12037 667 12273 903
rect 12358 667 12594 903
rect 12679 667 12915 903
rect 13000 667 13236 903
rect 13321 667 13557 903
rect 13642 667 13878 903
rect 13963 667 14199 903
rect 14284 667 14520 903
rect 14605 667 14841 903
rect 143 285 379 521
rect 465 285 701 521
rect 787 285 1023 521
rect 1109 285 1345 521
rect 1431 285 1667 521
rect 1753 285 1989 521
rect 2075 285 2311 521
rect 2397 285 2633 521
rect 2719 285 2955 521
rect 3041 285 3277 521
rect 3363 285 3599 521
rect 3685 285 3921 521
rect 4007 285 4243 521
rect 4329 285 4565 521
rect 4651 285 4887 521
rect 4973 285 5209 521
rect 5295 285 5531 521
rect 5617 285 5853 521
rect 5938 285 6174 521
rect 6259 285 6495 521
rect 6580 285 6816 521
rect 6901 285 7137 521
rect 7222 285 7458 521
rect 7543 285 7779 521
rect 7864 285 8100 521
rect 8185 285 8421 521
rect 8506 285 8742 521
rect 8827 285 9063 521
rect 9148 285 9384 521
rect 9469 285 9705 521
rect 9790 285 10026 521
rect 10111 285 10347 521
rect 10432 285 10668 521
rect 10753 285 10989 521
rect 11074 285 11310 521
rect 11395 285 11631 521
rect 11716 285 11952 521
rect 12037 285 12273 521
rect 12358 285 12594 521
rect 12679 285 12915 521
rect 13000 285 13236 521
rect 13321 285 13557 521
rect 13642 285 13878 521
rect 13963 285 14199 521
rect 14284 285 14520 521
rect 14605 285 14841 521
rect 143 -97 379 139
rect 465 -97 701 139
rect 787 -97 1023 139
rect 1109 -97 1345 139
rect 1431 -97 1667 139
rect 1753 -97 1989 139
rect 2075 -97 2311 139
rect 2397 -97 2633 139
rect 2719 -97 2955 139
rect 3041 -97 3277 139
rect 3363 -97 3599 139
rect 3685 -97 3921 139
rect 4007 -97 4243 139
rect 4329 -97 4565 139
rect 4651 -97 4887 139
rect 4973 -97 5209 139
rect 5295 -97 5531 139
rect 5617 -97 5853 139
rect 5938 -97 6174 139
rect 6259 -97 6495 139
rect 6580 -97 6816 139
rect 6901 -97 7137 139
rect 7222 -97 7458 139
rect 7543 -97 7779 139
rect 7864 -97 8100 139
rect 8185 -97 8421 139
rect 8506 -97 8742 139
rect 8827 -97 9063 139
rect 9148 -97 9384 139
rect 9469 -97 9705 139
rect 9790 -97 10026 139
rect 10111 -97 10347 139
rect 10432 -97 10668 139
rect 10753 -97 10989 139
rect 11074 -97 11310 139
rect 11395 -97 11631 139
rect 11716 -97 11952 139
rect 12037 -97 12273 139
rect 12358 -97 12594 139
rect 12679 -97 12915 139
rect 13000 -97 13236 139
rect 13321 -97 13557 139
rect 13642 -97 13878 139
rect 13963 -97 14199 139
rect 14284 -97 14520 139
rect 14605 -97 14841 139
<< metal5 >>
rect 0 39416 15000 39451
rect 0 39180 241 39416
rect 477 39180 568 39416
rect 804 39180 895 39416
rect 1131 39180 1222 39416
rect 1458 39180 1549 39416
rect 1785 39180 1876 39416
rect 2112 39180 2203 39416
rect 2439 39180 2530 39416
rect 2766 39180 2857 39416
rect 3093 39180 3184 39416
rect 3420 39180 3511 39416
rect 3747 39180 3838 39416
rect 4074 39180 4165 39416
rect 4401 39180 4492 39416
rect 4728 39180 4819 39416
rect 5055 39180 5146 39416
rect 5382 39180 5473 39416
rect 5709 39180 5800 39416
rect 6036 39180 6127 39416
rect 6363 39180 6454 39416
rect 6690 39180 6781 39416
rect 7017 39180 7108 39416
rect 7344 39180 7435 39416
rect 7671 39180 7762 39416
rect 7998 39180 8089 39416
rect 8325 39180 8415 39416
rect 8651 39180 8741 39416
rect 8977 39180 9067 39416
rect 9303 39180 9393 39416
rect 9629 39180 9719 39416
rect 9955 39180 10045 39416
rect 10281 39180 10371 39416
rect 10607 39180 10697 39416
rect 10933 39180 11023 39416
rect 11259 39180 11349 39416
rect 11585 39180 11675 39416
rect 11911 39180 12001 39416
rect 12237 39180 12327 39416
rect 12563 39180 12653 39416
rect 12889 39180 12979 39416
rect 13215 39180 13305 39416
rect 13541 39180 13631 39416
rect 13867 39180 13957 39416
rect 14193 39180 14283 39416
rect 14519 39180 14609 39416
rect 14845 39180 15000 39416
rect 0 39092 15000 39180
rect 0 38856 241 39092
rect 477 38856 568 39092
rect 804 38856 895 39092
rect 1131 38856 1222 39092
rect 1458 38856 1549 39092
rect 1785 38856 1876 39092
rect 2112 38856 2203 39092
rect 2439 38856 2530 39092
rect 2766 38856 2857 39092
rect 3093 38856 3184 39092
rect 3420 38856 3511 39092
rect 3747 38856 3838 39092
rect 4074 38856 4165 39092
rect 4401 38856 4492 39092
rect 4728 38856 4819 39092
rect 5055 38856 5146 39092
rect 5382 38856 5473 39092
rect 5709 38856 5800 39092
rect 6036 38856 6127 39092
rect 6363 38856 6454 39092
rect 6690 38856 6781 39092
rect 7017 38856 7108 39092
rect 7344 38856 7435 39092
rect 7671 38856 7762 39092
rect 7998 38856 8089 39092
rect 8325 38856 8415 39092
rect 8651 38856 8741 39092
rect 8977 38856 9067 39092
rect 9303 38856 9393 39092
rect 9629 38856 9719 39092
rect 9955 38856 10045 39092
rect 10281 38856 10371 39092
rect 10607 38856 10697 39092
rect 10933 38856 11023 39092
rect 11259 38856 11349 39092
rect 11585 38856 11675 39092
rect 11911 38856 12001 39092
rect 12237 38856 12327 39092
rect 12563 38856 12653 39092
rect 12889 38856 12979 39092
rect 13215 38856 13305 39092
rect 13541 38856 13631 39092
rect 13867 38856 13957 39092
rect 14193 38856 14283 39092
rect 14519 38856 14609 39092
rect 14845 38856 15000 39092
rect 0 38768 15000 38856
rect 0 38532 241 38768
rect 477 38532 568 38768
rect 804 38532 895 38768
rect 1131 38532 1222 38768
rect 1458 38532 1549 38768
rect 1785 38532 1876 38768
rect 2112 38532 2203 38768
rect 2439 38532 2530 38768
rect 2766 38532 2857 38768
rect 3093 38532 3184 38768
rect 3420 38532 3511 38768
rect 3747 38532 3838 38768
rect 4074 38532 4165 38768
rect 4401 38532 4492 38768
rect 4728 38532 4819 38768
rect 5055 38532 5146 38768
rect 5382 38532 5473 38768
rect 5709 38532 5800 38768
rect 6036 38532 6127 38768
rect 6363 38532 6454 38768
rect 6690 38532 6781 38768
rect 7017 38532 7108 38768
rect 7344 38532 7435 38768
rect 7671 38532 7762 38768
rect 7998 38532 8089 38768
rect 8325 38532 8415 38768
rect 8651 38532 8741 38768
rect 8977 38532 9067 38768
rect 9303 38532 9393 38768
rect 9629 38532 9719 38768
rect 9955 38532 10045 38768
rect 10281 38532 10371 38768
rect 10607 38532 10697 38768
rect 10933 38532 11023 38768
rect 11259 38532 11349 38768
rect 11585 38532 11675 38768
rect 11911 38532 12001 38768
rect 12237 38532 12327 38768
rect 12563 38532 12653 38768
rect 12889 38532 12979 38768
rect 13215 38532 13305 38768
rect 13541 38532 13631 38768
rect 13867 38532 13957 38768
rect 14193 38532 14283 38768
rect 14519 38532 14609 38768
rect 14845 38532 15000 38768
rect 0 38444 15000 38532
rect 0 38208 241 38444
rect 477 38208 568 38444
rect 804 38208 895 38444
rect 1131 38208 1222 38444
rect 1458 38208 1549 38444
rect 1785 38208 1876 38444
rect 2112 38208 2203 38444
rect 2439 38208 2530 38444
rect 2766 38208 2857 38444
rect 3093 38208 3184 38444
rect 3420 38208 3511 38444
rect 3747 38208 3838 38444
rect 4074 38208 4165 38444
rect 4401 38208 4492 38444
rect 4728 38208 4819 38444
rect 5055 38208 5146 38444
rect 5382 38208 5473 38444
rect 5709 38208 5800 38444
rect 6036 38208 6127 38444
rect 6363 38208 6454 38444
rect 6690 38208 6781 38444
rect 7017 38208 7108 38444
rect 7344 38208 7435 38444
rect 7671 38208 7762 38444
rect 7998 38208 8089 38444
rect 8325 38208 8415 38444
rect 8651 38208 8741 38444
rect 8977 38208 9067 38444
rect 9303 38208 9393 38444
rect 9629 38208 9719 38444
rect 9955 38208 10045 38444
rect 10281 38208 10371 38444
rect 10607 38208 10697 38444
rect 10933 38208 11023 38444
rect 11259 38208 11349 38444
rect 11585 38208 11675 38444
rect 11911 38208 12001 38444
rect 12237 38208 12327 38444
rect 12563 38208 12653 38444
rect 12889 38208 12979 38444
rect 13215 38208 13305 38444
rect 13541 38208 13631 38444
rect 13867 38208 13957 38444
rect 14193 38208 14283 38444
rect 14519 38208 14609 38444
rect 14845 38208 15000 38444
rect 0 38120 15000 38208
rect 0 37884 241 38120
rect 477 37884 568 38120
rect 804 37884 895 38120
rect 1131 37884 1222 38120
rect 1458 37884 1549 38120
rect 1785 37884 1876 38120
rect 2112 37884 2203 38120
rect 2439 37884 2530 38120
rect 2766 37884 2857 38120
rect 3093 37884 3184 38120
rect 3420 37884 3511 38120
rect 3747 37884 3838 38120
rect 4074 37884 4165 38120
rect 4401 37884 4492 38120
rect 4728 37884 4819 38120
rect 5055 37884 5146 38120
rect 5382 37884 5473 38120
rect 5709 37884 5800 38120
rect 6036 37884 6127 38120
rect 6363 37884 6454 38120
rect 6690 37884 6781 38120
rect 7017 37884 7108 38120
rect 7344 37884 7435 38120
rect 7671 37884 7762 38120
rect 7998 37884 8089 38120
rect 8325 37884 8415 38120
rect 8651 37884 8741 38120
rect 8977 37884 9067 38120
rect 9303 37884 9393 38120
rect 9629 37884 9719 38120
rect 9955 37884 10045 38120
rect 10281 37884 10371 38120
rect 10607 37884 10697 38120
rect 10933 37884 11023 38120
rect 11259 37884 11349 38120
rect 11585 37884 11675 38120
rect 11911 37884 12001 38120
rect 12237 37884 12327 38120
rect 12563 37884 12653 38120
rect 12889 37884 12979 38120
rect 13215 37884 13305 38120
rect 13541 37884 13631 38120
rect 13867 37884 13957 38120
rect 14193 37884 14283 38120
rect 14519 37884 14609 38120
rect 14845 37884 15000 38120
rect 0 37796 15000 37884
rect 0 37560 241 37796
rect 477 37560 568 37796
rect 804 37560 895 37796
rect 1131 37560 1222 37796
rect 1458 37560 1549 37796
rect 1785 37560 1876 37796
rect 2112 37560 2203 37796
rect 2439 37560 2530 37796
rect 2766 37560 2857 37796
rect 3093 37560 3184 37796
rect 3420 37560 3511 37796
rect 3747 37560 3838 37796
rect 4074 37560 4165 37796
rect 4401 37560 4492 37796
rect 4728 37560 4819 37796
rect 5055 37560 5146 37796
rect 5382 37560 5473 37796
rect 5709 37560 5800 37796
rect 6036 37560 6127 37796
rect 6363 37560 6454 37796
rect 6690 37560 6781 37796
rect 7017 37560 7108 37796
rect 7344 37560 7435 37796
rect 7671 37560 7762 37796
rect 7998 37560 8089 37796
rect 8325 37560 8415 37796
rect 8651 37560 8741 37796
rect 8977 37560 9067 37796
rect 9303 37560 9393 37796
rect 9629 37560 9719 37796
rect 9955 37560 10045 37796
rect 10281 37560 10371 37796
rect 10607 37560 10697 37796
rect 10933 37560 11023 37796
rect 11259 37560 11349 37796
rect 11585 37560 11675 37796
rect 11911 37560 12001 37796
rect 12237 37560 12327 37796
rect 12563 37560 12653 37796
rect 12889 37560 12979 37796
rect 13215 37560 13305 37796
rect 13541 37560 13631 37796
rect 13867 37560 13957 37796
rect 14193 37560 14283 37796
rect 14519 37560 14609 37796
rect 14845 37560 15000 37796
rect 0 37472 15000 37560
rect 0 37236 241 37472
rect 477 37236 568 37472
rect 804 37236 895 37472
rect 1131 37236 1222 37472
rect 1458 37236 1549 37472
rect 1785 37236 1876 37472
rect 2112 37236 2203 37472
rect 2439 37236 2530 37472
rect 2766 37236 2857 37472
rect 3093 37236 3184 37472
rect 3420 37236 3511 37472
rect 3747 37236 3838 37472
rect 4074 37236 4165 37472
rect 4401 37236 4492 37472
rect 4728 37236 4819 37472
rect 5055 37236 5146 37472
rect 5382 37236 5473 37472
rect 5709 37236 5800 37472
rect 6036 37236 6127 37472
rect 6363 37236 6454 37472
rect 6690 37236 6781 37472
rect 7017 37236 7108 37472
rect 7344 37236 7435 37472
rect 7671 37236 7762 37472
rect 7998 37236 8089 37472
rect 8325 37236 8415 37472
rect 8651 37236 8741 37472
rect 8977 37236 9067 37472
rect 9303 37236 9393 37472
rect 9629 37236 9719 37472
rect 9955 37236 10045 37472
rect 10281 37236 10371 37472
rect 10607 37236 10697 37472
rect 10933 37236 11023 37472
rect 11259 37236 11349 37472
rect 11585 37236 11675 37472
rect 11911 37236 12001 37472
rect 12237 37236 12327 37472
rect 12563 37236 12653 37472
rect 12889 37236 12979 37472
rect 13215 37236 13305 37472
rect 13541 37236 13631 37472
rect 13867 37236 13957 37472
rect 14193 37236 14283 37472
rect 14519 37236 14609 37472
rect 14845 37236 15000 37472
rect 0 37148 15000 37236
rect 0 36912 241 37148
rect 477 36912 568 37148
rect 804 36912 895 37148
rect 1131 36912 1222 37148
rect 1458 36912 1549 37148
rect 1785 36912 1876 37148
rect 2112 36912 2203 37148
rect 2439 36912 2530 37148
rect 2766 36912 2857 37148
rect 3093 36912 3184 37148
rect 3420 36912 3511 37148
rect 3747 36912 3838 37148
rect 4074 36912 4165 37148
rect 4401 36912 4492 37148
rect 4728 36912 4819 37148
rect 5055 36912 5146 37148
rect 5382 36912 5473 37148
rect 5709 36912 5800 37148
rect 6036 36912 6127 37148
rect 6363 36912 6454 37148
rect 6690 36912 6781 37148
rect 7017 36912 7108 37148
rect 7344 36912 7435 37148
rect 7671 36912 7762 37148
rect 7998 36912 8089 37148
rect 8325 36912 8415 37148
rect 8651 36912 8741 37148
rect 8977 36912 9067 37148
rect 9303 36912 9393 37148
rect 9629 36912 9719 37148
rect 9955 36912 10045 37148
rect 10281 36912 10371 37148
rect 10607 36912 10697 37148
rect 10933 36912 11023 37148
rect 11259 36912 11349 37148
rect 11585 36912 11675 37148
rect 11911 36912 12001 37148
rect 12237 36912 12327 37148
rect 12563 36912 12653 37148
rect 12889 36912 12979 37148
rect 13215 36912 13305 37148
rect 13541 36912 13631 37148
rect 13867 36912 13957 37148
rect 14193 36912 14283 37148
rect 14519 36912 14609 37148
rect 14845 36912 15000 37148
rect 0 36824 15000 36912
rect 0 36588 241 36824
rect 477 36588 568 36824
rect 804 36588 895 36824
rect 1131 36588 1222 36824
rect 1458 36588 1549 36824
rect 1785 36588 1876 36824
rect 2112 36588 2203 36824
rect 2439 36588 2530 36824
rect 2766 36588 2857 36824
rect 3093 36588 3184 36824
rect 3420 36588 3511 36824
rect 3747 36588 3838 36824
rect 4074 36588 4165 36824
rect 4401 36588 4492 36824
rect 4728 36588 4819 36824
rect 5055 36588 5146 36824
rect 5382 36588 5473 36824
rect 5709 36588 5800 36824
rect 6036 36588 6127 36824
rect 6363 36588 6454 36824
rect 6690 36588 6781 36824
rect 7017 36588 7108 36824
rect 7344 36588 7435 36824
rect 7671 36588 7762 36824
rect 7998 36588 8089 36824
rect 8325 36588 8415 36824
rect 8651 36588 8741 36824
rect 8977 36588 9067 36824
rect 9303 36588 9393 36824
rect 9629 36588 9719 36824
rect 9955 36588 10045 36824
rect 10281 36588 10371 36824
rect 10607 36588 10697 36824
rect 10933 36588 11023 36824
rect 11259 36588 11349 36824
rect 11585 36588 11675 36824
rect 11911 36588 12001 36824
rect 12237 36588 12327 36824
rect 12563 36588 12653 36824
rect 12889 36588 12979 36824
rect 13215 36588 13305 36824
rect 13541 36588 13631 36824
rect 13867 36588 13957 36824
rect 14193 36588 14283 36824
rect 14519 36588 14609 36824
rect 14845 36588 15000 36824
rect 0 36500 15000 36588
rect 0 36264 241 36500
rect 477 36264 568 36500
rect 804 36264 895 36500
rect 1131 36264 1222 36500
rect 1458 36264 1549 36500
rect 1785 36264 1876 36500
rect 2112 36264 2203 36500
rect 2439 36264 2530 36500
rect 2766 36264 2857 36500
rect 3093 36264 3184 36500
rect 3420 36264 3511 36500
rect 3747 36264 3838 36500
rect 4074 36264 4165 36500
rect 4401 36264 4492 36500
rect 4728 36264 4819 36500
rect 5055 36264 5146 36500
rect 5382 36264 5473 36500
rect 5709 36264 5800 36500
rect 6036 36264 6127 36500
rect 6363 36264 6454 36500
rect 6690 36264 6781 36500
rect 7017 36264 7108 36500
rect 7344 36264 7435 36500
rect 7671 36264 7762 36500
rect 7998 36264 8089 36500
rect 8325 36264 8415 36500
rect 8651 36264 8741 36500
rect 8977 36264 9067 36500
rect 9303 36264 9393 36500
rect 9629 36264 9719 36500
rect 9955 36264 10045 36500
rect 10281 36264 10371 36500
rect 10607 36264 10697 36500
rect 10933 36264 11023 36500
rect 11259 36264 11349 36500
rect 11585 36264 11675 36500
rect 11911 36264 12001 36500
rect 12237 36264 12327 36500
rect 12563 36264 12653 36500
rect 12889 36264 12979 36500
rect 13215 36264 13305 36500
rect 13541 36264 13631 36500
rect 13867 36264 13957 36500
rect 14193 36264 14283 36500
rect 14519 36264 14609 36500
rect 14845 36264 15000 36500
rect 0 36176 15000 36264
rect 0 35940 241 36176
rect 477 35940 568 36176
rect 804 35940 895 36176
rect 1131 35940 1222 36176
rect 1458 35940 1549 36176
rect 1785 35940 1876 36176
rect 2112 35940 2203 36176
rect 2439 35940 2530 36176
rect 2766 35940 2857 36176
rect 3093 35940 3184 36176
rect 3420 35940 3511 36176
rect 3747 35940 3838 36176
rect 4074 35940 4165 36176
rect 4401 35940 4492 36176
rect 4728 35940 4819 36176
rect 5055 35940 5146 36176
rect 5382 35940 5473 36176
rect 5709 35940 5800 36176
rect 6036 35940 6127 36176
rect 6363 35940 6454 36176
rect 6690 35940 6781 36176
rect 7017 35940 7108 36176
rect 7344 35940 7435 36176
rect 7671 35940 7762 36176
rect 7998 35940 8089 36176
rect 8325 35940 8415 36176
rect 8651 35940 8741 36176
rect 8977 35940 9067 36176
rect 9303 35940 9393 36176
rect 9629 35940 9719 36176
rect 9955 35940 10045 36176
rect 10281 35940 10371 36176
rect 10607 35940 10697 36176
rect 10933 35940 11023 36176
rect 11259 35940 11349 36176
rect 11585 35940 11675 36176
rect 11911 35940 12001 36176
rect 12237 35940 12327 36176
rect 12563 35940 12653 36176
rect 12889 35940 12979 36176
rect 13215 35940 13305 36176
rect 13541 35940 13631 36176
rect 13867 35940 13957 36176
rect 14193 35940 14283 36176
rect 14519 35940 14609 36176
rect 14845 35940 15000 36176
rect 0 35852 15000 35940
rect 0 35616 241 35852
rect 477 35616 568 35852
rect 804 35616 895 35852
rect 1131 35616 1222 35852
rect 1458 35616 1549 35852
rect 1785 35616 1876 35852
rect 2112 35616 2203 35852
rect 2439 35616 2530 35852
rect 2766 35616 2857 35852
rect 3093 35616 3184 35852
rect 3420 35616 3511 35852
rect 3747 35616 3838 35852
rect 4074 35616 4165 35852
rect 4401 35616 4492 35852
rect 4728 35616 4819 35852
rect 5055 35616 5146 35852
rect 5382 35616 5473 35852
rect 5709 35616 5800 35852
rect 6036 35616 6127 35852
rect 6363 35616 6454 35852
rect 6690 35616 6781 35852
rect 7017 35616 7108 35852
rect 7344 35616 7435 35852
rect 7671 35616 7762 35852
rect 7998 35616 8089 35852
rect 8325 35616 8415 35852
rect 8651 35616 8741 35852
rect 8977 35616 9067 35852
rect 9303 35616 9393 35852
rect 9629 35616 9719 35852
rect 9955 35616 10045 35852
rect 10281 35616 10371 35852
rect 10607 35616 10697 35852
rect 10933 35616 11023 35852
rect 11259 35616 11349 35852
rect 11585 35616 11675 35852
rect 11911 35616 12001 35852
rect 12237 35616 12327 35852
rect 12563 35616 12653 35852
rect 12889 35616 12979 35852
rect 13215 35616 13305 35852
rect 13541 35616 13631 35852
rect 13867 35616 13957 35852
rect 14193 35616 14283 35852
rect 14519 35616 14609 35852
rect 14845 35616 15000 35852
rect 0 35528 15000 35616
rect 0 35292 241 35528
rect 477 35292 568 35528
rect 804 35292 895 35528
rect 1131 35292 1222 35528
rect 1458 35292 1549 35528
rect 1785 35292 1876 35528
rect 2112 35292 2203 35528
rect 2439 35292 2530 35528
rect 2766 35292 2857 35528
rect 3093 35292 3184 35528
rect 3420 35292 3511 35528
rect 3747 35292 3838 35528
rect 4074 35292 4165 35528
rect 4401 35292 4492 35528
rect 4728 35292 4819 35528
rect 5055 35292 5146 35528
rect 5382 35292 5473 35528
rect 5709 35292 5800 35528
rect 6036 35292 6127 35528
rect 6363 35292 6454 35528
rect 6690 35292 6781 35528
rect 7017 35292 7108 35528
rect 7344 35292 7435 35528
rect 7671 35292 7762 35528
rect 7998 35292 8089 35528
rect 8325 35292 8415 35528
rect 8651 35292 8741 35528
rect 8977 35292 9067 35528
rect 9303 35292 9393 35528
rect 9629 35292 9719 35528
rect 9955 35292 10045 35528
rect 10281 35292 10371 35528
rect 10607 35292 10697 35528
rect 10933 35292 11023 35528
rect 11259 35292 11349 35528
rect 11585 35292 11675 35528
rect 11911 35292 12001 35528
rect 12237 35292 12327 35528
rect 12563 35292 12653 35528
rect 12889 35292 12979 35528
rect 13215 35292 13305 35528
rect 13541 35292 13631 35528
rect 13867 35292 13957 35528
rect 14193 35292 14283 35528
rect 14519 35292 14609 35528
rect 14845 35292 15000 35528
rect 0 35204 15000 35292
rect 0 34968 241 35204
rect 477 34968 568 35204
rect 804 34968 895 35204
rect 1131 34968 1222 35204
rect 1458 34968 1549 35204
rect 1785 34968 1876 35204
rect 2112 34968 2203 35204
rect 2439 34968 2530 35204
rect 2766 34968 2857 35204
rect 3093 34968 3184 35204
rect 3420 34968 3511 35204
rect 3747 34968 3838 35204
rect 4074 34968 4165 35204
rect 4401 34968 4492 35204
rect 4728 34968 4819 35204
rect 5055 34968 5146 35204
rect 5382 34968 5473 35204
rect 5709 34968 5800 35204
rect 6036 34968 6127 35204
rect 6363 34968 6454 35204
rect 6690 34968 6781 35204
rect 7017 34968 7108 35204
rect 7344 34968 7435 35204
rect 7671 34968 7762 35204
rect 7998 34968 8089 35204
rect 8325 34968 8415 35204
rect 8651 34968 8741 35204
rect 8977 34968 9067 35204
rect 9303 34968 9393 35204
rect 9629 34968 9719 35204
rect 9955 34968 10045 35204
rect 10281 34968 10371 35204
rect 10607 34968 10697 35204
rect 10933 34968 11023 35204
rect 11259 34968 11349 35204
rect 11585 34968 11675 35204
rect 11911 34968 12001 35204
rect 12237 34968 12327 35204
rect 12563 34968 12653 35204
rect 12889 34968 12979 35204
rect 13215 34968 13305 35204
rect 13541 34968 13631 35204
rect 13867 34968 13957 35204
rect 14193 34968 14283 35204
rect 14519 34968 14609 35204
rect 14845 34968 15000 35204
rect 0 34880 15000 34968
rect 0 34644 241 34880
rect 477 34644 568 34880
rect 804 34644 895 34880
rect 1131 34644 1222 34880
rect 1458 34644 1549 34880
rect 1785 34644 1876 34880
rect 2112 34644 2203 34880
rect 2439 34644 2530 34880
rect 2766 34644 2857 34880
rect 3093 34644 3184 34880
rect 3420 34644 3511 34880
rect 3747 34644 3838 34880
rect 4074 34644 4165 34880
rect 4401 34644 4492 34880
rect 4728 34644 4819 34880
rect 5055 34644 5146 34880
rect 5382 34644 5473 34880
rect 5709 34644 5800 34880
rect 6036 34644 6127 34880
rect 6363 34644 6454 34880
rect 6690 34644 6781 34880
rect 7017 34644 7108 34880
rect 7344 34644 7435 34880
rect 7671 34644 7762 34880
rect 7998 34644 8089 34880
rect 8325 34644 8415 34880
rect 8651 34644 8741 34880
rect 8977 34644 9067 34880
rect 9303 34644 9393 34880
rect 9629 34644 9719 34880
rect 9955 34644 10045 34880
rect 10281 34644 10371 34880
rect 10607 34644 10697 34880
rect 10933 34644 11023 34880
rect 11259 34644 11349 34880
rect 11585 34644 11675 34880
rect 11911 34644 12001 34880
rect 12237 34644 12327 34880
rect 12563 34644 12653 34880
rect 12889 34644 12979 34880
rect 13215 34644 13305 34880
rect 13541 34644 13631 34880
rect 13867 34644 13957 34880
rect 14193 34644 14283 34880
rect 14519 34644 14609 34880
rect 14845 34644 15000 34880
rect 0 34609 15000 34644
rect 0 34608 254 34609
rect 14746 34608 15000 34609
rect 0 18423 15000 18448
rect 0 18187 143 18423
rect 379 18187 465 18423
rect 701 18187 787 18423
rect 1023 18187 1109 18423
rect 1345 18187 1431 18423
rect 1667 18187 1753 18423
rect 1989 18187 2075 18423
rect 2311 18187 2397 18423
rect 2633 18187 2719 18423
rect 2955 18187 3041 18423
rect 3277 18187 3363 18423
rect 3599 18187 3685 18423
rect 3921 18187 4007 18423
rect 4243 18187 4329 18423
rect 4565 18187 4651 18423
rect 4887 18187 4973 18423
rect 5209 18187 5295 18423
rect 5531 18187 5617 18423
rect 5853 18187 5938 18423
rect 6174 18187 6259 18423
rect 6495 18187 6580 18423
rect 6816 18187 6901 18423
rect 7137 18187 7222 18423
rect 7458 18187 7543 18423
rect 7779 18187 7864 18423
rect 8100 18187 8185 18423
rect 8421 18187 8506 18423
rect 8742 18187 8827 18423
rect 9063 18187 9148 18423
rect 9384 18187 9469 18423
rect 9705 18187 9790 18423
rect 10026 18187 10111 18423
rect 10347 18187 10432 18423
rect 10668 18187 10753 18423
rect 10989 18187 11074 18423
rect 11310 18187 11395 18423
rect 11631 18187 11716 18423
rect 11952 18187 12037 18423
rect 12273 18187 12358 18423
rect 12594 18187 12679 18423
rect 12915 18187 13000 18423
rect 13236 18187 13321 18423
rect 13557 18187 13642 18423
rect 13878 18187 13963 18423
rect 14199 18187 14284 18423
rect 14520 18187 14605 18423
rect 14841 18187 15000 18423
rect 0 18087 15000 18187
rect 0 17851 143 18087
rect 379 17851 465 18087
rect 701 17851 787 18087
rect 1023 17851 1109 18087
rect 1345 17851 1431 18087
rect 1667 17851 1753 18087
rect 1989 17851 2075 18087
rect 2311 17851 2397 18087
rect 2633 17851 2719 18087
rect 2955 17851 3041 18087
rect 3277 17851 3363 18087
rect 3599 17851 3685 18087
rect 3921 17851 4007 18087
rect 4243 17851 4329 18087
rect 4565 17851 4651 18087
rect 4887 17851 4973 18087
rect 5209 17851 5295 18087
rect 5531 17851 5617 18087
rect 5853 17851 5938 18087
rect 6174 17851 6259 18087
rect 6495 17851 6580 18087
rect 6816 17851 6901 18087
rect 7137 17851 7222 18087
rect 7458 17851 7543 18087
rect 7779 17851 7864 18087
rect 8100 17851 8185 18087
rect 8421 17851 8506 18087
rect 8742 17851 8827 18087
rect 9063 17851 9148 18087
rect 9384 17851 9469 18087
rect 9705 17851 9790 18087
rect 10026 17851 10111 18087
rect 10347 17851 10432 18087
rect 10668 17851 10753 18087
rect 10989 17851 11074 18087
rect 11310 17851 11395 18087
rect 11631 17851 11716 18087
rect 11952 17851 12037 18087
rect 12273 17851 12358 18087
rect 12594 17851 12679 18087
rect 12915 17851 13000 18087
rect 13236 17851 13321 18087
rect 13557 17851 13642 18087
rect 13878 17851 13963 18087
rect 14199 17851 14284 18087
rect 14520 17851 14605 18087
rect 14841 17851 15000 18087
rect 0 17751 15000 17851
rect 0 17515 143 17751
rect 379 17515 465 17751
rect 701 17515 787 17751
rect 1023 17515 1109 17751
rect 1345 17515 1431 17751
rect 1667 17515 1753 17751
rect 1989 17515 2075 17751
rect 2311 17515 2397 17751
rect 2633 17515 2719 17751
rect 2955 17515 3041 17751
rect 3277 17515 3363 17751
rect 3599 17515 3685 17751
rect 3921 17515 4007 17751
rect 4243 17515 4329 17751
rect 4565 17515 4651 17751
rect 4887 17515 4973 17751
rect 5209 17515 5295 17751
rect 5531 17515 5617 17751
rect 5853 17515 5938 17751
rect 6174 17515 6259 17751
rect 6495 17515 6580 17751
rect 6816 17515 6901 17751
rect 7137 17515 7222 17751
rect 7458 17515 7543 17751
rect 7779 17515 7864 17751
rect 8100 17515 8185 17751
rect 8421 17515 8506 17751
rect 8742 17515 8827 17751
rect 9063 17515 9148 17751
rect 9384 17515 9469 17751
rect 9705 17515 9790 17751
rect 10026 17515 10111 17751
rect 10347 17515 10432 17751
rect 10668 17515 10753 17751
rect 10989 17515 11074 17751
rect 11310 17515 11395 17751
rect 11631 17515 11716 17751
rect 11952 17515 12037 17751
rect 12273 17515 12358 17751
rect 12594 17515 12679 17751
rect 12915 17515 13000 17751
rect 13236 17515 13321 17751
rect 13557 17515 13642 17751
rect 13878 17515 13963 17751
rect 14199 17515 14284 17751
rect 14520 17515 14605 17751
rect 14841 17515 15000 17751
rect 0 17415 15000 17515
rect 0 17179 143 17415
rect 379 17179 465 17415
rect 701 17179 787 17415
rect 1023 17179 1109 17415
rect 1345 17179 1431 17415
rect 1667 17179 1753 17415
rect 1989 17179 2075 17415
rect 2311 17179 2397 17415
rect 2633 17179 2719 17415
rect 2955 17179 3041 17415
rect 3277 17179 3363 17415
rect 3599 17179 3685 17415
rect 3921 17179 4007 17415
rect 4243 17179 4329 17415
rect 4565 17179 4651 17415
rect 4887 17179 4973 17415
rect 5209 17179 5295 17415
rect 5531 17179 5617 17415
rect 5853 17179 5938 17415
rect 6174 17179 6259 17415
rect 6495 17179 6580 17415
rect 6816 17179 6901 17415
rect 7137 17179 7222 17415
rect 7458 17179 7543 17415
rect 7779 17179 7864 17415
rect 8100 17179 8185 17415
rect 8421 17179 8506 17415
rect 8742 17179 8827 17415
rect 9063 17179 9148 17415
rect 9384 17179 9469 17415
rect 9705 17179 9790 17415
rect 10026 17179 10111 17415
rect 10347 17179 10432 17415
rect 10668 17179 10753 17415
rect 10989 17179 11074 17415
rect 11310 17179 11395 17415
rect 11631 17179 11716 17415
rect 11952 17179 12037 17415
rect 12273 17179 12358 17415
rect 12594 17179 12679 17415
rect 12915 17179 13000 17415
rect 13236 17179 13321 17415
rect 13557 17179 13642 17415
rect 13878 17179 13963 17415
rect 14199 17179 14284 17415
rect 14520 17179 14605 17415
rect 14841 17179 15000 17415
rect 0 17079 15000 17179
rect 0 16843 143 17079
rect 379 16843 465 17079
rect 701 16843 787 17079
rect 1023 16843 1109 17079
rect 1345 16843 1431 17079
rect 1667 16843 1753 17079
rect 1989 16843 2075 17079
rect 2311 16843 2397 17079
rect 2633 16843 2719 17079
rect 2955 16843 3041 17079
rect 3277 16843 3363 17079
rect 3599 16843 3685 17079
rect 3921 16843 4007 17079
rect 4243 16843 4329 17079
rect 4565 16843 4651 17079
rect 4887 16843 4973 17079
rect 5209 16843 5295 17079
rect 5531 16843 5617 17079
rect 5853 16843 5938 17079
rect 6174 16843 6259 17079
rect 6495 16843 6580 17079
rect 6816 16843 6901 17079
rect 7137 16843 7222 17079
rect 7458 16843 7543 17079
rect 7779 16843 7864 17079
rect 8100 16843 8185 17079
rect 8421 16843 8506 17079
rect 8742 16843 8827 17079
rect 9063 16843 9148 17079
rect 9384 16843 9469 17079
rect 9705 16843 9790 17079
rect 10026 16843 10111 17079
rect 10347 16843 10432 17079
rect 10668 16843 10753 17079
rect 10989 16843 11074 17079
rect 11310 16843 11395 17079
rect 11631 16843 11716 17079
rect 11952 16843 12037 17079
rect 12273 16843 12358 17079
rect 12594 16843 12679 17079
rect 12915 16843 13000 17079
rect 13236 16843 13321 17079
rect 13557 16843 13642 17079
rect 13878 16843 13963 17079
rect 14199 16843 14284 17079
rect 14520 16843 14605 17079
rect 14841 16843 15000 17079
rect 0 16743 15000 16843
rect 0 16507 143 16743
rect 379 16507 465 16743
rect 701 16507 787 16743
rect 1023 16507 1109 16743
rect 1345 16507 1431 16743
rect 1667 16507 1753 16743
rect 1989 16507 2075 16743
rect 2311 16507 2397 16743
rect 2633 16507 2719 16743
rect 2955 16507 3041 16743
rect 3277 16507 3363 16743
rect 3599 16507 3685 16743
rect 3921 16507 4007 16743
rect 4243 16507 4329 16743
rect 4565 16507 4651 16743
rect 4887 16507 4973 16743
rect 5209 16507 5295 16743
rect 5531 16507 5617 16743
rect 5853 16507 5938 16743
rect 6174 16507 6259 16743
rect 6495 16507 6580 16743
rect 6816 16507 6901 16743
rect 7137 16507 7222 16743
rect 7458 16507 7543 16743
rect 7779 16507 7864 16743
rect 8100 16507 8185 16743
rect 8421 16507 8506 16743
rect 8742 16507 8827 16743
rect 9063 16507 9148 16743
rect 9384 16507 9469 16743
rect 9705 16507 9790 16743
rect 10026 16507 10111 16743
rect 10347 16507 10432 16743
rect 10668 16507 10753 16743
rect 10989 16507 11074 16743
rect 11310 16507 11395 16743
rect 11631 16507 11716 16743
rect 11952 16507 12037 16743
rect 12273 16507 12358 16743
rect 12594 16507 12679 16743
rect 12915 16507 13000 16743
rect 13236 16507 13321 16743
rect 13557 16507 13642 16743
rect 13878 16507 13963 16743
rect 14199 16507 14284 16743
rect 14520 16507 14605 16743
rect 14841 16507 15000 16743
rect 0 16407 15000 16507
rect 0 16171 143 16407
rect 379 16171 465 16407
rect 701 16171 787 16407
rect 1023 16171 1109 16407
rect 1345 16171 1431 16407
rect 1667 16171 1753 16407
rect 1989 16171 2075 16407
rect 2311 16171 2397 16407
rect 2633 16171 2719 16407
rect 2955 16171 3041 16407
rect 3277 16171 3363 16407
rect 3599 16171 3685 16407
rect 3921 16171 4007 16407
rect 4243 16171 4329 16407
rect 4565 16171 4651 16407
rect 4887 16171 4973 16407
rect 5209 16171 5295 16407
rect 5531 16171 5617 16407
rect 5853 16171 5938 16407
rect 6174 16171 6259 16407
rect 6495 16171 6580 16407
rect 6816 16171 6901 16407
rect 7137 16171 7222 16407
rect 7458 16171 7543 16407
rect 7779 16171 7864 16407
rect 8100 16171 8185 16407
rect 8421 16171 8506 16407
rect 8742 16171 8827 16407
rect 9063 16171 9148 16407
rect 9384 16171 9469 16407
rect 9705 16171 9790 16407
rect 10026 16171 10111 16407
rect 10347 16171 10432 16407
rect 10668 16171 10753 16407
rect 10989 16171 11074 16407
rect 11310 16171 11395 16407
rect 11631 16171 11716 16407
rect 11952 16171 12037 16407
rect 12273 16171 12358 16407
rect 12594 16171 12679 16407
rect 12915 16171 13000 16407
rect 13236 16171 13321 16407
rect 13557 16171 13642 16407
rect 13878 16171 13963 16407
rect 14199 16171 14284 16407
rect 14520 16171 14605 16407
rect 14841 16171 15000 16407
rect 0 16071 15000 16171
rect 0 15835 143 16071
rect 379 15835 465 16071
rect 701 15835 787 16071
rect 1023 15835 1109 16071
rect 1345 15835 1431 16071
rect 1667 15835 1753 16071
rect 1989 15835 2075 16071
rect 2311 15835 2397 16071
rect 2633 15835 2719 16071
rect 2955 15835 3041 16071
rect 3277 15835 3363 16071
rect 3599 15835 3685 16071
rect 3921 15835 4007 16071
rect 4243 15835 4329 16071
rect 4565 15835 4651 16071
rect 4887 15835 4973 16071
rect 5209 15835 5295 16071
rect 5531 15835 5617 16071
rect 5853 15835 5938 16071
rect 6174 15835 6259 16071
rect 6495 15835 6580 16071
rect 6816 15835 6901 16071
rect 7137 15835 7222 16071
rect 7458 15835 7543 16071
rect 7779 15835 7864 16071
rect 8100 15835 8185 16071
rect 8421 15835 8506 16071
rect 8742 15835 8827 16071
rect 9063 15835 9148 16071
rect 9384 15835 9469 16071
rect 9705 15835 9790 16071
rect 10026 15835 10111 16071
rect 10347 15835 10432 16071
rect 10668 15835 10753 16071
rect 10989 15835 11074 16071
rect 11310 15835 11395 16071
rect 11631 15835 11716 16071
rect 11952 15835 12037 16071
rect 12273 15835 12358 16071
rect 12594 15835 12679 16071
rect 12915 15835 13000 16071
rect 13236 15835 13321 16071
rect 13557 15835 13642 16071
rect 13878 15835 13963 16071
rect 14199 15835 14284 16071
rect 14520 15835 14605 16071
rect 14841 15835 15000 16071
rect 0 15735 15000 15835
rect 0 15499 143 15735
rect 379 15499 465 15735
rect 701 15499 787 15735
rect 1023 15499 1109 15735
rect 1345 15499 1431 15735
rect 1667 15499 1753 15735
rect 1989 15499 2075 15735
rect 2311 15499 2397 15735
rect 2633 15499 2719 15735
rect 2955 15499 3041 15735
rect 3277 15499 3363 15735
rect 3599 15499 3685 15735
rect 3921 15499 4007 15735
rect 4243 15499 4329 15735
rect 4565 15499 4651 15735
rect 4887 15499 4973 15735
rect 5209 15499 5295 15735
rect 5531 15499 5617 15735
rect 5853 15499 5938 15735
rect 6174 15499 6259 15735
rect 6495 15499 6580 15735
rect 6816 15499 6901 15735
rect 7137 15499 7222 15735
rect 7458 15499 7543 15735
rect 7779 15499 7864 15735
rect 8100 15499 8185 15735
rect 8421 15499 8506 15735
rect 8742 15499 8827 15735
rect 9063 15499 9148 15735
rect 9384 15499 9469 15735
rect 9705 15499 9790 15735
rect 10026 15499 10111 15735
rect 10347 15499 10432 15735
rect 10668 15499 10753 15735
rect 10989 15499 11074 15735
rect 11310 15499 11395 15735
rect 11631 15499 11716 15735
rect 11952 15499 12037 15735
rect 12273 15499 12358 15735
rect 12594 15499 12679 15735
rect 12915 15499 13000 15735
rect 13236 15499 13321 15735
rect 13557 15499 13642 15735
rect 13878 15499 13963 15735
rect 14199 15499 14284 15735
rect 14520 15499 14605 15735
rect 14841 15499 15000 15735
rect 0 15399 15000 15499
rect 0 15163 143 15399
rect 379 15163 465 15399
rect 701 15163 787 15399
rect 1023 15163 1109 15399
rect 1345 15163 1431 15399
rect 1667 15163 1753 15399
rect 1989 15163 2075 15399
rect 2311 15163 2397 15399
rect 2633 15163 2719 15399
rect 2955 15163 3041 15399
rect 3277 15163 3363 15399
rect 3599 15163 3685 15399
rect 3921 15163 4007 15399
rect 4243 15163 4329 15399
rect 4565 15163 4651 15399
rect 4887 15163 4973 15399
rect 5209 15163 5295 15399
rect 5531 15163 5617 15399
rect 5853 15163 5938 15399
rect 6174 15163 6259 15399
rect 6495 15163 6580 15399
rect 6816 15163 6901 15399
rect 7137 15163 7222 15399
rect 7458 15163 7543 15399
rect 7779 15163 7864 15399
rect 8100 15163 8185 15399
rect 8421 15163 8506 15399
rect 8742 15163 8827 15399
rect 9063 15163 9148 15399
rect 9384 15163 9469 15399
rect 9705 15163 9790 15399
rect 10026 15163 10111 15399
rect 10347 15163 10432 15399
rect 10668 15163 10753 15399
rect 10989 15163 11074 15399
rect 11310 15163 11395 15399
rect 11631 15163 11716 15399
rect 11952 15163 12037 15399
rect 12273 15163 12358 15399
rect 12594 15163 12679 15399
rect 12915 15163 13000 15399
rect 13236 15163 13321 15399
rect 13557 15163 13642 15399
rect 13878 15163 13963 15399
rect 14199 15163 14284 15399
rect 14520 15163 14605 15399
rect 14841 15163 15000 15399
rect 0 15063 15000 15163
rect 0 14827 143 15063
rect 379 14827 465 15063
rect 701 14827 787 15063
rect 1023 14827 1109 15063
rect 1345 14827 1431 15063
rect 1667 14827 1753 15063
rect 1989 14827 2075 15063
rect 2311 14827 2397 15063
rect 2633 14827 2719 15063
rect 2955 14827 3041 15063
rect 3277 14827 3363 15063
rect 3599 14827 3685 15063
rect 3921 14827 4007 15063
rect 4243 14827 4329 15063
rect 4565 14827 4651 15063
rect 4887 14827 4973 15063
rect 5209 14827 5295 15063
rect 5531 14827 5617 15063
rect 5853 14827 5938 15063
rect 6174 14827 6259 15063
rect 6495 14827 6580 15063
rect 6816 14827 6901 15063
rect 7137 14827 7222 15063
rect 7458 14827 7543 15063
rect 7779 14827 7864 15063
rect 8100 14827 8185 15063
rect 8421 14827 8506 15063
rect 8742 14827 8827 15063
rect 9063 14827 9148 15063
rect 9384 14827 9469 15063
rect 9705 14827 9790 15063
rect 10026 14827 10111 15063
rect 10347 14827 10432 15063
rect 10668 14827 10753 15063
rect 10989 14827 11074 15063
rect 11310 14827 11395 15063
rect 11631 14827 11716 15063
rect 11952 14827 12037 15063
rect 12273 14827 12358 15063
rect 12594 14827 12679 15063
rect 12915 14827 13000 15063
rect 13236 14827 13321 15063
rect 13557 14827 13642 15063
rect 13878 14827 13963 15063
rect 14199 14827 14284 15063
rect 14520 14827 14605 15063
rect 14841 14827 15000 15063
rect 0 14727 15000 14827
rect 0 14491 143 14727
rect 379 14491 465 14727
rect 701 14491 787 14727
rect 1023 14491 1109 14727
rect 1345 14491 1431 14727
rect 1667 14491 1753 14727
rect 1989 14491 2075 14727
rect 2311 14491 2397 14727
rect 2633 14491 2719 14727
rect 2955 14491 3041 14727
rect 3277 14491 3363 14727
rect 3599 14491 3685 14727
rect 3921 14491 4007 14727
rect 4243 14491 4329 14727
rect 4565 14491 4651 14727
rect 4887 14491 4973 14727
rect 5209 14491 5295 14727
rect 5531 14491 5617 14727
rect 5853 14491 5938 14727
rect 6174 14491 6259 14727
rect 6495 14491 6580 14727
rect 6816 14491 6901 14727
rect 7137 14491 7222 14727
rect 7458 14491 7543 14727
rect 7779 14491 7864 14727
rect 8100 14491 8185 14727
rect 8421 14491 8506 14727
rect 8742 14491 8827 14727
rect 9063 14491 9148 14727
rect 9384 14491 9469 14727
rect 9705 14491 9790 14727
rect 10026 14491 10111 14727
rect 10347 14491 10432 14727
rect 10668 14491 10753 14727
rect 10989 14491 11074 14727
rect 11310 14491 11395 14727
rect 11631 14491 11716 14727
rect 11952 14491 12037 14727
rect 12273 14491 12358 14727
rect 12594 14491 12679 14727
rect 12915 14491 13000 14727
rect 13236 14491 13321 14727
rect 13557 14491 13642 14727
rect 13878 14491 13963 14727
rect 14199 14491 14284 14727
rect 14520 14491 14605 14727
rect 14841 14491 15000 14727
rect 0 14391 15000 14491
rect 0 14155 143 14391
rect 379 14155 465 14391
rect 701 14155 787 14391
rect 1023 14155 1109 14391
rect 1345 14155 1431 14391
rect 1667 14155 1753 14391
rect 1989 14155 2075 14391
rect 2311 14155 2397 14391
rect 2633 14155 2719 14391
rect 2955 14155 3041 14391
rect 3277 14155 3363 14391
rect 3599 14155 3685 14391
rect 3921 14155 4007 14391
rect 4243 14155 4329 14391
rect 4565 14155 4651 14391
rect 4887 14155 4973 14391
rect 5209 14155 5295 14391
rect 5531 14155 5617 14391
rect 5853 14155 5938 14391
rect 6174 14155 6259 14391
rect 6495 14155 6580 14391
rect 6816 14155 6901 14391
rect 7137 14155 7222 14391
rect 7458 14155 7543 14391
rect 7779 14155 7864 14391
rect 8100 14155 8185 14391
rect 8421 14155 8506 14391
rect 8742 14155 8827 14391
rect 9063 14155 9148 14391
rect 9384 14155 9469 14391
rect 9705 14155 9790 14391
rect 10026 14155 10111 14391
rect 10347 14155 10432 14391
rect 10668 14155 10753 14391
rect 10989 14155 11074 14391
rect 11310 14155 11395 14391
rect 11631 14155 11716 14391
rect 11952 14155 12037 14391
rect 12273 14155 12358 14391
rect 12594 14155 12679 14391
rect 12915 14155 13000 14391
rect 13236 14155 13321 14391
rect 13557 14155 13642 14391
rect 13878 14155 13963 14391
rect 14199 14155 14284 14391
rect 14520 14155 14605 14391
rect 14841 14155 15000 14391
rect 0 14055 15000 14155
rect 0 13819 143 14055
rect 379 13819 465 14055
rect 701 13819 787 14055
rect 1023 13819 1109 14055
rect 1345 13819 1431 14055
rect 1667 13819 1753 14055
rect 1989 13819 2075 14055
rect 2311 13819 2397 14055
rect 2633 13819 2719 14055
rect 2955 13819 3041 14055
rect 3277 13819 3363 14055
rect 3599 13819 3685 14055
rect 3921 13819 4007 14055
rect 4243 13819 4329 14055
rect 4565 13819 4651 14055
rect 4887 13819 4973 14055
rect 5209 13819 5295 14055
rect 5531 13819 5617 14055
rect 5853 13819 5938 14055
rect 6174 13819 6259 14055
rect 6495 13819 6580 14055
rect 6816 13819 6901 14055
rect 7137 13819 7222 14055
rect 7458 13819 7543 14055
rect 7779 13819 7864 14055
rect 8100 13819 8185 14055
rect 8421 13819 8506 14055
rect 8742 13819 8827 14055
rect 9063 13819 9148 14055
rect 9384 13819 9469 14055
rect 9705 13819 9790 14055
rect 10026 13819 10111 14055
rect 10347 13819 10432 14055
rect 10668 13819 10753 14055
rect 10989 13819 11074 14055
rect 11310 13819 11395 14055
rect 11631 13819 11716 14055
rect 11952 13819 12037 14055
rect 12273 13819 12358 14055
rect 12594 13819 12679 14055
rect 12915 13819 13000 14055
rect 13236 13819 13321 14055
rect 13557 13819 13642 14055
rect 13878 13819 13963 14055
rect 14199 13819 14284 14055
rect 14520 13819 14605 14055
rect 14841 13819 15000 14055
rect 0 13719 15000 13819
rect 0 13483 143 13719
rect 379 13483 465 13719
rect 701 13483 787 13719
rect 1023 13483 1109 13719
rect 1345 13483 1431 13719
rect 1667 13483 1753 13719
rect 1989 13483 2075 13719
rect 2311 13483 2397 13719
rect 2633 13483 2719 13719
rect 2955 13483 3041 13719
rect 3277 13483 3363 13719
rect 3599 13483 3685 13719
rect 3921 13483 4007 13719
rect 4243 13483 4329 13719
rect 4565 13483 4651 13719
rect 4887 13483 4973 13719
rect 5209 13483 5295 13719
rect 5531 13483 5617 13719
rect 5853 13483 5938 13719
rect 6174 13483 6259 13719
rect 6495 13483 6580 13719
rect 6816 13483 6901 13719
rect 7137 13483 7222 13719
rect 7458 13483 7543 13719
rect 7779 13483 7864 13719
rect 8100 13483 8185 13719
rect 8421 13483 8506 13719
rect 8742 13483 8827 13719
rect 9063 13483 9148 13719
rect 9384 13483 9469 13719
rect 9705 13483 9790 13719
rect 10026 13483 10111 13719
rect 10347 13483 10432 13719
rect 10668 13483 10753 13719
rect 10989 13483 11074 13719
rect 11310 13483 11395 13719
rect 11631 13483 11716 13719
rect 11952 13483 12037 13719
rect 12273 13483 12358 13719
rect 12594 13483 12679 13719
rect 12915 13483 13000 13719
rect 13236 13483 13321 13719
rect 13557 13483 13642 13719
rect 13878 13483 13963 13719
rect 14199 13483 14284 13719
rect 14520 13483 14605 13719
rect 14841 13483 15000 13719
rect 0 13458 15000 13483
rect 0 13114 15000 13138
rect 0 12878 143 13114
rect 379 12878 465 13114
rect 701 12878 787 13114
rect 1023 12878 1109 13114
rect 1345 12878 1431 13114
rect 1667 12878 1753 13114
rect 1989 12878 2075 13114
rect 2311 12878 2397 13114
rect 2633 12878 2719 13114
rect 2955 12878 3041 13114
rect 3277 12878 3363 13114
rect 3599 12878 3685 13114
rect 3921 12878 4007 13114
rect 4243 12878 4329 13114
rect 4565 12878 4651 13114
rect 4887 12878 4973 13114
rect 5209 12878 5294 13114
rect 5530 12878 5615 13114
rect 5851 12878 5936 13114
rect 6172 12878 6257 13114
rect 6493 12878 6578 13114
rect 6814 12878 6899 13114
rect 7135 12878 7220 13114
rect 7456 12878 7541 13114
rect 7777 12878 7862 13114
rect 8098 12878 8183 13114
rect 8419 12878 8504 13114
rect 8740 12878 8825 13114
rect 9061 12878 9146 13114
rect 9382 12878 9467 13114
rect 9703 12878 9788 13114
rect 10024 12878 10109 13114
rect 10345 12878 10430 13114
rect 10666 12878 10751 13114
rect 10987 12878 11072 13114
rect 11308 12878 11393 13114
rect 11629 12878 11714 13114
rect 11950 12878 12035 13114
rect 12271 12878 12356 13114
rect 12592 12878 12677 13114
rect 12913 12878 12998 13114
rect 13234 12878 13319 13114
rect 13555 12878 13640 13114
rect 13876 12878 13961 13114
rect 14197 12878 14282 13114
rect 14518 12878 14603 13114
rect 14839 12878 15000 13114
rect 0 12548 15000 12878
rect 0 12312 143 12548
rect 379 12312 465 12548
rect 701 12312 787 12548
rect 1023 12312 1109 12548
rect 1345 12312 1431 12548
rect 1667 12312 1753 12548
rect 1989 12312 2075 12548
rect 2311 12312 2397 12548
rect 2633 12312 2719 12548
rect 2955 12312 3041 12548
rect 3277 12312 3363 12548
rect 3599 12312 3685 12548
rect 3921 12312 4007 12548
rect 4243 12312 4329 12548
rect 4565 12312 4651 12548
rect 4887 12312 4973 12548
rect 5209 12312 5294 12548
rect 5530 12312 5615 12548
rect 5851 12312 5936 12548
rect 6172 12312 6257 12548
rect 6493 12312 6578 12548
rect 6814 12312 6899 12548
rect 7135 12312 7220 12548
rect 7456 12312 7541 12548
rect 7777 12312 7862 12548
rect 8098 12312 8183 12548
rect 8419 12312 8504 12548
rect 8740 12312 8825 12548
rect 9061 12312 9146 12548
rect 9382 12312 9467 12548
rect 9703 12312 9788 12548
rect 10024 12312 10109 12548
rect 10345 12312 10430 12548
rect 10666 12312 10751 12548
rect 10987 12312 11072 12548
rect 11308 12312 11393 12548
rect 11629 12312 11714 12548
rect 11950 12312 12035 12548
rect 12271 12312 12356 12548
rect 12592 12312 12677 12548
rect 12913 12312 12998 12548
rect 13234 12312 13319 12548
rect 13555 12312 13640 12548
rect 13876 12312 13961 12548
rect 14197 12312 14282 12548
rect 14518 12312 14603 12548
rect 14839 12312 15000 12548
rect 0 12288 15000 12312
rect 0 11944 15000 11968
rect 0 11708 143 11944
rect 379 11708 465 11944
rect 701 11708 787 11944
rect 1023 11708 1109 11944
rect 1345 11708 1431 11944
rect 1667 11708 1753 11944
rect 1989 11708 2075 11944
rect 2311 11708 2397 11944
rect 2633 11708 2719 11944
rect 2955 11708 3041 11944
rect 3277 11708 3363 11944
rect 3599 11708 3685 11944
rect 3921 11708 4007 11944
rect 4243 11708 4329 11944
rect 4565 11708 4651 11944
rect 4887 11708 4973 11944
rect 5209 11708 5294 11944
rect 5530 11708 5615 11944
rect 5851 11708 5936 11944
rect 6172 11708 6257 11944
rect 6493 11708 6578 11944
rect 6814 11708 6899 11944
rect 7135 11708 7220 11944
rect 7456 11708 7541 11944
rect 7777 11708 7862 11944
rect 8098 11708 8183 11944
rect 8419 11708 8504 11944
rect 8740 11708 8825 11944
rect 9061 11708 9146 11944
rect 9382 11708 9467 11944
rect 9703 11708 9788 11944
rect 10024 11708 10109 11944
rect 10345 11708 10430 11944
rect 10666 11708 10751 11944
rect 10987 11708 11072 11944
rect 11308 11708 11393 11944
rect 11629 11708 11714 11944
rect 11950 11708 12035 11944
rect 12271 11708 12356 11944
rect 12592 11708 12677 11944
rect 12913 11708 12998 11944
rect 13234 11708 13319 11944
rect 13555 11708 13640 11944
rect 13876 11708 13961 11944
rect 14197 11708 14282 11944
rect 14518 11708 14603 11944
rect 14839 11708 15000 11944
rect 0 11378 15000 11708
rect 0 11142 143 11378
rect 379 11142 465 11378
rect 701 11142 787 11378
rect 1023 11142 1109 11378
rect 1345 11142 1431 11378
rect 1667 11142 1753 11378
rect 1989 11142 2075 11378
rect 2311 11142 2397 11378
rect 2633 11142 2719 11378
rect 2955 11142 3041 11378
rect 3277 11142 3363 11378
rect 3599 11142 3685 11378
rect 3921 11142 4007 11378
rect 4243 11142 4329 11378
rect 4565 11142 4651 11378
rect 4887 11142 4973 11378
rect 5209 11142 5294 11378
rect 5530 11142 5615 11378
rect 5851 11142 5936 11378
rect 6172 11142 6257 11378
rect 6493 11142 6578 11378
rect 6814 11142 6899 11378
rect 7135 11142 7220 11378
rect 7456 11142 7541 11378
rect 7777 11142 7862 11378
rect 8098 11142 8183 11378
rect 8419 11142 8504 11378
rect 8740 11142 8825 11378
rect 9061 11142 9146 11378
rect 9382 11142 9467 11378
rect 9703 11142 9788 11378
rect 10024 11142 10109 11378
rect 10345 11142 10430 11378
rect 10666 11142 10751 11378
rect 10987 11142 11072 11378
rect 11308 11142 11393 11378
rect 11629 11142 11714 11378
rect 11950 11142 12035 11378
rect 12271 11142 12356 11378
rect 12592 11142 12677 11378
rect 12913 11142 12998 11378
rect 13234 11142 13319 11378
rect 13555 11142 13640 11378
rect 13876 11142 13961 11378
rect 14197 11142 14282 11378
rect 14518 11142 14603 11378
rect 14839 11142 15000 11378
rect 0 11118 15000 11142
rect 0 8998 254 10798
rect 14746 8998 15000 10798
rect 0 8654 15000 8678
rect 0 8418 143 8654
rect 379 8418 465 8654
rect 701 8418 787 8654
rect 1023 8418 1109 8654
rect 1345 8418 1431 8654
rect 1667 8418 1753 8654
rect 1989 8418 2075 8654
rect 2311 8418 2397 8654
rect 2633 8418 2719 8654
rect 2955 8418 3041 8654
rect 3277 8418 3363 8654
rect 3599 8418 3685 8654
rect 3921 8418 4007 8654
rect 4243 8418 4329 8654
rect 4565 8418 4651 8654
rect 4887 8418 4973 8654
rect 5209 8418 5295 8654
rect 5531 8418 5617 8654
rect 5853 8418 5938 8654
rect 6174 8418 6259 8654
rect 6495 8418 6580 8654
rect 6816 8418 6901 8654
rect 7137 8418 7222 8654
rect 7458 8418 7543 8654
rect 7779 8418 7864 8654
rect 8100 8418 8185 8654
rect 8421 8418 8506 8654
rect 8742 8418 8827 8654
rect 9063 8418 9148 8654
rect 9384 8418 9469 8654
rect 9705 8418 9790 8654
rect 10026 8418 10111 8654
rect 10347 8418 10432 8654
rect 10668 8418 10753 8654
rect 10989 8418 11074 8654
rect 11310 8418 11395 8654
rect 11631 8418 11716 8654
rect 11952 8418 12037 8654
rect 12273 8418 12358 8654
rect 12594 8418 12679 8654
rect 12915 8418 13000 8654
rect 13236 8418 13321 8654
rect 13557 8418 13642 8654
rect 13878 8418 13963 8654
rect 14199 8418 14284 8654
rect 14520 8418 14605 8654
rect 14841 8418 15000 8654
rect 0 8048 15000 8418
rect 0 7812 143 8048
rect 379 7812 465 8048
rect 701 7812 787 8048
rect 1023 7812 1109 8048
rect 1345 7812 1431 8048
rect 1667 7812 1753 8048
rect 1989 7812 2075 8048
rect 2311 7812 2397 8048
rect 2633 7812 2719 8048
rect 2955 7812 3041 8048
rect 3277 7812 3363 8048
rect 3599 7812 3685 8048
rect 3921 7812 4007 8048
rect 4243 7812 4329 8048
rect 4565 7812 4651 8048
rect 4887 7812 4973 8048
rect 5209 7812 5295 8048
rect 5531 7812 5617 8048
rect 5853 7812 5938 8048
rect 6174 7812 6259 8048
rect 6495 7812 6580 8048
rect 6816 7812 6901 8048
rect 7137 7812 7222 8048
rect 7458 7812 7543 8048
rect 7779 7812 7864 8048
rect 8100 7812 8185 8048
rect 8421 7812 8506 8048
rect 8742 7812 8827 8048
rect 9063 7812 9148 8048
rect 9384 7812 9469 8048
rect 9705 7812 9790 8048
rect 10026 7812 10111 8048
rect 10347 7812 10432 8048
rect 10668 7812 10753 8048
rect 10989 7812 11074 8048
rect 11310 7812 11395 8048
rect 11631 7812 11716 8048
rect 11952 7812 12037 8048
rect 12273 7812 12358 8048
rect 12594 7812 12679 8048
rect 12915 7812 13000 8048
rect 13236 7812 13321 8048
rect 13557 7812 13642 8048
rect 13878 7812 13963 8048
rect 14199 7812 14284 8048
rect 14520 7812 14605 8048
rect 14841 7812 15000 8048
rect 0 7788 15000 7812
rect 0 7444 15000 7468
rect 0 7208 143 7444
rect 379 7208 465 7444
rect 701 7208 787 7444
rect 1023 7208 1109 7444
rect 1345 7208 1431 7444
rect 1667 7208 1753 7444
rect 1989 7208 2075 7444
rect 2311 7208 2397 7444
rect 2633 7208 2719 7444
rect 2955 7208 3041 7444
rect 3277 7208 3363 7444
rect 3599 7208 3685 7444
rect 3921 7208 4007 7444
rect 4243 7208 4329 7444
rect 4565 7208 4651 7444
rect 4887 7208 4973 7444
rect 5209 7208 5295 7444
rect 5531 7208 5617 7444
rect 5853 7208 5938 7444
rect 6174 7208 6259 7444
rect 6495 7208 6580 7444
rect 6816 7208 6901 7444
rect 7137 7208 7222 7444
rect 7458 7208 7543 7444
rect 7779 7208 7864 7444
rect 8100 7208 8185 7444
rect 8421 7208 8506 7444
rect 8742 7208 8827 7444
rect 9063 7208 9148 7444
rect 9384 7208 9469 7444
rect 9705 7208 9790 7444
rect 10026 7208 10111 7444
rect 10347 7208 10432 7444
rect 10668 7208 10753 7444
rect 10989 7208 11074 7444
rect 11310 7208 11395 7444
rect 11631 7208 11716 7444
rect 11952 7208 12037 7444
rect 12273 7208 12358 7444
rect 12594 7208 12679 7444
rect 12915 7208 13000 7444
rect 13236 7208 13321 7444
rect 13557 7208 13642 7444
rect 13878 7208 13963 7444
rect 14199 7208 14284 7444
rect 14520 7208 14605 7444
rect 14841 7208 15000 7444
rect 0 7078 15000 7208
rect 0 6842 143 7078
rect 379 6842 465 7078
rect 701 6842 787 7078
rect 1023 6842 1109 7078
rect 1345 6842 1431 7078
rect 1667 6842 1753 7078
rect 1989 6842 2075 7078
rect 2311 6842 2397 7078
rect 2633 6842 2719 7078
rect 2955 6842 3041 7078
rect 3277 6842 3363 7078
rect 3599 6842 3685 7078
rect 3921 6842 4007 7078
rect 4243 6842 4329 7078
rect 4565 6842 4651 7078
rect 4887 6842 4973 7078
rect 5209 6842 5295 7078
rect 5531 6842 5617 7078
rect 5853 6842 5938 7078
rect 6174 6842 6259 7078
rect 6495 6842 6580 7078
rect 6816 6842 6901 7078
rect 7137 6842 7222 7078
rect 7458 6842 7543 7078
rect 7779 6842 7864 7078
rect 8100 6842 8185 7078
rect 8421 6842 8506 7078
rect 8742 6842 8827 7078
rect 9063 6842 9148 7078
rect 9384 6842 9469 7078
rect 9705 6842 9790 7078
rect 10026 6842 10111 7078
rect 10347 6842 10432 7078
rect 10668 6842 10753 7078
rect 10989 6842 11074 7078
rect 11310 6842 11395 7078
rect 11631 6842 11716 7078
rect 11952 6842 12037 7078
rect 12273 6842 12358 7078
rect 12594 6842 12679 7078
rect 12915 6842 13000 7078
rect 13236 6842 13321 7078
rect 13557 6842 13642 7078
rect 13878 6842 13963 7078
rect 14199 6842 14284 7078
rect 14520 6842 14605 7078
rect 14841 6842 15000 7078
rect 0 6819 15000 6842
rect 119 6818 14865 6819
rect 0 6474 15000 6498
rect 0 6238 143 6474
rect 379 6238 465 6474
rect 701 6238 787 6474
rect 1023 6238 1109 6474
rect 1345 6238 1431 6474
rect 1667 6238 1753 6474
rect 1989 6238 2075 6474
rect 2311 6238 2397 6474
rect 2633 6238 2719 6474
rect 2955 6238 3041 6474
rect 3277 6238 3363 6474
rect 3599 6238 3685 6474
rect 3921 6238 4007 6474
rect 4243 6238 4329 6474
rect 4565 6238 4651 6474
rect 4887 6238 4973 6474
rect 5209 6238 5295 6474
rect 5531 6238 5617 6474
rect 5853 6238 5938 6474
rect 6174 6238 6259 6474
rect 6495 6238 6580 6474
rect 6816 6238 6901 6474
rect 7137 6238 7222 6474
rect 7458 6238 7543 6474
rect 7779 6238 7864 6474
rect 8100 6238 8185 6474
rect 8421 6238 8506 6474
rect 8742 6238 8827 6474
rect 9063 6238 9148 6474
rect 9384 6238 9469 6474
rect 9705 6238 9790 6474
rect 10026 6238 10111 6474
rect 10347 6238 10432 6474
rect 10668 6238 10753 6474
rect 10989 6238 11074 6474
rect 11310 6238 11395 6474
rect 11631 6238 11716 6474
rect 11952 6238 12037 6474
rect 12273 6238 12358 6474
rect 12594 6238 12679 6474
rect 12915 6238 13000 6474
rect 13236 6238 13321 6474
rect 13557 6238 13642 6474
rect 13878 6238 13963 6474
rect 14199 6238 14284 6474
rect 14520 6238 14605 6474
rect 14841 6238 15000 6474
rect 0 6108 15000 6238
rect 0 5872 143 6108
rect 379 5872 465 6108
rect 701 5872 787 6108
rect 1023 5872 1109 6108
rect 1345 5872 1431 6108
rect 1667 5872 1753 6108
rect 1989 5872 2075 6108
rect 2311 5872 2397 6108
rect 2633 5872 2719 6108
rect 2955 5872 3041 6108
rect 3277 5872 3363 6108
rect 3599 5872 3685 6108
rect 3921 5872 4007 6108
rect 4243 5872 4329 6108
rect 4565 5872 4651 6108
rect 4887 5872 4973 6108
rect 5209 5872 5295 6108
rect 5531 5872 5617 6108
rect 5853 5872 5938 6108
rect 6174 5872 6259 6108
rect 6495 5872 6580 6108
rect 6816 5872 6901 6108
rect 7137 5872 7222 6108
rect 7458 5872 7543 6108
rect 7779 5872 7864 6108
rect 8100 5872 8185 6108
rect 8421 5872 8506 6108
rect 8742 5872 8827 6108
rect 9063 5872 9148 6108
rect 9384 5872 9469 6108
rect 9705 5872 9790 6108
rect 10026 5872 10111 6108
rect 10347 5872 10432 6108
rect 10668 5872 10753 6108
rect 10989 5872 11074 6108
rect 11310 5872 11395 6108
rect 11631 5872 11716 6108
rect 11952 5872 12037 6108
rect 12273 5872 12358 6108
rect 12594 5872 12679 6108
rect 12915 5872 13000 6108
rect 13236 5872 13321 6108
rect 13557 5872 13642 6108
rect 13878 5872 13963 6108
rect 14199 5872 14284 6108
rect 14520 5872 14605 6108
rect 14841 5872 15000 6108
rect 0 5848 15000 5872
rect 0 5504 15000 5528
rect 0 5268 143 5504
rect 379 5268 465 5504
rect 701 5268 787 5504
rect 1023 5268 1109 5504
rect 1345 5268 1431 5504
rect 1667 5268 1753 5504
rect 1989 5268 2075 5504
rect 2311 5268 2397 5504
rect 2633 5268 2719 5504
rect 2955 5268 3041 5504
rect 3277 5268 3363 5504
rect 3599 5268 3685 5504
rect 3921 5268 4007 5504
rect 4243 5268 4329 5504
rect 4565 5268 4651 5504
rect 4887 5268 4973 5504
rect 5209 5268 5295 5504
rect 5531 5268 5617 5504
rect 5853 5268 5938 5504
rect 6174 5268 6259 5504
rect 6495 5268 6580 5504
rect 6816 5268 6901 5504
rect 7137 5268 7222 5504
rect 7458 5268 7543 5504
rect 7779 5268 7864 5504
rect 8100 5268 8185 5504
rect 8421 5268 8506 5504
rect 8742 5268 8827 5504
rect 9063 5268 9148 5504
rect 9384 5268 9469 5504
rect 9705 5268 9790 5504
rect 10026 5268 10111 5504
rect 10347 5268 10432 5504
rect 10668 5268 10753 5504
rect 10989 5268 11074 5504
rect 11310 5268 11395 5504
rect 11631 5268 11716 5504
rect 11952 5268 12037 5504
rect 12273 5268 12358 5504
rect 12594 5268 12679 5504
rect 12915 5268 13000 5504
rect 13236 5268 13321 5504
rect 13557 5268 13642 5504
rect 13878 5268 13963 5504
rect 14199 5268 14284 5504
rect 14520 5268 14605 5504
rect 14841 5268 15000 5504
rect 0 4898 15000 5268
rect 0 4662 143 4898
rect 379 4662 465 4898
rect 701 4662 787 4898
rect 1023 4662 1109 4898
rect 1345 4662 1431 4898
rect 1667 4662 1753 4898
rect 1989 4662 2075 4898
rect 2311 4662 2397 4898
rect 2633 4662 2719 4898
rect 2955 4662 3041 4898
rect 3277 4662 3363 4898
rect 3599 4662 3685 4898
rect 3921 4662 4007 4898
rect 4243 4662 4329 4898
rect 4565 4662 4651 4898
rect 4887 4662 4973 4898
rect 5209 4662 5295 4898
rect 5531 4662 5617 4898
rect 5853 4662 5938 4898
rect 6174 4662 6259 4898
rect 6495 4662 6580 4898
rect 6816 4662 6901 4898
rect 7137 4662 7222 4898
rect 7458 4662 7543 4898
rect 7779 4662 7864 4898
rect 8100 4662 8185 4898
rect 8421 4662 8506 4898
rect 8742 4662 8827 4898
rect 9063 4662 9148 4898
rect 9384 4662 9469 4898
rect 9705 4662 9790 4898
rect 10026 4662 10111 4898
rect 10347 4662 10432 4898
rect 10668 4662 10753 4898
rect 10989 4662 11074 4898
rect 11310 4662 11395 4898
rect 11631 4662 11716 4898
rect 11952 4662 12037 4898
rect 12273 4662 12358 4898
rect 12594 4662 12679 4898
rect 12915 4662 13000 4898
rect 13236 4662 13321 4898
rect 13557 4662 13642 4898
rect 13878 4662 13963 4898
rect 14199 4662 14284 4898
rect 14520 4662 14605 4898
rect 14841 4662 15000 4898
rect 0 4638 15000 4662
rect 0 4294 15000 4318
rect 0 4058 143 4294
rect 379 4058 465 4294
rect 701 4058 787 4294
rect 1023 4058 1109 4294
rect 1345 4058 1431 4294
rect 1667 4058 1753 4294
rect 1989 4058 2075 4294
rect 2311 4058 2397 4294
rect 2633 4058 2719 4294
rect 2955 4058 3041 4294
rect 3277 4058 3363 4294
rect 3599 4058 3685 4294
rect 3921 4058 4007 4294
rect 4243 4058 4329 4294
rect 4565 4058 4651 4294
rect 4887 4058 4973 4294
rect 5209 4058 5295 4294
rect 5531 4058 5617 4294
rect 5853 4058 5938 4294
rect 6174 4058 6259 4294
rect 6495 4058 6580 4294
rect 6816 4058 6901 4294
rect 7137 4058 7222 4294
rect 7458 4058 7543 4294
rect 7779 4058 7864 4294
rect 8100 4058 8185 4294
rect 8421 4058 8506 4294
rect 8742 4058 8827 4294
rect 9063 4058 9148 4294
rect 9384 4058 9469 4294
rect 9705 4058 9790 4294
rect 10026 4058 10111 4294
rect 10347 4058 10432 4294
rect 10668 4058 10753 4294
rect 10989 4058 11074 4294
rect 11310 4058 11395 4294
rect 11631 4058 11716 4294
rect 11952 4058 12037 4294
rect 12273 4058 12358 4294
rect 12594 4058 12679 4294
rect 12915 4058 13000 4294
rect 13236 4058 13321 4294
rect 13557 4058 13642 4294
rect 13878 4058 13963 4294
rect 14199 4058 14284 4294
rect 14520 4058 14605 4294
rect 14841 4058 15000 4294
rect 0 3688 15000 4058
rect 0 3452 143 3688
rect 379 3452 465 3688
rect 701 3452 787 3688
rect 1023 3452 1109 3688
rect 1345 3452 1431 3688
rect 1667 3452 1753 3688
rect 1989 3452 2075 3688
rect 2311 3452 2397 3688
rect 2633 3452 2719 3688
rect 2955 3452 3041 3688
rect 3277 3452 3363 3688
rect 3599 3452 3685 3688
rect 3921 3452 4007 3688
rect 4243 3452 4329 3688
rect 4565 3452 4651 3688
rect 4887 3452 4973 3688
rect 5209 3452 5295 3688
rect 5531 3452 5617 3688
rect 5853 3452 5938 3688
rect 6174 3452 6259 3688
rect 6495 3452 6580 3688
rect 6816 3452 6901 3688
rect 7137 3452 7222 3688
rect 7458 3452 7543 3688
rect 7779 3452 7864 3688
rect 8100 3452 8185 3688
rect 8421 3452 8506 3688
rect 8742 3452 8827 3688
rect 9063 3452 9148 3688
rect 9384 3452 9469 3688
rect 9705 3452 9790 3688
rect 10026 3452 10111 3688
rect 10347 3452 10432 3688
rect 10668 3452 10753 3688
rect 10989 3452 11074 3688
rect 11310 3452 11395 3688
rect 11631 3452 11716 3688
rect 11952 3452 12037 3688
rect 12273 3452 12358 3688
rect 12594 3452 12679 3688
rect 12915 3452 13000 3688
rect 13236 3452 13321 3688
rect 13557 3452 13642 3688
rect 13878 3452 13963 3688
rect 14199 3452 14284 3688
rect 14520 3452 14605 3688
rect 14841 3452 15000 3688
rect 0 3428 15000 3452
rect 0 3084 15000 3108
rect 0 2848 143 3084
rect 379 2848 465 3084
rect 701 2848 787 3084
rect 1023 2848 1109 3084
rect 1345 2848 1431 3084
rect 1667 2848 1753 3084
rect 1989 2848 2075 3084
rect 2311 2848 2397 3084
rect 2633 2848 2719 3084
rect 2955 2848 3041 3084
rect 3277 2848 3363 3084
rect 3599 2848 3685 3084
rect 3921 2848 4007 3084
rect 4243 2848 4329 3084
rect 4565 2848 4651 3084
rect 4887 2848 4973 3084
rect 5209 2848 5295 3084
rect 5531 2848 5617 3084
rect 5853 2848 5938 3084
rect 6174 2848 6259 3084
rect 6495 2848 6580 3084
rect 6816 2848 6901 3084
rect 7137 2848 7222 3084
rect 7458 2848 7543 3084
rect 7779 2848 7864 3084
rect 8100 2848 8185 3084
rect 8421 2848 8506 3084
rect 8742 2848 8827 3084
rect 9063 2848 9148 3084
rect 9384 2848 9469 3084
rect 9705 2848 9790 3084
rect 10026 2848 10111 3084
rect 10347 2848 10432 3084
rect 10668 2848 10753 3084
rect 10989 2848 11074 3084
rect 11310 2848 11395 3084
rect 11631 2848 11716 3084
rect 11952 2848 12037 3084
rect 12273 2848 12358 3084
rect 12594 2848 12679 3084
rect 12915 2848 13000 3084
rect 13236 2848 13321 3084
rect 13557 2848 13642 3084
rect 13878 2848 13963 3084
rect 14199 2848 14284 3084
rect 14520 2848 14605 3084
rect 14841 2848 15000 3084
rect 0 2718 15000 2848
rect 0 2482 143 2718
rect 379 2482 465 2718
rect 701 2482 787 2718
rect 1023 2482 1109 2718
rect 1345 2482 1431 2718
rect 1667 2482 1753 2718
rect 1989 2482 2075 2718
rect 2311 2482 2397 2718
rect 2633 2482 2719 2718
rect 2955 2482 3041 2718
rect 3277 2482 3363 2718
rect 3599 2482 3685 2718
rect 3921 2482 4007 2718
rect 4243 2482 4329 2718
rect 4565 2482 4651 2718
rect 4887 2482 4973 2718
rect 5209 2482 5295 2718
rect 5531 2482 5617 2718
rect 5853 2482 5938 2718
rect 6174 2482 6259 2718
rect 6495 2482 6580 2718
rect 6816 2482 6901 2718
rect 7137 2482 7222 2718
rect 7458 2482 7543 2718
rect 7779 2482 7864 2718
rect 8100 2482 8185 2718
rect 8421 2482 8506 2718
rect 8742 2482 8827 2718
rect 9063 2482 9148 2718
rect 9384 2482 9469 2718
rect 9705 2482 9790 2718
rect 10026 2482 10111 2718
rect 10347 2482 10432 2718
rect 10668 2482 10753 2718
rect 10989 2482 11074 2718
rect 11310 2482 11395 2718
rect 11631 2482 11716 2718
rect 11952 2482 12037 2718
rect 12273 2482 12358 2718
rect 12594 2482 12679 2718
rect 12915 2482 13000 2718
rect 13236 2482 13321 2718
rect 13557 2482 13642 2718
rect 13878 2482 13963 2718
rect 14199 2482 14284 2718
rect 14520 2482 14605 2718
rect 14841 2482 15000 2718
rect 0 2458 15000 2482
rect 0 2114 15000 2138
rect 0 1878 143 2114
rect 379 1878 465 2114
rect 701 1878 787 2114
rect 1023 1878 1109 2114
rect 1345 1878 1431 2114
rect 1667 1878 1753 2114
rect 1989 1878 2075 2114
rect 2311 1878 2397 2114
rect 2633 1878 2719 2114
rect 2955 1878 3041 2114
rect 3277 1878 3363 2114
rect 3599 1878 3685 2114
rect 3921 1878 4007 2114
rect 4243 1878 4329 2114
rect 4565 1878 4651 2114
rect 4887 1878 4973 2114
rect 5209 1878 5295 2114
rect 5531 1878 5617 2114
rect 5853 1878 5938 2114
rect 6174 1878 6259 2114
rect 6495 1878 6580 2114
rect 6816 1878 6901 2114
rect 7137 1878 7222 2114
rect 7458 1878 7543 2114
rect 7779 1878 7864 2114
rect 8100 1878 8185 2114
rect 8421 1878 8506 2114
rect 8742 1878 8827 2114
rect 9063 1878 9148 2114
rect 9384 1878 9469 2114
rect 9705 1878 9790 2114
rect 10026 1878 10111 2114
rect 10347 1878 10432 2114
rect 10668 1878 10753 2114
rect 10989 1878 11074 2114
rect 11310 1878 11395 2114
rect 11631 1878 11716 2114
rect 11952 1878 12037 2114
rect 12273 1878 12358 2114
rect 12594 1878 12679 2114
rect 12915 1878 13000 2114
rect 13236 1878 13321 2114
rect 13557 1878 13642 2114
rect 13878 1878 13963 2114
rect 14199 1878 14284 2114
rect 14520 1878 14605 2114
rect 14841 1878 15000 2114
rect 0 1508 15000 1878
rect 0 1272 143 1508
rect 379 1272 465 1508
rect 701 1272 787 1508
rect 1023 1272 1109 1508
rect 1345 1272 1431 1508
rect 1667 1272 1753 1508
rect 1989 1272 2075 1508
rect 2311 1272 2397 1508
rect 2633 1272 2719 1508
rect 2955 1272 3041 1508
rect 3277 1272 3363 1508
rect 3599 1272 3685 1508
rect 3921 1272 4007 1508
rect 4243 1272 4329 1508
rect 4565 1272 4651 1508
rect 4887 1272 4973 1508
rect 5209 1272 5295 1508
rect 5531 1272 5617 1508
rect 5853 1272 5938 1508
rect 6174 1272 6259 1508
rect 6495 1272 6580 1508
rect 6816 1272 6901 1508
rect 7137 1272 7222 1508
rect 7458 1272 7543 1508
rect 7779 1272 7864 1508
rect 8100 1272 8185 1508
rect 8421 1272 8506 1508
rect 8742 1272 8827 1508
rect 9063 1272 9148 1508
rect 9384 1272 9469 1508
rect 9705 1272 9790 1508
rect 10026 1272 10111 1508
rect 10347 1272 10432 1508
rect 10668 1272 10753 1508
rect 10989 1272 11074 1508
rect 11310 1272 11395 1508
rect 11631 1272 11716 1508
rect 11952 1272 12037 1508
rect 12273 1272 12358 1508
rect 12594 1272 12679 1508
rect 12915 1272 13000 1508
rect 13236 1272 13321 1508
rect 13557 1272 13642 1508
rect 13878 1272 13963 1508
rect 14199 1272 14284 1508
rect 14520 1272 14605 1508
rect 14841 1272 15000 1508
rect 0 1248 15000 1272
rect 0 903 15000 928
rect 0 667 143 903
rect 379 667 465 903
rect 701 667 787 903
rect 1023 667 1109 903
rect 1345 667 1431 903
rect 1667 667 1753 903
rect 1989 667 2075 903
rect 2311 667 2397 903
rect 2633 667 2719 903
rect 2955 667 3041 903
rect 3277 667 3363 903
rect 3599 667 3685 903
rect 3921 667 4007 903
rect 4243 667 4329 903
rect 4565 667 4651 903
rect 4887 667 4973 903
rect 5209 667 5295 903
rect 5531 667 5617 903
rect 5853 667 5938 903
rect 6174 667 6259 903
rect 6495 667 6580 903
rect 6816 667 6901 903
rect 7137 667 7222 903
rect 7458 667 7543 903
rect 7779 667 7864 903
rect 8100 667 8185 903
rect 8421 667 8506 903
rect 8742 667 8827 903
rect 9063 667 9148 903
rect 9384 667 9469 903
rect 9705 667 9790 903
rect 10026 667 10111 903
rect 10347 667 10432 903
rect 10668 667 10753 903
rect 10989 667 11074 903
rect 11310 667 11395 903
rect 11631 667 11716 903
rect 11952 667 12037 903
rect 12273 667 12358 903
rect 12594 667 12679 903
rect 12915 667 13000 903
rect 13236 667 13321 903
rect 13557 667 13642 903
rect 13878 667 13963 903
rect 14199 667 14284 903
rect 14520 667 14605 903
rect 14841 667 15000 903
rect 0 521 15000 667
rect 0 285 143 521
rect 379 285 465 521
rect 701 285 787 521
rect 1023 285 1109 521
rect 1345 285 1431 521
rect 1667 285 1753 521
rect 1989 285 2075 521
rect 2311 285 2397 521
rect 2633 285 2719 521
rect 2955 285 3041 521
rect 3277 285 3363 521
rect 3599 285 3685 521
rect 3921 285 4007 521
rect 4243 285 4329 521
rect 4565 285 4651 521
rect 4887 285 4973 521
rect 5209 285 5295 521
rect 5531 285 5617 521
rect 5853 285 5938 521
rect 6174 285 6259 521
rect 6495 285 6580 521
rect 6816 285 6901 521
rect 7137 285 7222 521
rect 7458 285 7543 521
rect 7779 285 7864 521
rect 8100 285 8185 521
rect 8421 285 8506 521
rect 8742 285 8827 521
rect 9063 285 9148 521
rect 9384 285 9469 521
rect 9705 285 9790 521
rect 10026 285 10111 521
rect 10347 285 10432 521
rect 10668 285 10753 521
rect 10989 285 11074 521
rect 11310 285 11395 521
rect 11631 285 11716 521
rect 11952 285 12037 521
rect 12273 285 12358 521
rect 12594 285 12679 521
rect 12915 285 13000 521
rect 13236 285 13321 521
rect 13557 285 13642 521
rect 13878 285 13963 521
rect 14199 285 14284 521
rect 14520 285 14605 521
rect 14841 285 15000 521
rect 0 139 15000 285
rect 0 -97 143 139
rect 379 -97 465 139
rect 701 -97 787 139
rect 1023 -97 1109 139
rect 1345 -97 1431 139
rect 1667 -97 1753 139
rect 1989 -97 2075 139
rect 2311 -97 2397 139
rect 2633 -97 2719 139
rect 2955 -97 3041 139
rect 3277 -97 3363 139
rect 3599 -97 3685 139
rect 3921 -97 4007 139
rect 4243 -97 4329 139
rect 4565 -97 4651 139
rect 4887 -97 4973 139
rect 5209 -97 5295 139
rect 5531 -97 5617 139
rect 5853 -97 5938 139
rect 6174 -97 6259 139
rect 6495 -97 6580 139
rect 6816 -97 6901 139
rect 7137 -97 7222 139
rect 7458 -97 7543 139
rect 7779 -97 7864 139
rect 8100 -97 8185 139
rect 8421 -97 8506 139
rect 8742 -97 8827 139
rect 9063 -97 9148 139
rect 9384 -97 9469 139
rect 9705 -97 9790 139
rect 10026 -97 10111 139
rect 10347 -97 10432 139
rect 10668 -97 10753 139
rect 10989 -97 11074 139
rect 11310 -97 11395 139
rect 11631 -97 11716 139
rect 11952 -97 12037 139
rect 12273 -97 12358 139
rect 12594 -97 12679 139
rect 12915 -97 13000 139
rect 13236 -97 13321 139
rect 13557 -97 13642 139
rect 13878 -97 13963 139
rect 14199 -97 14284 139
rect 14520 -97 14605 139
rect 14841 -97 15000 139
rect 0 -122 15000 -97
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_0
timestamp 1666464484
transform 1 0 0 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_1
timestamp 1666464484
transform 1 0 1000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_2
timestamp 1666464484
transform 1 0 2000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_3
timestamp 1666464484
transform 1 0 3000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_4
timestamp 1666464484
transform 1 0 4000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_5
timestamp 1666464484
transform 1 0 5000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_6
timestamp 1666464484
transform 1 0 6000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_7
timestamp 1666464484
transform 1 0 7000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_8
timestamp 1666464484
transform 1 0 8000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_9
timestamp 1666464484
transform 1 0 9000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_10
timestamp 1666464484
transform 1 0 14000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_11
timestamp 1666464484
transform 1 0 13000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_12
timestamp 1666464484
transform 1 0 12000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_13
timestamp 1666464484
transform 1 0 11000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_14
timestamp 1666464484
transform 1 0 10000 0 1 -6457
box 0 6315 1000 45908
<< labels >>
flabel metal5 s 14746 34608 15000 39451 3 FreeSans 520 180 0 0 VSSIO
port 1 nsew
flabel metal5 s 14746 8998 15000 10798 3 FreeSans 520 180 0 0 VSSA
port 2 nsew
flabel metal5 s 14807 2458 15000 3108 3 FreeSans 520 180 0 0 VDDA
port 3 nsew
flabel metal5 s 14746 7788 15000 8678 3 FreeSans 520 180 0 0 VSSD
port 4 nsew
flabel metal5 s 14746 11118 15000 11968 3 FreeSans 520 180 0 0 VSSIO_Q
port 5 nsew
flabel metal5 s 14746 4638 15000 5528 3 FreeSans 520 180 0 0 VSSIO
port 1 nsew
flabel metal5 s 14746 5848 15000 6498 3 FreeSans 520 180 0 0 VSWITCH
port 6 nsew
flabel metal5 s 14746 6819 15000 7468 3 FreeSans 520 180 0 0 VSSA
port 2 nsew
flabel metal5 s 14746 1248 15000 2138 3 FreeSans 520 180 0 0 VCCD
port 7 nsew
flabel metal5 s 14746 12288 15000 13138 3 FreeSans 520 180 0 0 VDDIO_Q
port 8 nsew
flabel metal5 s 14746 13458 15000 18448 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew
flabel metal5 s 14746 -122 15000 928 3 FreeSans 520 180 0 0 VCCHIB
port 10 nsew
flabel metal5 s 14746 3428 15000 4318 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew
flabel metal5 s 0 34608 254 39451 3 FreeSans 520 0 0 0 VSSIO
port 1 nsew
flabel metal5 s 0 13458 254 18448 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew
flabel metal5 s 0 7788 254 8678 3 FreeSans 520 0 0 0 VSSD
port 4 nsew
flabel metal5 s 0 11118 254 11968 3 FreeSans 520 0 0 0 VSSIO_Q
port 5 nsew
flabel metal5 s 0 5848 254 6498 3 FreeSans 520 0 0 0 VSWITCH
port 6 nsew
flabel metal5 s 0 4638 254 5528 3 FreeSans 520 0 0 0 VSSIO
port 1 nsew
flabel metal5 s 0 2458 193 3108 3 FreeSans 520 0 0 0 VDDA
port 3 nsew
flabel metal5 s 0 3428 254 4318 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew
flabel metal5 s 0 1248 254 2138 3 FreeSans 520 0 0 0 VCCD
port 7 nsew
flabel metal5 s 0 12288 254 13138 3 FreeSans 520 0 0 0 VDDIO_Q
port 8 nsew
flabel metal5 s 0 8998 254 10798 3 FreeSans 520 0 0 0 VSSA
port 2 nsew
flabel metal5 s 0 6819 254 7468 3 FreeSans 520 0 0 0 VSSA
port 2 nsew
flabel metal5 s 0 -122 254 928 3 FreeSans 520 0 0 0 VCCHIB
port 10 nsew
flabel metal4 s 14746 7768 15000 8698 3 FreeSans 520 180 0 0 VSSD
port 4 nsew
flabel metal4 s 14807 2438 15000 3128 3 FreeSans 520 180 0 0 VDDA
port 3 nsew
flabel metal4 s 14746 11098 15000 11988 3 FreeSans 520 180 0 0 VSSIO_Q
port 5 nsew
flabel metal4 s 14746 4618 15000 5548 3 FreeSans 520 180 0 0 VSSIO
port 1 nsew
flabel metal4 s 14746 5828 15000 6518 3 FreeSans 520 180 0 0 VSWITCH
port 6 nsew
flabel metal4 s 14746 9780 15000 10016 3 FreeSans 520 180 0 0 VSSA
port 2 nsew
flabel metal4 s 14746 10732 15000 10798 3 FreeSans 520 180 0 0 VSSA
port 2 nsew
flabel metal4 s 14746 -142 15000 948 3 FreeSans 520 180 0 0 VCCHIB
port 10 nsew
flabel metal4 s 14746 3408 15000 4338 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew
flabel metal4 s 14746 8998 15000 9064 3 FreeSans 520 180 0 0 VSSA
port 2 nsew
flabel metal4 s 14746 6798 15000 7488 3 FreeSans 520 180 0 0 VSSA
port 2 nsew
flabel metal4 s 14746 12268 15000 13158 3 FreeSans 520 180 0 0 VDDIO_Q
port 8 nsew
flabel metal4 s 14746 1228 15000 2158 3 FreeSans 520 180 0 0 VCCD
port 7 nsew
flabel metal4 s 14746 9124 15000 9720 3 FreeSans 520 180 0 0 AMUXBUS_B
port 11 nsew
flabel metal4 s 14746 34608 15000 39451 3 FreeSans 520 180 0 0 VSSIO
port 1 nsew
flabel metal4 s 14746 10076 15000 10672 3 FreeSans 520 180 0 0 AMUXBUS_A
port 12 nsew
flabel metal4 s 14746 13458 15000 18451 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew
flabel metal4 s 0 34608 254 39451 3 FreeSans 520 0 0 0 VSSIO
port 1 nsew
flabel metal4 s 0 3408 254 4338 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew
flabel metal4 s 0 12268 254 13158 3 FreeSans 520 0 0 0 VDDIO_Q
port 8 nsew
flabel metal4 s 0 13458 254 18451 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew
flabel metal4 s 0 1228 254 2158 3 FreeSans 520 0 0 0 VCCD
port 7 nsew
flabel metal4 s 0 8998 254 9064 3 FreeSans 520 0 0 0 VSSA
port 2 nsew
flabel metal4 s 0 5828 254 6518 3 FreeSans 520 0 0 0 VSWITCH
port 6 nsew
flabel metal4 s 0 -142 254 948 3 FreeSans 520 0 0 0 VCCHIB
port 10 nsew
flabel metal4 s 0 9780 254 10016 3 FreeSans 520 0 0 0 VSSA
port 2 nsew
flabel metal4 s 0 11098 254 11988 3 FreeSans 520 0 0 0 VSSIO_Q
port 5 nsew
flabel metal4 s 0 4618 254 5548 3 FreeSans 520 0 0 0 VSSIO
port 1 nsew
flabel metal4 s 0 2438 193 3128 3 FreeSans 520 0 0 0 VDDA
port 3 nsew
flabel metal4 s 0 10076 254 10672 3 FreeSans 520 0 0 0 AMUXBUS_A
port 12 nsew
flabel metal4 s 0 10732 254 10798 3 FreeSans 520 0 0 0 VSSA
port 2 nsew
flabel metal4 s 0 6798 254 7488 3 FreeSans 520 0 0 0 VSSA
port 2 nsew
flabel metal4 s 0 7768 254 8698 3 FreeSans 520 0 0 0 VSSD
port 4 nsew
flabel metal4 s 0 9124 254 9720 3 FreeSans 520 0 0 0 AMUXBUS_B
port 11 nsew
<< properties >>
string GDS_END 179026
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 19010
<< end >>
