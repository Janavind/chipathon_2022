magic
tech sky130B
magscale 1 2
timestamp 1666464484
use sky130_fd_pr__dfm1sd__example_55959141808169  sky130_fd_pr__dfm1sd__example_55959141808169_0
timestamp 1666464484
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfm1sd__example_55959141808169  sky130_fd_pr__dfm1sd__example_55959141808169_1
timestamp 1666464484
transform 1 0 100 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 35440366
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35439316
<< end >>
