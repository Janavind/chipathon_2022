magic
tech sky130B
timestamp 1666199351
<< properties >>
string GDS_END 31970976
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31970524
<< end >>
