magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 133 157 919 203
rect 36 21 919 157
rect 36 17 58 21
rect 24 -17 58 17
<< scnmos >>
rect 114 47 144 131
rect 209 47 239 177
rect 433 47 463 131
rect 528 47 558 177
rect 716 47 746 131
rect 811 47 841 177
<< scpmoshvt >>
rect 114 413 144 497
rect 209 297 239 497
rect 433 413 463 497
rect 528 297 558 497
rect 716 413 746 497
rect 811 297 841 497
<< ndiff >>
rect 159 131 209 177
rect 62 106 114 131
rect 62 72 70 106
rect 104 72 114 106
rect 62 47 114 72
rect 144 93 209 131
rect 144 59 159 93
rect 193 59 209 93
rect 144 47 209 59
rect 239 105 291 177
rect 478 131 528 177
rect 239 71 249 105
rect 283 71 291 105
rect 239 47 291 71
rect 381 105 433 131
rect 381 71 389 105
rect 423 71 433 105
rect 381 47 433 71
rect 463 93 528 131
rect 463 59 478 93
rect 512 59 528 93
rect 463 47 528 59
rect 558 105 610 177
rect 761 131 811 177
rect 558 71 568 105
rect 602 71 610 105
rect 558 47 610 71
rect 664 105 716 131
rect 664 71 672 105
rect 706 71 716 105
rect 664 47 716 71
rect 746 93 811 131
rect 746 59 761 93
rect 795 59 811 93
rect 746 47 811 59
rect 841 105 893 177
rect 841 71 851 105
rect 885 71 893 105
rect 841 47 893 71
<< pdiff >>
rect 62 472 114 497
rect 62 438 70 472
rect 104 438 114 472
rect 62 413 114 438
rect 144 489 209 497
rect 144 455 160 489
rect 194 455 209 489
rect 144 413 209 455
rect 159 297 209 413
rect 239 477 291 497
rect 239 443 249 477
rect 283 443 291 477
rect 239 409 291 443
rect 381 472 433 497
rect 381 438 389 472
rect 423 438 433 472
rect 381 413 433 438
rect 463 489 528 497
rect 463 455 479 489
rect 513 455 528 489
rect 463 413 528 455
rect 239 375 249 409
rect 283 375 291 409
rect 239 297 291 375
rect 478 297 528 413
rect 558 477 610 497
rect 558 443 568 477
rect 602 443 610 477
rect 558 409 610 443
rect 664 472 716 497
rect 664 438 672 472
rect 706 438 716 472
rect 664 413 716 438
rect 746 489 811 497
rect 746 455 762 489
rect 796 455 811 489
rect 746 413 811 455
rect 558 375 568 409
rect 602 375 610 409
rect 558 297 610 375
rect 761 297 811 413
rect 841 477 893 497
rect 841 443 851 477
rect 885 443 893 477
rect 841 409 893 443
rect 841 375 851 409
rect 885 375 893 409
rect 841 297 893 375
<< ndiffc >>
rect 70 72 104 106
rect 159 59 193 93
rect 249 71 283 105
rect 389 71 423 105
rect 478 59 512 93
rect 568 71 602 105
rect 672 71 706 105
rect 761 59 795 93
rect 851 71 885 105
<< pdiffc >>
rect 70 438 104 472
rect 160 455 194 489
rect 249 443 283 477
rect 389 438 423 472
rect 479 455 513 489
rect 249 375 283 409
rect 568 443 602 477
rect 672 438 706 472
rect 762 455 796 489
rect 568 375 602 409
rect 851 443 885 477
rect 851 375 885 409
<< poly >>
rect 114 497 144 523
rect 209 497 239 523
rect 433 497 463 523
rect 528 497 558 523
rect 716 497 746 523
rect 811 497 841 523
rect 114 265 144 413
rect 209 265 239 297
rect 433 265 463 413
rect 528 265 558 297
rect 716 265 746 413
rect 811 265 841 297
rect 57 249 144 265
rect 57 215 67 249
rect 101 215 144 249
rect 57 199 144 215
rect 186 249 240 265
rect 186 215 196 249
rect 230 215 240 249
rect 186 199 240 215
rect 376 249 463 265
rect 376 215 386 249
rect 420 215 463 249
rect 376 199 463 215
rect 505 249 559 265
rect 505 215 515 249
rect 549 215 559 249
rect 505 199 559 215
rect 659 249 746 265
rect 659 215 669 249
rect 703 215 746 249
rect 659 199 746 215
rect 788 249 842 265
rect 788 215 798 249
rect 832 215 842 249
rect 788 199 842 215
rect 114 131 144 199
rect 209 177 239 199
rect 433 131 463 199
rect 528 177 558 199
rect 716 131 746 199
rect 811 177 841 199
rect 114 21 144 47
rect 209 21 239 47
rect 433 21 463 47
rect 528 21 558 47
rect 716 21 746 47
rect 811 21 841 47
<< polycont >>
rect 67 215 101 249
rect 196 215 230 249
rect 386 215 420 249
rect 515 215 549 249
rect 669 215 703 249
rect 798 215 832 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 472 104 493
rect 17 438 70 472
rect 138 489 215 527
rect 138 455 160 489
rect 194 455 215 489
rect 138 442 215 455
rect 249 477 334 493
rect 283 443 334 477
rect 17 408 104 438
rect 249 409 334 443
rect 17 374 215 408
rect 17 249 114 340
rect 17 215 67 249
rect 101 215 114 249
rect 17 199 114 215
rect 148 265 215 374
rect 283 375 334 409
rect 249 335 334 375
rect 368 472 423 493
rect 368 438 389 472
rect 457 489 534 527
rect 457 455 479 489
rect 513 455 534 489
rect 457 442 534 455
rect 568 477 617 493
rect 602 443 617 477
rect 368 408 423 438
rect 568 409 617 443
rect 368 369 534 408
rect 249 299 430 335
rect 148 249 230 265
rect 148 215 196 249
rect 148 199 230 215
rect 264 249 430 299
rect 264 215 386 249
rect 420 215 430 249
rect 264 199 430 215
rect 464 265 534 369
rect 602 375 617 409
rect 568 335 617 375
rect 655 472 706 493
rect 655 438 672 472
rect 740 489 817 527
rect 740 455 762 489
rect 796 455 817 489
rect 740 442 817 455
rect 851 477 903 493
rect 885 443 903 477
rect 655 408 706 438
rect 851 409 903 443
rect 655 369 817 408
rect 568 299 713 335
rect 464 249 549 265
rect 464 215 515 249
rect 464 199 549 215
rect 583 249 713 299
rect 583 215 669 249
rect 703 215 713 249
rect 583 199 713 215
rect 747 265 817 369
rect 885 375 903 409
rect 851 299 903 375
rect 747 249 832 265
rect 747 215 798 249
rect 747 199 832 215
rect 148 165 215 199
rect 264 165 334 199
rect 464 165 534 199
rect 583 165 617 199
rect 747 165 817 199
rect 866 165 903 299
rect 17 131 215 165
rect 17 106 104 131
rect 17 72 70 106
rect 249 105 334 165
rect 17 51 104 72
rect 138 93 215 97
rect 138 59 159 93
rect 193 59 215 93
rect 138 17 215 59
rect 283 71 334 105
rect 249 51 334 71
rect 372 131 534 165
rect 372 105 423 131
rect 372 71 389 105
rect 568 105 617 165
rect 372 51 423 71
rect 457 93 534 97
rect 457 59 478 93
rect 512 59 534 93
rect 457 17 534 59
rect 602 71 617 105
rect 568 51 617 71
rect 655 131 817 165
rect 655 105 706 131
rect 655 71 672 105
rect 851 105 903 165
rect 655 51 706 71
rect 740 93 817 97
rect 740 59 761 93
rect 795 59 817 93
rect 740 17 817 59
rect 885 71 903 105
rect 851 51 903 71
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel metal1 s 24 527 58 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 24 -17 58 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel nwell s 24 527 58 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 24 -17 58 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel locali s 24 221 58 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 300 289 334 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 24 289 58 323 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 300 357 334 391 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 300 425 334 459 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 300 221 334 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 300 153 334 187 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 300 85 334 119 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 392 221 426 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 392 289 426 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
rlabel comment s 0 0 0 0 4 dlymetal6s2s_1
rlabel metal1 s 0 -48 920 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 2917254
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2909478
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 23.000 13.600 
<< end >>
