magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< metal1 >>
rect 1465 2168 1471 2220
rect 1523 2168 1529 2220
rect 1570 1130 1604 2256
rect 1646 1142 1674 2256
rect 6457 2168 6463 2220
rect 6515 2168 6521 2220
rect 1793 2016 1799 2068
rect 1851 2016 1857 2068
rect 1711 1242 1717 1294
rect 1769 1242 1775 1294
rect 6562 1130 6596 2256
rect 6638 1142 6666 2256
rect 11449 2168 11455 2220
rect 11507 2168 11513 2220
rect 6785 2016 6791 2068
rect 6843 2016 6849 2068
rect 6703 1242 6709 1294
rect 6761 1242 6767 1294
rect 11554 1130 11588 2256
rect 11630 1142 11658 2256
rect 16441 2168 16447 2220
rect 16499 2168 16505 2220
rect 11777 2016 11783 2068
rect 11835 2016 11841 2068
rect 11695 1242 11701 1294
rect 11753 1242 11759 1294
rect 16546 1130 16580 2256
rect 16622 1142 16650 2256
rect 21433 2168 21439 2220
rect 21491 2168 21497 2220
rect 16769 2016 16775 2068
rect 16827 2016 16833 2068
rect 16687 1242 16693 1294
rect 16745 1242 16751 1294
rect 21538 1130 21572 2256
rect 21614 1142 21642 2256
rect 26425 2168 26431 2220
rect 26483 2168 26489 2220
rect 21761 2016 21767 2068
rect 21819 2016 21825 2068
rect 21679 1242 21685 1294
rect 21737 1242 21743 1294
rect 26530 1130 26564 2256
rect 26606 1142 26634 2256
rect 31417 2168 31423 2220
rect 31475 2168 31481 2220
rect 26753 2016 26759 2068
rect 26811 2016 26817 2068
rect 26671 1242 26677 1294
rect 26729 1242 26735 1294
rect 31522 1130 31556 2256
rect 31598 1142 31626 2256
rect 36409 2168 36415 2220
rect 36467 2168 36473 2220
rect 31745 2016 31751 2068
rect 31803 2016 31809 2068
rect 31663 1242 31669 1294
rect 31721 1242 31727 1294
rect 36514 1130 36548 2256
rect 36590 1142 36618 2256
rect 36737 2016 36743 2068
rect 36795 2016 36801 2068
rect 36655 1242 36661 1294
rect 36713 1242 36719 1294
rect 1723 404 1729 456
rect 1781 404 1787 456
rect 6715 404 6721 456
rect 6773 404 6779 456
rect 11707 404 11713 456
rect 11765 404 11771 456
rect 16699 404 16705 456
rect 16757 404 16763 456
rect 21691 404 21697 456
rect 21749 404 21755 456
rect 26683 404 26689 456
rect 26741 404 26747 456
rect 31675 404 31681 456
rect 31733 404 31739 456
rect 36667 404 36673 456
rect 36725 404 36731 456
rect 1478 0 1524 254
rect 1723 82 1729 134
rect 1781 82 1787 134
rect 6470 0 6516 254
rect 6715 82 6721 134
rect 6773 82 6779 134
rect 11462 0 11508 254
rect 11707 82 11713 134
rect 11765 82 11771 134
rect 16454 0 16500 254
rect 16699 82 16705 134
rect 16757 82 16763 134
rect 21446 0 21492 254
rect 21691 82 21697 134
rect 21749 82 21755 134
rect 26438 0 26484 254
rect 26683 82 26689 134
rect 26741 82 26747 134
rect 31430 0 31476 254
rect 31675 82 31681 134
rect 31733 82 31739 134
rect 36422 0 36468 254
rect 36667 82 36673 134
rect 36725 82 36731 134
<< via1 >>
rect 1471 2168 1523 2220
rect 6463 2168 6515 2220
rect 1799 2016 1851 2068
rect 1717 1242 1769 1294
rect 11455 2168 11507 2220
rect 6791 2016 6843 2068
rect 6709 1242 6761 1294
rect 16447 2168 16499 2220
rect 11783 2016 11835 2068
rect 11701 1242 11753 1294
rect 21439 2168 21491 2220
rect 16775 2016 16827 2068
rect 16693 1242 16745 1294
rect 26431 2168 26483 2220
rect 21767 2016 21819 2068
rect 21685 1242 21737 1294
rect 31423 2168 31475 2220
rect 26759 2016 26811 2068
rect 26677 1242 26729 1294
rect 36415 2168 36467 2220
rect 31751 2016 31803 2068
rect 31669 1242 31721 1294
rect 36743 2016 36795 2068
rect 36661 1242 36713 1294
rect 1729 404 1781 456
rect 6721 404 6773 456
rect 11713 404 11765 456
rect 16705 404 16757 456
rect 21697 404 21749 456
rect 26689 404 26741 456
rect 31681 404 31733 456
rect 36673 404 36725 456
rect 1729 82 1781 134
rect 6721 82 6773 134
rect 11713 82 11765 134
rect 16705 82 16757 134
rect 21697 82 21749 134
rect 26689 82 26741 134
rect 31681 82 31733 134
rect 36673 82 36725 134
<< metal2 >>
rect 1469 2222 1525 2231
rect 1469 2157 1525 2166
rect 6461 2222 6517 2231
rect 6461 2157 6517 2166
rect 11453 2222 11509 2231
rect 11453 2157 11509 2166
rect 16445 2222 16501 2231
rect 16445 2157 16501 2166
rect 21437 2222 21493 2231
rect 21437 2157 21493 2166
rect 26429 2222 26485 2231
rect 26429 2157 26485 2166
rect 31421 2222 31477 2231
rect 31421 2157 31477 2166
rect 36413 2222 36469 2231
rect 36413 2157 36469 2166
rect 1797 2070 1853 2079
rect 1797 2005 1853 2014
rect 6789 2070 6845 2079
rect 6789 2005 6845 2014
rect 11781 2070 11837 2079
rect 11781 2005 11837 2014
rect 16773 2070 16829 2079
rect 16773 2005 16829 2014
rect 21765 2070 21821 2079
rect 21765 2005 21821 2014
rect 26757 2070 26813 2079
rect 26757 2005 26813 2014
rect 31749 2070 31805 2079
rect 31749 2005 31805 2014
rect 36741 2070 36797 2079
rect 36741 2005 36797 2014
rect 1715 1296 1771 1305
rect 1715 1231 1771 1240
rect 6707 1296 6763 1305
rect 6707 1231 6763 1240
rect 11699 1296 11755 1305
rect 11699 1231 11755 1240
rect 16691 1296 16747 1305
rect 16691 1231 16747 1240
rect 21683 1296 21739 1305
rect 21683 1231 21739 1240
rect 26675 1296 26731 1305
rect 26675 1231 26731 1240
rect 31667 1296 31723 1305
rect 31667 1231 31723 1240
rect 36659 1296 36715 1305
rect 36659 1231 36715 1240
rect 1727 458 1783 467
rect 1727 393 1783 402
rect 6719 458 6775 467
rect 6719 393 6775 402
rect 11711 458 11767 467
rect 11711 393 11767 402
rect 16703 458 16759 467
rect 16703 393 16759 402
rect 21695 458 21751 467
rect 21695 393 21751 402
rect 26687 458 26743 467
rect 26687 393 26743 402
rect 31679 458 31735 467
rect 31679 393 31735 402
rect 36671 458 36727 467
rect 36671 393 36727 402
rect 1727 136 1783 145
rect 1727 71 1783 80
rect 6719 136 6775 145
rect 6719 71 6775 80
rect 11711 136 11767 145
rect 11711 71 11767 80
rect 16703 136 16759 145
rect 16703 71 16759 80
rect 21695 136 21751 145
rect 21695 71 21751 80
rect 26687 136 26743 145
rect 26687 71 26743 80
rect 31679 136 31735 145
rect 31679 71 31735 80
rect 36671 136 36727 145
rect 36671 71 36727 80
<< via2 >>
rect 1469 2220 1525 2222
rect 1469 2168 1471 2220
rect 1471 2168 1523 2220
rect 1523 2168 1525 2220
rect 1469 2166 1525 2168
rect 6461 2220 6517 2222
rect 6461 2168 6463 2220
rect 6463 2168 6515 2220
rect 6515 2168 6517 2220
rect 6461 2166 6517 2168
rect 11453 2220 11509 2222
rect 11453 2168 11455 2220
rect 11455 2168 11507 2220
rect 11507 2168 11509 2220
rect 11453 2166 11509 2168
rect 16445 2220 16501 2222
rect 16445 2168 16447 2220
rect 16447 2168 16499 2220
rect 16499 2168 16501 2220
rect 16445 2166 16501 2168
rect 21437 2220 21493 2222
rect 21437 2168 21439 2220
rect 21439 2168 21491 2220
rect 21491 2168 21493 2220
rect 21437 2166 21493 2168
rect 26429 2220 26485 2222
rect 26429 2168 26431 2220
rect 26431 2168 26483 2220
rect 26483 2168 26485 2220
rect 26429 2166 26485 2168
rect 31421 2220 31477 2222
rect 31421 2168 31423 2220
rect 31423 2168 31475 2220
rect 31475 2168 31477 2220
rect 31421 2166 31477 2168
rect 36413 2220 36469 2222
rect 36413 2168 36415 2220
rect 36415 2168 36467 2220
rect 36467 2168 36469 2220
rect 36413 2166 36469 2168
rect 1797 2068 1853 2070
rect 1797 2016 1799 2068
rect 1799 2016 1851 2068
rect 1851 2016 1853 2068
rect 1797 2014 1853 2016
rect 6789 2068 6845 2070
rect 6789 2016 6791 2068
rect 6791 2016 6843 2068
rect 6843 2016 6845 2068
rect 6789 2014 6845 2016
rect 11781 2068 11837 2070
rect 11781 2016 11783 2068
rect 11783 2016 11835 2068
rect 11835 2016 11837 2068
rect 11781 2014 11837 2016
rect 16773 2068 16829 2070
rect 16773 2016 16775 2068
rect 16775 2016 16827 2068
rect 16827 2016 16829 2068
rect 16773 2014 16829 2016
rect 21765 2068 21821 2070
rect 21765 2016 21767 2068
rect 21767 2016 21819 2068
rect 21819 2016 21821 2068
rect 21765 2014 21821 2016
rect 26757 2068 26813 2070
rect 26757 2016 26759 2068
rect 26759 2016 26811 2068
rect 26811 2016 26813 2068
rect 26757 2014 26813 2016
rect 31749 2068 31805 2070
rect 31749 2016 31751 2068
rect 31751 2016 31803 2068
rect 31803 2016 31805 2068
rect 31749 2014 31805 2016
rect 36741 2068 36797 2070
rect 36741 2016 36743 2068
rect 36743 2016 36795 2068
rect 36795 2016 36797 2068
rect 36741 2014 36797 2016
rect 1715 1294 1771 1296
rect 1715 1242 1717 1294
rect 1717 1242 1769 1294
rect 1769 1242 1771 1294
rect 1715 1240 1771 1242
rect 6707 1294 6763 1296
rect 6707 1242 6709 1294
rect 6709 1242 6761 1294
rect 6761 1242 6763 1294
rect 6707 1240 6763 1242
rect 11699 1294 11755 1296
rect 11699 1242 11701 1294
rect 11701 1242 11753 1294
rect 11753 1242 11755 1294
rect 11699 1240 11755 1242
rect 16691 1294 16747 1296
rect 16691 1242 16693 1294
rect 16693 1242 16745 1294
rect 16745 1242 16747 1294
rect 16691 1240 16747 1242
rect 21683 1294 21739 1296
rect 21683 1242 21685 1294
rect 21685 1242 21737 1294
rect 21737 1242 21739 1294
rect 21683 1240 21739 1242
rect 26675 1294 26731 1296
rect 26675 1242 26677 1294
rect 26677 1242 26729 1294
rect 26729 1242 26731 1294
rect 26675 1240 26731 1242
rect 31667 1294 31723 1296
rect 31667 1242 31669 1294
rect 31669 1242 31721 1294
rect 31721 1242 31723 1294
rect 31667 1240 31723 1242
rect 36659 1294 36715 1296
rect 36659 1242 36661 1294
rect 36661 1242 36713 1294
rect 36713 1242 36715 1294
rect 36659 1240 36715 1242
rect 1727 456 1783 458
rect 1727 404 1729 456
rect 1729 404 1781 456
rect 1781 404 1783 456
rect 1727 402 1783 404
rect 6719 456 6775 458
rect 6719 404 6721 456
rect 6721 404 6773 456
rect 6773 404 6775 456
rect 6719 402 6775 404
rect 11711 456 11767 458
rect 11711 404 11713 456
rect 11713 404 11765 456
rect 11765 404 11767 456
rect 11711 402 11767 404
rect 16703 456 16759 458
rect 16703 404 16705 456
rect 16705 404 16757 456
rect 16757 404 16759 456
rect 16703 402 16759 404
rect 21695 456 21751 458
rect 21695 404 21697 456
rect 21697 404 21749 456
rect 21749 404 21751 456
rect 21695 402 21751 404
rect 26687 456 26743 458
rect 26687 404 26689 456
rect 26689 404 26741 456
rect 26741 404 26743 456
rect 26687 402 26743 404
rect 31679 456 31735 458
rect 31679 404 31681 456
rect 31681 404 31733 456
rect 31733 404 31735 456
rect 31679 402 31735 404
rect 36671 456 36727 458
rect 36671 404 36673 456
rect 36673 404 36725 456
rect 36725 404 36727 456
rect 36671 402 36727 404
rect 1727 134 1783 136
rect 1727 82 1729 134
rect 1729 82 1781 134
rect 1781 82 1783 134
rect 1727 80 1783 82
rect 6719 134 6775 136
rect 6719 82 6721 134
rect 6721 82 6773 134
rect 6773 82 6775 134
rect 6719 80 6775 82
rect 11711 134 11767 136
rect 11711 82 11713 134
rect 11713 82 11765 134
rect 11765 82 11767 134
rect 11711 80 11767 82
rect 16703 134 16759 136
rect 16703 82 16705 134
rect 16705 82 16757 134
rect 16757 82 16759 134
rect 16703 80 16759 82
rect 21695 134 21751 136
rect 21695 82 21697 134
rect 21697 82 21749 134
rect 21749 82 21751 134
rect 21695 80 21751 82
rect 26687 134 26743 136
rect 26687 82 26689 134
rect 26689 82 26741 134
rect 26741 82 26743 134
rect 26687 80 26743 82
rect 31679 134 31735 136
rect 31679 82 31681 134
rect 31681 82 31733 134
rect 31733 82 31735 134
rect 31679 80 31735 82
rect 36671 134 36727 136
rect 36671 82 36673 134
rect 36673 82 36725 134
rect 36725 82 36727 134
rect 36671 80 36727 82
<< metal3 >>
rect 1464 2224 1530 2227
rect 6456 2224 6522 2227
rect 11448 2224 11514 2227
rect 16440 2224 16506 2227
rect 21432 2224 21498 2227
rect 26424 2224 26490 2227
rect 31416 2224 31482 2227
rect 36408 2224 36474 2227
rect 0 2222 36818 2224
rect 0 2166 1469 2222
rect 1525 2166 6461 2222
rect 6517 2166 11453 2222
rect 11509 2166 16445 2222
rect 16501 2166 21437 2222
rect 21493 2166 26429 2222
rect 26485 2166 31421 2222
rect 31477 2166 36413 2222
rect 36469 2166 36818 2222
rect 0 2164 36818 2166
rect 1464 2161 1530 2164
rect 6456 2161 6522 2164
rect 11448 2161 11514 2164
rect 16440 2161 16506 2164
rect 21432 2161 21498 2164
rect 26424 2161 26490 2164
rect 31416 2161 31482 2164
rect 36408 2161 36474 2164
rect 1776 2070 1874 2091
rect 1776 2014 1797 2070
rect 1853 2014 1874 2070
rect 1776 1993 1874 2014
rect 6768 2070 6866 2091
rect 6768 2014 6789 2070
rect 6845 2014 6866 2070
rect 6768 1993 6866 2014
rect 11760 2070 11858 2091
rect 11760 2014 11781 2070
rect 11837 2014 11858 2070
rect 11760 1993 11858 2014
rect 16752 2070 16850 2091
rect 16752 2014 16773 2070
rect 16829 2014 16850 2070
rect 16752 1993 16850 2014
rect 21744 2070 21842 2091
rect 21744 2014 21765 2070
rect 21821 2014 21842 2070
rect 21744 1993 21842 2014
rect 26736 2070 26834 2091
rect 26736 2014 26757 2070
rect 26813 2014 26834 2070
rect 26736 1993 26834 2014
rect 31728 2070 31826 2091
rect 31728 2014 31749 2070
rect 31805 2014 31826 2070
rect 31728 1993 31826 2014
rect 36720 2070 36818 2091
rect 36720 2014 36741 2070
rect 36797 2014 36818 2070
rect 36720 1993 36818 2014
rect 1694 1296 1792 1317
rect 1694 1240 1715 1296
rect 1771 1240 1792 1296
rect 1694 1219 1792 1240
rect 6686 1296 6784 1317
rect 6686 1240 6707 1296
rect 6763 1240 6784 1296
rect 6686 1219 6784 1240
rect 11678 1296 11776 1317
rect 11678 1240 11699 1296
rect 11755 1240 11776 1296
rect 11678 1219 11776 1240
rect 16670 1296 16768 1317
rect 16670 1240 16691 1296
rect 16747 1240 16768 1296
rect 16670 1219 16768 1240
rect 21662 1296 21760 1317
rect 21662 1240 21683 1296
rect 21739 1240 21760 1296
rect 21662 1219 21760 1240
rect 26654 1296 26752 1317
rect 26654 1240 26675 1296
rect 26731 1240 26752 1296
rect 26654 1219 26752 1240
rect 31646 1296 31744 1317
rect 31646 1240 31667 1296
rect 31723 1240 31744 1296
rect 31646 1219 31744 1240
rect 36638 1296 36736 1317
rect 36638 1240 36659 1296
rect 36715 1240 36736 1296
rect 36638 1219 36736 1240
rect 1706 458 1804 479
rect 1706 402 1727 458
rect 1783 402 1804 458
rect 1706 381 1804 402
rect 6698 458 6796 479
rect 6698 402 6719 458
rect 6775 402 6796 458
rect 6698 381 6796 402
rect 11690 458 11788 479
rect 11690 402 11711 458
rect 11767 402 11788 458
rect 11690 381 11788 402
rect 16682 458 16780 479
rect 16682 402 16703 458
rect 16759 402 16780 458
rect 16682 381 16780 402
rect 21674 458 21772 479
rect 21674 402 21695 458
rect 21751 402 21772 458
rect 21674 381 21772 402
rect 26666 458 26764 479
rect 26666 402 26687 458
rect 26743 402 26764 458
rect 26666 381 26764 402
rect 31658 458 31756 479
rect 31658 402 31679 458
rect 31735 402 31756 458
rect 31658 381 31756 402
rect 36650 458 36748 479
rect 36650 402 36671 458
rect 36727 402 36748 458
rect 36650 381 36748 402
rect 1706 136 1804 157
rect 1706 80 1727 136
rect 1783 80 1804 136
rect 1706 59 1804 80
rect 6698 136 6796 157
rect 6698 80 6719 136
rect 6775 80 6796 136
rect 6698 59 6796 80
rect 11690 136 11788 157
rect 11690 80 11711 136
rect 11767 80 11788 136
rect 11690 59 11788 80
rect 16682 136 16780 157
rect 16682 80 16703 136
rect 16759 80 16780 136
rect 16682 59 16780 80
rect 21674 136 21772 157
rect 21674 80 21695 136
rect 21751 80 21772 136
rect 21674 59 21772 80
rect 26666 136 26764 157
rect 26666 80 26687 136
rect 26743 80 26764 136
rect 26666 59 26764 80
rect 31658 136 31756 157
rect 31658 80 31679 136
rect 31735 80 31756 136
rect 31658 59 31756 80
rect 36650 136 36748 157
rect 36650 80 36671 136
rect 36727 80 36748 136
rect 36650 59 36748 80
use sky130_fd_bd_sram__openram_sense_amp_1  sky130_fd_bd_sram__openram_sense_amp_0
timestamp 1666464484
transform 1 0 36318 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_1  sky130_fd_bd_sram__openram_sense_amp_1
timestamp 1666464484
transform 1 0 31326 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_1  sky130_fd_bd_sram__openram_sense_amp_2
timestamp 1666464484
transform 1 0 26334 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_1  sky130_fd_bd_sram__openram_sense_amp_3
timestamp 1666464484
transform 1 0 21342 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_1  sky130_fd_bd_sram__openram_sense_amp_4
timestamp 1666464484
transform 1 0 16350 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_1  sky130_fd_bd_sram__openram_sense_amp_5
timestamp 1666464484
transform 1 0 11358 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_1  sky130_fd_bd_sram__openram_sense_amp_6
timestamp 1666464484
transform 1 0 6366 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_1  sky130_fd_bd_sram__openram_sense_amp_7
timestamp 1666464484
transform 1 0 1374 0 1 0
box -541 0 937 2256
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_0
timestamp 1666464484
transform 1 0 36408 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_1
timestamp 1666464484
transform 1 0 31416 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_2
timestamp 1666464484
transform 1 0 26424 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_3
timestamp 1666464484
transform 1 0 21432 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_4
timestamp 1666464484
transform 1 0 16440 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_5
timestamp 1666464484
transform 1 0 11448 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_6
timestamp 1666464484
transform 1 0 6456 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_7
timestamp 1666464484
transform 1 0 1464 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_8
timestamp 1666464484
transform 1 0 36666 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_9
timestamp 1666464484
transform 1 0 36654 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_10
timestamp 1666464484
transform 1 0 36666 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_11
timestamp 1666464484
transform 1 0 36736 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_12
timestamp 1666464484
transform 1 0 31674 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_13
timestamp 1666464484
transform 1 0 31662 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_14
timestamp 1666464484
transform 1 0 31674 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_15
timestamp 1666464484
transform 1 0 31744 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_16
timestamp 1666464484
transform 1 0 26682 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_17
timestamp 1666464484
transform 1 0 26670 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_18
timestamp 1666464484
transform 1 0 26682 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_19
timestamp 1666464484
transform 1 0 26752 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_20
timestamp 1666464484
transform 1 0 21690 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_21
timestamp 1666464484
transform 1 0 21678 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_22
timestamp 1666464484
transform 1 0 21690 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_23
timestamp 1666464484
transform 1 0 21760 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_24
timestamp 1666464484
transform 1 0 16698 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_25
timestamp 1666464484
transform 1 0 16686 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_26
timestamp 1666464484
transform 1 0 16698 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_27
timestamp 1666464484
transform 1 0 16768 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_28
timestamp 1666464484
transform 1 0 11706 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_29
timestamp 1666464484
transform 1 0 11694 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_30
timestamp 1666464484
transform 1 0 11706 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_31
timestamp 1666464484
transform 1 0 11776 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_32
timestamp 1666464484
transform 1 0 6714 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_33
timestamp 1666464484
transform 1 0 6702 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_34
timestamp 1666464484
transform 1 0 6714 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_35
timestamp 1666464484
transform 1 0 6784 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_36
timestamp 1666464484
transform 1 0 1722 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_37
timestamp 1666464484
transform 1 0 1710 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_38
timestamp 1666464484
transform 1 0 1722 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_39
timestamp 1666464484
transform 1 0 1792 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_0
timestamp 1666464484
transform 1 0 36409 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_1
timestamp 1666464484
transform 1 0 31417 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_2
timestamp 1666464484
transform 1 0 26425 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_3
timestamp 1666464484
transform 1 0 21433 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_4
timestamp 1666464484
transform 1 0 16441 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_5
timestamp 1666464484
transform 1 0 11449 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_6
timestamp 1666464484
transform 1 0 6457 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_7
timestamp 1666464484
transform 1 0 1465 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_8
timestamp 1666464484
transform 1 0 36667 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_9
timestamp 1666464484
transform 1 0 36655 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_10
timestamp 1666464484
transform 1 0 36667 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_11
timestamp 1666464484
transform 1 0 36737 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_12
timestamp 1666464484
transform 1 0 31675 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_13
timestamp 1666464484
transform 1 0 31663 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_14
timestamp 1666464484
transform 1 0 31675 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_15
timestamp 1666464484
transform 1 0 31745 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_16
timestamp 1666464484
transform 1 0 26683 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_17
timestamp 1666464484
transform 1 0 26671 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_18
timestamp 1666464484
transform 1 0 26683 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_19
timestamp 1666464484
transform 1 0 26753 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_20
timestamp 1666464484
transform 1 0 21691 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_21
timestamp 1666464484
transform 1 0 21679 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_22
timestamp 1666464484
transform 1 0 21691 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_23
timestamp 1666464484
transform 1 0 21761 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_24
timestamp 1666464484
transform 1 0 16699 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_25
timestamp 1666464484
transform 1 0 16687 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_26
timestamp 1666464484
transform 1 0 16699 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_27
timestamp 1666464484
transform 1 0 16769 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_28
timestamp 1666464484
transform 1 0 11707 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_29
timestamp 1666464484
transform 1 0 11695 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_30
timestamp 1666464484
transform 1 0 11707 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_31
timestamp 1666464484
transform 1 0 11777 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_32
timestamp 1666464484
transform 1 0 6715 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_33
timestamp 1666464484
transform 1 0 6703 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_34
timestamp 1666464484
transform 1 0 6715 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_35
timestamp 1666464484
transform 1 0 6785 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_36
timestamp 1666464484
transform 1 0 1723 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_37
timestamp 1666464484
transform 1 0 1711 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_38
timestamp 1666464484
transform 1 0 1723 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_39
timestamp 1666464484
transform 1 0 1793 0 1 2010
box 0 0 1 1
<< labels >>
rlabel metal3 s 26736 1993 26834 2091 4 gnd
port 1 nsew
rlabel metal3 s 31728 1993 31826 2091 4 gnd
port 1 nsew
rlabel metal3 s 1776 1993 1874 2091 4 gnd
port 1 nsew
rlabel metal3 s 11690 59 11788 157 4 gnd
port 1 nsew
rlabel metal3 s 11760 1993 11858 2091 4 gnd
port 1 nsew
rlabel metal3 s 21674 59 21772 157 4 gnd
port 1 nsew
rlabel metal3 s 21744 1993 21842 2091 4 gnd
port 1 nsew
rlabel metal3 s 26666 59 26764 157 4 gnd
port 1 nsew
rlabel metal3 s 16682 59 16780 157 4 gnd
port 1 nsew
rlabel metal3 s 36650 59 36748 157 4 gnd
port 1 nsew
rlabel metal3 s 6698 59 6796 157 4 gnd
port 1 nsew
rlabel metal3 s 1706 59 1804 157 4 gnd
port 1 nsew
rlabel metal3 s 36720 1993 36818 2091 4 gnd
port 1 nsew
rlabel metal3 s 6768 1993 6866 2091 4 gnd
port 1 nsew
rlabel metal3 s 31658 59 31756 157 4 gnd
port 1 nsew
rlabel metal3 s 16752 1993 16850 2091 4 gnd
port 1 nsew
rlabel metal3 s 16682 381 16780 479 4 vdd
port 2 nsew
rlabel metal3 s 21662 1219 21760 1317 4 vdd
port 2 nsew
rlabel metal3 s 26666 381 26764 479 4 vdd
port 2 nsew
rlabel metal3 s 36650 381 36748 479 4 vdd
port 2 nsew
rlabel metal3 s 31646 1219 31744 1317 4 vdd
port 2 nsew
rlabel metal3 s 36638 1219 36736 1317 4 vdd
port 2 nsew
rlabel metal3 s 11678 1219 11776 1317 4 vdd
port 2 nsew
rlabel metal3 s 6686 1219 6784 1317 4 vdd
port 2 nsew
rlabel metal3 s 21674 381 21772 479 4 vdd
port 2 nsew
rlabel metal3 s 26654 1219 26752 1317 4 vdd
port 2 nsew
rlabel metal3 s 1706 381 1804 479 4 vdd
port 2 nsew
rlabel metal3 s 11690 381 11788 479 4 vdd
port 2 nsew
rlabel metal3 s 6698 381 6796 479 4 vdd
port 2 nsew
rlabel metal3 s 16670 1219 16768 1317 4 vdd
port 2 nsew
rlabel metal3 s 1694 1219 1792 1317 4 vdd
port 2 nsew
rlabel metal3 s 31658 381 31756 479 4 vdd
port 2 nsew
rlabel metal3 s 0 2164 36818 2224 4 en
port 3 nsew
rlabel metal1 s 1570 1130 1604 2256 4 bl_0
port 4 nsew
rlabel metal1 s 1646 1142 1674 2256 4 br_0
port 5 nsew
rlabel metal1 s 1478 0 1524 254 4 data_0
port 6 nsew
rlabel metal1 s 6562 1130 6596 2256 4 bl_1
port 7 nsew
rlabel metal1 s 6638 1142 6666 2256 4 br_1
port 8 nsew
rlabel metal1 s 6470 0 6516 254 4 data_1
port 9 nsew
rlabel metal1 s 11554 1130 11588 2256 4 bl_2
port 10 nsew
rlabel metal1 s 11630 1142 11658 2256 4 br_2
port 11 nsew
rlabel metal1 s 11462 0 11508 254 4 data_2
port 12 nsew
rlabel metal1 s 16546 1130 16580 2256 4 bl_3
port 13 nsew
rlabel metal1 s 16622 1142 16650 2256 4 br_3
port 14 nsew
rlabel metal1 s 16454 0 16500 254 4 data_3
port 15 nsew
rlabel metal1 s 21538 1130 21572 2256 4 bl_4
port 16 nsew
rlabel metal1 s 21614 1142 21642 2256 4 br_4
port 17 nsew
rlabel metal1 s 21446 0 21492 254 4 data_4
port 18 nsew
rlabel metal1 s 26530 1130 26564 2256 4 bl_5
port 19 nsew
rlabel metal1 s 26606 1142 26634 2256 4 br_5
port 20 nsew
rlabel metal1 s 26438 0 26484 254 4 data_5
port 21 nsew
rlabel metal1 s 31522 1130 31556 2256 4 bl_6
port 22 nsew
rlabel metal1 s 31598 1142 31626 2256 4 br_6
port 23 nsew
rlabel metal1 s 31430 0 31476 254 4 data_6
port 24 nsew
rlabel metal1 s 36514 1130 36548 2256 4 bl_7
port 25 nsew
rlabel metal1 s 36590 1142 36618 2256 4 br_7
port 26 nsew
rlabel metal1 s 36422 0 36468 254 4 data_7
port 27 nsew
<< properties >>
string FIXED_BBOX 0 0 36818 2256
string GDS_END 1091860
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 1072788
<< end >>
