magic
tech sky130B
magscale 1 2
timestamp 1666199351
use sky130_fd_pr__hvdfl1sd__example_55959141808137  sky130_fd_pr__hvdfl1sd__example_55959141808137_0
timestamp 1666199351
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808449  sky130_fd_pr__hvdfm1sd2__example_55959141808449_0
timestamp 1666199351
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808200  sky130_fd_pr__hvdfm1sd__example_55959141808200_0
timestamp 1666199351
transform 1 0 296 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 30063970
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30062398
<< end >>
