magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< pwell >>
rect 15 163 1347 1633
<< mvnmos >>
rect 241 189 341 1607
rect 397 189 497 1607
rect 553 189 653 1607
rect 709 189 809 1607
rect 865 189 965 1607
rect 1021 189 1121 1607
<< mvndiff >>
rect 181 1595 241 1607
rect 181 1561 196 1595
rect 230 1561 241 1595
rect 181 1527 241 1561
rect 181 1493 196 1527
rect 230 1493 241 1527
rect 181 1459 241 1493
rect 181 1425 196 1459
rect 230 1425 241 1459
rect 181 1391 241 1425
rect 181 1357 196 1391
rect 230 1357 241 1391
rect 181 1323 241 1357
rect 181 1289 196 1323
rect 230 1289 241 1323
rect 181 1255 241 1289
rect 181 1221 196 1255
rect 230 1221 241 1255
rect 181 1187 241 1221
rect 181 1153 196 1187
rect 230 1153 241 1187
rect 181 1119 241 1153
rect 181 1085 196 1119
rect 230 1085 241 1119
rect 181 1051 241 1085
rect 181 1017 196 1051
rect 230 1017 241 1051
rect 181 983 241 1017
rect 181 949 196 983
rect 230 949 241 983
rect 181 915 241 949
rect 181 881 196 915
rect 230 881 241 915
rect 181 847 241 881
rect 181 813 196 847
rect 230 813 241 847
rect 181 779 241 813
rect 181 745 196 779
rect 230 745 241 779
rect 181 711 241 745
rect 181 677 196 711
rect 230 677 241 711
rect 181 643 241 677
rect 181 609 196 643
rect 230 609 241 643
rect 181 575 241 609
rect 181 541 196 575
rect 230 541 241 575
rect 181 507 241 541
rect 181 473 196 507
rect 230 473 241 507
rect 181 439 241 473
rect 181 405 196 439
rect 230 405 241 439
rect 181 371 241 405
rect 181 337 196 371
rect 230 337 241 371
rect 181 303 241 337
rect 181 269 196 303
rect 230 269 241 303
rect 181 235 241 269
rect 181 201 196 235
rect 230 201 241 235
rect 181 189 241 201
rect 341 1595 397 1607
rect 341 1561 352 1595
rect 386 1561 397 1595
rect 341 1527 397 1561
rect 341 1493 352 1527
rect 386 1493 397 1527
rect 341 1459 397 1493
rect 341 1425 352 1459
rect 386 1425 397 1459
rect 341 1391 397 1425
rect 341 1357 352 1391
rect 386 1357 397 1391
rect 341 1323 397 1357
rect 341 1289 352 1323
rect 386 1289 397 1323
rect 341 1255 397 1289
rect 341 1221 352 1255
rect 386 1221 397 1255
rect 341 1187 397 1221
rect 341 1153 352 1187
rect 386 1153 397 1187
rect 341 1119 397 1153
rect 341 1085 352 1119
rect 386 1085 397 1119
rect 341 1051 397 1085
rect 341 1017 352 1051
rect 386 1017 397 1051
rect 341 983 397 1017
rect 341 949 352 983
rect 386 949 397 983
rect 341 915 397 949
rect 341 881 352 915
rect 386 881 397 915
rect 341 847 397 881
rect 341 813 352 847
rect 386 813 397 847
rect 341 779 397 813
rect 341 745 352 779
rect 386 745 397 779
rect 341 711 397 745
rect 341 677 352 711
rect 386 677 397 711
rect 341 643 397 677
rect 341 609 352 643
rect 386 609 397 643
rect 341 575 397 609
rect 341 541 352 575
rect 386 541 397 575
rect 341 507 397 541
rect 341 473 352 507
rect 386 473 397 507
rect 341 439 397 473
rect 341 405 352 439
rect 386 405 397 439
rect 341 371 397 405
rect 341 337 352 371
rect 386 337 397 371
rect 341 303 397 337
rect 341 269 352 303
rect 386 269 397 303
rect 341 235 397 269
rect 341 201 352 235
rect 386 201 397 235
rect 341 189 397 201
rect 497 1595 553 1607
rect 497 1561 508 1595
rect 542 1561 553 1595
rect 497 1527 553 1561
rect 497 1493 508 1527
rect 542 1493 553 1527
rect 497 1459 553 1493
rect 497 1425 508 1459
rect 542 1425 553 1459
rect 497 1391 553 1425
rect 497 1357 508 1391
rect 542 1357 553 1391
rect 497 1323 553 1357
rect 497 1289 508 1323
rect 542 1289 553 1323
rect 497 1255 553 1289
rect 497 1221 508 1255
rect 542 1221 553 1255
rect 497 1187 553 1221
rect 497 1153 508 1187
rect 542 1153 553 1187
rect 497 1119 553 1153
rect 497 1085 508 1119
rect 542 1085 553 1119
rect 497 1051 553 1085
rect 497 1017 508 1051
rect 542 1017 553 1051
rect 497 983 553 1017
rect 497 949 508 983
rect 542 949 553 983
rect 497 915 553 949
rect 497 881 508 915
rect 542 881 553 915
rect 497 847 553 881
rect 497 813 508 847
rect 542 813 553 847
rect 497 779 553 813
rect 497 745 508 779
rect 542 745 553 779
rect 497 711 553 745
rect 497 677 508 711
rect 542 677 553 711
rect 497 643 553 677
rect 497 609 508 643
rect 542 609 553 643
rect 497 575 553 609
rect 497 541 508 575
rect 542 541 553 575
rect 497 507 553 541
rect 497 473 508 507
rect 542 473 553 507
rect 497 439 553 473
rect 497 405 508 439
rect 542 405 553 439
rect 497 371 553 405
rect 497 337 508 371
rect 542 337 553 371
rect 497 303 553 337
rect 497 269 508 303
rect 542 269 553 303
rect 497 235 553 269
rect 497 201 508 235
rect 542 201 553 235
rect 497 189 553 201
rect 653 1595 709 1607
rect 653 1561 664 1595
rect 698 1561 709 1595
rect 653 1527 709 1561
rect 653 1493 664 1527
rect 698 1493 709 1527
rect 653 1459 709 1493
rect 653 1425 664 1459
rect 698 1425 709 1459
rect 653 1391 709 1425
rect 653 1357 664 1391
rect 698 1357 709 1391
rect 653 1323 709 1357
rect 653 1289 664 1323
rect 698 1289 709 1323
rect 653 1255 709 1289
rect 653 1221 664 1255
rect 698 1221 709 1255
rect 653 1187 709 1221
rect 653 1153 664 1187
rect 698 1153 709 1187
rect 653 1119 709 1153
rect 653 1085 664 1119
rect 698 1085 709 1119
rect 653 1051 709 1085
rect 653 1017 664 1051
rect 698 1017 709 1051
rect 653 983 709 1017
rect 653 949 664 983
rect 698 949 709 983
rect 653 915 709 949
rect 653 881 664 915
rect 698 881 709 915
rect 653 847 709 881
rect 653 813 664 847
rect 698 813 709 847
rect 653 779 709 813
rect 653 745 664 779
rect 698 745 709 779
rect 653 711 709 745
rect 653 677 664 711
rect 698 677 709 711
rect 653 643 709 677
rect 653 609 664 643
rect 698 609 709 643
rect 653 575 709 609
rect 653 541 664 575
rect 698 541 709 575
rect 653 507 709 541
rect 653 473 664 507
rect 698 473 709 507
rect 653 439 709 473
rect 653 405 664 439
rect 698 405 709 439
rect 653 371 709 405
rect 653 337 664 371
rect 698 337 709 371
rect 653 303 709 337
rect 653 269 664 303
rect 698 269 709 303
rect 653 235 709 269
rect 653 201 664 235
rect 698 201 709 235
rect 653 189 709 201
rect 809 1595 865 1607
rect 809 1561 820 1595
rect 854 1561 865 1595
rect 809 1527 865 1561
rect 809 1493 820 1527
rect 854 1493 865 1527
rect 809 1459 865 1493
rect 809 1425 820 1459
rect 854 1425 865 1459
rect 809 1391 865 1425
rect 809 1357 820 1391
rect 854 1357 865 1391
rect 809 1323 865 1357
rect 809 1289 820 1323
rect 854 1289 865 1323
rect 809 1255 865 1289
rect 809 1221 820 1255
rect 854 1221 865 1255
rect 809 1187 865 1221
rect 809 1153 820 1187
rect 854 1153 865 1187
rect 809 1119 865 1153
rect 809 1085 820 1119
rect 854 1085 865 1119
rect 809 1051 865 1085
rect 809 1017 820 1051
rect 854 1017 865 1051
rect 809 983 865 1017
rect 809 949 820 983
rect 854 949 865 983
rect 809 915 865 949
rect 809 881 820 915
rect 854 881 865 915
rect 809 847 865 881
rect 809 813 820 847
rect 854 813 865 847
rect 809 779 865 813
rect 809 745 820 779
rect 854 745 865 779
rect 809 711 865 745
rect 809 677 820 711
rect 854 677 865 711
rect 809 643 865 677
rect 809 609 820 643
rect 854 609 865 643
rect 809 575 865 609
rect 809 541 820 575
rect 854 541 865 575
rect 809 507 865 541
rect 809 473 820 507
rect 854 473 865 507
rect 809 439 865 473
rect 809 405 820 439
rect 854 405 865 439
rect 809 371 865 405
rect 809 337 820 371
rect 854 337 865 371
rect 809 303 865 337
rect 809 269 820 303
rect 854 269 865 303
rect 809 235 865 269
rect 809 201 820 235
rect 854 201 865 235
rect 809 189 865 201
rect 965 1595 1021 1607
rect 965 1561 976 1595
rect 1010 1561 1021 1595
rect 965 1527 1021 1561
rect 965 1493 976 1527
rect 1010 1493 1021 1527
rect 965 1459 1021 1493
rect 965 1425 976 1459
rect 1010 1425 1021 1459
rect 965 1391 1021 1425
rect 965 1357 976 1391
rect 1010 1357 1021 1391
rect 965 1323 1021 1357
rect 965 1289 976 1323
rect 1010 1289 1021 1323
rect 965 1255 1021 1289
rect 965 1221 976 1255
rect 1010 1221 1021 1255
rect 965 1187 1021 1221
rect 965 1153 976 1187
rect 1010 1153 1021 1187
rect 965 1119 1021 1153
rect 965 1085 976 1119
rect 1010 1085 1021 1119
rect 965 1051 1021 1085
rect 965 1017 976 1051
rect 1010 1017 1021 1051
rect 965 983 1021 1017
rect 965 949 976 983
rect 1010 949 1021 983
rect 965 915 1021 949
rect 965 881 976 915
rect 1010 881 1021 915
rect 965 847 1021 881
rect 965 813 976 847
rect 1010 813 1021 847
rect 965 779 1021 813
rect 965 745 976 779
rect 1010 745 1021 779
rect 965 711 1021 745
rect 965 677 976 711
rect 1010 677 1021 711
rect 965 643 1021 677
rect 965 609 976 643
rect 1010 609 1021 643
rect 965 575 1021 609
rect 965 541 976 575
rect 1010 541 1021 575
rect 965 507 1021 541
rect 965 473 976 507
rect 1010 473 1021 507
rect 965 439 1021 473
rect 965 405 976 439
rect 1010 405 1021 439
rect 965 371 1021 405
rect 965 337 976 371
rect 1010 337 1021 371
rect 965 303 1021 337
rect 965 269 976 303
rect 1010 269 1021 303
rect 965 235 1021 269
rect 965 201 976 235
rect 1010 201 1021 235
rect 965 189 1021 201
rect 1121 1595 1181 1607
rect 1121 1561 1132 1595
rect 1166 1561 1181 1595
rect 1121 1527 1181 1561
rect 1121 1493 1132 1527
rect 1166 1493 1181 1527
rect 1121 1459 1181 1493
rect 1121 1425 1132 1459
rect 1166 1425 1181 1459
rect 1121 1391 1181 1425
rect 1121 1357 1132 1391
rect 1166 1357 1181 1391
rect 1121 1323 1181 1357
rect 1121 1289 1132 1323
rect 1166 1289 1181 1323
rect 1121 1255 1181 1289
rect 1121 1221 1132 1255
rect 1166 1221 1181 1255
rect 1121 1187 1181 1221
rect 1121 1153 1132 1187
rect 1166 1153 1181 1187
rect 1121 1119 1181 1153
rect 1121 1085 1132 1119
rect 1166 1085 1181 1119
rect 1121 1051 1181 1085
rect 1121 1017 1132 1051
rect 1166 1017 1181 1051
rect 1121 983 1181 1017
rect 1121 949 1132 983
rect 1166 949 1181 983
rect 1121 915 1181 949
rect 1121 881 1132 915
rect 1166 881 1181 915
rect 1121 847 1181 881
rect 1121 813 1132 847
rect 1166 813 1181 847
rect 1121 779 1181 813
rect 1121 745 1132 779
rect 1166 745 1181 779
rect 1121 711 1181 745
rect 1121 677 1132 711
rect 1166 677 1181 711
rect 1121 643 1181 677
rect 1121 609 1132 643
rect 1166 609 1181 643
rect 1121 575 1181 609
rect 1121 541 1132 575
rect 1166 541 1181 575
rect 1121 507 1181 541
rect 1121 473 1132 507
rect 1166 473 1181 507
rect 1121 439 1181 473
rect 1121 405 1132 439
rect 1166 405 1181 439
rect 1121 371 1181 405
rect 1121 337 1132 371
rect 1166 337 1181 371
rect 1121 303 1181 337
rect 1121 269 1132 303
rect 1166 269 1181 303
rect 1121 235 1181 269
rect 1121 201 1132 235
rect 1166 201 1181 235
rect 1121 189 1181 201
<< mvndiffc >>
rect 196 1561 230 1595
rect 196 1493 230 1527
rect 196 1425 230 1459
rect 196 1357 230 1391
rect 196 1289 230 1323
rect 196 1221 230 1255
rect 196 1153 230 1187
rect 196 1085 230 1119
rect 196 1017 230 1051
rect 196 949 230 983
rect 196 881 230 915
rect 196 813 230 847
rect 196 745 230 779
rect 196 677 230 711
rect 196 609 230 643
rect 196 541 230 575
rect 196 473 230 507
rect 196 405 230 439
rect 196 337 230 371
rect 196 269 230 303
rect 196 201 230 235
rect 352 1561 386 1595
rect 352 1493 386 1527
rect 352 1425 386 1459
rect 352 1357 386 1391
rect 352 1289 386 1323
rect 352 1221 386 1255
rect 352 1153 386 1187
rect 352 1085 386 1119
rect 352 1017 386 1051
rect 352 949 386 983
rect 352 881 386 915
rect 352 813 386 847
rect 352 745 386 779
rect 352 677 386 711
rect 352 609 386 643
rect 352 541 386 575
rect 352 473 386 507
rect 352 405 386 439
rect 352 337 386 371
rect 352 269 386 303
rect 352 201 386 235
rect 508 1561 542 1595
rect 508 1493 542 1527
rect 508 1425 542 1459
rect 508 1357 542 1391
rect 508 1289 542 1323
rect 508 1221 542 1255
rect 508 1153 542 1187
rect 508 1085 542 1119
rect 508 1017 542 1051
rect 508 949 542 983
rect 508 881 542 915
rect 508 813 542 847
rect 508 745 542 779
rect 508 677 542 711
rect 508 609 542 643
rect 508 541 542 575
rect 508 473 542 507
rect 508 405 542 439
rect 508 337 542 371
rect 508 269 542 303
rect 508 201 542 235
rect 664 1561 698 1595
rect 664 1493 698 1527
rect 664 1425 698 1459
rect 664 1357 698 1391
rect 664 1289 698 1323
rect 664 1221 698 1255
rect 664 1153 698 1187
rect 664 1085 698 1119
rect 664 1017 698 1051
rect 664 949 698 983
rect 664 881 698 915
rect 664 813 698 847
rect 664 745 698 779
rect 664 677 698 711
rect 664 609 698 643
rect 664 541 698 575
rect 664 473 698 507
rect 664 405 698 439
rect 664 337 698 371
rect 664 269 698 303
rect 664 201 698 235
rect 820 1561 854 1595
rect 820 1493 854 1527
rect 820 1425 854 1459
rect 820 1357 854 1391
rect 820 1289 854 1323
rect 820 1221 854 1255
rect 820 1153 854 1187
rect 820 1085 854 1119
rect 820 1017 854 1051
rect 820 949 854 983
rect 820 881 854 915
rect 820 813 854 847
rect 820 745 854 779
rect 820 677 854 711
rect 820 609 854 643
rect 820 541 854 575
rect 820 473 854 507
rect 820 405 854 439
rect 820 337 854 371
rect 820 269 854 303
rect 820 201 854 235
rect 976 1561 1010 1595
rect 976 1493 1010 1527
rect 976 1425 1010 1459
rect 976 1357 1010 1391
rect 976 1289 1010 1323
rect 976 1221 1010 1255
rect 976 1153 1010 1187
rect 976 1085 1010 1119
rect 976 1017 1010 1051
rect 976 949 1010 983
rect 976 881 1010 915
rect 976 813 1010 847
rect 976 745 1010 779
rect 976 677 1010 711
rect 976 609 1010 643
rect 976 541 1010 575
rect 976 473 1010 507
rect 976 405 1010 439
rect 976 337 1010 371
rect 976 269 1010 303
rect 976 201 1010 235
rect 1132 1561 1166 1595
rect 1132 1493 1166 1527
rect 1132 1425 1166 1459
rect 1132 1357 1166 1391
rect 1132 1289 1166 1323
rect 1132 1221 1166 1255
rect 1132 1153 1166 1187
rect 1132 1085 1166 1119
rect 1132 1017 1166 1051
rect 1132 949 1166 983
rect 1132 881 1166 915
rect 1132 813 1166 847
rect 1132 745 1166 779
rect 1132 677 1166 711
rect 1132 609 1166 643
rect 1132 541 1166 575
rect 1132 473 1166 507
rect 1132 405 1166 439
rect 1132 337 1166 371
rect 1132 269 1166 303
rect 1132 201 1166 235
<< mvpsubdiff >>
rect 41 1595 181 1607
rect 41 201 60 1595
rect 162 201 181 1595
rect 41 189 181 201
rect 1181 1595 1321 1607
rect 1181 201 1200 1595
rect 1302 201 1321 1595
rect 1181 189 1321 201
<< mvpsubdiffcont >>
rect 60 201 162 1595
rect 1200 201 1302 1595
<< poly >>
rect 383 1775 979 1796
rect 190 1683 341 1699
rect 190 1649 206 1683
rect 240 1649 341 1683
rect 383 1673 426 1775
rect 936 1673 979 1775
rect 383 1657 979 1673
rect 1021 1683 1172 1699
rect 190 1633 341 1649
rect 241 1607 341 1633
rect 397 1607 497 1657
rect 553 1607 653 1657
rect 709 1607 809 1657
rect 865 1607 965 1657
rect 1021 1649 1122 1683
rect 1156 1649 1172 1683
rect 1021 1633 1172 1649
rect 1021 1607 1121 1633
rect 241 163 341 189
rect 190 147 341 163
rect 190 113 206 147
rect 240 113 341 147
rect 397 139 497 189
rect 553 139 653 189
rect 709 139 809 189
rect 865 139 965 189
rect 1021 163 1121 189
rect 1021 147 1172 163
rect 190 97 341 113
rect 383 123 979 139
rect 383 21 426 123
rect 936 21 979 123
rect 1021 113 1122 147
rect 1156 113 1172 147
rect 1021 97 1172 113
rect 383 0 979 21
<< polycont >>
rect 206 1649 240 1683
rect 426 1673 936 1775
rect 1122 1649 1156 1683
rect 206 113 240 147
rect 426 21 936 123
rect 1122 113 1156 147
<< locali >>
rect 400 1777 962 1796
rect 190 1683 256 1699
rect 190 1649 206 1683
rect 240 1649 256 1683
rect 400 1671 412 1777
rect 950 1671 962 1777
rect 400 1659 962 1671
rect 1106 1683 1172 1699
rect 190 1633 256 1649
rect 1106 1649 1122 1683
rect 1156 1649 1172 1683
rect 1106 1633 1172 1649
rect 190 1611 230 1633
rect 1132 1611 1172 1633
rect 41 1595 230 1611
rect 41 201 60 1595
rect 162 1561 196 1595
rect 162 1527 230 1561
rect 162 1493 196 1527
rect 162 1459 230 1493
rect 162 1425 196 1459
rect 162 1391 230 1425
rect 162 1357 196 1391
rect 162 1323 230 1357
rect 162 1289 196 1323
rect 162 1255 230 1289
rect 162 1221 196 1255
rect 162 1187 230 1221
rect 162 1153 196 1187
rect 162 1119 230 1153
rect 162 1085 196 1119
rect 162 1051 230 1085
rect 162 1017 196 1051
rect 162 983 230 1017
rect 162 949 196 983
rect 162 915 230 949
rect 162 881 196 915
rect 162 847 230 881
rect 162 813 196 847
rect 162 779 230 813
rect 162 745 196 779
rect 162 711 230 745
rect 162 677 196 711
rect 162 643 230 677
rect 162 609 196 643
rect 162 575 230 609
rect 162 541 196 575
rect 162 507 230 541
rect 162 473 196 507
rect 162 439 230 473
rect 162 405 196 439
rect 162 371 230 405
rect 162 337 196 371
rect 162 303 230 337
rect 162 269 196 303
rect 162 235 230 269
rect 162 201 196 235
rect 41 185 230 201
rect 352 1595 386 1611
rect 352 1527 386 1529
rect 352 1491 386 1493
rect 352 1419 386 1425
rect 352 1347 386 1357
rect 352 1275 386 1289
rect 352 1203 386 1221
rect 352 1131 386 1153
rect 352 1059 386 1085
rect 352 987 386 1017
rect 352 915 386 949
rect 352 847 386 881
rect 352 779 386 809
rect 352 711 386 737
rect 352 643 386 665
rect 352 575 386 593
rect 352 507 386 521
rect 352 439 386 449
rect 352 371 386 377
rect 352 303 386 305
rect 352 267 386 269
rect 352 185 386 201
rect 508 1595 542 1611
rect 508 1527 542 1529
rect 508 1491 542 1493
rect 508 1419 542 1425
rect 508 1347 542 1357
rect 508 1275 542 1289
rect 508 1203 542 1221
rect 508 1131 542 1153
rect 508 1059 542 1085
rect 508 987 542 1017
rect 508 915 542 949
rect 508 847 542 881
rect 508 779 542 809
rect 508 711 542 737
rect 508 643 542 665
rect 508 575 542 593
rect 508 507 542 521
rect 508 439 542 449
rect 508 371 542 377
rect 508 303 542 305
rect 508 267 542 269
rect 508 185 542 201
rect 664 1595 698 1611
rect 664 1527 698 1529
rect 664 1491 698 1493
rect 664 1419 698 1425
rect 664 1347 698 1357
rect 664 1275 698 1289
rect 664 1203 698 1221
rect 664 1131 698 1153
rect 664 1059 698 1085
rect 664 987 698 1017
rect 664 915 698 949
rect 664 847 698 881
rect 664 779 698 809
rect 664 711 698 737
rect 664 643 698 665
rect 664 575 698 593
rect 664 507 698 521
rect 664 439 698 449
rect 664 371 698 377
rect 664 303 698 305
rect 664 267 698 269
rect 664 185 698 201
rect 820 1595 854 1611
rect 820 1527 854 1529
rect 820 1491 854 1493
rect 820 1419 854 1425
rect 820 1347 854 1357
rect 820 1275 854 1289
rect 820 1203 854 1221
rect 820 1131 854 1153
rect 820 1059 854 1085
rect 820 987 854 1017
rect 820 915 854 949
rect 820 847 854 881
rect 820 779 854 809
rect 820 711 854 737
rect 820 643 854 665
rect 820 575 854 593
rect 820 507 854 521
rect 820 439 854 449
rect 820 371 854 377
rect 820 303 854 305
rect 820 267 854 269
rect 820 185 854 201
rect 976 1595 1010 1611
rect 976 1527 1010 1529
rect 976 1491 1010 1493
rect 976 1419 1010 1425
rect 976 1347 1010 1357
rect 976 1275 1010 1289
rect 976 1203 1010 1221
rect 976 1131 1010 1153
rect 976 1059 1010 1085
rect 976 987 1010 1017
rect 976 915 1010 949
rect 976 847 1010 881
rect 976 779 1010 809
rect 976 711 1010 737
rect 976 643 1010 665
rect 976 575 1010 593
rect 976 507 1010 521
rect 976 439 1010 449
rect 976 371 1010 377
rect 976 303 1010 305
rect 976 267 1010 269
rect 976 185 1010 201
rect 1132 1595 1321 1611
rect 1166 1561 1200 1595
rect 1132 1527 1200 1561
rect 1166 1493 1200 1527
rect 1132 1459 1200 1493
rect 1166 1425 1200 1459
rect 1132 1391 1200 1425
rect 1166 1357 1200 1391
rect 1132 1323 1200 1357
rect 1166 1289 1200 1323
rect 1132 1255 1200 1289
rect 1166 1221 1200 1255
rect 1132 1187 1200 1221
rect 1166 1153 1200 1187
rect 1132 1119 1200 1153
rect 1166 1085 1200 1119
rect 1132 1051 1200 1085
rect 1166 1017 1200 1051
rect 1132 983 1200 1017
rect 1166 949 1200 983
rect 1132 915 1200 949
rect 1166 881 1200 915
rect 1132 847 1200 881
rect 1166 813 1200 847
rect 1132 779 1200 813
rect 1166 745 1200 779
rect 1132 711 1200 745
rect 1166 677 1200 711
rect 1132 643 1200 677
rect 1166 609 1200 643
rect 1132 575 1200 609
rect 1166 541 1200 575
rect 1132 507 1200 541
rect 1166 473 1200 507
rect 1132 439 1200 473
rect 1166 405 1200 439
rect 1132 371 1200 405
rect 1166 337 1200 371
rect 1132 303 1200 337
rect 1166 269 1200 303
rect 1132 235 1200 269
rect 1166 201 1200 235
rect 1302 201 1321 1595
rect 1132 185 1321 201
rect 190 163 230 185
rect 1132 163 1172 185
rect 190 147 256 163
rect 190 113 206 147
rect 240 113 256 147
rect 1106 147 1172 163
rect 190 97 256 113
rect 400 125 962 137
rect 400 19 412 125
rect 950 19 962 125
rect 1106 113 1122 147
rect 1156 113 1172 147
rect 1106 97 1172 113
rect 400 0 962 19
<< viali >>
rect 412 1775 950 1777
rect 412 1673 426 1775
rect 426 1673 936 1775
rect 936 1673 950 1775
rect 412 1671 950 1673
rect 60 1529 94 1563
rect 60 1457 94 1491
rect 60 1385 94 1419
rect 60 1313 94 1347
rect 60 1241 94 1275
rect 60 1169 94 1203
rect 60 1097 94 1131
rect 60 1025 94 1059
rect 60 953 94 987
rect 60 881 94 915
rect 60 809 94 843
rect 60 737 94 771
rect 60 665 94 699
rect 60 593 94 627
rect 60 521 94 555
rect 60 449 94 483
rect 60 377 94 411
rect 60 305 94 339
rect 60 233 94 267
rect 352 1561 386 1563
rect 352 1529 386 1561
rect 352 1459 386 1491
rect 352 1457 386 1459
rect 352 1391 386 1419
rect 352 1385 386 1391
rect 352 1323 386 1347
rect 352 1313 386 1323
rect 352 1255 386 1275
rect 352 1241 386 1255
rect 352 1187 386 1203
rect 352 1169 386 1187
rect 352 1119 386 1131
rect 352 1097 386 1119
rect 352 1051 386 1059
rect 352 1025 386 1051
rect 352 983 386 987
rect 352 953 386 983
rect 352 881 386 915
rect 352 813 386 843
rect 352 809 386 813
rect 352 745 386 771
rect 352 737 386 745
rect 352 677 386 699
rect 352 665 386 677
rect 352 609 386 627
rect 352 593 386 609
rect 352 541 386 555
rect 352 521 386 541
rect 352 473 386 483
rect 352 449 386 473
rect 352 405 386 411
rect 352 377 386 405
rect 352 337 386 339
rect 352 305 386 337
rect 352 235 386 267
rect 352 233 386 235
rect 508 1561 542 1563
rect 508 1529 542 1561
rect 508 1459 542 1491
rect 508 1457 542 1459
rect 508 1391 542 1419
rect 508 1385 542 1391
rect 508 1323 542 1347
rect 508 1313 542 1323
rect 508 1255 542 1275
rect 508 1241 542 1255
rect 508 1187 542 1203
rect 508 1169 542 1187
rect 508 1119 542 1131
rect 508 1097 542 1119
rect 508 1051 542 1059
rect 508 1025 542 1051
rect 508 983 542 987
rect 508 953 542 983
rect 508 881 542 915
rect 508 813 542 843
rect 508 809 542 813
rect 508 745 542 771
rect 508 737 542 745
rect 508 677 542 699
rect 508 665 542 677
rect 508 609 542 627
rect 508 593 542 609
rect 508 541 542 555
rect 508 521 542 541
rect 508 473 542 483
rect 508 449 542 473
rect 508 405 542 411
rect 508 377 542 405
rect 508 337 542 339
rect 508 305 542 337
rect 508 235 542 267
rect 508 233 542 235
rect 664 1561 698 1563
rect 664 1529 698 1561
rect 664 1459 698 1491
rect 664 1457 698 1459
rect 664 1391 698 1419
rect 664 1385 698 1391
rect 664 1323 698 1347
rect 664 1313 698 1323
rect 664 1255 698 1275
rect 664 1241 698 1255
rect 664 1187 698 1203
rect 664 1169 698 1187
rect 664 1119 698 1131
rect 664 1097 698 1119
rect 664 1051 698 1059
rect 664 1025 698 1051
rect 664 983 698 987
rect 664 953 698 983
rect 664 881 698 915
rect 664 813 698 843
rect 664 809 698 813
rect 664 745 698 771
rect 664 737 698 745
rect 664 677 698 699
rect 664 665 698 677
rect 664 609 698 627
rect 664 593 698 609
rect 664 541 698 555
rect 664 521 698 541
rect 664 473 698 483
rect 664 449 698 473
rect 664 405 698 411
rect 664 377 698 405
rect 664 337 698 339
rect 664 305 698 337
rect 664 235 698 267
rect 664 233 698 235
rect 820 1561 854 1563
rect 820 1529 854 1561
rect 820 1459 854 1491
rect 820 1457 854 1459
rect 820 1391 854 1419
rect 820 1385 854 1391
rect 820 1323 854 1347
rect 820 1313 854 1323
rect 820 1255 854 1275
rect 820 1241 854 1255
rect 820 1187 854 1203
rect 820 1169 854 1187
rect 820 1119 854 1131
rect 820 1097 854 1119
rect 820 1051 854 1059
rect 820 1025 854 1051
rect 820 983 854 987
rect 820 953 854 983
rect 820 881 854 915
rect 820 813 854 843
rect 820 809 854 813
rect 820 745 854 771
rect 820 737 854 745
rect 820 677 854 699
rect 820 665 854 677
rect 820 609 854 627
rect 820 593 854 609
rect 820 541 854 555
rect 820 521 854 541
rect 820 473 854 483
rect 820 449 854 473
rect 820 405 854 411
rect 820 377 854 405
rect 820 337 854 339
rect 820 305 854 337
rect 820 235 854 267
rect 820 233 854 235
rect 976 1561 1010 1563
rect 976 1529 1010 1561
rect 976 1459 1010 1491
rect 976 1457 1010 1459
rect 976 1391 1010 1419
rect 976 1385 1010 1391
rect 976 1323 1010 1347
rect 976 1313 1010 1323
rect 976 1255 1010 1275
rect 976 1241 1010 1255
rect 976 1187 1010 1203
rect 976 1169 1010 1187
rect 976 1119 1010 1131
rect 976 1097 1010 1119
rect 976 1051 1010 1059
rect 976 1025 1010 1051
rect 976 983 1010 987
rect 976 953 1010 983
rect 976 881 1010 915
rect 976 813 1010 843
rect 976 809 1010 813
rect 976 745 1010 771
rect 976 737 1010 745
rect 976 677 1010 699
rect 976 665 1010 677
rect 976 609 1010 627
rect 976 593 1010 609
rect 976 541 1010 555
rect 976 521 1010 541
rect 976 473 1010 483
rect 976 449 1010 473
rect 976 405 1010 411
rect 976 377 1010 405
rect 976 337 1010 339
rect 976 305 1010 337
rect 976 235 1010 267
rect 976 233 1010 235
rect 1268 1529 1302 1563
rect 1268 1457 1302 1491
rect 1268 1385 1302 1419
rect 1268 1313 1302 1347
rect 1268 1241 1302 1275
rect 1268 1169 1302 1203
rect 1268 1097 1302 1131
rect 1268 1025 1302 1059
rect 1268 953 1302 987
rect 1268 881 1302 915
rect 1268 809 1302 843
rect 1268 737 1302 771
rect 1268 665 1302 699
rect 1268 593 1302 627
rect 1268 521 1302 555
rect 1268 449 1302 483
rect 1268 377 1302 411
rect 1268 305 1302 339
rect 1268 233 1302 267
rect 412 123 950 125
rect 412 21 426 123
rect 426 21 936 123
rect 936 21 950 123
rect 412 19 950 21
<< metal1 >>
rect 400 1777 962 1796
rect 400 1671 412 1777
rect 950 1671 962 1777
rect 400 1659 962 1671
rect 41 1563 100 1594
rect 41 1529 60 1563
rect 94 1529 100 1563
rect 41 1491 100 1529
rect 41 1457 60 1491
rect 94 1457 100 1491
rect 41 1419 100 1457
rect 41 1385 60 1419
rect 94 1385 100 1419
rect 41 1347 100 1385
rect 41 1313 60 1347
rect 94 1313 100 1347
rect 41 1275 100 1313
rect 41 1241 60 1275
rect 94 1241 100 1275
rect 41 1203 100 1241
rect 41 1169 60 1203
rect 94 1169 100 1203
rect 41 1131 100 1169
rect 41 1097 60 1131
rect 94 1097 100 1131
rect 41 1059 100 1097
rect 41 1025 60 1059
rect 94 1025 100 1059
rect 41 987 100 1025
rect 41 953 60 987
rect 94 953 100 987
rect 41 915 100 953
rect 41 881 60 915
rect 94 881 100 915
rect 41 843 100 881
rect 41 809 60 843
rect 94 809 100 843
rect 41 771 100 809
rect 41 737 60 771
rect 94 737 100 771
rect 41 699 100 737
rect 41 665 60 699
rect 94 665 100 699
rect 41 627 100 665
rect 41 593 60 627
rect 94 593 100 627
rect 41 555 100 593
rect 41 521 60 555
rect 94 521 100 555
rect 41 483 100 521
rect 41 449 60 483
rect 94 449 100 483
rect 41 411 100 449
rect 41 377 60 411
rect 94 377 100 411
rect 41 339 100 377
rect 41 305 60 339
rect 94 305 100 339
rect 41 267 100 305
rect 41 233 60 267
rect 94 233 100 267
rect 41 202 100 233
rect 343 1588 395 1594
rect 343 1529 352 1536
rect 386 1529 395 1536
rect 343 1524 395 1529
rect 343 1460 352 1472
rect 386 1460 395 1472
rect 343 1396 352 1408
rect 386 1396 395 1408
rect 343 1332 352 1344
rect 386 1332 395 1344
rect 343 1275 395 1280
rect 343 1241 352 1275
rect 386 1241 395 1275
rect 343 1203 395 1241
rect 343 1169 352 1203
rect 386 1169 395 1203
rect 343 1131 395 1169
rect 343 1097 352 1131
rect 386 1097 395 1131
rect 343 1059 395 1097
rect 343 1025 352 1059
rect 386 1025 395 1059
rect 343 987 395 1025
rect 343 953 352 987
rect 386 953 395 987
rect 343 915 395 953
rect 343 881 352 915
rect 386 881 395 915
rect 343 843 395 881
rect 343 809 352 843
rect 386 809 395 843
rect 343 771 395 809
rect 343 737 352 771
rect 386 737 395 771
rect 343 699 395 737
rect 343 665 352 699
rect 386 665 395 699
rect 343 627 395 665
rect 343 593 352 627
rect 386 593 395 627
rect 343 555 395 593
rect 343 521 352 555
rect 386 521 395 555
rect 343 516 395 521
rect 343 452 352 464
rect 386 452 395 464
rect 343 388 352 400
rect 386 388 395 400
rect 343 324 352 336
rect 386 324 395 336
rect 343 267 395 272
rect 343 260 352 267
rect 386 260 395 267
rect 343 202 395 208
rect 499 1563 551 1594
rect 499 1529 508 1563
rect 542 1529 551 1563
rect 499 1491 551 1529
rect 499 1457 508 1491
rect 542 1457 551 1491
rect 499 1419 551 1457
rect 499 1385 508 1419
rect 542 1385 551 1419
rect 499 1347 551 1385
rect 499 1313 508 1347
rect 542 1313 551 1347
rect 499 1275 551 1313
rect 499 1241 508 1275
rect 542 1241 551 1275
rect 499 1212 551 1241
rect 499 1148 551 1160
rect 499 1084 551 1096
rect 499 1025 508 1032
rect 542 1025 551 1032
rect 499 1020 551 1025
rect 499 956 508 968
rect 542 956 551 968
rect 499 892 508 904
rect 542 892 551 904
rect 499 828 508 840
rect 542 828 551 840
rect 499 771 551 776
rect 499 764 508 771
rect 542 764 551 771
rect 499 700 551 712
rect 499 636 551 648
rect 499 555 551 584
rect 499 521 508 555
rect 542 521 551 555
rect 499 483 551 521
rect 499 449 508 483
rect 542 449 551 483
rect 499 411 551 449
rect 499 377 508 411
rect 542 377 551 411
rect 499 339 551 377
rect 499 305 508 339
rect 542 305 551 339
rect 499 267 551 305
rect 499 233 508 267
rect 542 233 551 267
rect 499 202 551 233
rect 655 1588 707 1594
rect 655 1529 664 1536
rect 698 1529 707 1536
rect 655 1524 707 1529
rect 655 1460 664 1472
rect 698 1460 707 1472
rect 655 1396 664 1408
rect 698 1396 707 1408
rect 655 1332 664 1344
rect 698 1332 707 1344
rect 655 1275 707 1280
rect 655 1241 664 1275
rect 698 1241 707 1275
rect 655 1203 707 1241
rect 655 1169 664 1203
rect 698 1169 707 1203
rect 655 1131 707 1169
rect 655 1097 664 1131
rect 698 1097 707 1131
rect 655 1059 707 1097
rect 655 1025 664 1059
rect 698 1025 707 1059
rect 655 987 707 1025
rect 655 953 664 987
rect 698 953 707 987
rect 655 915 707 953
rect 655 881 664 915
rect 698 881 707 915
rect 655 843 707 881
rect 655 809 664 843
rect 698 809 707 843
rect 655 771 707 809
rect 655 737 664 771
rect 698 737 707 771
rect 655 699 707 737
rect 655 665 664 699
rect 698 665 707 699
rect 655 627 707 665
rect 655 593 664 627
rect 698 593 707 627
rect 655 555 707 593
rect 655 521 664 555
rect 698 521 707 555
rect 655 516 707 521
rect 655 452 664 464
rect 698 452 707 464
rect 655 388 664 400
rect 698 388 707 400
rect 655 324 664 336
rect 698 324 707 336
rect 655 267 707 272
rect 655 260 664 267
rect 698 260 707 267
rect 655 202 707 208
rect 811 1563 863 1594
rect 811 1529 820 1563
rect 854 1529 863 1563
rect 811 1491 863 1529
rect 811 1457 820 1491
rect 854 1457 863 1491
rect 811 1419 863 1457
rect 811 1385 820 1419
rect 854 1385 863 1419
rect 811 1347 863 1385
rect 811 1313 820 1347
rect 854 1313 863 1347
rect 811 1275 863 1313
rect 811 1241 820 1275
rect 854 1241 863 1275
rect 811 1212 863 1241
rect 811 1148 863 1160
rect 811 1084 863 1096
rect 811 1025 820 1032
rect 854 1025 863 1032
rect 811 1020 863 1025
rect 811 956 820 968
rect 854 956 863 968
rect 811 892 820 904
rect 854 892 863 904
rect 811 828 820 840
rect 854 828 863 840
rect 811 771 863 776
rect 811 764 820 771
rect 854 764 863 771
rect 811 700 863 712
rect 811 636 863 648
rect 811 555 863 584
rect 811 521 820 555
rect 854 521 863 555
rect 811 483 863 521
rect 811 449 820 483
rect 854 449 863 483
rect 811 411 863 449
rect 811 377 820 411
rect 854 377 863 411
rect 811 339 863 377
rect 811 305 820 339
rect 854 305 863 339
rect 811 267 863 305
rect 811 233 820 267
rect 854 233 863 267
rect 811 202 863 233
rect 967 1588 1019 1594
rect 967 1529 976 1536
rect 1010 1529 1019 1536
rect 967 1524 1019 1529
rect 967 1460 976 1472
rect 1010 1460 1019 1472
rect 967 1396 976 1408
rect 1010 1396 1019 1408
rect 967 1332 976 1344
rect 1010 1332 1019 1344
rect 967 1275 1019 1280
rect 967 1241 976 1275
rect 1010 1241 1019 1275
rect 967 1203 1019 1241
rect 967 1169 976 1203
rect 1010 1169 1019 1203
rect 967 1131 1019 1169
rect 967 1097 976 1131
rect 1010 1097 1019 1131
rect 967 1059 1019 1097
rect 967 1025 976 1059
rect 1010 1025 1019 1059
rect 967 987 1019 1025
rect 967 953 976 987
rect 1010 953 1019 987
rect 967 915 1019 953
rect 967 881 976 915
rect 1010 881 1019 915
rect 967 843 1019 881
rect 967 809 976 843
rect 1010 809 1019 843
rect 967 771 1019 809
rect 967 737 976 771
rect 1010 737 1019 771
rect 967 699 1019 737
rect 967 665 976 699
rect 1010 665 1019 699
rect 967 627 1019 665
rect 967 593 976 627
rect 1010 593 1019 627
rect 967 555 1019 593
rect 967 521 976 555
rect 1010 521 1019 555
rect 967 516 1019 521
rect 967 452 976 464
rect 1010 452 1019 464
rect 967 388 976 400
rect 1010 388 1019 400
rect 967 324 976 336
rect 1010 324 1019 336
rect 967 267 1019 272
rect 967 260 976 267
rect 1010 260 1019 267
rect 967 202 1019 208
rect 1262 1563 1321 1594
rect 1262 1529 1268 1563
rect 1302 1529 1321 1563
rect 1262 1491 1321 1529
rect 1262 1457 1268 1491
rect 1302 1457 1321 1491
rect 1262 1419 1321 1457
rect 1262 1385 1268 1419
rect 1302 1385 1321 1419
rect 1262 1347 1321 1385
rect 1262 1313 1268 1347
rect 1302 1313 1321 1347
rect 1262 1275 1321 1313
rect 1262 1241 1268 1275
rect 1302 1241 1321 1275
rect 1262 1203 1321 1241
rect 1262 1169 1268 1203
rect 1302 1169 1321 1203
rect 1262 1131 1321 1169
rect 1262 1097 1268 1131
rect 1302 1097 1321 1131
rect 1262 1059 1321 1097
rect 1262 1025 1268 1059
rect 1302 1025 1321 1059
rect 1262 987 1321 1025
rect 1262 953 1268 987
rect 1302 953 1321 987
rect 1262 915 1321 953
rect 1262 881 1268 915
rect 1302 881 1321 915
rect 1262 843 1321 881
rect 1262 809 1268 843
rect 1302 809 1321 843
rect 1262 771 1321 809
rect 1262 737 1268 771
rect 1302 737 1321 771
rect 1262 699 1321 737
rect 1262 665 1268 699
rect 1302 665 1321 699
rect 1262 627 1321 665
rect 1262 593 1268 627
rect 1302 593 1321 627
rect 1262 555 1321 593
rect 1262 521 1268 555
rect 1302 521 1321 555
rect 1262 483 1321 521
rect 1262 449 1268 483
rect 1302 449 1321 483
rect 1262 411 1321 449
rect 1262 377 1268 411
rect 1302 377 1321 411
rect 1262 339 1321 377
rect 1262 305 1268 339
rect 1302 305 1321 339
rect 1262 267 1321 305
rect 1262 233 1268 267
rect 1302 233 1321 267
rect 1262 202 1321 233
rect 400 125 962 137
rect 400 19 412 125
rect 950 19 962 125
rect 400 0 962 19
<< via1 >>
rect 343 1563 395 1588
rect 343 1536 352 1563
rect 352 1536 386 1563
rect 386 1536 395 1563
rect 343 1491 395 1524
rect 343 1472 352 1491
rect 352 1472 386 1491
rect 386 1472 395 1491
rect 343 1457 352 1460
rect 352 1457 386 1460
rect 386 1457 395 1460
rect 343 1419 395 1457
rect 343 1408 352 1419
rect 352 1408 386 1419
rect 386 1408 395 1419
rect 343 1385 352 1396
rect 352 1385 386 1396
rect 386 1385 395 1396
rect 343 1347 395 1385
rect 343 1344 352 1347
rect 352 1344 386 1347
rect 386 1344 395 1347
rect 343 1313 352 1332
rect 352 1313 386 1332
rect 386 1313 395 1332
rect 343 1280 395 1313
rect 343 483 395 516
rect 343 464 352 483
rect 352 464 386 483
rect 386 464 395 483
rect 343 449 352 452
rect 352 449 386 452
rect 386 449 395 452
rect 343 411 395 449
rect 343 400 352 411
rect 352 400 386 411
rect 386 400 395 411
rect 343 377 352 388
rect 352 377 386 388
rect 386 377 395 388
rect 343 339 395 377
rect 343 336 352 339
rect 352 336 386 339
rect 386 336 395 339
rect 343 305 352 324
rect 352 305 386 324
rect 386 305 395 324
rect 343 272 395 305
rect 343 233 352 260
rect 352 233 386 260
rect 386 233 395 260
rect 343 208 395 233
rect 499 1203 551 1212
rect 499 1169 508 1203
rect 508 1169 542 1203
rect 542 1169 551 1203
rect 499 1160 551 1169
rect 499 1131 551 1148
rect 499 1097 508 1131
rect 508 1097 542 1131
rect 542 1097 551 1131
rect 499 1096 551 1097
rect 499 1059 551 1084
rect 499 1032 508 1059
rect 508 1032 542 1059
rect 542 1032 551 1059
rect 499 987 551 1020
rect 499 968 508 987
rect 508 968 542 987
rect 542 968 551 987
rect 499 953 508 956
rect 508 953 542 956
rect 542 953 551 956
rect 499 915 551 953
rect 499 904 508 915
rect 508 904 542 915
rect 542 904 551 915
rect 499 881 508 892
rect 508 881 542 892
rect 542 881 551 892
rect 499 843 551 881
rect 499 840 508 843
rect 508 840 542 843
rect 542 840 551 843
rect 499 809 508 828
rect 508 809 542 828
rect 542 809 551 828
rect 499 776 551 809
rect 499 737 508 764
rect 508 737 542 764
rect 542 737 551 764
rect 499 712 551 737
rect 499 699 551 700
rect 499 665 508 699
rect 508 665 542 699
rect 542 665 551 699
rect 499 648 551 665
rect 499 627 551 636
rect 499 593 508 627
rect 508 593 542 627
rect 542 593 551 627
rect 499 584 551 593
rect 655 1563 707 1588
rect 655 1536 664 1563
rect 664 1536 698 1563
rect 698 1536 707 1563
rect 655 1491 707 1524
rect 655 1472 664 1491
rect 664 1472 698 1491
rect 698 1472 707 1491
rect 655 1457 664 1460
rect 664 1457 698 1460
rect 698 1457 707 1460
rect 655 1419 707 1457
rect 655 1408 664 1419
rect 664 1408 698 1419
rect 698 1408 707 1419
rect 655 1385 664 1396
rect 664 1385 698 1396
rect 698 1385 707 1396
rect 655 1347 707 1385
rect 655 1344 664 1347
rect 664 1344 698 1347
rect 698 1344 707 1347
rect 655 1313 664 1332
rect 664 1313 698 1332
rect 698 1313 707 1332
rect 655 1280 707 1313
rect 655 483 707 516
rect 655 464 664 483
rect 664 464 698 483
rect 698 464 707 483
rect 655 449 664 452
rect 664 449 698 452
rect 698 449 707 452
rect 655 411 707 449
rect 655 400 664 411
rect 664 400 698 411
rect 698 400 707 411
rect 655 377 664 388
rect 664 377 698 388
rect 698 377 707 388
rect 655 339 707 377
rect 655 336 664 339
rect 664 336 698 339
rect 698 336 707 339
rect 655 305 664 324
rect 664 305 698 324
rect 698 305 707 324
rect 655 272 707 305
rect 655 233 664 260
rect 664 233 698 260
rect 698 233 707 260
rect 655 208 707 233
rect 811 1203 863 1212
rect 811 1169 820 1203
rect 820 1169 854 1203
rect 854 1169 863 1203
rect 811 1160 863 1169
rect 811 1131 863 1148
rect 811 1097 820 1131
rect 820 1097 854 1131
rect 854 1097 863 1131
rect 811 1096 863 1097
rect 811 1059 863 1084
rect 811 1032 820 1059
rect 820 1032 854 1059
rect 854 1032 863 1059
rect 811 987 863 1020
rect 811 968 820 987
rect 820 968 854 987
rect 854 968 863 987
rect 811 953 820 956
rect 820 953 854 956
rect 854 953 863 956
rect 811 915 863 953
rect 811 904 820 915
rect 820 904 854 915
rect 854 904 863 915
rect 811 881 820 892
rect 820 881 854 892
rect 854 881 863 892
rect 811 843 863 881
rect 811 840 820 843
rect 820 840 854 843
rect 854 840 863 843
rect 811 809 820 828
rect 820 809 854 828
rect 854 809 863 828
rect 811 776 863 809
rect 811 737 820 764
rect 820 737 854 764
rect 854 737 863 764
rect 811 712 863 737
rect 811 699 863 700
rect 811 665 820 699
rect 820 665 854 699
rect 854 665 863 699
rect 811 648 863 665
rect 811 627 863 636
rect 811 593 820 627
rect 820 593 854 627
rect 854 593 863 627
rect 811 584 863 593
rect 967 1563 1019 1588
rect 967 1536 976 1563
rect 976 1536 1010 1563
rect 1010 1536 1019 1563
rect 967 1491 1019 1524
rect 967 1472 976 1491
rect 976 1472 1010 1491
rect 1010 1472 1019 1491
rect 967 1457 976 1460
rect 976 1457 1010 1460
rect 1010 1457 1019 1460
rect 967 1419 1019 1457
rect 967 1408 976 1419
rect 976 1408 1010 1419
rect 1010 1408 1019 1419
rect 967 1385 976 1396
rect 976 1385 1010 1396
rect 1010 1385 1019 1396
rect 967 1347 1019 1385
rect 967 1344 976 1347
rect 976 1344 1010 1347
rect 1010 1344 1019 1347
rect 967 1313 976 1332
rect 976 1313 1010 1332
rect 1010 1313 1019 1332
rect 967 1280 1019 1313
rect 967 483 1019 516
rect 967 464 976 483
rect 976 464 1010 483
rect 1010 464 1019 483
rect 967 449 976 452
rect 976 449 1010 452
rect 1010 449 1019 452
rect 967 411 1019 449
rect 967 400 976 411
rect 976 400 1010 411
rect 1010 400 1019 411
rect 967 377 976 388
rect 976 377 1010 388
rect 1010 377 1019 388
rect 967 339 1019 377
rect 967 336 976 339
rect 976 336 1010 339
rect 1010 336 1019 339
rect 967 305 976 324
rect 976 305 1010 324
rect 1010 305 1019 324
rect 967 272 1019 305
rect 967 233 976 260
rect 976 233 1010 260
rect 1010 233 1019 260
rect 967 208 1019 233
<< metal2 >>
rect 14 1588 1348 1594
rect 14 1536 343 1588
rect 395 1536 655 1588
rect 707 1536 967 1588
rect 1019 1536 1348 1588
rect 14 1524 1348 1536
rect 14 1472 343 1524
rect 395 1472 655 1524
rect 707 1472 967 1524
rect 1019 1472 1348 1524
rect 14 1460 1348 1472
rect 14 1408 343 1460
rect 395 1408 655 1460
rect 707 1408 967 1460
rect 1019 1408 1348 1460
rect 14 1396 1348 1408
rect 14 1344 343 1396
rect 395 1344 655 1396
rect 707 1344 967 1396
rect 1019 1344 1348 1396
rect 14 1332 1348 1344
rect 14 1280 343 1332
rect 395 1280 655 1332
rect 707 1280 967 1332
rect 1019 1280 1348 1332
rect 14 1274 1348 1280
rect 14 1212 1348 1218
rect 14 1160 499 1212
rect 551 1160 811 1212
rect 863 1160 1348 1212
rect 14 1148 1348 1160
rect 14 1096 499 1148
rect 551 1096 811 1148
rect 863 1096 1348 1148
rect 14 1084 1348 1096
rect 14 1032 499 1084
rect 551 1032 811 1084
rect 863 1032 1348 1084
rect 14 1020 1348 1032
rect 14 968 499 1020
rect 551 968 811 1020
rect 863 968 1348 1020
rect 14 956 1348 968
rect 14 904 499 956
rect 551 904 811 956
rect 863 904 1348 956
rect 14 892 1348 904
rect 14 840 499 892
rect 551 840 811 892
rect 863 840 1348 892
rect 14 828 1348 840
rect 14 776 499 828
rect 551 776 811 828
rect 863 776 1348 828
rect 14 764 1348 776
rect 14 712 499 764
rect 551 712 811 764
rect 863 712 1348 764
rect 14 700 1348 712
rect 14 648 499 700
rect 551 648 811 700
rect 863 648 1348 700
rect 14 636 1348 648
rect 14 584 499 636
rect 551 584 811 636
rect 863 584 1348 636
rect 14 578 1348 584
rect 14 516 1348 522
rect 14 464 343 516
rect 395 464 655 516
rect 707 464 967 516
rect 1019 464 1348 516
rect 14 452 1348 464
rect 14 400 343 452
rect 395 400 655 452
rect 707 400 967 452
rect 1019 400 1348 452
rect 14 388 1348 400
rect 14 336 343 388
rect 395 336 655 388
rect 707 336 967 388
rect 1019 336 1348 388
rect 14 324 1348 336
rect 14 272 343 324
rect 395 272 655 324
rect 707 272 967 324
rect 1019 272 1348 324
rect 14 260 1348 272
rect 14 208 343 260
rect 395 208 655 260
rect 707 208 967 260
rect 1019 208 1348 260
rect 14 202 1348 208
<< labels >>
flabel metal2 s 216 250 258 446 0 FreeSans 200 90 0 0 SOURCE
port 3 nsew
flabel metal2 s 219 1356 255 1517 0 FreeSans 200 90 0 0 SOURCE
port 3 nsew
flabel metal2 s 276 780 317 1016 0 FreeSans 200 90 0 0 DRAIN
port 1 nsew
flabel metal1 s 628 1669 729 1709 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel metal1 s 628 17 729 57 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel comment s 837 898 837 898 0 FreeSans 300 0 0 0 S
flabel comment s 993 898 993 898 0 FreeSans 300 0 0 0 S
flabel comment s 837 898 837 898 0 FreeSans 300 0 0 0 D
flabel comment s 681 898 681 898 0 FreeSans 300 0 0 0 S
flabel comment s 681 898 681 898 0 FreeSans 300 0 0 0 S
flabel comment s 525 898 525 898 0 FreeSans 300 0 0 0 S
flabel comment s 525 898 525 898 0 FreeSans 300 0 0 0 D
flabel comment s 369 898 369 898 0 FreeSans 300 0 0 0 S
flabel comment s 369 898 369 898 0 FreeSans 300 0 0 0 S
flabel comment s 1062 932 1062 932 0 FreeSans 400 90 0 0 dummy_poly
flabel comment s 286 919 286 919 0 FreeSans 400 90 0 0 dummy_poly
flabel metal1 s 41 1231 100 1261 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 1262 1221 1321 1251 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
<< properties >>
string GDS_END 8554414
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8516230
string device primitive
<< end >>
