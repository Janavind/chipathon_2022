magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -1543 3178 -413 3394
rect -1543 3062 -1049 3178
<< pwell >>
rect 577 923 991 1175
rect 293 97 1611 749
rect 1164 70 1611 97
rect 1164 -16 1692 70
<< mvnmos >>
rect 656 949 756 1149
rect 812 949 912 1149
rect 372 123 472 723
rect 528 123 628 723
rect 684 123 784 723
rect 840 123 940 723
rect 996 123 1096 723
rect 1152 123 1252 723
rect 1432 123 1532 723
<< mvpmos >>
rect -1424 3128 -1324 3328
rect -1268 3128 -1168 3328
rect -988 3244 -788 3328
rect -732 3244 -532 3328
<< mvndiff >>
rect 603 1131 656 1149
rect 603 1097 611 1131
rect 645 1097 656 1131
rect 603 1063 656 1097
rect 603 1029 611 1063
rect 645 1029 656 1063
rect 603 995 656 1029
rect 603 961 611 995
rect 645 961 656 995
rect 603 949 656 961
rect 756 1131 812 1149
rect 756 1097 767 1131
rect 801 1097 812 1131
rect 756 1063 812 1097
rect 756 1029 767 1063
rect 801 1029 812 1063
rect 756 995 812 1029
rect 756 961 767 995
rect 801 961 812 995
rect 756 949 812 961
rect 912 1131 965 1149
rect 912 1097 923 1131
rect 957 1097 965 1131
rect 912 1063 965 1097
rect 912 1029 923 1063
rect 957 1029 965 1063
rect 912 995 965 1029
rect 912 961 923 995
rect 957 961 965 995
rect 912 949 965 961
rect 319 645 372 723
rect 319 611 327 645
rect 361 611 372 645
rect 319 577 372 611
rect 319 543 327 577
rect 361 543 372 577
rect 319 509 372 543
rect 319 475 327 509
rect 361 475 372 509
rect 319 441 372 475
rect 319 407 327 441
rect 361 407 372 441
rect 319 373 372 407
rect 319 339 327 373
rect 361 339 372 373
rect 319 305 372 339
rect 319 271 327 305
rect 361 271 372 305
rect 319 237 372 271
rect 319 203 327 237
rect 361 203 372 237
rect 319 169 372 203
rect 319 135 327 169
rect 361 135 372 169
rect 319 123 372 135
rect 472 645 528 723
rect 472 611 483 645
rect 517 611 528 645
rect 472 577 528 611
rect 472 543 483 577
rect 517 543 528 577
rect 472 509 528 543
rect 472 475 483 509
rect 517 475 528 509
rect 472 441 528 475
rect 472 407 483 441
rect 517 407 528 441
rect 472 373 528 407
rect 472 339 483 373
rect 517 339 528 373
rect 472 305 528 339
rect 472 271 483 305
rect 517 271 528 305
rect 472 237 528 271
rect 472 203 483 237
rect 517 203 528 237
rect 472 169 528 203
rect 472 135 483 169
rect 517 135 528 169
rect 472 123 528 135
rect 628 645 684 723
rect 628 611 639 645
rect 673 611 684 645
rect 628 577 684 611
rect 628 543 639 577
rect 673 543 684 577
rect 628 509 684 543
rect 628 475 639 509
rect 673 475 684 509
rect 628 441 684 475
rect 628 407 639 441
rect 673 407 684 441
rect 628 373 684 407
rect 628 339 639 373
rect 673 339 684 373
rect 628 305 684 339
rect 628 271 639 305
rect 673 271 684 305
rect 628 237 684 271
rect 628 203 639 237
rect 673 203 684 237
rect 628 169 684 203
rect 628 135 639 169
rect 673 135 684 169
rect 628 123 684 135
rect 784 645 840 723
rect 784 611 795 645
rect 829 611 840 645
rect 784 577 840 611
rect 784 543 795 577
rect 829 543 840 577
rect 784 509 840 543
rect 784 475 795 509
rect 829 475 840 509
rect 784 441 840 475
rect 784 407 795 441
rect 829 407 840 441
rect 784 373 840 407
rect 784 339 795 373
rect 829 339 840 373
rect 784 305 840 339
rect 784 271 795 305
rect 829 271 840 305
rect 784 237 840 271
rect 784 203 795 237
rect 829 203 840 237
rect 784 169 840 203
rect 784 135 795 169
rect 829 135 840 169
rect 784 123 840 135
rect 940 645 996 723
rect 940 611 951 645
rect 985 611 996 645
rect 940 577 996 611
rect 940 543 951 577
rect 985 543 996 577
rect 940 509 996 543
rect 940 475 951 509
rect 985 475 996 509
rect 940 441 996 475
rect 940 407 951 441
rect 985 407 996 441
rect 940 373 996 407
rect 940 339 951 373
rect 985 339 996 373
rect 940 305 996 339
rect 940 271 951 305
rect 985 271 996 305
rect 940 237 996 271
rect 940 203 951 237
rect 985 203 996 237
rect 940 169 996 203
rect 940 135 951 169
rect 985 135 996 169
rect 940 123 996 135
rect 1096 645 1152 723
rect 1096 611 1107 645
rect 1141 611 1152 645
rect 1096 577 1152 611
rect 1096 543 1107 577
rect 1141 543 1152 577
rect 1096 509 1152 543
rect 1096 475 1107 509
rect 1141 475 1152 509
rect 1096 441 1152 475
rect 1096 407 1107 441
rect 1141 407 1152 441
rect 1096 373 1152 407
rect 1096 339 1107 373
rect 1141 339 1152 373
rect 1096 305 1152 339
rect 1096 271 1107 305
rect 1141 271 1152 305
rect 1096 237 1152 271
rect 1096 203 1107 237
rect 1141 203 1152 237
rect 1096 169 1152 203
rect 1096 135 1107 169
rect 1141 135 1152 169
rect 1096 123 1152 135
rect 1252 645 1305 723
rect 1252 611 1263 645
rect 1297 611 1305 645
rect 1252 577 1305 611
rect 1252 543 1263 577
rect 1297 543 1305 577
rect 1252 509 1305 543
rect 1252 475 1263 509
rect 1297 475 1305 509
rect 1252 441 1305 475
rect 1252 407 1263 441
rect 1297 407 1305 441
rect 1252 373 1305 407
rect 1252 339 1263 373
rect 1297 339 1305 373
rect 1252 305 1305 339
rect 1252 271 1263 305
rect 1297 271 1305 305
rect 1252 237 1305 271
rect 1252 203 1263 237
rect 1297 203 1305 237
rect 1252 169 1305 203
rect 1252 135 1263 169
rect 1297 135 1305 169
rect 1252 123 1305 135
rect 1379 645 1432 723
rect 1379 611 1387 645
rect 1421 611 1432 645
rect 1379 577 1432 611
rect 1379 543 1387 577
rect 1421 543 1432 577
rect 1379 509 1432 543
rect 1379 475 1387 509
rect 1421 475 1432 509
rect 1379 441 1432 475
rect 1379 407 1387 441
rect 1421 407 1432 441
rect 1379 373 1432 407
rect 1379 339 1387 373
rect 1421 339 1432 373
rect 1379 305 1432 339
rect 1379 271 1387 305
rect 1421 271 1432 305
rect 1379 237 1432 271
rect 1379 203 1387 237
rect 1421 203 1432 237
rect 1379 169 1432 203
rect 1379 135 1387 169
rect 1421 135 1432 169
rect 1379 123 1432 135
rect 1532 645 1585 723
rect 1532 611 1543 645
rect 1577 611 1585 645
rect 1532 577 1585 611
rect 1532 543 1543 577
rect 1577 543 1585 577
rect 1532 509 1585 543
rect 1532 475 1543 509
rect 1577 475 1585 509
rect 1532 441 1585 475
rect 1532 407 1543 441
rect 1577 407 1585 441
rect 1532 373 1585 407
rect 1532 339 1543 373
rect 1577 339 1585 373
rect 1532 305 1585 339
rect 1532 271 1543 305
rect 1577 271 1585 305
rect 1532 237 1585 271
rect 1532 203 1543 237
rect 1577 203 1585 237
rect 1532 169 1585 203
rect 1532 135 1543 169
rect 1577 135 1585 169
rect 1532 123 1585 135
<< mvpdiff >>
rect -1477 3310 -1424 3328
rect -1477 3276 -1469 3310
rect -1435 3276 -1424 3310
rect -1477 3242 -1424 3276
rect -1477 3208 -1469 3242
rect -1435 3208 -1424 3242
rect -1477 3174 -1424 3208
rect -1477 3140 -1469 3174
rect -1435 3140 -1424 3174
rect -1477 3128 -1424 3140
rect -1324 3310 -1268 3328
rect -1324 3276 -1313 3310
rect -1279 3276 -1268 3310
rect -1324 3242 -1268 3276
rect -1324 3208 -1313 3242
rect -1279 3208 -1268 3242
rect -1324 3174 -1268 3208
rect -1324 3140 -1313 3174
rect -1279 3140 -1268 3174
rect -1324 3128 -1268 3140
rect -1168 3310 -1115 3328
rect -1168 3276 -1157 3310
rect -1123 3276 -1115 3310
rect -1168 3242 -1115 3276
rect -1041 3316 -988 3328
rect -1041 3282 -1033 3316
rect -999 3282 -988 3316
rect -1041 3244 -988 3282
rect -788 3316 -732 3328
rect -788 3282 -777 3316
rect -743 3282 -732 3316
rect -788 3244 -732 3282
rect -532 3316 -479 3328
rect -532 3282 -521 3316
rect -487 3282 -479 3316
rect -532 3244 -479 3282
rect -1168 3208 -1157 3242
rect -1123 3208 -1115 3242
rect -1168 3174 -1115 3208
rect -1168 3140 -1157 3174
rect -1123 3140 -1115 3174
rect -1168 3128 -1115 3140
<< mvndiffc >>
rect 611 1097 645 1131
rect 611 1029 645 1063
rect 611 961 645 995
rect 767 1097 801 1131
rect 767 1029 801 1063
rect 767 961 801 995
rect 923 1097 957 1131
rect 923 1029 957 1063
rect 923 961 957 995
rect 327 611 361 645
rect 327 543 361 577
rect 327 475 361 509
rect 327 407 361 441
rect 327 339 361 373
rect 327 271 361 305
rect 327 203 361 237
rect 327 135 361 169
rect 483 611 517 645
rect 483 543 517 577
rect 483 475 517 509
rect 483 407 517 441
rect 483 339 517 373
rect 483 271 517 305
rect 483 203 517 237
rect 483 135 517 169
rect 639 611 673 645
rect 639 543 673 577
rect 639 475 673 509
rect 639 407 673 441
rect 639 339 673 373
rect 639 271 673 305
rect 639 203 673 237
rect 639 135 673 169
rect 795 611 829 645
rect 795 543 829 577
rect 795 475 829 509
rect 795 407 829 441
rect 795 339 829 373
rect 795 271 829 305
rect 795 203 829 237
rect 795 135 829 169
rect 951 611 985 645
rect 951 543 985 577
rect 951 475 985 509
rect 951 407 985 441
rect 951 339 985 373
rect 951 271 985 305
rect 951 203 985 237
rect 951 135 985 169
rect 1107 611 1141 645
rect 1107 543 1141 577
rect 1107 475 1141 509
rect 1107 407 1141 441
rect 1107 339 1141 373
rect 1107 271 1141 305
rect 1107 203 1141 237
rect 1107 135 1141 169
rect 1263 611 1297 645
rect 1263 543 1297 577
rect 1263 475 1297 509
rect 1263 407 1297 441
rect 1263 339 1297 373
rect 1263 271 1297 305
rect 1263 203 1297 237
rect 1263 135 1297 169
rect 1387 611 1421 645
rect 1387 543 1421 577
rect 1387 475 1421 509
rect 1387 407 1421 441
rect 1387 339 1421 373
rect 1387 271 1421 305
rect 1387 203 1421 237
rect 1387 135 1421 169
rect 1543 611 1577 645
rect 1543 543 1577 577
rect 1543 475 1577 509
rect 1543 407 1577 441
rect 1543 339 1577 373
rect 1543 271 1577 305
rect 1543 203 1577 237
rect 1543 135 1577 169
<< mvpdiffc >>
rect -1469 3276 -1435 3310
rect -1469 3208 -1435 3242
rect -1469 3140 -1435 3174
rect -1313 3276 -1279 3310
rect -1313 3208 -1279 3242
rect -1313 3140 -1279 3174
rect -1157 3276 -1123 3310
rect -1033 3282 -999 3316
rect -777 3282 -743 3316
rect -521 3282 -487 3316
rect -1157 3208 -1123 3242
rect -1157 3140 -1123 3174
<< psubdiff >>
rect 1190 10 1224 44
rect 1258 10 1318 44
rect 1352 10 1412 44
rect 1446 10 1505 44
rect 1539 10 1598 44
rect 1632 10 1666 44
<< psubdiffcont >>
rect 1224 10 1258 44
rect 1318 10 1352 44
rect 1412 10 1446 44
rect 1505 10 1539 44
rect 1598 10 1632 44
<< poly >>
rect -1424 3328 -1324 3360
rect -1268 3328 -1168 3360
rect -988 3328 -788 3360
rect -732 3328 -532 3360
rect -988 3196 -788 3244
rect -988 3162 -972 3196
rect -938 3162 -838 3196
rect -804 3162 -788 3196
rect -988 3146 -788 3162
rect -732 3196 -532 3244
rect -732 3162 -716 3196
rect -682 3162 -582 3196
rect -548 3162 -532 3196
rect -732 3146 -532 3162
rect -1424 3096 -1324 3128
rect -1268 3096 -1168 3128
rect -1424 3080 -1168 3096
rect -1424 3046 -1408 3080
rect -1374 3046 -1313 3080
rect -1279 3046 -1218 3080
rect -1184 3046 -1168 3080
rect -1424 3030 -1168 3046
rect 656 1149 756 1175
rect 812 1149 912 1175
rect 656 923 756 949
rect 622 907 756 923
rect 622 873 638 907
rect 672 873 706 907
rect 740 873 756 907
rect 622 857 756 873
rect 812 923 912 949
rect 812 907 946 923
rect 812 873 828 907
rect 862 873 896 907
rect 930 873 946 907
rect 812 857 946 873
rect 372 799 784 815
rect 372 765 388 799
rect 422 765 458 799
rect 492 765 527 799
rect 561 765 596 799
rect 630 765 665 799
rect 699 765 734 799
rect 768 765 784 799
rect 372 749 784 765
rect 372 723 472 749
rect 528 723 628 749
rect 684 723 784 749
rect 840 799 1252 815
rect 840 765 856 799
rect 890 765 925 799
rect 959 765 994 799
rect 1028 765 1063 799
rect 1097 765 1132 799
rect 1166 765 1202 799
rect 1236 765 1252 799
rect 840 749 1252 765
rect 1410 799 1544 815
rect 1410 765 1426 799
rect 1460 765 1494 799
rect 1528 765 1544 799
rect 1410 749 1544 765
rect 840 723 940 749
rect 996 723 1096 749
rect 1152 723 1252 749
rect 1432 723 1532 749
rect 372 97 472 123
rect 528 97 628 123
rect 684 97 784 123
rect 840 97 940 123
rect 996 97 1096 123
rect 1152 97 1252 123
rect 1432 97 1532 123
<< polycont >>
rect -972 3162 -938 3196
rect -838 3162 -804 3196
rect -716 3162 -682 3196
rect -582 3162 -548 3196
rect -1408 3046 -1374 3080
rect -1313 3046 -1279 3080
rect -1218 3046 -1184 3080
rect 638 873 672 907
rect 706 873 740 907
rect 828 873 862 907
rect 896 873 930 907
rect 388 765 422 799
rect 458 765 492 799
rect 527 765 561 799
rect 596 765 630 799
rect 665 765 699 799
rect 734 765 768 799
rect 856 765 890 799
rect 925 765 959 799
rect 994 765 1028 799
rect 1063 765 1097 799
rect 1132 765 1166 799
rect 1202 765 1236 799
rect 1426 765 1460 799
rect 1494 765 1528 799
<< locali >>
rect -1469 3310 -1435 3330
rect -1469 3242 -1435 3258
rect -1469 3174 -1435 3208
rect -1313 3310 -1279 3326
rect -1313 3242 -1279 3276
rect -1313 3174 -1279 3208
rect -1469 3124 -1435 3140
rect -1314 3140 -1313 3160
rect -1157 3310 -1123 3330
rect -1157 3242 -1123 3258
rect -1157 3174 -1123 3208
rect -1279 3140 -1276 3160
rect -1314 3126 -1276 3140
rect -1313 3124 -1279 3126
rect -1157 3124 -1123 3140
rect -1089 3316 -999 3332
rect -1089 3282 -1033 3316
rect -1089 3266 -999 3282
rect -777 3316 -743 3330
rect -1089 3115 -1022 3266
rect -521 3316 -388 3332
rect -487 3282 -388 3316
rect -521 3266 -388 3282
rect -498 3196 -388 3266
rect -988 3162 -972 3196
rect -938 3162 -923 3196
rect -889 3162 -851 3196
rect -804 3162 -788 3196
rect -732 3162 -716 3196
rect -682 3162 -582 3196
rect -548 3162 -532 3196
rect -460 3162 -422 3196
rect -732 3122 -532 3162
rect -732 3115 -653 3122
rect -1089 3088 -653 3115
rect -619 3088 -581 3122
rect -547 3088 -532 3122
rect -1089 3080 -532 3088
rect -1425 3046 -1408 3080
rect -1374 3046 -1313 3080
rect -1279 3046 -1218 3080
rect -1184 3046 -532 3080
rect -1425 2982 -532 3046
rect 611 1131 645 1147
rect 611 1087 645 1097
rect 767 1131 801 1147
rect 767 1069 801 1097
rect 923 1131 957 1147
rect 923 1078 957 1097
rect 764 1063 802 1069
rect 764 1035 767 1063
rect 611 1015 645 1029
rect 611 945 645 961
rect 801 1035 802 1063
rect 923 1063 924 1078
rect 767 995 801 1029
rect 767 945 801 961
rect 957 1029 958 1044
rect 923 1006 958 1029
rect 923 995 924 1006
rect 923 945 957 961
rect 622 901 638 907
rect 672 901 706 907
rect 622 873 633 901
rect 672 873 705 901
rect 740 873 756 907
rect 812 901 828 907
rect 812 873 826 901
rect 862 873 896 907
rect 930 901 946 907
rect 932 873 946 901
rect 667 867 705 873
rect 860 867 898 873
rect 372 765 388 799
rect 422 765 458 799
rect 492 765 510 799
rect 561 765 582 799
rect 630 765 665 799
rect 699 765 734 799
rect 768 765 784 799
rect 840 765 856 799
rect 897 765 925 799
rect 969 765 994 799
rect 1028 765 1063 799
rect 1097 765 1132 799
rect 1166 765 1202 799
rect 1236 765 1252 799
rect 1410 765 1424 799
rect 1460 765 1494 799
rect 1530 765 1544 799
rect 327 645 361 661
rect 327 593 361 611
rect 483 645 517 661
rect 325 577 363 593
rect 325 559 327 577
rect 361 559 363 577
rect 483 577 517 611
rect 639 645 673 661
rect 639 593 673 611
rect 795 645 829 661
rect 327 509 361 543
rect 635 577 673 593
rect 635 559 639 577
rect 483 519 517 543
rect 795 577 829 611
rect 951 645 985 661
rect 951 593 985 611
rect 1107 645 1141 661
rect 484 509 522 519
rect 517 485 522 509
rect 639 509 673 543
rect 949 577 987 593
rect 949 559 951 577
rect 795 519 829 543
rect 985 559 987 577
rect 1107 577 1141 611
rect 1263 645 1297 661
rect 1263 593 1297 611
rect 1387 645 1421 661
rect 327 441 361 475
rect 327 373 361 407
rect 327 305 361 339
rect 327 237 361 271
rect 327 169 361 203
rect 327 119 361 135
rect 483 441 517 475
rect 483 373 517 407
rect 483 305 517 339
rect 483 237 517 271
rect 483 169 517 203
rect 483 119 517 135
rect 794 509 832 519
rect 794 485 795 509
rect 639 441 673 475
rect 639 373 673 407
rect 639 305 673 339
rect 639 237 673 271
rect 639 169 673 203
rect 639 119 673 135
rect 829 485 832 509
rect 951 509 985 543
rect 1260 577 1298 593
rect 1260 559 1263 577
rect 1107 519 1141 543
rect 1297 559 1298 577
rect 1387 577 1421 611
rect 795 441 829 475
rect 795 373 829 407
rect 795 305 829 339
rect 795 237 829 271
rect 795 169 829 203
rect 795 119 829 135
rect 1075 509 1113 519
rect 1075 485 1107 509
rect 1263 509 1297 543
rect 1387 519 1421 543
rect 1543 645 1577 661
rect 1543 577 1577 611
rect 951 441 985 475
rect 951 373 985 407
rect 951 305 985 339
rect 951 237 985 271
rect 951 169 985 203
rect 951 119 985 135
rect 1107 441 1141 475
rect 1107 373 1141 407
rect 1107 305 1141 339
rect 1107 237 1141 271
rect 1107 169 1141 203
rect 1107 119 1141 135
rect 1385 509 1423 519
rect 1385 485 1387 509
rect 1263 441 1297 475
rect 1263 373 1297 407
rect 1263 305 1297 339
rect 1263 237 1297 271
rect 1263 169 1297 203
rect 1263 119 1297 135
rect 1421 485 1423 509
rect 1543 509 1577 543
rect 1387 441 1421 475
rect 1387 373 1421 407
rect 1387 305 1421 339
rect 1387 237 1421 271
rect 1387 169 1421 203
rect 1387 119 1421 135
rect 1543 441 1577 475
rect 1543 373 1577 407
rect 1543 305 1577 339
rect 1543 237 1577 271
rect 1543 189 1577 203
rect 1543 117 1577 135
rect 1190 10 1198 44
rect 1258 10 1276 44
rect 1310 10 1318 44
rect 1352 10 1353 44
rect 1387 10 1412 44
rect 1464 10 1505 44
rect 1541 10 1584 44
rect 1632 10 1666 44
<< viali >>
rect -1469 3330 -1435 3364
rect -1157 3330 -1123 3364
rect -1469 3276 -1435 3292
rect -1469 3258 -1435 3276
rect -1348 3126 -1314 3160
rect -1157 3276 -1123 3292
rect -1157 3258 -1123 3276
rect -1276 3126 -1242 3160
rect -777 3330 -743 3364
rect -777 3282 -743 3292
rect -777 3258 -743 3282
rect -923 3162 -889 3196
rect -851 3162 -838 3196
rect -838 3162 -817 3196
rect -494 3162 -460 3196
rect -422 3162 -388 3196
rect -653 3088 -619 3122
rect -581 3088 -547 3122
rect 611 1063 645 1087
rect 611 1053 645 1063
rect 730 1035 764 1069
rect 611 995 645 1015
rect 611 981 645 995
rect 802 1035 836 1069
rect 924 1063 958 1078
rect 924 1044 957 1063
rect 957 1044 958 1063
rect 924 995 958 1006
rect 924 972 957 995
rect 957 972 958 995
rect 633 873 638 901
rect 638 873 667 901
rect 705 873 706 901
rect 706 873 739 901
rect 826 873 828 901
rect 828 873 860 901
rect 898 873 930 901
rect 930 873 932 901
rect 633 867 667 873
rect 705 867 739 873
rect 826 867 860 873
rect 898 867 932 873
rect 510 765 527 799
rect 527 765 544 799
rect 582 765 596 799
rect 596 765 616 799
rect 863 765 890 799
rect 890 765 897 799
rect 935 765 959 799
rect 959 765 969 799
rect 1424 765 1426 799
rect 1426 765 1458 799
rect 1496 765 1528 799
rect 1528 765 1530 799
rect 291 559 325 593
rect 363 559 397 593
rect 601 559 635 593
rect 673 559 707 593
rect 450 509 484 519
rect 450 485 483 509
rect 483 485 484 509
rect 522 485 556 519
rect 915 559 949 593
rect 987 559 1021 593
rect 760 485 794 519
rect 832 485 866 519
rect 1226 559 1260 593
rect 1298 559 1332 593
rect 1041 485 1075 519
rect 1113 509 1147 519
rect 1113 485 1141 509
rect 1141 485 1147 509
rect 1351 485 1385 519
rect 1423 485 1457 519
rect 1543 169 1577 189
rect 1543 155 1577 169
rect 1543 83 1577 117
rect 1198 10 1224 44
rect 1224 10 1232 44
rect 1276 10 1310 44
rect 1353 10 1387 44
rect 1430 10 1446 44
rect 1446 10 1464 44
rect 1507 10 1539 44
rect 1539 10 1541 44
rect 1584 10 1598 44
rect 1598 10 1618 44
<< metal1 >>
rect -1475 3364 -737 3442
rect -1475 3330 -1469 3364
rect -1435 3330 -1157 3364
rect -1123 3330 -777 3364
rect -743 3330 -737 3364
rect -1475 3292 -737 3330
rect -1475 3258 -1469 3292
rect -1435 3258 -1157 3292
rect -1123 3258 -777 3292
rect -743 3258 -737 3292
rect -1475 3246 -737 3258
rect -935 3196 -203 3202
rect -1360 3160 -1230 3166
rect -1360 3126 -1348 3160
rect -1314 3126 -1276 3160
rect -1242 3126 -1230 3160
rect -935 3162 -923 3196
rect -889 3162 -851 3196
rect -817 3162 -494 3196
rect -460 3162 -422 3196
rect -388 3162 -203 3196
rect -935 3156 -203 3162
tri -289 3128 -261 3156 ne
rect -261 3128 -203 3156
rect -1360 3088 -1230 3126
rect -665 3122 -303 3128
tri -303 3122 -297 3128 sw
tri -261 3122 -255 3128 ne
tri -1230 3088 -1198 3120 sw
rect -665 3088 -653 3122
rect -619 3088 -581 3122
rect -547 3108 -297 3122
tri -297 3108 -283 3122 sw
rect -547 3094 -283 3108
rect -547 3088 -535 3094
rect -1360 3082 -1198 3088
tri -1198 3082 -1192 3088 sw
rect -665 3082 -535 3088
tri -535 3082 -523 3094 nw
tri -365 3082 -353 3094 ne
rect -353 3082 -283 3094
rect -1360 3064 -1192 3082
tri -1192 3064 -1174 3082 sw
tri -353 3064 -335 3082 ne
rect -1360 3050 -1174 3064
tri -1174 3050 -1160 3064 sw
rect -1360 3044 -363 3050
rect -1360 3016 -415 3044
rect -415 2980 -363 2992
rect -415 2922 -363 2928
rect -335 3044 -283 3082
rect -335 2980 -283 2992
rect -335 2922 -283 2928
rect -255 3044 -203 3128
rect -255 2980 -203 2992
rect -255 2922 -203 2928
rect -335 1249 -283 1255
rect -335 1185 -283 1197
rect -415 1173 -363 1179
tri -283 1161 -249 1195 sw
rect -237 1189 -231 1241
rect -179 1189 -167 1241
rect -115 1235 -109 1241
tri -109 1235 -103 1241 sw
rect -115 1189 1057 1235
rect -283 1138 941 1161
tri 941 1138 964 1161 sw
rect -283 1133 964 1138
rect -335 1127 964 1133
rect -415 1109 -363 1121
tri -363 1099 -347 1115 sw
rect -363 1087 -347 1099
tri -347 1087 -335 1099 sw
tri 587 1087 599 1099 se
rect -363 1085 -335 1087
tri -335 1085 -333 1087 sw
tri 585 1085 587 1087 se
rect 587 1085 599 1087
rect 605 1087 651 1099
rect 605 1085 611 1087
rect -363 1057 611 1085
rect -415 1053 611 1057
rect 645 1053 651 1087
rect 918 1078 964 1127
rect -415 1051 651 1053
tri 565 1035 581 1051 ne
rect 581 1035 599 1051
tri 581 1017 599 1035 ne
rect 605 1015 651 1051
rect 718 1069 848 1078
rect 718 1035 730 1069
rect 764 1035 802 1069
rect 836 1035 848 1069
rect 718 1026 848 1035
rect 918 1044 924 1078
rect 958 1044 964 1078
tri 917 1026 918 1027 se
rect 918 1026 964 1044
rect 605 981 611 1015
rect 645 981 651 1015
tri 897 1006 917 1026 se
rect 917 1006 964 1026
tri 885 994 897 1006 se
rect 897 994 924 1006
rect 605 971 651 981
rect 599 969 651 971
rect 697 972 924 994
rect 958 972 964 1006
rect 697 960 964 972
tri 663 907 697 941 se
rect 697 907 751 960
tri 751 922 789 960 nw
rect 621 901 751 907
rect 621 867 633 901
rect 667 867 705 901
rect 739 867 751 901
rect 621 861 751 867
tri 671 829 703 861 ne
rect 703 829 751 861
rect 814 901 959 907
rect 814 867 826 901
rect 860 867 898 901
rect 932 867 959 901
rect 814 854 959 867
tri 597 827 599 829 se
tri 703 827 705 829 ne
tri 575 805 597 827 se
rect 597 805 599 827
rect 498 799 628 805
rect 498 765 510 799
rect 544 765 582 799
rect 616 765 628 799
rect 498 759 628 765
tri 565 725 599 759 ne
tri 671 599 705 633 se
rect 705 599 751 829
rect 851 799 981 805
rect 851 765 863 799
rect 897 765 935 799
rect 969 765 981 799
rect 851 759 981 765
tri 851 725 885 759 nw
tri 977 599 1011 633 se
rect 1011 599 1057 1189
rect 1412 799 1542 805
rect 1412 765 1424 799
rect 1458 765 1496 799
rect 1530 765 1542 799
rect 1412 759 1542 765
tri 1057 599 1091 633 sw
rect 279 593 751 599
rect 279 559 291 593
rect 325 559 363 593
rect 397 559 601 593
rect 635 559 673 593
rect 707 559 751 593
rect 279 553 751 559
rect 903 593 1344 599
rect 903 559 915 593
rect 949 559 987 593
rect 1021 559 1226 593
rect 1260 559 1298 593
rect 1332 559 1344 593
rect 903 553 1344 559
rect 438 519 1469 525
rect 438 485 450 519
rect 484 485 522 519
rect 556 485 760 519
rect 794 485 832 519
rect 866 485 1041 519
rect 1075 485 1113 519
rect 1147 485 1351 519
rect 1385 485 1423 519
rect 1457 485 1469 519
rect 438 479 1469 485
rect 1362 189 1583 201
rect 1362 155 1543 189
rect 1577 155 1583 189
rect 1362 117 1583 155
rect 1362 83 1543 117
rect 1577 83 1583 117
rect 1362 50 1583 83
rect 1186 44 1630 50
rect 1186 10 1198 44
rect 1232 10 1276 44
rect 1310 10 1353 44
rect 1387 10 1430 44
rect 1464 10 1507 44
rect 1541 10 1584 44
rect 1618 10 1630 44
rect 1186 4 1630 10
<< via1 >>
rect -415 2992 -363 3044
rect -415 2928 -363 2980
rect -335 2992 -283 3044
rect -335 2928 -283 2980
rect -255 2992 -203 3044
rect -255 2928 -203 2980
rect -335 1197 -283 1249
rect -415 1121 -363 1173
rect -335 1133 -283 1185
rect -231 1189 -179 1241
rect -167 1189 -115 1241
rect -415 1057 -363 1109
<< metal2 >>
rect -415 3044 -363 3050
rect -415 2980 -363 2992
rect -415 1173 -363 2928
rect -335 3044 -283 3050
rect -335 2980 -283 2992
rect -335 1249 -283 2928
rect -335 1185 -283 1197
rect -255 3044 -203 3050
rect -255 2980 -203 2992
rect -255 1241 -203 2928
rect -255 1189 -231 1241
rect -179 1189 -167 1241
rect -115 1189 -109 1241
rect -335 1127 -283 1133
rect -415 1109 -363 1121
rect -415 1051 -363 1057
use sky130_fd_pr__nfet_01v8__example_55959141808568  sky130_fd_pr__nfet_01v8__example_55959141808568_0
timestamp 1666199351
transform -1 0 1532 0 1 123
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808569  sky130_fd_pr__nfet_01v8__example_55959141808569_0
timestamp 1666199351
transform -1 0 784 0 1 123
box -1 0 413 1
use sky130_fd_pr__nfet_01v8__example_55959141808569  sky130_fd_pr__nfet_01v8__example_55959141808569_1
timestamp 1666199351
transform 1 0 840 0 1 123
box -1 0 413 1
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_0
timestamp 1666199351
transform 1 0 812 0 1 949
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_1
timestamp 1666199351
transform -1 0 756 0 1 949
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_0
timestamp 1666199351
transform 1 0 -732 0 -1 3328
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_1
timestamp 1666199351
transform -1 0 -788 0 -1 3328
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808567  sky130_fd_pr__pfet_01v8__example_55959141808567_0
timestamp 1666199351
transform 1 0 -1424 0 1 3128
box -1 0 257 1
<< labels >>
flabel metal1 s -1310 3348 -1282 3376 3 FreeSans 520 0 0 0 VPWR_HV
port 1 nsew
flabel metal1 s 894 771 922 799 3 FreeSans 520 0 0 0 IN
port 2 nsew
flabel metal1 s 1452 126 1480 154 3 FreeSans 520 0 0 0 VGND
port 3 nsew
flabel metal1 s 848 866 876 894 3 FreeSans 520 0 0 0 RST_H
port 4 nsew
flabel metal1 s 1468 768 1496 796 3 FreeSans 520 0 0 0 HLD_H_N
port 5 nsew
flabel metal1 s 552 770 580 798 3 FreeSans 520 0 0 0 IN_B
port 6 nsew
flabel metal1 s 614 1026 642 1054 3 FreeSans 520 0 0 0 OUT_H_N
port 7 nsew
flabel metal1 s 765 1038 793 1066 3 FreeSans 520 0 0 0 VGND
port 3 nsew
<< properties >>
string GDS_END 43568498
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43552564
<< end >>
