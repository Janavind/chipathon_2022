magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect 12570 14777 14442 15721
rect 8293 8874 15173 8875
rect -32 6931 15173 8874
<< pwell >>
rect -973 8935 15143 9711
rect 18 6661 7134 6869
rect 12467 6661 15143 6869
rect 18 6025 15143 6661
rect 14891 5962 15143 6025
rect 14951 1314 15143 5962
rect 7018 1308 15143 1314
rect 42 1225 15143 1308
rect 6996 962 15143 1225
rect 6996 395 7780 962
rect 9661 702 15143 962
rect 9661 395 11682 702
rect 14439 395 15143 702
rect 6996 -7 15143 395
<< mvpsubdiff >>
rect -947 9680 15117 9685
rect -947 9647 -723 9680
rect -947 9613 -932 9647
rect -898 9613 -864 9647
rect -830 9613 -796 9647
rect -762 9646 -723 9647
rect -689 9646 -654 9680
rect -620 9646 -585 9680
rect -551 9646 -516 9680
rect -482 9646 -447 9680
rect -413 9646 -378 9680
rect -344 9646 -309 9680
rect -275 9646 -240 9680
rect -206 9646 -171 9680
rect -137 9646 -102 9680
rect -68 9646 -33 9680
rect -762 9613 -33 9646
rect -947 9612 -33 9613
rect -947 9578 -723 9612
rect -689 9578 -654 9612
rect -620 9578 -585 9612
rect -551 9578 -516 9612
rect -482 9578 -447 9612
rect -413 9578 -378 9612
rect -344 9578 -309 9612
rect -275 9578 -240 9612
rect -206 9578 -171 9612
rect -137 9578 -102 9612
rect -68 9578 -33 9612
rect -947 9571 -33 9578
rect -947 9537 -932 9571
rect -898 9537 -864 9571
rect -830 9537 -796 9571
rect -762 9544 -33 9571
rect -762 9537 -723 9544
rect -947 9510 -723 9537
rect -689 9510 -654 9544
rect -620 9510 -585 9544
rect -551 9510 -516 9544
rect -482 9510 -447 9544
rect -413 9510 -378 9544
rect -344 9510 -309 9544
rect -275 9510 -240 9544
rect -206 9510 -171 9544
rect -137 9510 -102 9544
rect -68 9510 -33 9544
rect -947 9495 -33 9510
rect -947 9461 -932 9495
rect -898 9461 -864 9495
rect -830 9461 -796 9495
rect -762 9476 -33 9495
rect -762 9461 -723 9476
rect -947 9442 -723 9461
rect -689 9442 -654 9476
rect -620 9442 -585 9476
rect -551 9442 -516 9476
rect -482 9442 -447 9476
rect -413 9442 -378 9476
rect -344 9442 -309 9476
rect -275 9442 -240 9476
rect -206 9442 -171 9476
rect -137 9442 -102 9476
rect -68 9442 -33 9476
rect -947 9418 -33 9442
rect -947 9384 -932 9418
rect -898 9384 -864 9418
rect -830 9384 -796 9418
rect -762 9408 -33 9418
rect -762 9384 -723 9408
rect -947 9374 -723 9384
rect -689 9374 -654 9408
rect -620 9374 -585 9408
rect -551 9374 -516 9408
rect -482 9374 -447 9408
rect -413 9374 -378 9408
rect -344 9374 -309 9408
rect -275 9374 -240 9408
rect -206 9374 -171 9408
rect -137 9374 -102 9408
rect -68 9374 -33 9408
rect -947 9341 -33 9374
rect -947 9307 -932 9341
rect -898 9307 -864 9341
rect -830 9307 -796 9341
rect -762 9340 -33 9341
rect -762 9307 -723 9340
rect -947 9306 -723 9307
rect -689 9306 -654 9340
rect -620 9306 -585 9340
rect -551 9306 -516 9340
rect -482 9306 -447 9340
rect -413 9306 -378 9340
rect -344 9306 -309 9340
rect -275 9306 -240 9340
rect -206 9306 -171 9340
rect -137 9306 -102 9340
rect -68 9306 -33 9340
rect -947 9272 -33 9306
rect -947 9264 -723 9272
rect -947 9230 -932 9264
rect -898 9230 -864 9264
rect -830 9230 -796 9264
rect -762 9238 -723 9264
rect -689 9238 -654 9272
rect -620 9238 -585 9272
rect -551 9238 -516 9272
rect -482 9238 -447 9272
rect -413 9238 -378 9272
rect -344 9238 -309 9272
rect -275 9238 -240 9272
rect -206 9238 -171 9272
rect -137 9238 -102 9272
rect -68 9238 -33 9272
rect -762 9230 -33 9238
rect -947 9204 -33 9230
rect -947 9187 -723 9204
rect -947 9153 -932 9187
rect -898 9153 -864 9187
rect -830 9153 -796 9187
rect -762 9170 -723 9187
rect -689 9170 -654 9204
rect -620 9170 -585 9204
rect -551 9170 -516 9204
rect -482 9170 -447 9204
rect -413 9170 -378 9204
rect -344 9170 -309 9204
rect -275 9170 -240 9204
rect -206 9170 -171 9204
rect -137 9170 -102 9204
rect -68 9170 -33 9204
rect -762 9153 -33 9170
rect -947 9136 -33 9153
rect -947 9110 -723 9136
rect -947 9076 -932 9110
rect -898 9076 -864 9110
rect -830 9076 -796 9110
rect -762 9102 -723 9110
rect -689 9102 -654 9136
rect -620 9102 -585 9136
rect -551 9102 -516 9136
rect -482 9102 -447 9136
rect -413 9102 -378 9136
rect -344 9102 -309 9136
rect -275 9102 -240 9136
rect -206 9102 -171 9136
rect -137 9102 -102 9136
rect -68 9102 -33 9136
rect -762 9076 -33 9102
rect -947 9068 -33 9076
rect -947 9034 -723 9068
rect -689 9034 -654 9068
rect -620 9034 -585 9068
rect -551 9034 -516 9068
rect -482 9034 -447 9068
rect -413 9034 -378 9068
rect -344 9034 -309 9068
rect -275 9034 -240 9068
rect -206 9034 -171 9068
rect -137 9034 -102 9068
rect -68 9034 -33 9068
rect -947 9033 -33 9034
rect -947 8999 -932 9033
rect -898 8999 -864 9033
rect -830 8999 -796 9033
rect -762 9000 -33 9033
rect -762 8999 -723 9000
rect -947 8966 -723 8999
rect -689 8966 -654 9000
rect -620 8966 -585 9000
rect -551 8966 -516 9000
rect -482 8966 -447 9000
rect -413 8966 -378 9000
rect -344 8966 -309 9000
rect -275 8966 -240 9000
rect -206 8966 -171 9000
rect -137 8966 -102 9000
rect -68 8966 -33 9000
rect 14893 9647 15117 9680
rect 14893 9613 14932 9647
rect 14966 9613 15000 9647
rect 15034 9613 15068 9647
rect 15102 9613 15117 9647
rect 14893 9571 15117 9613
rect 14893 9537 14932 9571
rect 14966 9537 15000 9571
rect 15034 9537 15068 9571
rect 15102 9537 15117 9571
rect 14893 9495 15117 9537
rect 14893 9461 14932 9495
rect 14966 9461 15000 9495
rect 15034 9461 15068 9495
rect 15102 9461 15117 9495
rect 14893 9418 15117 9461
rect 14893 9384 14932 9418
rect 14966 9384 15000 9418
rect 15034 9384 15068 9418
rect 15102 9384 15117 9418
rect 14893 9341 15117 9384
rect 14893 9307 14932 9341
rect 14966 9307 15000 9341
rect 15034 9307 15068 9341
rect 15102 9307 15117 9341
rect 14893 9264 15117 9307
rect 14893 9230 14932 9264
rect 14966 9230 15000 9264
rect 15034 9230 15068 9264
rect 15102 9230 15117 9264
rect 14893 9187 15117 9230
rect 14893 9153 14932 9187
rect 14966 9153 15000 9187
rect 15034 9153 15068 9187
rect 15102 9153 15117 9187
rect 14893 9110 15117 9153
rect 14893 9076 14932 9110
rect 14966 9076 15000 9110
rect 15034 9076 15068 9110
rect 15102 9076 15117 9110
rect 14893 9033 15117 9076
rect 14893 8999 14932 9033
rect 14966 8999 15000 9033
rect 15034 8999 15068 9033
rect 15102 8999 15117 9033
rect 14893 8966 15117 8999
rect -947 8961 15117 8966
rect 44 6809 68 6843
rect 102 6809 137 6843
rect 171 6809 206 6843
rect 240 6809 275 6843
rect 309 6809 344 6843
rect 378 6809 413 6843
rect 447 6809 482 6843
rect 516 6809 551 6843
rect 585 6809 620 6843
rect 654 6809 689 6843
rect 723 6809 758 6843
rect 792 6809 827 6843
rect 861 6809 896 6843
rect 930 6809 965 6843
rect 999 6809 1034 6843
rect 1068 6809 1103 6843
rect 1137 6809 1172 6843
rect 1206 6809 1241 6843
rect 1275 6809 1310 6843
rect 1344 6809 1379 6843
rect 1413 6809 1448 6843
rect 1482 6809 1517 6843
rect 1551 6809 1586 6843
rect 1620 6809 1655 6843
rect 1689 6809 1724 6843
rect 1758 6809 1793 6843
rect 1827 6809 1862 6843
rect 1896 6809 1931 6843
rect 1965 6809 2000 6843
rect 2034 6809 2069 6843
rect 2103 6809 2138 6843
rect 2172 6809 2207 6843
rect 2241 6809 2276 6843
rect 2310 6809 2345 6843
rect 2379 6809 2414 6843
rect 2448 6809 2483 6843
rect 2517 6809 2552 6843
rect 2586 6809 2621 6843
rect 2655 6809 2690 6843
rect 2724 6809 2759 6843
rect 2793 6809 2828 6843
rect 2862 6809 2897 6843
rect 2931 6809 2966 6843
rect 3000 6809 3035 6843
rect 3069 6809 3104 6843
rect 3138 6809 3173 6843
rect 3207 6809 3242 6843
rect 3276 6809 3310 6843
rect 3344 6809 3378 6843
rect 3412 6809 3446 6843
rect 3480 6809 3514 6843
rect 3548 6809 3582 6843
rect 3616 6809 3650 6843
rect 3684 6809 3718 6843
rect 3752 6809 3786 6843
rect 3820 6809 3854 6843
rect 3888 6809 3922 6843
rect 3956 6809 3990 6843
rect 4024 6809 4058 6843
rect 4092 6809 4126 6843
rect 4160 6809 4194 6843
rect 4228 6809 4262 6843
rect 4296 6809 4330 6843
rect 4364 6809 4398 6843
rect 4432 6809 4466 6843
rect 4500 6809 4534 6843
rect 4568 6809 4602 6843
rect 4636 6809 4670 6843
rect 4704 6809 4738 6843
rect 4772 6809 4806 6843
rect 4840 6809 4874 6843
rect 4908 6809 4942 6843
rect 4976 6809 5010 6843
rect 5044 6809 5078 6843
rect 5112 6809 5146 6843
rect 5180 6809 5214 6843
rect 5248 6809 5282 6843
rect 5316 6809 5350 6843
rect 5384 6809 5418 6843
rect 5452 6809 5486 6843
rect 5520 6809 5554 6843
rect 5588 6809 5622 6843
rect 5656 6809 5690 6843
rect 5724 6809 5758 6843
rect 5792 6809 5826 6843
rect 5860 6809 5894 6843
rect 5928 6809 5962 6843
rect 5996 6809 6030 6843
rect 6064 6809 6098 6843
rect 6132 6809 6166 6843
rect 6200 6809 6234 6843
rect 6268 6809 6302 6843
rect 6336 6809 6370 6843
rect 6404 6809 6438 6843
rect 6472 6809 6506 6843
rect 6540 6809 6574 6843
rect 6608 6809 6642 6843
rect 6676 6809 6710 6843
rect 6744 6809 6778 6843
rect 6812 6809 6846 6843
rect 6880 6809 6914 6843
rect 6948 6809 6982 6843
rect 7016 6809 7050 6843
rect 7084 6809 7108 6843
rect 44 6756 7108 6809
rect 44 6722 68 6756
rect 102 6722 137 6756
rect 171 6722 206 6756
rect 240 6722 275 6756
rect 309 6722 344 6756
rect 378 6722 413 6756
rect 447 6722 482 6756
rect 516 6722 551 6756
rect 585 6722 620 6756
rect 654 6722 689 6756
rect 723 6722 758 6756
rect 792 6722 827 6756
rect 861 6722 896 6756
rect 930 6722 965 6756
rect 999 6722 1034 6756
rect 1068 6722 1103 6756
rect 1137 6722 1172 6756
rect 1206 6722 1241 6756
rect 1275 6722 1310 6756
rect 1344 6722 1379 6756
rect 1413 6722 1448 6756
rect 1482 6722 1517 6756
rect 1551 6722 1586 6756
rect 1620 6722 1655 6756
rect 1689 6722 1724 6756
rect 1758 6722 1793 6756
rect 1827 6722 1862 6756
rect 1896 6722 1931 6756
rect 1965 6722 2000 6756
rect 2034 6722 2069 6756
rect 2103 6722 2138 6756
rect 2172 6722 2207 6756
rect 2241 6722 2276 6756
rect 2310 6722 2345 6756
rect 2379 6722 2414 6756
rect 2448 6722 2483 6756
rect 2517 6722 2552 6756
rect 2586 6722 2621 6756
rect 2655 6722 2690 6756
rect 2724 6722 2759 6756
rect 2793 6722 2828 6756
rect 2862 6722 2897 6756
rect 2931 6722 2966 6756
rect 3000 6722 3035 6756
rect 3069 6722 3104 6756
rect 3138 6722 3173 6756
rect 3207 6722 3242 6756
rect 3276 6722 3310 6756
rect 3344 6722 3378 6756
rect 3412 6722 3446 6756
rect 3480 6722 3514 6756
rect 3548 6722 3582 6756
rect 3616 6722 3650 6756
rect 3684 6722 3718 6756
rect 3752 6722 3786 6756
rect 3820 6722 3854 6756
rect 3888 6722 3922 6756
rect 3956 6722 3990 6756
rect 4024 6722 4058 6756
rect 4092 6722 4126 6756
rect 4160 6722 4194 6756
rect 4228 6722 4262 6756
rect 4296 6722 4330 6756
rect 4364 6722 4398 6756
rect 4432 6722 4466 6756
rect 4500 6722 4534 6756
rect 4568 6722 4602 6756
rect 4636 6722 4670 6756
rect 4704 6722 4738 6756
rect 4772 6722 4806 6756
rect 4840 6722 4874 6756
rect 4908 6722 4942 6756
rect 4976 6722 5010 6756
rect 5044 6722 5078 6756
rect 5112 6722 5146 6756
rect 5180 6722 5214 6756
rect 5248 6722 5282 6756
rect 5316 6722 5350 6756
rect 5384 6722 5418 6756
rect 5452 6722 5486 6756
rect 5520 6722 5554 6756
rect 5588 6722 5622 6756
rect 5656 6722 5690 6756
rect 5724 6722 5758 6756
rect 5792 6722 5826 6756
rect 5860 6722 5894 6756
rect 5928 6722 5962 6756
rect 5996 6722 6030 6756
rect 6064 6722 6098 6756
rect 6132 6722 6166 6756
rect 6200 6722 6234 6756
rect 6268 6722 6302 6756
rect 6336 6722 6370 6756
rect 6404 6722 6438 6756
rect 6472 6722 6506 6756
rect 6540 6722 6574 6756
rect 6608 6722 6642 6756
rect 6676 6722 6710 6756
rect 6744 6722 6778 6756
rect 6812 6722 6846 6756
rect 6880 6722 6914 6756
rect 6948 6722 6982 6756
rect 7016 6722 7050 6756
rect 7084 6722 7108 6756
rect 44 6669 7108 6722
rect 44 6635 68 6669
rect 102 6635 137 6669
rect 171 6635 206 6669
rect 240 6635 275 6669
rect 309 6635 344 6669
rect 378 6635 413 6669
rect 447 6635 482 6669
rect 516 6635 551 6669
rect 585 6635 620 6669
rect 654 6635 689 6669
rect 723 6635 758 6669
rect 792 6635 827 6669
rect 861 6635 896 6669
rect 930 6635 965 6669
rect 999 6635 1034 6669
rect 1068 6635 1103 6669
rect 1137 6635 1172 6669
rect 1206 6635 1241 6669
rect 1275 6635 1310 6669
rect 1344 6635 1379 6669
rect 1413 6635 1448 6669
rect 1482 6635 1517 6669
rect 1551 6635 1586 6669
rect 1620 6635 1655 6669
rect 1689 6635 1724 6669
rect 1758 6635 1793 6669
rect 1827 6635 1862 6669
rect 1896 6635 1931 6669
rect 1965 6635 2000 6669
rect 2034 6635 2069 6669
rect 2103 6635 2138 6669
rect 2172 6635 2207 6669
rect 2241 6635 2276 6669
rect 2310 6635 2345 6669
rect 2379 6635 2414 6669
rect 2448 6635 2483 6669
rect 2517 6635 2552 6669
rect 2586 6635 2621 6669
rect 2655 6635 2690 6669
rect 2724 6635 2759 6669
rect 2793 6635 2828 6669
rect 2862 6635 2897 6669
rect 2931 6635 2966 6669
rect 3000 6635 3035 6669
rect 3069 6635 3104 6669
rect 3138 6635 3173 6669
rect 3207 6635 3242 6669
rect 3276 6635 3310 6669
rect 3344 6635 3378 6669
rect 3412 6635 3446 6669
rect 3480 6635 3514 6669
rect 3548 6635 3582 6669
rect 3616 6635 3650 6669
rect 3684 6635 3718 6669
rect 3752 6635 3786 6669
rect 3820 6635 3854 6669
rect 3888 6635 3922 6669
rect 3956 6635 3990 6669
rect 4024 6635 4058 6669
rect 4092 6635 4126 6669
rect 4160 6635 4194 6669
rect 4228 6635 4262 6669
rect 4296 6635 4330 6669
rect 4364 6635 4398 6669
rect 4432 6635 4466 6669
rect 4500 6635 4534 6669
rect 4568 6635 4602 6669
rect 4636 6635 4670 6669
rect 4704 6635 4738 6669
rect 4772 6635 4806 6669
rect 4840 6635 4874 6669
rect 4908 6635 4942 6669
rect 4976 6635 5010 6669
rect 5044 6635 5078 6669
rect 5112 6635 5146 6669
rect 5180 6635 5214 6669
rect 5248 6635 5282 6669
rect 5316 6635 5350 6669
rect 5384 6635 5418 6669
rect 5452 6635 5486 6669
rect 5520 6635 5554 6669
rect 5588 6635 5622 6669
rect 5656 6635 5690 6669
rect 5724 6635 5758 6669
rect 5792 6635 5826 6669
rect 5860 6635 5894 6669
rect 5928 6635 5962 6669
rect 5996 6635 6030 6669
rect 6064 6635 6098 6669
rect 6132 6635 6166 6669
rect 6200 6635 6234 6669
rect 6268 6635 6302 6669
rect 6336 6635 6370 6669
rect 6404 6635 6438 6669
rect 6472 6635 6506 6669
rect 6540 6635 6574 6669
rect 6608 6635 6642 6669
rect 6676 6635 6710 6669
rect 6744 6635 6778 6669
rect 6812 6635 6846 6669
rect 6880 6635 6914 6669
rect 6948 6635 6982 6669
rect 7016 6635 7050 6669
rect 7084 6635 7108 6669
rect 12493 6809 12517 6843
rect 12551 6809 12586 6843
rect 12620 6809 12655 6843
rect 12689 6809 12724 6843
rect 12758 6809 12793 6843
rect 12827 6809 12862 6843
rect 12896 6809 12931 6843
rect 12965 6809 13000 6843
rect 13034 6809 13069 6843
rect 13103 6809 13138 6843
rect 13172 6809 13207 6843
rect 13241 6809 13276 6843
rect 13310 6809 13345 6843
rect 13379 6809 13414 6843
rect 13448 6809 13483 6843
rect 13517 6809 13552 6843
rect 13586 6809 13621 6843
rect 13655 6809 13690 6843
rect 13724 6809 13759 6843
rect 13793 6809 13828 6843
rect 13862 6809 13897 6843
rect 13931 6809 13966 6843
rect 14000 6809 14035 6843
rect 14069 6809 14104 6843
rect 14138 6809 14173 6843
rect 14207 6809 14242 6843
rect 14276 6809 14311 6843
rect 14345 6809 14380 6843
rect 14414 6809 14449 6843
rect 14483 6809 14518 6843
rect 14552 6809 14587 6843
rect 14621 6809 14655 6843
rect 14689 6809 14723 6843
rect 14757 6809 14791 6843
rect 14825 6809 14859 6843
rect 14893 6809 15117 6843
rect 12493 6805 15117 6809
rect 12493 6771 14932 6805
rect 14966 6771 15000 6805
rect 15034 6771 15068 6805
rect 15102 6771 15117 6805
rect 12493 6756 15117 6771
rect 12493 6722 12517 6756
rect 12551 6722 12586 6756
rect 12620 6722 12655 6756
rect 12689 6722 12724 6756
rect 12758 6722 12793 6756
rect 12827 6722 12862 6756
rect 12896 6722 12931 6756
rect 12965 6722 13000 6756
rect 13034 6722 13069 6756
rect 13103 6722 13138 6756
rect 13172 6722 13207 6756
rect 13241 6722 13276 6756
rect 13310 6722 13345 6756
rect 13379 6722 13414 6756
rect 13448 6722 13483 6756
rect 13517 6722 13552 6756
rect 13586 6722 13621 6756
rect 13655 6722 13690 6756
rect 13724 6722 13759 6756
rect 13793 6722 13828 6756
rect 13862 6722 13897 6756
rect 13931 6722 13966 6756
rect 14000 6722 14035 6756
rect 14069 6722 14104 6756
rect 14138 6722 14173 6756
rect 14207 6722 14242 6756
rect 14276 6722 14311 6756
rect 14345 6722 14380 6756
rect 14414 6722 14449 6756
rect 14483 6722 14518 6756
rect 14552 6722 14587 6756
rect 14621 6722 14655 6756
rect 14689 6722 14723 6756
rect 14757 6722 14791 6756
rect 14825 6722 14859 6756
rect 14893 6731 15117 6756
rect 14893 6722 14932 6731
rect 12493 6697 14932 6722
rect 14966 6697 15000 6731
rect 15034 6697 15068 6731
rect 15102 6697 15117 6731
rect 12493 6669 15117 6697
rect 12493 6635 12517 6669
rect 12551 6635 12586 6669
rect 12620 6635 12655 6669
rect 12689 6635 12724 6669
rect 12758 6635 12793 6669
rect 12827 6635 12862 6669
rect 12896 6635 12931 6669
rect 12965 6635 13000 6669
rect 13034 6635 13069 6669
rect 13103 6635 13138 6669
rect 13172 6635 13207 6669
rect 13241 6635 13276 6669
rect 13310 6635 13345 6669
rect 13379 6635 13414 6669
rect 13448 6635 13483 6669
rect 13517 6635 13552 6669
rect 13586 6635 13621 6669
rect 13655 6635 13690 6669
rect 13724 6635 13759 6669
rect 13793 6635 13828 6669
rect 13862 6635 13897 6669
rect 13931 6635 13966 6669
rect 14000 6635 14035 6669
rect 14069 6635 14104 6669
rect 14138 6635 14173 6669
rect 14207 6635 14242 6669
rect 14276 6635 14311 6669
rect 14345 6635 14380 6669
rect 14414 6635 14449 6669
rect 14483 6635 14518 6669
rect 14552 6635 14587 6669
rect 14621 6635 14655 6669
rect 14689 6635 14723 6669
rect 14757 6635 14791 6669
rect 14825 6635 14859 6669
rect 14893 6657 15117 6669
rect 14893 6635 14932 6657
rect 44 6623 14932 6635
rect 14966 6623 15000 6657
rect 15034 6623 15068 6657
rect 15102 6623 15117 6657
rect 44 6583 15117 6623
rect 44 6582 14932 6583
rect 44 6548 68 6582
rect 102 6548 137 6582
rect 171 6548 206 6582
rect 240 6548 275 6582
rect 309 6548 344 6582
rect 378 6548 413 6582
rect 447 6548 482 6582
rect 516 6548 551 6582
rect 585 6548 620 6582
rect 654 6548 689 6582
rect 723 6548 758 6582
rect 792 6548 827 6582
rect 861 6548 896 6582
rect 930 6548 965 6582
rect 999 6548 1034 6582
rect 1068 6548 1103 6582
rect 1137 6548 1172 6582
rect 1206 6548 1241 6582
rect 1275 6548 1310 6582
rect 1344 6548 1379 6582
rect 1413 6548 1448 6582
rect 1482 6548 1517 6582
rect 1551 6548 1586 6582
rect 1620 6548 1655 6582
rect 1689 6548 1724 6582
rect 1758 6548 1793 6582
rect 1827 6548 1862 6582
rect 1896 6548 1931 6582
rect 1965 6548 2000 6582
rect 2034 6548 2069 6582
rect 2103 6548 2138 6582
rect 2172 6548 2207 6582
rect 2241 6548 2276 6582
rect 2310 6548 2345 6582
rect 2379 6548 2414 6582
rect 2448 6548 2483 6582
rect 2517 6548 2551 6582
rect 2585 6548 2619 6582
rect 2653 6548 2687 6582
rect 2721 6548 2755 6582
rect 2789 6548 2823 6582
rect 2857 6548 2891 6582
rect 2925 6548 2959 6582
rect 2993 6548 3027 6582
rect 3061 6548 3095 6582
rect 3129 6548 3163 6582
rect 3197 6548 3231 6582
rect 3265 6548 3299 6582
rect 3333 6548 3367 6582
rect 3401 6548 3435 6582
rect 3469 6548 3503 6582
rect 3537 6548 3571 6582
rect 3605 6548 3639 6582
rect 3673 6548 3707 6582
rect 3741 6548 3775 6582
rect 3809 6548 3843 6582
rect 3877 6548 3911 6582
rect 3945 6548 3979 6582
rect 4013 6548 4047 6582
rect 4081 6548 4115 6582
rect 4149 6548 4183 6582
rect 4217 6548 4251 6582
rect 4285 6548 4319 6582
rect 4353 6548 4387 6582
rect 4421 6548 4455 6582
rect 4489 6548 4523 6582
rect 4557 6548 4591 6582
rect 4625 6548 4659 6582
rect 4693 6548 4727 6582
rect 4761 6548 4795 6582
rect 4829 6548 4863 6582
rect 4897 6548 4931 6582
rect 4965 6548 4999 6582
rect 5033 6548 5067 6582
rect 5101 6548 5135 6582
rect 5169 6548 5203 6582
rect 5237 6548 5271 6582
rect 5305 6548 5339 6582
rect 5373 6548 5407 6582
rect 5441 6548 5475 6582
rect 5509 6548 5543 6582
rect 5577 6548 5611 6582
rect 5645 6548 5679 6582
rect 5713 6548 5747 6582
rect 5781 6548 5815 6582
rect 5849 6548 5883 6582
rect 5917 6548 5951 6582
rect 5985 6548 6019 6582
rect 6053 6548 6087 6582
rect 6121 6548 6155 6582
rect 6189 6548 6223 6582
rect 6257 6548 6291 6582
rect 6325 6548 6359 6582
rect 6393 6548 6427 6582
rect 6461 6548 6495 6582
rect 6529 6548 6563 6582
rect 6597 6548 6631 6582
rect 6665 6548 6699 6582
rect 6733 6548 6767 6582
rect 6801 6548 6835 6582
rect 6869 6548 6903 6582
rect 6937 6548 6971 6582
rect 7005 6548 7039 6582
rect 7073 6548 7107 6582
rect 7141 6548 7175 6582
rect 7209 6548 7243 6582
rect 7277 6548 7311 6582
rect 7345 6548 7379 6582
rect 7413 6548 7447 6582
rect 7481 6548 7515 6582
rect 7549 6548 7583 6582
rect 7617 6548 7651 6582
rect 7685 6548 7719 6582
rect 7753 6548 7787 6582
rect 7821 6548 7855 6582
rect 7889 6548 7923 6582
rect 7957 6548 7991 6582
rect 8025 6548 8059 6582
rect 8093 6548 8127 6582
rect 8161 6548 8195 6582
rect 8229 6548 8263 6582
rect 8297 6548 8331 6582
rect 8365 6548 8399 6582
rect 8433 6548 8467 6582
rect 8501 6548 8535 6582
rect 8569 6548 8603 6582
rect 8637 6548 8671 6582
rect 8705 6548 8739 6582
rect 8773 6548 8807 6582
rect 8841 6548 8875 6582
rect 8909 6548 8943 6582
rect 8977 6548 9011 6582
rect 9045 6548 9079 6582
rect 9113 6548 9147 6582
rect 9181 6548 9215 6582
rect 9249 6548 9283 6582
rect 9317 6548 9351 6582
rect 9385 6548 9419 6582
rect 9453 6548 9487 6582
rect 9521 6548 9555 6582
rect 9589 6548 9623 6582
rect 9657 6548 9691 6582
rect 9725 6548 9759 6582
rect 9793 6548 9827 6582
rect 9861 6548 9895 6582
rect 9929 6548 9963 6582
rect 9997 6548 10031 6582
rect 10065 6548 10099 6582
rect 10133 6548 10167 6582
rect 10201 6548 10235 6582
rect 10269 6548 10303 6582
rect 10337 6548 10371 6582
rect 10405 6548 10439 6582
rect 10473 6548 10507 6582
rect 10541 6548 10575 6582
rect 10609 6548 10643 6582
rect 10677 6548 10711 6582
rect 10745 6548 10779 6582
rect 10813 6548 10847 6582
rect 10881 6548 10915 6582
rect 10949 6548 10983 6582
rect 11017 6548 11051 6582
rect 11085 6548 11119 6582
rect 11153 6548 11187 6582
rect 11221 6548 11255 6582
rect 11289 6548 11323 6582
rect 11357 6548 11391 6582
rect 11425 6548 11459 6582
rect 11493 6548 11527 6582
rect 11561 6548 11595 6582
rect 11629 6548 11663 6582
rect 11697 6548 11731 6582
rect 11765 6548 11799 6582
rect 11833 6548 11867 6582
rect 11901 6548 11935 6582
rect 11969 6548 12003 6582
rect 12037 6548 12071 6582
rect 12105 6548 12139 6582
rect 12173 6548 12207 6582
rect 12241 6548 12275 6582
rect 12309 6548 12343 6582
rect 12377 6548 12411 6582
rect 12445 6548 12479 6582
rect 12513 6548 12547 6582
rect 12581 6548 12615 6582
rect 12649 6548 12683 6582
rect 12717 6548 12751 6582
rect 12785 6548 12819 6582
rect 12853 6548 12887 6582
rect 12921 6548 12955 6582
rect 12989 6548 13023 6582
rect 13057 6548 13091 6582
rect 13125 6548 13159 6582
rect 13193 6548 13227 6582
rect 13261 6548 13295 6582
rect 13329 6548 13363 6582
rect 13397 6548 13431 6582
rect 13465 6548 13499 6582
rect 13533 6548 13567 6582
rect 13601 6548 13635 6582
rect 13669 6548 13703 6582
rect 13737 6548 13771 6582
rect 13805 6548 13839 6582
rect 13873 6548 13907 6582
rect 13941 6548 13975 6582
rect 14009 6548 14043 6582
rect 14077 6548 14111 6582
rect 14145 6548 14179 6582
rect 14213 6548 14247 6582
rect 14281 6548 14315 6582
rect 14349 6548 14383 6582
rect 14417 6548 14451 6582
rect 14485 6548 14519 6582
rect 14553 6548 14587 6582
rect 14621 6548 14655 6582
rect 14689 6548 14723 6582
rect 14757 6548 14791 6582
rect 14825 6548 14859 6582
rect 14893 6549 14932 6582
rect 14966 6549 15000 6583
rect 15034 6549 15068 6583
rect 15102 6549 15117 6583
rect 14893 6548 15117 6549
rect 44 6509 15117 6548
rect 44 6508 14932 6509
rect 44 6474 68 6508
rect 102 6474 137 6508
rect 171 6474 206 6508
rect 240 6474 275 6508
rect 309 6474 344 6508
rect 378 6474 413 6508
rect 447 6474 482 6508
rect 516 6474 551 6508
rect 585 6474 620 6508
rect 654 6474 689 6508
rect 723 6474 758 6508
rect 792 6474 827 6508
rect 861 6474 896 6508
rect 930 6474 965 6508
rect 999 6474 1034 6508
rect 1068 6474 1103 6508
rect 1137 6474 1172 6508
rect 1206 6474 1241 6508
rect 1275 6474 1310 6508
rect 1344 6474 1379 6508
rect 1413 6474 1448 6508
rect 1482 6474 1517 6508
rect 1551 6474 1586 6508
rect 1620 6474 1655 6508
rect 1689 6474 1724 6508
rect 1758 6474 1793 6508
rect 1827 6474 1862 6508
rect 1896 6474 1931 6508
rect 1965 6474 2000 6508
rect 2034 6474 2069 6508
rect 2103 6474 2138 6508
rect 2172 6474 2207 6508
rect 2241 6474 2276 6508
rect 2310 6474 2345 6508
rect 2379 6474 2414 6508
rect 2448 6474 2483 6508
rect 2517 6474 2551 6508
rect 2585 6474 2619 6508
rect 2653 6474 2687 6508
rect 2721 6474 2755 6508
rect 2789 6474 2823 6508
rect 2857 6474 2891 6508
rect 2925 6474 2959 6508
rect 2993 6474 3027 6508
rect 3061 6474 3095 6508
rect 3129 6474 3163 6508
rect 3197 6474 3231 6508
rect 3265 6474 3299 6508
rect 3333 6474 3367 6508
rect 3401 6474 3435 6508
rect 3469 6474 3503 6508
rect 3537 6474 3571 6508
rect 3605 6474 3639 6508
rect 3673 6474 3707 6508
rect 3741 6474 3775 6508
rect 3809 6474 3843 6508
rect 3877 6474 3911 6508
rect 3945 6474 3979 6508
rect 4013 6474 4047 6508
rect 4081 6474 4115 6508
rect 4149 6474 4183 6508
rect 4217 6474 4251 6508
rect 4285 6474 4319 6508
rect 4353 6474 4387 6508
rect 4421 6474 4455 6508
rect 4489 6474 4523 6508
rect 4557 6474 4591 6508
rect 4625 6474 4659 6508
rect 4693 6474 4727 6508
rect 4761 6474 4795 6508
rect 4829 6474 4863 6508
rect 4897 6474 4931 6508
rect 4965 6474 4999 6508
rect 5033 6474 5067 6508
rect 5101 6474 5135 6508
rect 5169 6474 5203 6508
rect 5237 6474 5271 6508
rect 5305 6474 5339 6508
rect 5373 6474 5407 6508
rect 5441 6474 5475 6508
rect 5509 6474 5543 6508
rect 5577 6474 5611 6508
rect 5645 6474 5679 6508
rect 5713 6474 5747 6508
rect 5781 6474 5815 6508
rect 5849 6474 5883 6508
rect 5917 6474 5951 6508
rect 5985 6474 6019 6508
rect 6053 6474 6087 6508
rect 6121 6474 6155 6508
rect 6189 6474 6223 6508
rect 6257 6474 6291 6508
rect 6325 6474 6359 6508
rect 6393 6474 6427 6508
rect 6461 6474 6495 6508
rect 6529 6474 6563 6508
rect 6597 6474 6631 6508
rect 6665 6474 6699 6508
rect 6733 6474 6767 6508
rect 6801 6474 6835 6508
rect 6869 6474 6903 6508
rect 6937 6474 6971 6508
rect 7005 6474 7039 6508
rect 7073 6474 7107 6508
rect 7141 6474 7175 6508
rect 7209 6474 7243 6508
rect 7277 6474 7311 6508
rect 7345 6474 7379 6508
rect 7413 6474 7447 6508
rect 7481 6474 7515 6508
rect 7549 6474 7583 6508
rect 7617 6474 7651 6508
rect 7685 6474 7719 6508
rect 7753 6474 7787 6508
rect 7821 6474 7855 6508
rect 7889 6474 7923 6508
rect 7957 6474 7991 6508
rect 8025 6474 8059 6508
rect 8093 6474 8127 6508
rect 8161 6474 8195 6508
rect 8229 6474 8263 6508
rect 8297 6474 8331 6508
rect 8365 6474 8399 6508
rect 8433 6474 8467 6508
rect 8501 6474 8535 6508
rect 8569 6474 8603 6508
rect 8637 6474 8671 6508
rect 8705 6474 8739 6508
rect 8773 6474 8807 6508
rect 8841 6474 8875 6508
rect 8909 6474 8943 6508
rect 8977 6474 9011 6508
rect 9045 6474 9079 6508
rect 9113 6474 9147 6508
rect 9181 6474 9215 6508
rect 9249 6474 9283 6508
rect 9317 6474 9351 6508
rect 9385 6474 9419 6508
rect 9453 6474 9487 6508
rect 9521 6474 9555 6508
rect 9589 6474 9623 6508
rect 9657 6474 9691 6508
rect 9725 6474 9759 6508
rect 9793 6474 9827 6508
rect 9861 6474 9895 6508
rect 9929 6474 9963 6508
rect 9997 6474 10031 6508
rect 10065 6474 10099 6508
rect 10133 6474 10167 6508
rect 10201 6474 10235 6508
rect 10269 6474 10303 6508
rect 10337 6474 10371 6508
rect 10405 6474 10439 6508
rect 10473 6474 10507 6508
rect 10541 6474 10575 6508
rect 10609 6474 10643 6508
rect 10677 6474 10711 6508
rect 10745 6474 10779 6508
rect 10813 6474 10847 6508
rect 10881 6474 10915 6508
rect 10949 6474 10983 6508
rect 11017 6474 11051 6508
rect 11085 6474 11119 6508
rect 11153 6474 11187 6508
rect 11221 6474 11255 6508
rect 11289 6474 11323 6508
rect 11357 6474 11391 6508
rect 11425 6474 11459 6508
rect 11493 6474 11527 6508
rect 11561 6474 11595 6508
rect 11629 6474 11663 6508
rect 11697 6474 11731 6508
rect 11765 6474 11799 6508
rect 11833 6474 11867 6508
rect 11901 6474 11935 6508
rect 11969 6474 12003 6508
rect 12037 6474 12071 6508
rect 12105 6474 12139 6508
rect 12173 6474 12207 6508
rect 12241 6474 12275 6508
rect 12309 6474 12343 6508
rect 12377 6474 12411 6508
rect 12445 6474 12479 6508
rect 12513 6474 12547 6508
rect 12581 6474 12615 6508
rect 12649 6474 12683 6508
rect 12717 6474 12751 6508
rect 12785 6474 12819 6508
rect 12853 6474 12887 6508
rect 12921 6474 12955 6508
rect 12989 6474 13023 6508
rect 13057 6474 13091 6508
rect 13125 6474 13159 6508
rect 13193 6474 13227 6508
rect 13261 6474 13295 6508
rect 13329 6474 13363 6508
rect 13397 6474 13431 6508
rect 13465 6474 13499 6508
rect 13533 6474 13567 6508
rect 13601 6474 13635 6508
rect 13669 6474 13703 6508
rect 13737 6474 13771 6508
rect 13805 6474 13839 6508
rect 13873 6474 13907 6508
rect 13941 6474 13975 6508
rect 14009 6474 14043 6508
rect 14077 6474 14111 6508
rect 14145 6474 14179 6508
rect 14213 6474 14247 6508
rect 14281 6474 14315 6508
rect 14349 6474 14383 6508
rect 14417 6474 14451 6508
rect 14485 6474 14519 6508
rect 14553 6474 14587 6508
rect 14621 6474 14655 6508
rect 14689 6474 14723 6508
rect 14757 6474 14791 6508
rect 14825 6474 14859 6508
rect 14893 6475 14932 6508
rect 14966 6475 15000 6509
rect 15034 6475 15068 6509
rect 15102 6475 15117 6509
rect 14893 6474 15117 6475
rect 44 6435 15117 6474
rect 44 6434 14932 6435
rect 44 6400 68 6434
rect 102 6400 137 6434
rect 171 6400 206 6434
rect 240 6400 275 6434
rect 309 6400 344 6434
rect 378 6400 413 6434
rect 447 6400 482 6434
rect 516 6400 551 6434
rect 585 6400 620 6434
rect 654 6400 689 6434
rect 723 6400 758 6434
rect 792 6400 827 6434
rect 861 6400 896 6434
rect 930 6400 965 6434
rect 999 6400 1034 6434
rect 1068 6400 1103 6434
rect 1137 6400 1172 6434
rect 1206 6400 1241 6434
rect 1275 6400 1310 6434
rect 1344 6400 1379 6434
rect 1413 6400 1448 6434
rect 1482 6400 1517 6434
rect 1551 6400 1586 6434
rect 1620 6400 1655 6434
rect 1689 6400 1724 6434
rect 1758 6400 1793 6434
rect 1827 6400 1862 6434
rect 1896 6400 1931 6434
rect 1965 6400 2000 6434
rect 2034 6400 2069 6434
rect 2103 6400 2138 6434
rect 2172 6400 2207 6434
rect 2241 6400 2276 6434
rect 2310 6400 2345 6434
rect 2379 6400 2414 6434
rect 2448 6400 2483 6434
rect 2517 6400 2551 6434
rect 2585 6400 2619 6434
rect 2653 6400 2687 6434
rect 2721 6400 2755 6434
rect 2789 6400 2823 6434
rect 2857 6400 2891 6434
rect 2925 6400 2959 6434
rect 2993 6400 3027 6434
rect 3061 6400 3095 6434
rect 3129 6400 3163 6434
rect 3197 6400 3231 6434
rect 3265 6400 3299 6434
rect 3333 6400 3367 6434
rect 3401 6400 3435 6434
rect 3469 6400 3503 6434
rect 3537 6400 3571 6434
rect 3605 6400 3639 6434
rect 3673 6400 3707 6434
rect 3741 6400 3775 6434
rect 3809 6400 3843 6434
rect 3877 6400 3911 6434
rect 3945 6400 3979 6434
rect 4013 6400 4047 6434
rect 4081 6400 4115 6434
rect 4149 6400 4183 6434
rect 4217 6400 4251 6434
rect 4285 6400 4319 6434
rect 4353 6400 4387 6434
rect 4421 6400 4455 6434
rect 4489 6400 4523 6434
rect 4557 6400 4591 6434
rect 4625 6400 4659 6434
rect 4693 6400 4727 6434
rect 4761 6400 4795 6434
rect 4829 6400 4863 6434
rect 4897 6400 4931 6434
rect 4965 6400 4999 6434
rect 5033 6400 5067 6434
rect 5101 6400 5135 6434
rect 5169 6400 5203 6434
rect 5237 6400 5271 6434
rect 5305 6400 5339 6434
rect 5373 6400 5407 6434
rect 5441 6400 5475 6434
rect 5509 6400 5543 6434
rect 5577 6400 5611 6434
rect 5645 6400 5679 6434
rect 5713 6400 5747 6434
rect 5781 6400 5815 6434
rect 5849 6400 5883 6434
rect 5917 6400 5951 6434
rect 5985 6400 6019 6434
rect 6053 6400 6087 6434
rect 6121 6400 6155 6434
rect 6189 6400 6223 6434
rect 6257 6400 6291 6434
rect 6325 6400 6359 6434
rect 6393 6400 6427 6434
rect 6461 6400 6495 6434
rect 6529 6400 6563 6434
rect 6597 6400 6631 6434
rect 6665 6400 6699 6434
rect 6733 6400 6767 6434
rect 6801 6400 6835 6434
rect 6869 6400 6903 6434
rect 6937 6400 6971 6434
rect 7005 6400 7039 6434
rect 7073 6400 7107 6434
rect 7141 6400 7175 6434
rect 7209 6400 7243 6434
rect 7277 6400 7311 6434
rect 7345 6400 7379 6434
rect 7413 6400 7447 6434
rect 7481 6400 7515 6434
rect 7549 6400 7583 6434
rect 7617 6400 7651 6434
rect 7685 6400 7719 6434
rect 7753 6400 7787 6434
rect 7821 6400 7855 6434
rect 7889 6400 7923 6434
rect 7957 6400 7991 6434
rect 8025 6400 8059 6434
rect 8093 6400 8127 6434
rect 8161 6400 8195 6434
rect 8229 6400 8263 6434
rect 8297 6400 8331 6434
rect 8365 6400 8399 6434
rect 8433 6400 8467 6434
rect 8501 6400 8535 6434
rect 8569 6400 8603 6434
rect 8637 6400 8671 6434
rect 8705 6400 8739 6434
rect 8773 6400 8807 6434
rect 8841 6400 8875 6434
rect 8909 6400 8943 6434
rect 8977 6400 9011 6434
rect 9045 6400 9079 6434
rect 9113 6400 9147 6434
rect 9181 6400 9215 6434
rect 9249 6400 9283 6434
rect 9317 6400 9351 6434
rect 9385 6400 9419 6434
rect 9453 6400 9487 6434
rect 9521 6400 9555 6434
rect 9589 6400 9623 6434
rect 9657 6400 9691 6434
rect 9725 6400 9759 6434
rect 9793 6400 9827 6434
rect 9861 6400 9895 6434
rect 9929 6400 9963 6434
rect 9997 6400 10031 6434
rect 10065 6400 10099 6434
rect 10133 6400 10167 6434
rect 10201 6400 10235 6434
rect 10269 6400 10303 6434
rect 10337 6400 10371 6434
rect 10405 6400 10439 6434
rect 10473 6400 10507 6434
rect 10541 6400 10575 6434
rect 10609 6400 10643 6434
rect 10677 6400 10711 6434
rect 10745 6400 10779 6434
rect 10813 6400 10847 6434
rect 10881 6400 10915 6434
rect 10949 6400 10983 6434
rect 11017 6400 11051 6434
rect 11085 6400 11119 6434
rect 11153 6400 11187 6434
rect 11221 6400 11255 6434
rect 11289 6400 11323 6434
rect 11357 6400 11391 6434
rect 11425 6400 11459 6434
rect 11493 6400 11527 6434
rect 11561 6400 11595 6434
rect 11629 6400 11663 6434
rect 11697 6400 11731 6434
rect 11765 6400 11799 6434
rect 11833 6400 11867 6434
rect 11901 6400 11935 6434
rect 11969 6400 12003 6434
rect 12037 6400 12071 6434
rect 12105 6400 12139 6434
rect 12173 6400 12207 6434
rect 12241 6400 12275 6434
rect 12309 6400 12343 6434
rect 12377 6400 12411 6434
rect 12445 6400 12479 6434
rect 12513 6400 12547 6434
rect 12581 6400 12615 6434
rect 12649 6400 12683 6434
rect 12717 6400 12751 6434
rect 12785 6400 12819 6434
rect 12853 6400 12887 6434
rect 12921 6400 12955 6434
rect 12989 6400 13023 6434
rect 13057 6400 13091 6434
rect 13125 6400 13159 6434
rect 13193 6400 13227 6434
rect 13261 6400 13295 6434
rect 13329 6400 13363 6434
rect 13397 6400 13431 6434
rect 13465 6400 13499 6434
rect 13533 6400 13567 6434
rect 13601 6400 13635 6434
rect 13669 6400 13703 6434
rect 13737 6400 13771 6434
rect 13805 6400 13839 6434
rect 13873 6400 13907 6434
rect 13941 6400 13975 6434
rect 14009 6400 14043 6434
rect 14077 6400 14111 6434
rect 14145 6400 14179 6434
rect 14213 6400 14247 6434
rect 14281 6400 14315 6434
rect 14349 6400 14383 6434
rect 14417 6400 14451 6434
rect 14485 6400 14519 6434
rect 14553 6400 14587 6434
rect 14621 6400 14655 6434
rect 14689 6400 14723 6434
rect 14757 6400 14791 6434
rect 14825 6400 14859 6434
rect 14893 6401 14932 6434
rect 14966 6401 15000 6435
rect 15034 6401 15068 6435
rect 15102 6401 15117 6435
rect 14893 6400 15117 6401
rect 44 6360 15117 6400
rect 44 6326 68 6360
rect 102 6326 137 6360
rect 171 6326 206 6360
rect 240 6326 275 6360
rect 309 6326 344 6360
rect 378 6326 413 6360
rect 447 6326 482 6360
rect 516 6326 551 6360
rect 585 6326 620 6360
rect 654 6326 689 6360
rect 723 6326 758 6360
rect 792 6326 827 6360
rect 861 6326 896 6360
rect 930 6326 965 6360
rect 999 6326 1034 6360
rect 1068 6326 1103 6360
rect 1137 6326 1172 6360
rect 1206 6326 1241 6360
rect 1275 6326 1310 6360
rect 1344 6326 1379 6360
rect 1413 6326 1448 6360
rect 1482 6326 1517 6360
rect 1551 6326 1586 6360
rect 1620 6326 1655 6360
rect 1689 6326 1724 6360
rect 1758 6326 1793 6360
rect 1827 6326 1862 6360
rect 1896 6326 1931 6360
rect 1965 6326 2000 6360
rect 2034 6326 2069 6360
rect 2103 6326 2138 6360
rect 2172 6326 2207 6360
rect 2241 6326 2276 6360
rect 2310 6326 2345 6360
rect 2379 6326 2414 6360
rect 2448 6326 2483 6360
rect 2517 6326 2551 6360
rect 2585 6326 2619 6360
rect 2653 6326 2687 6360
rect 2721 6326 2755 6360
rect 2789 6326 2823 6360
rect 2857 6326 2891 6360
rect 2925 6326 2959 6360
rect 2993 6326 3027 6360
rect 3061 6326 3095 6360
rect 3129 6326 3163 6360
rect 3197 6326 3231 6360
rect 3265 6326 3299 6360
rect 3333 6326 3367 6360
rect 3401 6326 3435 6360
rect 3469 6326 3503 6360
rect 3537 6326 3571 6360
rect 3605 6326 3639 6360
rect 3673 6326 3707 6360
rect 3741 6326 3775 6360
rect 3809 6326 3843 6360
rect 3877 6326 3911 6360
rect 3945 6326 3979 6360
rect 4013 6326 4047 6360
rect 4081 6326 4115 6360
rect 4149 6326 4183 6360
rect 4217 6326 4251 6360
rect 4285 6326 4319 6360
rect 4353 6326 4387 6360
rect 4421 6326 4455 6360
rect 4489 6326 4523 6360
rect 4557 6326 4591 6360
rect 4625 6326 4659 6360
rect 4693 6326 4727 6360
rect 4761 6326 4795 6360
rect 4829 6326 4863 6360
rect 4897 6326 4931 6360
rect 4965 6326 4999 6360
rect 5033 6326 5067 6360
rect 5101 6326 5135 6360
rect 5169 6326 5203 6360
rect 5237 6326 5271 6360
rect 5305 6326 5339 6360
rect 5373 6326 5407 6360
rect 5441 6326 5475 6360
rect 5509 6326 5543 6360
rect 5577 6326 5611 6360
rect 5645 6326 5679 6360
rect 5713 6326 5747 6360
rect 5781 6326 5815 6360
rect 5849 6326 5883 6360
rect 5917 6326 5951 6360
rect 5985 6326 6019 6360
rect 6053 6326 6087 6360
rect 6121 6326 6155 6360
rect 6189 6326 6223 6360
rect 6257 6326 6291 6360
rect 6325 6326 6359 6360
rect 6393 6326 6427 6360
rect 6461 6326 6495 6360
rect 6529 6326 6563 6360
rect 6597 6326 6631 6360
rect 6665 6326 6699 6360
rect 6733 6326 6767 6360
rect 6801 6326 6835 6360
rect 6869 6326 6903 6360
rect 6937 6326 6971 6360
rect 7005 6326 7039 6360
rect 7073 6326 7107 6360
rect 7141 6326 7175 6360
rect 7209 6326 7243 6360
rect 7277 6326 7311 6360
rect 7345 6326 7379 6360
rect 7413 6326 7447 6360
rect 7481 6326 7515 6360
rect 7549 6326 7583 6360
rect 7617 6326 7651 6360
rect 7685 6326 7719 6360
rect 7753 6326 7787 6360
rect 7821 6326 7855 6360
rect 7889 6326 7923 6360
rect 7957 6326 7991 6360
rect 8025 6326 8059 6360
rect 8093 6326 8127 6360
rect 8161 6326 8195 6360
rect 8229 6326 8263 6360
rect 8297 6326 8331 6360
rect 8365 6326 8399 6360
rect 8433 6326 8467 6360
rect 8501 6326 8535 6360
rect 8569 6326 8603 6360
rect 8637 6326 8671 6360
rect 8705 6326 8739 6360
rect 8773 6326 8807 6360
rect 8841 6326 8875 6360
rect 8909 6326 8943 6360
rect 8977 6326 9011 6360
rect 9045 6326 9079 6360
rect 9113 6326 9147 6360
rect 9181 6326 9215 6360
rect 9249 6326 9283 6360
rect 9317 6326 9351 6360
rect 9385 6326 9419 6360
rect 9453 6326 9487 6360
rect 9521 6326 9555 6360
rect 9589 6326 9623 6360
rect 9657 6326 9691 6360
rect 9725 6326 9759 6360
rect 9793 6326 9827 6360
rect 9861 6326 9895 6360
rect 9929 6326 9963 6360
rect 9997 6326 10031 6360
rect 10065 6326 10099 6360
rect 10133 6326 10167 6360
rect 10201 6326 10235 6360
rect 10269 6326 10303 6360
rect 10337 6326 10371 6360
rect 10405 6326 10439 6360
rect 10473 6326 10507 6360
rect 10541 6326 10575 6360
rect 10609 6326 10643 6360
rect 10677 6326 10711 6360
rect 10745 6326 10779 6360
rect 10813 6326 10847 6360
rect 10881 6326 10915 6360
rect 10949 6326 10983 6360
rect 11017 6326 11051 6360
rect 11085 6326 11119 6360
rect 11153 6326 11187 6360
rect 11221 6326 11255 6360
rect 11289 6326 11323 6360
rect 11357 6326 11391 6360
rect 11425 6326 11459 6360
rect 11493 6326 11527 6360
rect 11561 6326 11595 6360
rect 11629 6326 11663 6360
rect 11697 6326 11731 6360
rect 11765 6326 11799 6360
rect 11833 6326 11867 6360
rect 11901 6326 11935 6360
rect 11969 6326 12003 6360
rect 12037 6326 12071 6360
rect 12105 6326 12139 6360
rect 12173 6326 12207 6360
rect 12241 6326 12275 6360
rect 12309 6326 12343 6360
rect 12377 6326 12411 6360
rect 12445 6326 12479 6360
rect 12513 6326 12547 6360
rect 12581 6326 12615 6360
rect 12649 6326 12683 6360
rect 12717 6326 12751 6360
rect 12785 6326 12819 6360
rect 12853 6326 12887 6360
rect 12921 6326 12955 6360
rect 12989 6326 13023 6360
rect 13057 6326 13091 6360
rect 13125 6326 13159 6360
rect 13193 6326 13227 6360
rect 13261 6326 13295 6360
rect 13329 6326 13363 6360
rect 13397 6326 13431 6360
rect 13465 6326 13499 6360
rect 13533 6326 13567 6360
rect 13601 6326 13635 6360
rect 13669 6326 13703 6360
rect 13737 6326 13771 6360
rect 13805 6326 13839 6360
rect 13873 6326 13907 6360
rect 13941 6326 13975 6360
rect 14009 6326 14043 6360
rect 14077 6326 14111 6360
rect 14145 6326 14179 6360
rect 14213 6326 14247 6360
rect 14281 6326 14315 6360
rect 14349 6326 14383 6360
rect 14417 6326 14451 6360
rect 14485 6326 14519 6360
rect 14553 6326 14587 6360
rect 14621 6326 14655 6360
rect 14689 6326 14723 6360
rect 14757 6326 14791 6360
rect 14825 6326 14859 6360
rect 14893 6326 14932 6360
rect 14966 6326 15000 6360
rect 15034 6326 15068 6360
rect 15102 6326 15117 6360
rect 44 6286 15117 6326
rect 44 6252 68 6286
rect 102 6252 137 6286
rect 171 6252 206 6286
rect 240 6252 275 6286
rect 309 6252 344 6286
rect 378 6252 413 6286
rect 447 6252 482 6286
rect 516 6252 551 6286
rect 585 6252 620 6286
rect 654 6252 689 6286
rect 723 6252 758 6286
rect 792 6252 827 6286
rect 861 6252 896 6286
rect 930 6252 965 6286
rect 999 6252 1034 6286
rect 1068 6252 1103 6286
rect 1137 6252 1172 6286
rect 1206 6252 1241 6286
rect 1275 6252 1310 6286
rect 1344 6252 1379 6286
rect 1413 6252 1448 6286
rect 1482 6252 1517 6286
rect 1551 6252 1586 6286
rect 1620 6252 1655 6286
rect 1689 6252 1724 6286
rect 1758 6252 1793 6286
rect 1827 6252 1862 6286
rect 1896 6252 1931 6286
rect 1965 6252 2000 6286
rect 2034 6252 2069 6286
rect 2103 6252 2138 6286
rect 2172 6252 2207 6286
rect 2241 6252 2276 6286
rect 2310 6252 2345 6286
rect 2379 6252 2414 6286
rect 2448 6252 2483 6286
rect 2517 6252 2551 6286
rect 2585 6252 2619 6286
rect 2653 6252 2687 6286
rect 2721 6252 2755 6286
rect 2789 6252 2823 6286
rect 2857 6252 2891 6286
rect 2925 6252 2959 6286
rect 2993 6252 3027 6286
rect 3061 6252 3095 6286
rect 3129 6252 3163 6286
rect 3197 6252 3231 6286
rect 3265 6252 3299 6286
rect 3333 6252 3367 6286
rect 3401 6252 3435 6286
rect 3469 6252 3503 6286
rect 3537 6252 3571 6286
rect 3605 6252 3639 6286
rect 3673 6252 3707 6286
rect 3741 6252 3775 6286
rect 3809 6252 3843 6286
rect 3877 6252 3911 6286
rect 3945 6252 3979 6286
rect 4013 6252 4047 6286
rect 4081 6252 4115 6286
rect 4149 6252 4183 6286
rect 4217 6252 4251 6286
rect 4285 6252 4319 6286
rect 4353 6252 4387 6286
rect 4421 6252 4455 6286
rect 4489 6252 4523 6286
rect 4557 6252 4591 6286
rect 4625 6252 4659 6286
rect 4693 6252 4727 6286
rect 4761 6252 4795 6286
rect 4829 6252 4863 6286
rect 4897 6252 4931 6286
rect 4965 6252 4999 6286
rect 5033 6252 5067 6286
rect 5101 6252 5135 6286
rect 5169 6252 5203 6286
rect 5237 6252 5271 6286
rect 5305 6252 5339 6286
rect 5373 6252 5407 6286
rect 5441 6252 5475 6286
rect 5509 6252 5543 6286
rect 5577 6252 5611 6286
rect 5645 6252 5679 6286
rect 5713 6252 5747 6286
rect 5781 6252 5815 6286
rect 5849 6252 5883 6286
rect 5917 6252 5951 6286
rect 5985 6252 6019 6286
rect 6053 6252 6087 6286
rect 6121 6252 6155 6286
rect 6189 6252 6223 6286
rect 6257 6252 6291 6286
rect 6325 6252 6359 6286
rect 6393 6252 6427 6286
rect 6461 6252 6495 6286
rect 6529 6252 6563 6286
rect 6597 6252 6631 6286
rect 6665 6252 6699 6286
rect 6733 6252 6767 6286
rect 6801 6252 6835 6286
rect 6869 6252 6903 6286
rect 6937 6252 6971 6286
rect 7005 6252 7039 6286
rect 7073 6252 7107 6286
rect 7141 6252 7175 6286
rect 7209 6252 7243 6286
rect 7277 6252 7311 6286
rect 7345 6252 7379 6286
rect 7413 6252 7447 6286
rect 7481 6252 7515 6286
rect 7549 6252 7583 6286
rect 7617 6252 7651 6286
rect 7685 6252 7719 6286
rect 7753 6252 7787 6286
rect 7821 6252 7855 6286
rect 7889 6252 7923 6286
rect 7957 6252 7991 6286
rect 8025 6252 8059 6286
rect 8093 6252 8127 6286
rect 8161 6252 8195 6286
rect 8229 6252 8263 6286
rect 8297 6252 8331 6286
rect 8365 6252 8399 6286
rect 8433 6252 8467 6286
rect 8501 6252 8535 6286
rect 8569 6252 8603 6286
rect 8637 6252 8671 6286
rect 8705 6252 8739 6286
rect 8773 6252 8807 6286
rect 8841 6252 8875 6286
rect 8909 6252 8943 6286
rect 8977 6252 9011 6286
rect 9045 6252 9079 6286
rect 9113 6252 9147 6286
rect 9181 6252 9215 6286
rect 9249 6252 9283 6286
rect 9317 6252 9351 6286
rect 9385 6252 9419 6286
rect 9453 6252 9487 6286
rect 9521 6252 9555 6286
rect 9589 6252 9623 6286
rect 9657 6252 9691 6286
rect 9725 6252 9759 6286
rect 9793 6252 9827 6286
rect 9861 6252 9895 6286
rect 9929 6252 9963 6286
rect 9997 6252 10031 6286
rect 10065 6252 10099 6286
rect 10133 6252 10167 6286
rect 10201 6252 10235 6286
rect 10269 6252 10303 6286
rect 10337 6252 10371 6286
rect 10405 6252 10439 6286
rect 10473 6252 10507 6286
rect 10541 6252 10575 6286
rect 10609 6252 10643 6286
rect 10677 6252 10711 6286
rect 10745 6252 10779 6286
rect 10813 6252 10847 6286
rect 10881 6252 10915 6286
rect 10949 6252 10983 6286
rect 11017 6252 11051 6286
rect 11085 6252 11119 6286
rect 11153 6252 11187 6286
rect 11221 6252 11255 6286
rect 11289 6252 11323 6286
rect 11357 6252 11391 6286
rect 11425 6252 11459 6286
rect 11493 6252 11527 6286
rect 11561 6252 11595 6286
rect 11629 6252 11663 6286
rect 11697 6252 11731 6286
rect 11765 6252 11799 6286
rect 11833 6252 11867 6286
rect 11901 6252 11935 6286
rect 11969 6252 12003 6286
rect 12037 6252 12071 6286
rect 12105 6252 12139 6286
rect 12173 6252 12207 6286
rect 12241 6252 12275 6286
rect 12309 6252 12343 6286
rect 12377 6252 12411 6286
rect 12445 6252 12479 6286
rect 12513 6252 12547 6286
rect 12581 6252 12615 6286
rect 12649 6252 12683 6286
rect 12717 6252 12751 6286
rect 12785 6252 12819 6286
rect 12853 6252 12887 6286
rect 12921 6252 12955 6286
rect 12989 6252 13023 6286
rect 13057 6252 13091 6286
rect 13125 6252 13159 6286
rect 13193 6252 13227 6286
rect 13261 6252 13295 6286
rect 13329 6252 13363 6286
rect 13397 6252 13431 6286
rect 13465 6252 13499 6286
rect 13533 6252 13567 6286
rect 13601 6252 13635 6286
rect 13669 6252 13703 6286
rect 13737 6252 13771 6286
rect 13805 6252 13839 6286
rect 13873 6252 13907 6286
rect 13941 6252 13975 6286
rect 14009 6252 14043 6286
rect 14077 6252 14111 6286
rect 14145 6252 14179 6286
rect 14213 6252 14247 6286
rect 14281 6252 14315 6286
rect 14349 6252 14383 6286
rect 14417 6252 14451 6286
rect 14485 6252 14519 6286
rect 14553 6252 14587 6286
rect 14621 6252 14655 6286
rect 14689 6252 14723 6286
rect 14757 6252 14791 6286
rect 14825 6252 14859 6286
rect 14893 6285 15117 6286
rect 14893 6252 14932 6285
rect 44 6251 14932 6252
rect 14966 6251 15000 6285
rect 15034 6251 15068 6285
rect 15102 6251 15117 6285
rect 44 6212 15117 6251
rect 44 6178 68 6212
rect 102 6178 137 6212
rect 171 6178 206 6212
rect 240 6178 275 6212
rect 309 6178 344 6212
rect 378 6178 413 6212
rect 447 6178 482 6212
rect 516 6178 551 6212
rect 585 6178 620 6212
rect 654 6178 689 6212
rect 723 6178 758 6212
rect 792 6178 827 6212
rect 861 6178 896 6212
rect 930 6178 965 6212
rect 999 6178 1034 6212
rect 1068 6178 1103 6212
rect 1137 6178 1172 6212
rect 1206 6178 1241 6212
rect 1275 6178 1310 6212
rect 1344 6178 1379 6212
rect 1413 6178 1448 6212
rect 1482 6178 1517 6212
rect 1551 6178 1586 6212
rect 1620 6178 1655 6212
rect 1689 6178 1724 6212
rect 1758 6178 1793 6212
rect 1827 6178 1862 6212
rect 1896 6178 1931 6212
rect 1965 6178 2000 6212
rect 2034 6178 2069 6212
rect 2103 6178 2138 6212
rect 2172 6178 2207 6212
rect 2241 6178 2276 6212
rect 2310 6178 2345 6212
rect 2379 6178 2414 6212
rect 2448 6178 2483 6212
rect 2517 6178 2551 6212
rect 2585 6178 2619 6212
rect 2653 6178 2687 6212
rect 2721 6178 2755 6212
rect 2789 6178 2823 6212
rect 2857 6178 2891 6212
rect 2925 6178 2959 6212
rect 2993 6178 3027 6212
rect 3061 6178 3095 6212
rect 3129 6178 3163 6212
rect 3197 6178 3231 6212
rect 3265 6178 3299 6212
rect 3333 6178 3367 6212
rect 3401 6178 3435 6212
rect 3469 6178 3503 6212
rect 3537 6178 3571 6212
rect 3605 6178 3639 6212
rect 3673 6178 3707 6212
rect 3741 6178 3775 6212
rect 3809 6178 3843 6212
rect 3877 6178 3911 6212
rect 3945 6178 3979 6212
rect 4013 6178 4047 6212
rect 4081 6178 4115 6212
rect 4149 6178 4183 6212
rect 4217 6178 4251 6212
rect 4285 6178 4319 6212
rect 4353 6178 4387 6212
rect 4421 6178 4455 6212
rect 4489 6178 4523 6212
rect 4557 6178 4591 6212
rect 4625 6178 4659 6212
rect 4693 6178 4727 6212
rect 4761 6178 4795 6212
rect 4829 6178 4863 6212
rect 4897 6178 4931 6212
rect 4965 6178 4999 6212
rect 5033 6178 5067 6212
rect 5101 6178 5135 6212
rect 5169 6178 5203 6212
rect 5237 6178 5271 6212
rect 5305 6178 5339 6212
rect 5373 6178 5407 6212
rect 5441 6178 5475 6212
rect 5509 6178 5543 6212
rect 5577 6178 5611 6212
rect 5645 6178 5679 6212
rect 5713 6178 5747 6212
rect 5781 6178 5815 6212
rect 5849 6178 5883 6212
rect 5917 6178 5951 6212
rect 5985 6178 6019 6212
rect 6053 6178 6087 6212
rect 6121 6178 6155 6212
rect 6189 6178 6223 6212
rect 6257 6178 6291 6212
rect 6325 6178 6359 6212
rect 6393 6178 6427 6212
rect 6461 6178 6495 6212
rect 6529 6178 6563 6212
rect 6597 6178 6631 6212
rect 6665 6178 6699 6212
rect 6733 6178 6767 6212
rect 6801 6178 6835 6212
rect 6869 6178 6903 6212
rect 6937 6178 6971 6212
rect 7005 6178 7039 6212
rect 7073 6178 7107 6212
rect 7141 6178 7175 6212
rect 7209 6178 7243 6212
rect 7277 6178 7311 6212
rect 7345 6178 7379 6212
rect 7413 6178 7447 6212
rect 7481 6178 7515 6212
rect 7549 6178 7583 6212
rect 7617 6178 7651 6212
rect 7685 6178 7719 6212
rect 7753 6178 7787 6212
rect 7821 6178 7855 6212
rect 7889 6178 7923 6212
rect 7957 6178 7991 6212
rect 8025 6178 8059 6212
rect 8093 6178 8127 6212
rect 8161 6178 8195 6212
rect 8229 6178 8263 6212
rect 8297 6178 8331 6212
rect 8365 6178 8399 6212
rect 8433 6178 8467 6212
rect 8501 6178 8535 6212
rect 8569 6178 8603 6212
rect 8637 6178 8671 6212
rect 8705 6178 8739 6212
rect 8773 6178 8807 6212
rect 8841 6178 8875 6212
rect 8909 6178 8943 6212
rect 8977 6178 9011 6212
rect 9045 6178 9079 6212
rect 9113 6178 9147 6212
rect 9181 6178 9215 6212
rect 9249 6178 9283 6212
rect 9317 6178 9351 6212
rect 9385 6178 9419 6212
rect 9453 6178 9487 6212
rect 9521 6178 9555 6212
rect 9589 6178 9623 6212
rect 9657 6178 9691 6212
rect 9725 6178 9759 6212
rect 9793 6178 9827 6212
rect 9861 6178 9895 6212
rect 9929 6178 9963 6212
rect 9997 6178 10031 6212
rect 10065 6178 10099 6212
rect 10133 6178 10167 6212
rect 10201 6178 10235 6212
rect 10269 6178 10303 6212
rect 10337 6178 10371 6212
rect 10405 6178 10439 6212
rect 10473 6178 10507 6212
rect 10541 6178 10575 6212
rect 10609 6178 10643 6212
rect 10677 6178 10711 6212
rect 10745 6178 10779 6212
rect 10813 6178 10847 6212
rect 10881 6178 10915 6212
rect 10949 6178 10983 6212
rect 11017 6178 11051 6212
rect 11085 6178 11119 6212
rect 11153 6178 11187 6212
rect 11221 6178 11255 6212
rect 11289 6178 11323 6212
rect 11357 6178 11391 6212
rect 11425 6178 11459 6212
rect 11493 6178 11527 6212
rect 11561 6178 11595 6212
rect 11629 6178 11663 6212
rect 11697 6178 11731 6212
rect 11765 6178 11799 6212
rect 11833 6178 11867 6212
rect 11901 6178 11935 6212
rect 11969 6178 12003 6212
rect 12037 6178 12071 6212
rect 12105 6178 12139 6212
rect 12173 6178 12207 6212
rect 12241 6178 12275 6212
rect 12309 6178 12343 6212
rect 12377 6178 12411 6212
rect 12445 6178 12479 6212
rect 12513 6178 12547 6212
rect 12581 6178 12615 6212
rect 12649 6178 12683 6212
rect 12717 6178 12751 6212
rect 12785 6178 12819 6212
rect 12853 6178 12887 6212
rect 12921 6178 12955 6212
rect 12989 6178 13023 6212
rect 13057 6178 13091 6212
rect 13125 6178 13159 6212
rect 13193 6178 13227 6212
rect 13261 6178 13295 6212
rect 13329 6178 13363 6212
rect 13397 6178 13431 6212
rect 13465 6178 13499 6212
rect 13533 6178 13567 6212
rect 13601 6178 13635 6212
rect 13669 6178 13703 6212
rect 13737 6178 13771 6212
rect 13805 6178 13839 6212
rect 13873 6178 13907 6212
rect 13941 6178 13975 6212
rect 14009 6178 14043 6212
rect 14077 6178 14111 6212
rect 14145 6178 14179 6212
rect 14213 6178 14247 6212
rect 14281 6178 14315 6212
rect 14349 6178 14383 6212
rect 14417 6178 14451 6212
rect 14485 6178 14519 6212
rect 14553 6178 14587 6212
rect 14621 6178 14655 6212
rect 14689 6178 14723 6212
rect 14757 6178 14791 6212
rect 14825 6178 14859 6212
rect 14893 6210 15117 6212
rect 14893 6178 14932 6210
rect 44 6176 14932 6178
rect 14966 6176 15000 6210
rect 15034 6176 15068 6210
rect 15102 6176 15117 6210
rect 44 6138 15117 6176
rect 44 6104 68 6138
rect 102 6104 137 6138
rect 171 6104 206 6138
rect 240 6104 275 6138
rect 309 6104 344 6138
rect 378 6104 413 6138
rect 447 6104 482 6138
rect 516 6104 551 6138
rect 585 6104 620 6138
rect 654 6104 689 6138
rect 723 6104 758 6138
rect 792 6104 827 6138
rect 861 6104 896 6138
rect 930 6104 965 6138
rect 999 6104 1034 6138
rect 1068 6104 1103 6138
rect 1137 6104 1172 6138
rect 1206 6104 1241 6138
rect 1275 6104 1310 6138
rect 1344 6104 1379 6138
rect 1413 6104 1448 6138
rect 1482 6104 1517 6138
rect 1551 6104 1586 6138
rect 1620 6104 1655 6138
rect 1689 6104 1724 6138
rect 1758 6104 1793 6138
rect 1827 6104 1862 6138
rect 1896 6104 1931 6138
rect 1965 6104 2000 6138
rect 2034 6104 2069 6138
rect 2103 6104 2138 6138
rect 2172 6104 2207 6138
rect 2241 6104 2276 6138
rect 2310 6104 2345 6138
rect 2379 6104 2414 6138
rect 2448 6104 2483 6138
rect 2517 6104 2551 6138
rect 2585 6104 2619 6138
rect 2653 6104 2687 6138
rect 2721 6104 2755 6138
rect 2789 6104 2823 6138
rect 2857 6104 2891 6138
rect 2925 6104 2959 6138
rect 2993 6104 3027 6138
rect 3061 6104 3095 6138
rect 3129 6104 3163 6138
rect 3197 6104 3231 6138
rect 3265 6104 3299 6138
rect 3333 6104 3367 6138
rect 3401 6104 3435 6138
rect 3469 6104 3503 6138
rect 3537 6104 3571 6138
rect 3605 6104 3639 6138
rect 3673 6104 3707 6138
rect 3741 6104 3775 6138
rect 3809 6104 3843 6138
rect 3877 6104 3911 6138
rect 3945 6104 3979 6138
rect 4013 6104 4047 6138
rect 4081 6104 4115 6138
rect 4149 6104 4183 6138
rect 4217 6104 4251 6138
rect 4285 6104 4319 6138
rect 4353 6104 4387 6138
rect 4421 6104 4455 6138
rect 4489 6104 4523 6138
rect 4557 6104 4591 6138
rect 4625 6104 4659 6138
rect 4693 6104 4727 6138
rect 4761 6104 4795 6138
rect 4829 6104 4863 6138
rect 4897 6104 4931 6138
rect 4965 6104 4999 6138
rect 5033 6104 5067 6138
rect 5101 6104 5135 6138
rect 5169 6104 5203 6138
rect 5237 6104 5271 6138
rect 5305 6104 5339 6138
rect 5373 6104 5407 6138
rect 5441 6104 5475 6138
rect 5509 6104 5543 6138
rect 5577 6104 5611 6138
rect 5645 6104 5679 6138
rect 5713 6104 5747 6138
rect 5781 6104 5815 6138
rect 5849 6104 5883 6138
rect 5917 6104 5951 6138
rect 5985 6104 6019 6138
rect 6053 6104 6087 6138
rect 6121 6104 6155 6138
rect 6189 6104 6223 6138
rect 6257 6104 6291 6138
rect 6325 6104 6359 6138
rect 6393 6104 6427 6138
rect 6461 6104 6495 6138
rect 6529 6104 6563 6138
rect 6597 6104 6631 6138
rect 6665 6104 6699 6138
rect 6733 6104 6767 6138
rect 6801 6104 6835 6138
rect 6869 6104 6903 6138
rect 6937 6104 6971 6138
rect 7005 6104 7039 6138
rect 7073 6104 7107 6138
rect 7141 6104 7175 6138
rect 7209 6104 7243 6138
rect 7277 6104 7311 6138
rect 7345 6104 7379 6138
rect 7413 6104 7447 6138
rect 7481 6104 7515 6138
rect 7549 6104 7583 6138
rect 7617 6104 7651 6138
rect 7685 6104 7719 6138
rect 7753 6104 7787 6138
rect 7821 6104 7855 6138
rect 7889 6104 7923 6138
rect 7957 6104 7991 6138
rect 8025 6104 8059 6138
rect 8093 6104 8127 6138
rect 8161 6104 8195 6138
rect 8229 6104 8263 6138
rect 8297 6104 8331 6138
rect 8365 6104 8399 6138
rect 8433 6104 8467 6138
rect 8501 6104 8535 6138
rect 8569 6104 8603 6138
rect 8637 6104 8671 6138
rect 8705 6104 8739 6138
rect 8773 6104 8807 6138
rect 8841 6104 8875 6138
rect 8909 6104 8943 6138
rect 8977 6104 9011 6138
rect 9045 6104 9079 6138
rect 9113 6104 9147 6138
rect 9181 6104 9215 6138
rect 9249 6104 9283 6138
rect 9317 6104 9351 6138
rect 9385 6104 9419 6138
rect 9453 6104 9487 6138
rect 9521 6104 9555 6138
rect 9589 6104 9623 6138
rect 9657 6104 9691 6138
rect 9725 6104 9759 6138
rect 9793 6104 9827 6138
rect 9861 6104 9895 6138
rect 9929 6104 9963 6138
rect 9997 6104 10031 6138
rect 10065 6104 10099 6138
rect 10133 6104 10167 6138
rect 10201 6104 10235 6138
rect 10269 6104 10303 6138
rect 10337 6104 10371 6138
rect 10405 6104 10439 6138
rect 10473 6104 10507 6138
rect 10541 6104 10575 6138
rect 10609 6104 10643 6138
rect 10677 6104 10711 6138
rect 10745 6104 10779 6138
rect 10813 6104 10847 6138
rect 10881 6104 10915 6138
rect 10949 6104 10983 6138
rect 11017 6104 11051 6138
rect 11085 6104 11119 6138
rect 11153 6104 11187 6138
rect 11221 6104 11255 6138
rect 11289 6104 11323 6138
rect 11357 6104 11391 6138
rect 11425 6104 11459 6138
rect 11493 6104 11527 6138
rect 11561 6104 11595 6138
rect 11629 6104 11663 6138
rect 11697 6104 11731 6138
rect 11765 6104 11799 6138
rect 11833 6104 11867 6138
rect 11901 6104 11935 6138
rect 11969 6104 12003 6138
rect 12037 6104 12071 6138
rect 12105 6104 12139 6138
rect 12173 6104 12207 6138
rect 12241 6104 12275 6138
rect 12309 6104 12343 6138
rect 12377 6104 12411 6138
rect 12445 6104 12479 6138
rect 12513 6104 12547 6138
rect 12581 6104 12615 6138
rect 12649 6104 12683 6138
rect 12717 6104 12751 6138
rect 12785 6104 12819 6138
rect 12853 6104 12887 6138
rect 12921 6104 12955 6138
rect 12989 6104 13023 6138
rect 13057 6104 13091 6138
rect 13125 6104 13159 6138
rect 13193 6104 13227 6138
rect 13261 6104 13295 6138
rect 13329 6104 13363 6138
rect 13397 6104 13431 6138
rect 13465 6104 13499 6138
rect 13533 6104 13567 6138
rect 13601 6104 13635 6138
rect 13669 6104 13703 6138
rect 13737 6104 13771 6138
rect 13805 6104 13839 6138
rect 13873 6104 13907 6138
rect 13941 6104 13975 6138
rect 14009 6104 14043 6138
rect 14077 6104 14111 6138
rect 14145 6104 14179 6138
rect 14213 6104 14247 6138
rect 14281 6104 14315 6138
rect 14349 6104 14383 6138
rect 14417 6104 14451 6138
rect 14485 6104 14519 6138
rect 14553 6104 14587 6138
rect 14621 6104 14655 6138
rect 14689 6104 14723 6138
rect 14757 6104 14791 6138
rect 14825 6104 14859 6138
rect 14893 6135 15117 6138
rect 14893 6104 14932 6135
rect 44 6101 14932 6104
rect 14966 6101 15000 6135
rect 15034 6101 15068 6135
rect 15102 6101 15117 6135
rect 44 6060 15117 6101
rect 44 6051 14932 6060
rect 14917 6026 14932 6051
rect 14966 6026 15000 6060
rect 15034 6026 15068 6060
rect 15102 6026 15117 6060
rect 14917 5988 15117 6026
rect 14977 5954 15117 5988
rect 14977 4628 15000 5954
rect 15102 4628 15117 5954
rect 14977 4593 15117 4628
rect 14977 4559 15000 4593
rect 15034 4559 15068 4593
rect 15102 4559 15117 4593
rect 14977 4524 15117 4559
rect 14977 4490 15000 4524
rect 15034 4490 15068 4524
rect 15102 4490 15117 4524
rect 14977 4455 15117 4490
rect 14977 4421 15000 4455
rect 15034 4421 15068 4455
rect 15102 4421 15117 4455
rect 14977 4386 15117 4421
rect 14977 4352 15000 4386
rect 15034 4352 15068 4386
rect 15102 4352 15117 4386
rect 14977 4317 15117 4352
rect 14977 4283 15000 4317
rect 15034 4283 15068 4317
rect 15102 4283 15117 4317
rect 14977 4248 15117 4283
rect 14977 4214 15000 4248
rect 15034 4214 15068 4248
rect 15102 4214 15117 4248
rect 14977 4179 15117 4214
rect 14977 4145 15000 4179
rect 15034 4145 15068 4179
rect 15102 4145 15117 4179
rect 14977 4110 15117 4145
rect 14977 4076 15000 4110
rect 15034 4076 15068 4110
rect 15102 4076 15117 4110
rect 14977 4041 15117 4076
rect 14977 4007 15000 4041
rect 15034 4007 15068 4041
rect 15102 4007 15117 4041
rect 14977 3972 15117 4007
rect 14977 3938 15000 3972
rect 15034 3938 15068 3972
rect 15102 3938 15117 3972
rect 14977 3903 15117 3938
rect 14977 3869 15000 3903
rect 15034 3869 15068 3903
rect 15102 3869 15117 3903
rect 14977 3834 15117 3869
rect 14977 3800 15000 3834
rect 15034 3800 15068 3834
rect 15102 3800 15117 3834
rect 14977 3765 15117 3800
rect 14977 3731 15000 3765
rect 15034 3731 15068 3765
rect 15102 3731 15117 3765
rect 14977 3696 15117 3731
rect 14977 3662 15000 3696
rect 15034 3662 15068 3696
rect 15102 3662 15117 3696
rect 14977 3627 15117 3662
rect 14977 3593 15000 3627
rect 15034 3593 15068 3627
rect 15102 3593 15117 3627
rect 14977 3558 15117 3593
rect 14977 3524 15000 3558
rect 15034 3524 15068 3558
rect 15102 3524 15117 3558
rect 14977 3489 15117 3524
rect 14977 3455 15000 3489
rect 15034 3455 15068 3489
rect 15102 3455 15117 3489
rect 14977 3420 15117 3455
rect 14977 3386 15000 3420
rect 15034 3386 15068 3420
rect 15102 3386 15117 3420
rect 14977 3351 15117 3386
rect 14977 3317 15000 3351
rect 15034 3317 15068 3351
rect 15102 3317 15117 3351
rect 14977 3282 15117 3317
rect 14977 3248 15000 3282
rect 15034 3248 15068 3282
rect 15102 3248 15117 3282
rect 14977 3213 15117 3248
rect 14977 3179 15000 3213
rect 15034 3179 15068 3213
rect 15102 3179 15117 3213
rect 14977 3144 15117 3179
rect 14977 3110 15000 3144
rect 15034 3110 15068 3144
rect 15102 3110 15117 3144
rect 14977 3075 15117 3110
rect 14977 3041 15000 3075
rect 15034 3041 15068 3075
rect 15102 3041 15117 3075
rect 14977 3006 15117 3041
rect 14977 2972 15000 3006
rect 15034 2972 15068 3006
rect 15102 2972 15117 3006
rect 14977 2937 15117 2972
rect 14977 2903 15000 2937
rect 15034 2903 15068 2937
rect 15102 2903 15117 2937
rect 14977 2868 15117 2903
rect 14977 2834 15000 2868
rect 15034 2834 15068 2868
rect 15102 2834 15117 2868
rect 14977 2799 15117 2834
rect 14977 2765 15000 2799
rect 15034 2765 15068 2799
rect 15102 2765 15117 2799
rect 14977 2730 15117 2765
rect 14977 2696 15000 2730
rect 15034 2696 15068 2730
rect 15102 2696 15117 2730
rect 14977 2661 15117 2696
rect 14977 2627 15000 2661
rect 15034 2627 15068 2661
rect 15102 2627 15117 2661
rect 14977 2592 15117 2627
rect 14977 2558 15000 2592
rect 15034 2558 15068 2592
rect 15102 2558 15117 2592
rect 14977 2523 15117 2558
rect 14977 2489 15000 2523
rect 15034 2489 15068 2523
rect 15102 2489 15117 2523
rect 14977 2454 15117 2489
rect 14977 2420 15000 2454
rect 15034 2420 15068 2454
rect 15102 2420 15117 2454
rect 14977 2385 15117 2420
rect 14977 2351 15000 2385
rect 15034 2351 15068 2385
rect 15102 2351 15117 2385
rect 14977 2316 15117 2351
rect 14977 2282 15000 2316
rect 15034 2282 15068 2316
rect 15102 2282 15117 2316
rect 14977 2247 15117 2282
rect 14977 2213 15000 2247
rect 15034 2213 15068 2247
rect 15102 2213 15117 2247
rect 14977 2178 15117 2213
rect 14977 2144 15000 2178
rect 15034 2144 15068 2178
rect 15102 2144 15117 2178
rect 14977 2109 15117 2144
rect 14977 2075 15000 2109
rect 15034 2075 15068 2109
rect 15102 2075 15117 2109
rect 14977 2040 15117 2075
rect 14977 2006 15000 2040
rect 15034 2006 15068 2040
rect 15102 2006 15117 2040
rect 14977 1971 15117 2006
rect 14977 1937 15000 1971
rect 15034 1937 15068 1971
rect 15102 1937 15117 1971
rect 14977 1902 15117 1937
rect 14977 1868 15000 1902
rect 15034 1868 15068 1902
rect 15102 1868 15117 1902
rect 14977 1833 15117 1868
rect 14977 1799 15000 1833
rect 15034 1799 15068 1833
rect 15102 1799 15117 1833
rect 14977 1764 15117 1799
rect 14977 1730 15000 1764
rect 15034 1730 15068 1764
rect 15102 1730 15117 1764
rect 14977 1695 15117 1730
rect 14977 1661 15000 1695
rect 15034 1661 15068 1695
rect 15102 1661 15117 1695
rect 14977 1626 15117 1661
rect 14977 1592 15000 1626
rect 15034 1592 15068 1626
rect 15102 1592 15117 1626
rect 14977 1557 15117 1592
rect 14977 1523 15000 1557
rect 15034 1523 15068 1557
rect 15102 1523 15117 1557
rect 14977 1488 15117 1523
rect 14977 1454 15000 1488
rect 15034 1454 15068 1488
rect 15102 1454 15117 1488
rect 14977 1419 15117 1454
rect 14977 1385 15000 1419
rect 15034 1385 15068 1419
rect 15102 1385 15117 1419
rect 14977 1350 15117 1385
rect 14977 1316 15000 1350
rect 15034 1316 15068 1350
rect 15102 1316 15117 1350
rect 7044 1282 14917 1288
rect 14977 1282 15117 1316
rect 7018 1257 15117 1282
rect 7018 1251 7068 1257
rect 7022 1223 7068 1251
rect 7102 1223 7137 1257
rect 7171 1223 7206 1257
rect 7240 1223 7275 1257
rect 7309 1223 7344 1257
rect 7378 1223 7413 1257
rect 7447 1223 7482 1257
rect 7516 1223 7551 1257
rect 7585 1223 7620 1257
rect 7654 1223 7689 1257
rect 7723 1223 7758 1257
rect 7792 1223 7827 1257
rect 7861 1223 7896 1257
rect 7930 1223 7965 1257
rect 7999 1223 8034 1257
rect 8068 1223 8103 1257
rect 8137 1223 8172 1257
rect 8206 1223 8241 1257
rect 8275 1223 8310 1257
rect 8344 1223 8379 1257
rect 8413 1223 8448 1257
rect 8482 1223 8517 1257
rect 8551 1223 8586 1257
rect 8620 1223 8655 1257
rect 8689 1223 8724 1257
rect 8758 1223 8793 1257
rect 8827 1223 8862 1257
rect 8896 1223 8931 1257
rect 8965 1223 9000 1257
rect 9034 1223 9069 1257
rect 9103 1223 9138 1257
rect 9172 1223 9207 1257
rect 9241 1223 9276 1257
rect 9310 1223 9345 1257
rect 9379 1223 9414 1257
rect 9448 1223 9483 1257
rect 9517 1223 9552 1257
rect 9586 1223 9621 1257
rect 9655 1223 9690 1257
rect 9724 1223 9759 1257
rect 7022 1189 9759 1223
rect 7022 1155 7068 1189
rect 7102 1155 7137 1189
rect 7171 1155 7206 1189
rect 7240 1155 7275 1189
rect 7309 1155 7344 1189
rect 7378 1155 7413 1189
rect 7447 1155 7482 1189
rect 7516 1155 7551 1189
rect 7585 1155 7620 1189
rect 7654 1155 7689 1189
rect 7723 1155 7758 1189
rect 7792 1155 7827 1189
rect 7861 1155 7896 1189
rect 7930 1155 7965 1189
rect 7999 1155 8034 1189
rect 8068 1155 8103 1189
rect 8137 1155 8172 1189
rect 8206 1155 8241 1189
rect 8275 1155 8310 1189
rect 8344 1155 8379 1189
rect 8413 1155 8448 1189
rect 8482 1155 8517 1189
rect 8551 1155 8586 1189
rect 8620 1155 8655 1189
rect 8689 1155 8724 1189
rect 8758 1155 8793 1189
rect 8827 1155 8862 1189
rect 8896 1155 8931 1189
rect 8965 1155 9000 1189
rect 9034 1155 9069 1189
rect 9103 1155 9138 1189
rect 9172 1155 9207 1189
rect 9241 1155 9276 1189
rect 9310 1155 9345 1189
rect 9379 1155 9414 1189
rect 9448 1155 9483 1189
rect 9517 1155 9552 1189
rect 9586 1155 9621 1189
rect 9655 1155 9690 1189
rect 9724 1155 9759 1189
rect 7022 1121 9759 1155
rect 7022 1087 7068 1121
rect 7102 1087 7137 1121
rect 7171 1087 7206 1121
rect 7240 1087 7275 1121
rect 7309 1087 7344 1121
rect 7378 1087 7413 1121
rect 7447 1087 7482 1121
rect 7516 1087 7551 1121
rect 7585 1087 7620 1121
rect 7654 1087 7689 1121
rect 7723 1087 7758 1121
rect 7792 1087 7827 1121
rect 7861 1087 7896 1121
rect 7930 1087 7965 1121
rect 7999 1087 8034 1121
rect 8068 1087 8103 1121
rect 8137 1087 8172 1121
rect 8206 1087 8241 1121
rect 8275 1087 8310 1121
rect 8344 1087 8379 1121
rect 8413 1087 8448 1121
rect 8482 1087 8517 1121
rect 8551 1087 8586 1121
rect 8620 1087 8655 1121
rect 8689 1087 8724 1121
rect 8758 1087 8793 1121
rect 8827 1087 8862 1121
rect 8896 1087 8931 1121
rect 8965 1087 9000 1121
rect 9034 1087 9069 1121
rect 9103 1087 9138 1121
rect 9172 1087 9207 1121
rect 9241 1087 9276 1121
rect 9310 1087 9345 1121
rect 9379 1087 9414 1121
rect 9448 1087 9483 1121
rect 9517 1087 9552 1121
rect 9586 1087 9621 1121
rect 9655 1087 9690 1121
rect 9724 1087 9759 1121
rect 7022 1053 9759 1087
rect 7022 1019 7068 1053
rect 7102 1019 7137 1053
rect 7171 1019 7206 1053
rect 7240 1019 7275 1053
rect 7309 1019 7344 1053
rect 7378 1019 7413 1053
rect 7447 1019 7482 1053
rect 7516 1019 7551 1053
rect 7585 1019 7620 1053
rect 7654 1019 7689 1053
rect 7723 1019 7758 1053
rect 7792 1019 7827 1053
rect 7861 1019 7896 1053
rect 7930 1019 7965 1053
rect 7999 1019 8034 1053
rect 8068 1019 8103 1053
rect 8137 1019 8172 1053
rect 8206 1019 8241 1053
rect 8275 1019 8310 1053
rect 8344 1019 8379 1053
rect 8413 1019 8448 1053
rect 8482 1019 8517 1053
rect 8551 1019 8586 1053
rect 8620 1019 8655 1053
rect 8689 1019 8724 1053
rect 8758 1019 8793 1053
rect 8827 1019 8862 1053
rect 8896 1019 8931 1053
rect 8965 1019 9000 1053
rect 9034 1019 9069 1053
rect 9103 1019 9138 1053
rect 9172 1019 9207 1053
rect 9241 1019 9276 1053
rect 9310 1019 9345 1053
rect 9379 1019 9414 1053
rect 9448 1019 9483 1053
rect 9517 1019 9552 1053
rect 9586 1019 9621 1053
rect 9655 1019 9690 1053
rect 9724 1019 9759 1053
rect 14893 1244 15117 1257
rect 14893 1210 14932 1244
rect 14966 1210 15000 1244
rect 15034 1210 15068 1244
rect 15102 1210 15117 1244
rect 14893 1172 15117 1210
rect 14893 1138 14932 1172
rect 14966 1138 15000 1172
rect 15034 1138 15068 1172
rect 15102 1138 15117 1172
rect 14893 1100 15117 1138
rect 14893 1066 14932 1100
rect 14966 1066 15000 1100
rect 15034 1066 15068 1100
rect 15102 1066 15117 1100
rect 14893 1028 15117 1066
rect 14893 1019 14932 1028
rect 7022 994 14932 1019
rect 14966 994 15000 1028
rect 15034 994 15068 1028
rect 15102 994 15117 1028
rect 7022 988 15117 994
rect 7022 947 7754 988
rect 7022 913 7067 947
rect 7101 913 7137 947
rect 7171 913 7207 947
rect 7241 913 7277 947
rect 7311 913 7347 947
rect 7381 913 7417 947
rect 7451 913 7487 947
rect 7521 913 7557 947
rect 7591 913 7627 947
rect 7661 913 7696 947
rect 7730 913 7754 947
rect 7022 875 7754 913
rect 7022 841 7067 875
rect 7101 841 7137 875
rect 7171 841 7207 875
rect 7241 841 7277 875
rect 7311 841 7347 875
rect 7381 841 7417 875
rect 7451 841 7487 875
rect 7521 841 7557 875
rect 7591 841 7627 875
rect 7661 841 7696 875
rect 7730 841 7754 875
rect 7022 803 7754 841
rect 7022 769 7067 803
rect 7101 769 7137 803
rect 7171 769 7207 803
rect 7241 769 7277 803
rect 7311 769 7347 803
rect 7381 769 7417 803
rect 7451 769 7487 803
rect 7521 769 7557 803
rect 7591 769 7627 803
rect 7661 769 7696 803
rect 7730 769 7754 803
rect 7022 731 7754 769
rect 7022 697 7067 731
rect 7101 697 7137 731
rect 7171 697 7207 731
rect 7241 697 7277 731
rect 7311 697 7347 731
rect 7381 697 7417 731
rect 7451 697 7487 731
rect 7521 697 7557 731
rect 7591 697 7627 731
rect 7661 697 7696 731
rect 7730 697 7754 731
rect 7022 659 7754 697
rect 7022 625 7067 659
rect 7101 625 7137 659
rect 7171 625 7207 659
rect 7241 625 7277 659
rect 7311 625 7347 659
rect 7381 625 7417 659
rect 7451 625 7487 659
rect 7521 625 7557 659
rect 7591 625 7627 659
rect 7661 625 7696 659
rect 7730 625 7754 659
rect 7022 587 7754 625
rect 7022 553 7067 587
rect 7101 553 7137 587
rect 7171 553 7207 587
rect 7241 553 7277 587
rect 7311 553 7347 587
rect 7381 553 7417 587
rect 7451 553 7487 587
rect 7521 553 7557 587
rect 7591 553 7627 587
rect 7661 553 7696 587
rect 7730 553 7754 587
rect 7022 515 7754 553
rect 7022 481 7067 515
rect 7101 481 7137 515
rect 7171 481 7207 515
rect 7241 481 7277 515
rect 7311 481 7347 515
rect 7381 481 7417 515
rect 7451 481 7487 515
rect 7521 481 7557 515
rect 7591 481 7627 515
rect 7661 481 7696 515
rect 7730 481 7754 515
rect 7022 443 7754 481
rect 7022 409 7067 443
rect 7101 409 7137 443
rect 7171 409 7207 443
rect 7241 409 7277 443
rect 7311 409 7347 443
rect 7381 409 7417 443
rect 7451 409 7487 443
rect 7521 409 7557 443
rect 7591 409 7627 443
rect 7661 409 7696 443
rect 7730 409 7754 443
rect 7022 369 7754 409
rect 9687 956 15117 988
rect 9687 955 14932 956
rect 9687 947 11680 955
rect 9687 913 9711 947
rect 9745 913 9781 947
rect 9815 913 9851 947
rect 9885 913 9921 947
rect 9955 913 9991 947
rect 10025 913 10061 947
rect 10095 913 10131 947
rect 10165 913 10201 947
rect 10235 913 10271 947
rect 10305 913 10341 947
rect 10375 913 10411 947
rect 10445 913 10481 947
rect 10515 913 10551 947
rect 10585 913 10621 947
rect 10655 913 10691 947
rect 10725 913 10761 947
rect 10795 913 10831 947
rect 10865 913 10901 947
rect 10935 913 10971 947
rect 11005 913 11041 947
rect 11075 913 11111 947
rect 11145 913 11181 947
rect 11215 913 11251 947
rect 11285 913 11321 947
rect 11355 913 11391 947
rect 11425 913 11460 947
rect 11494 913 11529 947
rect 11563 913 11598 947
rect 11632 921 11680 947
rect 11714 921 11750 955
rect 11784 921 11820 955
rect 11854 921 11890 955
rect 11924 921 11960 955
rect 11994 921 12030 955
rect 12064 921 12099 955
rect 12133 921 12168 955
rect 12202 921 12237 955
rect 12271 921 12306 955
rect 12340 921 12375 955
rect 12409 921 12444 955
rect 12478 921 12513 955
rect 12547 921 12582 955
rect 12616 921 12651 955
rect 12685 921 12720 955
rect 12754 921 12789 955
rect 12823 921 12858 955
rect 12892 921 12927 955
rect 12961 921 12996 955
rect 13030 921 13065 955
rect 13099 921 13134 955
rect 13168 921 13203 955
rect 13237 921 13272 955
rect 13306 921 13341 955
rect 13375 921 13410 955
rect 13444 921 13479 955
rect 13513 921 13548 955
rect 13582 921 13617 955
rect 13651 921 13686 955
rect 13720 921 13755 955
rect 13789 921 13824 955
rect 13858 921 13893 955
rect 13927 921 13962 955
rect 13996 921 14031 955
rect 14065 921 14100 955
rect 14134 921 14169 955
rect 14203 921 14238 955
rect 14272 921 14307 955
rect 14341 921 14376 955
rect 14410 921 14445 955
rect 14479 921 14514 955
rect 14548 921 14583 955
rect 14617 921 14652 955
rect 14686 921 14721 955
rect 14755 921 14790 955
rect 14824 921 14859 955
rect 14893 922 14932 955
rect 14966 922 15000 956
rect 15034 922 15068 956
rect 15102 922 15117 956
rect 14893 921 15117 922
rect 11632 913 15117 921
rect 9687 884 15117 913
rect 9687 875 14932 884
rect 9687 841 9711 875
rect 9745 841 9781 875
rect 9815 841 9851 875
rect 9885 841 9921 875
rect 9955 841 9991 875
rect 10025 841 10061 875
rect 10095 841 10131 875
rect 10165 841 10201 875
rect 10235 841 10271 875
rect 10305 841 10341 875
rect 10375 841 10411 875
rect 10445 841 10481 875
rect 10515 841 10551 875
rect 10585 841 10621 875
rect 10655 841 10691 875
rect 10725 841 10761 875
rect 10795 841 10831 875
rect 10865 841 10901 875
rect 10935 841 10971 875
rect 11005 841 11041 875
rect 11075 841 11111 875
rect 11145 841 11181 875
rect 11215 841 11251 875
rect 11285 841 11321 875
rect 11355 841 11391 875
rect 11425 841 11460 875
rect 11494 841 11529 875
rect 11563 841 11598 875
rect 11632 841 11680 875
rect 11714 841 11750 875
rect 11784 841 11820 875
rect 11854 841 11890 875
rect 11924 841 11960 875
rect 11994 841 12030 875
rect 12064 841 12099 875
rect 12133 841 12168 875
rect 12202 841 12237 875
rect 12271 841 12306 875
rect 12340 841 12375 875
rect 12409 841 12444 875
rect 12478 841 12513 875
rect 12547 841 12582 875
rect 12616 841 12651 875
rect 12685 841 12720 875
rect 12754 841 12789 875
rect 12823 841 12858 875
rect 12892 841 12927 875
rect 12961 841 12996 875
rect 13030 841 13065 875
rect 13099 841 13134 875
rect 13168 841 13203 875
rect 13237 841 13272 875
rect 13306 841 13341 875
rect 13375 841 13410 875
rect 13444 841 13479 875
rect 13513 841 13548 875
rect 13582 841 13617 875
rect 13651 841 13686 875
rect 13720 841 13755 875
rect 13789 841 13824 875
rect 13858 841 13893 875
rect 13927 841 13962 875
rect 13996 841 14031 875
rect 14065 841 14100 875
rect 14134 841 14169 875
rect 14203 841 14238 875
rect 14272 841 14307 875
rect 14341 841 14376 875
rect 14410 841 14445 875
rect 14479 841 14514 875
rect 14548 841 14583 875
rect 14617 841 14652 875
rect 14686 841 14721 875
rect 14755 841 14790 875
rect 14824 841 14859 875
rect 14893 850 14932 875
rect 14966 850 15000 884
rect 15034 850 15068 884
rect 15102 850 15117 884
rect 14893 841 15117 850
rect 9687 812 15117 841
rect 9687 803 14932 812
rect 9687 769 9711 803
rect 9745 769 9781 803
rect 9815 769 9851 803
rect 9885 769 9921 803
rect 9955 769 9991 803
rect 10025 769 10061 803
rect 10095 769 10131 803
rect 10165 769 10201 803
rect 10235 769 10271 803
rect 10305 769 10341 803
rect 10375 769 10411 803
rect 10445 769 10481 803
rect 10515 769 10551 803
rect 10585 769 10621 803
rect 10655 769 10691 803
rect 10725 769 10761 803
rect 10795 769 10831 803
rect 10865 769 10901 803
rect 10935 769 10971 803
rect 11005 769 11041 803
rect 11075 769 11111 803
rect 11145 769 11181 803
rect 11215 769 11251 803
rect 11285 769 11321 803
rect 11355 769 11391 803
rect 11425 769 11460 803
rect 11494 769 11529 803
rect 11563 769 11598 803
rect 11632 795 14932 803
rect 11632 769 11680 795
rect 9687 761 11680 769
rect 11714 761 11750 795
rect 11784 761 11820 795
rect 11854 761 11890 795
rect 11924 761 11960 795
rect 11994 761 12030 795
rect 12064 761 12099 795
rect 12133 761 12168 795
rect 12202 761 12237 795
rect 12271 761 12306 795
rect 12340 761 12375 795
rect 12409 761 12444 795
rect 12478 761 12513 795
rect 12547 761 12582 795
rect 12616 761 12651 795
rect 12685 761 12720 795
rect 12754 761 12789 795
rect 12823 761 12858 795
rect 12892 761 12927 795
rect 12961 761 12996 795
rect 13030 761 13065 795
rect 13099 761 13134 795
rect 13168 761 13203 795
rect 13237 761 13272 795
rect 13306 761 13341 795
rect 13375 761 13410 795
rect 13444 761 13479 795
rect 13513 761 13548 795
rect 13582 761 13617 795
rect 13651 761 13686 795
rect 13720 761 13755 795
rect 13789 761 13824 795
rect 13858 761 13893 795
rect 13927 761 13962 795
rect 13996 761 14031 795
rect 14065 761 14100 795
rect 14134 761 14169 795
rect 14203 761 14238 795
rect 14272 761 14307 795
rect 14341 761 14376 795
rect 14410 761 14445 795
rect 14479 761 14514 795
rect 14548 761 14583 795
rect 14617 761 14652 795
rect 14686 761 14721 795
rect 14755 761 14790 795
rect 14824 761 14859 795
rect 14893 778 14932 795
rect 14966 778 15000 812
rect 15034 778 15068 812
rect 15102 778 15117 812
rect 14893 761 15117 778
rect 9687 740 15117 761
rect 9687 731 14932 740
rect 9687 697 9711 731
rect 9745 697 9781 731
rect 9815 697 9851 731
rect 9885 697 9921 731
rect 9955 697 9991 731
rect 10025 697 10061 731
rect 10095 697 10131 731
rect 10165 697 10201 731
rect 10235 697 10271 731
rect 10305 697 10341 731
rect 10375 697 10411 731
rect 10445 697 10481 731
rect 10515 697 10551 731
rect 10585 697 10621 731
rect 10655 697 10691 731
rect 10725 697 10761 731
rect 10795 697 10831 731
rect 10865 697 10901 731
rect 10935 697 10971 731
rect 11005 697 11041 731
rect 11075 697 11111 731
rect 11145 697 11181 731
rect 11215 697 11251 731
rect 11285 697 11321 731
rect 11355 697 11391 731
rect 11425 697 11460 731
rect 11494 697 11529 731
rect 11563 697 11598 731
rect 11632 728 14932 731
rect 11632 697 11656 728
rect 9687 659 11656 697
rect 9687 625 9711 659
rect 9745 625 9781 659
rect 9815 625 9851 659
rect 9885 625 9921 659
rect 9955 625 9991 659
rect 10025 625 10061 659
rect 10095 625 10131 659
rect 10165 625 10201 659
rect 10235 625 10271 659
rect 10305 625 10341 659
rect 10375 625 10411 659
rect 10445 625 10481 659
rect 10515 625 10551 659
rect 10585 625 10621 659
rect 10655 625 10691 659
rect 10725 625 10761 659
rect 10795 625 10831 659
rect 10865 625 10901 659
rect 10935 625 10971 659
rect 11005 625 11041 659
rect 11075 625 11111 659
rect 11145 625 11181 659
rect 11215 625 11251 659
rect 11285 625 11321 659
rect 11355 625 11391 659
rect 11425 625 11460 659
rect 11494 625 11529 659
rect 11563 625 11598 659
rect 11632 625 11656 659
rect 9687 587 11656 625
rect 9687 553 9711 587
rect 9745 553 9781 587
rect 9815 553 9851 587
rect 9885 553 9921 587
rect 9955 553 9991 587
rect 10025 553 10061 587
rect 10095 553 10131 587
rect 10165 553 10201 587
rect 10235 553 10271 587
rect 10305 553 10341 587
rect 10375 553 10411 587
rect 10445 553 10481 587
rect 10515 553 10551 587
rect 10585 553 10621 587
rect 10655 553 10691 587
rect 10725 553 10761 587
rect 10795 553 10831 587
rect 10865 553 10901 587
rect 10935 553 10971 587
rect 11005 553 11041 587
rect 11075 553 11111 587
rect 11145 553 11181 587
rect 11215 553 11251 587
rect 11285 553 11321 587
rect 11355 553 11391 587
rect 11425 553 11460 587
rect 11494 553 11529 587
rect 11563 553 11598 587
rect 11632 553 11656 587
rect 9687 515 11656 553
rect 9687 481 9711 515
rect 9745 481 9781 515
rect 9815 481 9851 515
rect 9885 481 9921 515
rect 9955 481 9991 515
rect 10025 481 10061 515
rect 10095 481 10131 515
rect 10165 481 10201 515
rect 10235 481 10271 515
rect 10305 481 10341 515
rect 10375 481 10411 515
rect 10445 481 10481 515
rect 10515 481 10551 515
rect 10585 481 10621 515
rect 10655 481 10691 515
rect 10725 481 10761 515
rect 10795 481 10831 515
rect 10865 481 10901 515
rect 10935 481 10971 515
rect 11005 481 11041 515
rect 11075 481 11111 515
rect 11145 481 11181 515
rect 11215 481 11251 515
rect 11285 481 11321 515
rect 11355 481 11391 515
rect 11425 481 11460 515
rect 11494 481 11529 515
rect 11563 481 11598 515
rect 11632 481 11656 515
rect 9687 443 11656 481
rect 9687 409 9711 443
rect 9745 409 9781 443
rect 9815 409 9851 443
rect 9885 409 9921 443
rect 9955 409 9991 443
rect 10025 409 10061 443
rect 10095 409 10131 443
rect 10165 409 10201 443
rect 10235 409 10271 443
rect 10305 409 10341 443
rect 10375 409 10411 443
rect 10445 409 10481 443
rect 10515 409 10551 443
rect 10585 409 10621 443
rect 10655 409 10691 443
rect 10725 409 10761 443
rect 10795 409 10831 443
rect 10865 409 10901 443
rect 10935 409 10971 443
rect 11005 409 11041 443
rect 11075 409 11111 443
rect 11145 409 11181 443
rect 11215 409 11251 443
rect 11285 409 11321 443
rect 11355 409 11391 443
rect 11425 409 11460 443
rect 11494 409 11529 443
rect 11563 409 11598 443
rect 11632 409 11656 443
rect 9687 369 11656 409
rect 14465 706 14932 728
rect 14966 706 15000 740
rect 15034 706 15068 740
rect 15102 706 15117 740
rect 14465 695 15117 706
rect 14499 661 14543 695
rect 14577 661 14621 695
rect 14655 661 14698 695
rect 14732 661 14775 695
rect 14809 661 14852 695
rect 14886 668 15117 695
rect 14886 661 14932 668
rect 14465 634 14932 661
rect 14966 634 15000 668
rect 15034 634 15068 668
rect 15102 634 15117 668
rect 14465 609 15117 634
rect 14499 575 14543 609
rect 14577 575 14621 609
rect 14655 575 14698 609
rect 14732 575 14775 609
rect 14809 575 14852 609
rect 14886 596 15117 609
rect 14886 575 14932 596
rect 14465 562 14932 575
rect 14966 562 15000 596
rect 15034 562 15068 596
rect 15102 562 15117 596
rect 14465 524 15117 562
rect 14465 523 14932 524
rect 14499 489 14543 523
rect 14577 489 14621 523
rect 14655 489 14698 523
rect 14732 489 14775 523
rect 14809 489 14852 523
rect 14886 490 14932 523
rect 14966 490 15000 524
rect 15034 490 15068 524
rect 15102 490 15117 524
rect 14886 489 15117 490
rect 14465 452 15117 489
rect 14465 437 14932 452
rect 14499 403 14543 437
rect 14577 403 14621 437
rect 14655 403 14698 437
rect 14732 403 14775 437
rect 14809 403 14852 437
rect 14886 418 14932 437
rect 14966 418 15000 452
rect 15034 418 15068 452
rect 15102 418 15117 452
rect 14886 403 15117 418
rect 14465 380 15117 403
rect 14465 369 14932 380
rect 7022 367 14932 369
rect 7022 333 7056 367
rect 7090 333 7125 367
rect 7159 333 7194 367
rect 7228 333 7263 367
rect 7297 333 7332 367
rect 7366 333 7401 367
rect 7435 333 7470 367
rect 7504 333 7539 367
rect 7573 333 7608 367
rect 7642 333 7677 367
rect 7711 333 7746 367
rect 7780 333 7815 367
rect 7849 333 7884 367
rect 7918 333 7953 367
rect 7987 333 8022 367
rect 8056 333 8091 367
rect 8125 333 8160 367
rect 8194 333 8229 367
rect 8263 333 8298 367
rect 8332 333 8367 367
rect 8401 333 8436 367
rect 8470 333 8505 367
rect 8539 333 8574 367
rect 8608 333 8643 367
rect 8677 333 8712 367
rect 8746 333 8781 367
rect 8815 333 8850 367
rect 8884 333 8919 367
rect 8953 333 8988 367
rect 9022 333 9057 367
rect 9091 333 9126 367
rect 9160 333 9195 367
rect 9229 333 9264 367
rect 9298 333 9333 367
rect 9367 333 9402 367
rect 9436 333 9471 367
rect 9505 333 9540 367
rect 9574 333 9609 367
rect 9643 333 9678 367
rect 9712 333 9747 367
rect 9781 333 9816 367
rect 9850 333 9885 367
rect 9919 333 9954 367
rect 9988 333 10023 367
rect 10057 333 10092 367
rect 10126 333 10161 367
rect 10195 333 10230 367
rect 10264 333 10299 367
rect 10333 333 10368 367
rect 10402 333 10437 367
rect 10471 333 10506 367
rect 10540 333 10575 367
rect 10609 333 10643 367
rect 10677 333 10711 367
rect 10745 333 10779 367
rect 10813 333 10847 367
rect 10881 333 10915 367
rect 10949 333 10983 367
rect 11017 333 11051 367
rect 11085 333 11119 367
rect 11153 333 11187 367
rect 11221 333 11255 367
rect 11289 333 11323 367
rect 11357 333 11391 367
rect 11425 333 11459 367
rect 11493 333 11527 367
rect 11561 333 11595 367
rect 11629 333 11663 367
rect 11697 333 11731 367
rect 11765 333 11799 367
rect 11833 333 11867 367
rect 11901 333 11935 367
rect 11969 333 12003 367
rect 12037 333 12071 367
rect 12105 333 12139 367
rect 12173 333 12207 367
rect 12241 333 12275 367
rect 12309 333 12343 367
rect 12377 333 12411 367
rect 12445 333 12479 367
rect 12513 333 12547 367
rect 12581 333 12615 367
rect 12649 333 12683 367
rect 12717 333 12751 367
rect 12785 333 12819 367
rect 12853 333 12887 367
rect 12921 333 12955 367
rect 12989 333 13023 367
rect 13057 333 13091 367
rect 13125 333 13159 367
rect 13193 333 13227 367
rect 13261 333 13295 367
rect 13329 333 13363 367
rect 13397 333 13431 367
rect 13465 333 13499 367
rect 13533 333 13567 367
rect 13601 333 13635 367
rect 13669 333 13703 367
rect 13737 333 13771 367
rect 13805 333 13839 367
rect 13873 333 13907 367
rect 13941 333 13975 367
rect 14009 333 14043 367
rect 14077 333 14111 367
rect 14145 333 14179 367
rect 14213 333 14247 367
rect 14281 333 14315 367
rect 14349 333 14383 367
rect 14417 333 14451 367
rect 14485 333 14519 367
rect 14553 333 14587 367
rect 14621 333 14655 367
rect 14689 333 14723 367
rect 14757 333 14791 367
rect 14825 333 14859 367
rect 14893 346 14932 367
rect 14966 346 15000 380
rect 15034 346 15068 380
rect 15102 346 15117 380
rect 14893 333 15117 346
rect 7022 308 15117 333
rect 7022 289 14932 308
rect 7022 255 7056 289
rect 7090 255 7125 289
rect 7159 255 7194 289
rect 7228 255 7263 289
rect 7297 255 7332 289
rect 7366 255 7401 289
rect 7435 255 7470 289
rect 7504 255 7539 289
rect 7573 255 7608 289
rect 7642 255 7677 289
rect 7711 255 7746 289
rect 7780 255 7815 289
rect 7849 255 7884 289
rect 7918 255 7953 289
rect 7987 255 8022 289
rect 8056 255 8091 289
rect 8125 255 8160 289
rect 8194 255 8229 289
rect 8263 255 8298 289
rect 8332 255 8367 289
rect 8401 255 8436 289
rect 8470 255 8505 289
rect 8539 255 8574 289
rect 8608 255 8643 289
rect 8677 255 8712 289
rect 8746 255 8781 289
rect 8815 255 8850 289
rect 8884 255 8919 289
rect 8953 255 8988 289
rect 9022 255 9057 289
rect 9091 255 9126 289
rect 9160 255 9195 289
rect 9229 255 9264 289
rect 9298 255 9333 289
rect 9367 255 9402 289
rect 9436 255 9471 289
rect 9505 255 9540 289
rect 9574 255 9609 289
rect 9643 255 9678 289
rect 9712 255 9747 289
rect 9781 255 9816 289
rect 9850 255 9885 289
rect 9919 255 9954 289
rect 9988 255 10023 289
rect 10057 255 10092 289
rect 10126 255 10161 289
rect 10195 255 10230 289
rect 10264 255 10299 289
rect 10333 255 10368 289
rect 10402 255 10437 289
rect 10471 255 10506 289
rect 10540 255 10575 289
rect 10609 255 10643 289
rect 10677 255 10711 289
rect 10745 255 10779 289
rect 10813 255 10847 289
rect 10881 255 10915 289
rect 10949 255 10983 289
rect 11017 255 11051 289
rect 11085 255 11119 289
rect 11153 255 11187 289
rect 11221 255 11255 289
rect 11289 255 11323 289
rect 11357 255 11391 289
rect 11425 255 11459 289
rect 11493 255 11527 289
rect 11561 255 11595 289
rect 11629 255 11663 289
rect 11697 255 11731 289
rect 11765 255 11799 289
rect 11833 255 11867 289
rect 11901 255 11935 289
rect 11969 255 12003 289
rect 12037 255 12071 289
rect 12105 255 12139 289
rect 12173 255 12207 289
rect 12241 255 12275 289
rect 12309 255 12343 289
rect 12377 255 12411 289
rect 12445 255 12479 289
rect 12513 255 12547 289
rect 12581 255 12615 289
rect 12649 255 12683 289
rect 12717 255 12751 289
rect 12785 255 12819 289
rect 12853 255 12887 289
rect 12921 255 12955 289
rect 12989 255 13023 289
rect 13057 255 13091 289
rect 13125 255 13159 289
rect 13193 255 13227 289
rect 13261 255 13295 289
rect 13329 255 13363 289
rect 13397 255 13431 289
rect 13465 255 13499 289
rect 13533 255 13567 289
rect 13601 255 13635 289
rect 13669 255 13703 289
rect 13737 255 13771 289
rect 13805 255 13839 289
rect 13873 255 13907 289
rect 13941 255 13975 289
rect 14009 255 14043 289
rect 14077 255 14111 289
rect 14145 255 14179 289
rect 14213 255 14247 289
rect 14281 255 14315 289
rect 14349 255 14383 289
rect 14417 255 14451 289
rect 14485 255 14519 289
rect 14553 255 14587 289
rect 14621 255 14655 289
rect 14689 255 14723 289
rect 14757 255 14791 289
rect 14825 255 14859 289
rect 14893 274 14932 289
rect 14966 274 15000 308
rect 15034 274 15068 308
rect 15102 274 15117 308
rect 14893 255 15117 274
rect 7022 236 15117 255
rect 7022 211 14932 236
rect 7022 177 7056 211
rect 7090 177 7125 211
rect 7159 177 7194 211
rect 7228 177 7263 211
rect 7297 177 7332 211
rect 7366 177 7401 211
rect 7435 177 7470 211
rect 7504 177 7539 211
rect 7573 177 7608 211
rect 7642 177 7677 211
rect 7711 177 7746 211
rect 7780 177 7815 211
rect 7849 177 7884 211
rect 7918 177 7953 211
rect 7987 177 8022 211
rect 8056 177 8091 211
rect 8125 177 8160 211
rect 8194 177 8229 211
rect 8263 177 8298 211
rect 8332 177 8367 211
rect 8401 177 8436 211
rect 8470 177 8505 211
rect 8539 177 8574 211
rect 8608 177 8643 211
rect 8677 177 8712 211
rect 8746 177 8781 211
rect 8815 177 8850 211
rect 8884 177 8919 211
rect 8953 177 8988 211
rect 9022 177 9057 211
rect 9091 177 9126 211
rect 9160 177 9195 211
rect 9229 177 9264 211
rect 9298 177 9333 211
rect 9367 177 9402 211
rect 9436 177 9471 211
rect 9505 177 9540 211
rect 9574 177 9609 211
rect 9643 177 9678 211
rect 9712 177 9747 211
rect 9781 177 9816 211
rect 9850 177 9885 211
rect 9919 177 9954 211
rect 9988 177 10023 211
rect 10057 177 10092 211
rect 10126 177 10161 211
rect 10195 177 10230 211
rect 10264 177 10299 211
rect 10333 177 10368 211
rect 10402 177 10437 211
rect 10471 177 10506 211
rect 10540 177 10575 211
rect 10609 177 10643 211
rect 10677 177 10711 211
rect 10745 177 10779 211
rect 10813 177 10847 211
rect 10881 177 10915 211
rect 10949 177 10983 211
rect 11017 177 11051 211
rect 11085 177 11119 211
rect 11153 177 11187 211
rect 11221 177 11255 211
rect 11289 177 11323 211
rect 11357 177 11391 211
rect 11425 177 11459 211
rect 11493 177 11527 211
rect 11561 177 11595 211
rect 11629 177 11663 211
rect 11697 177 11731 211
rect 11765 177 11799 211
rect 11833 177 11867 211
rect 11901 177 11935 211
rect 11969 177 12003 211
rect 12037 177 12071 211
rect 12105 177 12139 211
rect 12173 177 12207 211
rect 12241 177 12275 211
rect 12309 177 12343 211
rect 12377 177 12411 211
rect 12445 177 12479 211
rect 12513 177 12547 211
rect 12581 177 12615 211
rect 12649 177 12683 211
rect 12717 177 12751 211
rect 12785 177 12819 211
rect 12853 177 12887 211
rect 12921 177 12955 211
rect 12989 177 13023 211
rect 13057 177 13091 211
rect 13125 177 13159 211
rect 13193 177 13227 211
rect 13261 177 13295 211
rect 13329 177 13363 211
rect 13397 177 13431 211
rect 13465 177 13499 211
rect 13533 177 13567 211
rect 13601 177 13635 211
rect 13669 177 13703 211
rect 13737 177 13771 211
rect 13805 177 13839 211
rect 13873 177 13907 211
rect 13941 177 13975 211
rect 14009 177 14043 211
rect 14077 177 14111 211
rect 14145 177 14179 211
rect 14213 177 14247 211
rect 14281 177 14315 211
rect 14349 177 14383 211
rect 14417 177 14451 211
rect 14485 177 14519 211
rect 14553 177 14587 211
rect 14621 177 14655 211
rect 14689 177 14723 211
rect 14757 177 14791 211
rect 14825 177 14859 211
rect 14893 202 14932 211
rect 14966 202 15000 236
rect 15034 202 15068 236
rect 15102 202 15117 236
rect 14893 177 15117 202
rect 7022 164 15117 177
rect 7022 133 14932 164
rect 7022 99 7056 133
rect 7090 99 7125 133
rect 7159 99 7194 133
rect 7228 99 7263 133
rect 7297 99 7332 133
rect 7366 99 7401 133
rect 7435 99 7470 133
rect 7504 99 7539 133
rect 7573 99 7608 133
rect 7642 99 7677 133
rect 7711 99 7746 133
rect 7780 99 7815 133
rect 7849 99 7884 133
rect 7918 99 7953 133
rect 7987 99 8022 133
rect 8056 99 8091 133
rect 8125 99 8160 133
rect 8194 99 8229 133
rect 8263 99 8298 133
rect 8332 99 8367 133
rect 8401 99 8436 133
rect 8470 99 8505 133
rect 8539 99 8574 133
rect 8608 99 8643 133
rect 8677 99 8712 133
rect 8746 99 8781 133
rect 8815 99 8850 133
rect 8884 99 8919 133
rect 8953 99 8988 133
rect 9022 99 9057 133
rect 9091 99 9126 133
rect 9160 99 9195 133
rect 9229 99 9264 133
rect 9298 99 9333 133
rect 9367 99 9402 133
rect 9436 99 9471 133
rect 9505 99 9540 133
rect 9574 99 9609 133
rect 9643 99 9678 133
rect 9712 99 9747 133
rect 9781 99 9816 133
rect 9850 99 9885 133
rect 9919 99 9954 133
rect 9988 99 10023 133
rect 10057 99 10092 133
rect 10126 99 10161 133
rect 10195 99 10230 133
rect 10264 99 10299 133
rect 10333 99 10368 133
rect 10402 99 10437 133
rect 10471 99 10506 133
rect 10540 99 10575 133
rect 10609 99 10643 133
rect 10677 99 10711 133
rect 10745 99 10779 133
rect 10813 99 10847 133
rect 10881 99 10915 133
rect 10949 99 10983 133
rect 11017 99 11051 133
rect 11085 99 11119 133
rect 11153 99 11187 133
rect 11221 99 11255 133
rect 11289 99 11323 133
rect 11357 99 11391 133
rect 11425 99 11459 133
rect 11493 99 11527 133
rect 11561 99 11595 133
rect 11629 99 11663 133
rect 11697 99 11731 133
rect 11765 99 11799 133
rect 11833 99 11867 133
rect 11901 99 11935 133
rect 11969 99 12003 133
rect 12037 99 12071 133
rect 12105 99 12139 133
rect 12173 99 12207 133
rect 12241 99 12275 133
rect 12309 99 12343 133
rect 12377 99 12411 133
rect 12445 99 12479 133
rect 12513 99 12547 133
rect 12581 99 12615 133
rect 12649 99 12683 133
rect 12717 99 12751 133
rect 12785 99 12819 133
rect 12853 99 12887 133
rect 12921 99 12955 133
rect 12989 99 13023 133
rect 13057 99 13091 133
rect 13125 99 13159 133
rect 13193 99 13227 133
rect 13261 99 13295 133
rect 13329 99 13363 133
rect 13397 99 13431 133
rect 13465 99 13499 133
rect 13533 99 13567 133
rect 13601 99 13635 133
rect 13669 99 13703 133
rect 13737 99 13771 133
rect 13805 99 13839 133
rect 13873 99 13907 133
rect 13941 99 13975 133
rect 14009 99 14043 133
rect 14077 99 14111 133
rect 14145 99 14179 133
rect 14213 99 14247 133
rect 14281 99 14315 133
rect 14349 99 14383 133
rect 14417 99 14451 133
rect 14485 99 14519 133
rect 14553 99 14587 133
rect 14621 99 14655 133
rect 14689 99 14723 133
rect 14757 99 14791 133
rect 14825 99 14859 133
rect 14893 130 14932 133
rect 14966 130 15000 164
rect 15034 130 15068 164
rect 15102 130 15117 164
rect 14893 99 15117 130
rect 7022 91 15117 99
rect 7022 57 14932 91
rect 14966 57 15000 91
rect 15034 57 15068 91
rect 15102 57 15117 91
rect 7022 55 15117 57
rect 7022 21 7056 55
rect 7090 21 7125 55
rect 7159 21 7194 55
rect 7228 21 7263 55
rect 7297 21 7332 55
rect 7366 21 7401 55
rect 7435 21 7470 55
rect 7504 21 7539 55
rect 7573 21 7608 55
rect 7642 21 7677 55
rect 7711 21 7746 55
rect 7780 21 7815 55
rect 7849 21 7884 55
rect 7918 21 7953 55
rect 7987 21 8022 55
rect 8056 21 8091 55
rect 8125 21 8160 55
rect 8194 21 8229 55
rect 8263 21 8298 55
rect 8332 21 8367 55
rect 8401 21 8436 55
rect 8470 21 8505 55
rect 8539 21 8574 55
rect 8608 21 8643 55
rect 8677 21 8712 55
rect 8746 21 8781 55
rect 8815 21 8850 55
rect 8884 21 8919 55
rect 8953 21 8988 55
rect 9022 21 9057 55
rect 9091 21 9126 55
rect 9160 21 9195 55
rect 9229 21 9264 55
rect 9298 21 9333 55
rect 9367 21 9402 55
rect 9436 21 9471 55
rect 9505 21 9540 55
rect 9574 21 9609 55
rect 9643 21 9678 55
rect 9712 21 9747 55
rect 9781 21 9816 55
rect 9850 21 9885 55
rect 9919 21 9954 55
rect 9988 21 10023 55
rect 10057 21 10092 55
rect 10126 21 10161 55
rect 10195 21 10230 55
rect 10264 21 10299 55
rect 10333 21 10368 55
rect 10402 21 10437 55
rect 10471 21 10506 55
rect 10540 21 10575 55
rect 10609 21 10643 55
rect 10677 21 10711 55
rect 10745 21 10779 55
rect 10813 21 10847 55
rect 10881 21 10915 55
rect 10949 21 10983 55
rect 11017 21 11051 55
rect 11085 21 11119 55
rect 11153 21 11187 55
rect 11221 21 11255 55
rect 11289 21 11323 55
rect 11357 21 11391 55
rect 11425 21 11459 55
rect 11493 21 11527 55
rect 11561 21 11595 55
rect 11629 21 11663 55
rect 11697 21 11731 55
rect 11765 21 11799 55
rect 11833 21 11867 55
rect 11901 21 11935 55
rect 11969 21 12003 55
rect 12037 21 12071 55
rect 12105 21 12139 55
rect 12173 21 12207 55
rect 12241 21 12275 55
rect 12309 21 12343 55
rect 12377 21 12411 55
rect 12445 21 12479 55
rect 12513 21 12547 55
rect 12581 21 12615 55
rect 12649 21 12683 55
rect 12717 21 12751 55
rect 12785 21 12819 55
rect 12853 21 12887 55
rect 12921 21 12955 55
rect 12989 21 13023 55
rect 13057 21 13091 55
rect 13125 21 13159 55
rect 13193 21 13227 55
rect 13261 21 13295 55
rect 13329 21 13363 55
rect 13397 21 13431 55
rect 13465 21 13499 55
rect 13533 21 13567 55
rect 13601 21 13635 55
rect 13669 21 13703 55
rect 13737 21 13771 55
rect 13805 21 13839 55
rect 13873 21 13907 55
rect 13941 21 13975 55
rect 14009 21 14043 55
rect 14077 21 14111 55
rect 14145 21 14179 55
rect 14213 21 14247 55
rect 14281 21 14315 55
rect 14349 21 14383 55
rect 14417 21 14451 55
rect 14485 21 14519 55
rect 14553 21 14587 55
rect 14621 21 14655 55
rect 14689 21 14723 55
rect 14757 21 14791 55
rect 14825 21 14859 55
rect 14893 21 15117 55
rect 7022 19 15117 21
<< mvnsubdiff >>
rect 12580 15655 12636 15661
rect 14376 15655 14416 15661
rect 12580 15651 14416 15655
rect 12580 15617 12660 15651
rect 12694 15617 12730 15651
rect 12764 15617 12800 15651
rect 12834 15617 12869 15651
rect 12903 15617 12938 15651
rect 12972 15617 13007 15651
rect 13041 15617 13076 15651
rect 13110 15617 13145 15651
rect 13179 15617 13214 15651
rect 13248 15617 13283 15651
rect 13317 15617 13352 15651
rect 13386 15617 13421 15651
rect 13455 15617 13490 15651
rect 13524 15617 13559 15651
rect 13593 15617 13628 15651
rect 13662 15617 13697 15651
rect 13731 15617 13766 15651
rect 13800 15617 13835 15651
rect 13869 15617 13904 15651
rect 13938 15617 13973 15651
rect 14007 15617 14042 15651
rect 14076 15617 14111 15651
rect 14145 15617 14180 15651
rect 14214 15617 14249 15651
rect 14283 15617 14318 15651
rect 14352 15617 14416 15651
rect 12580 15581 14416 15617
rect 12580 15547 12660 15581
rect 12694 15547 12730 15581
rect 12764 15547 12800 15581
rect 12834 15547 12869 15581
rect 12903 15547 12938 15581
rect 12972 15547 13007 15581
rect 13041 15547 13076 15581
rect 13110 15547 13145 15581
rect 13179 15547 13214 15581
rect 13248 15547 13283 15581
rect 13317 15547 13352 15581
rect 13386 15547 13421 15581
rect 13455 15547 13490 15581
rect 13524 15547 13559 15581
rect 13593 15547 13628 15581
rect 13662 15547 13697 15581
rect 13731 15547 13766 15581
rect 13800 15547 13835 15581
rect 13869 15547 13904 15581
rect 13938 15547 13973 15581
rect 14007 15547 14042 15581
rect 14076 15547 14111 15581
rect 14145 15547 14180 15581
rect 14214 15547 14249 15581
rect 14283 15547 14318 15581
rect 14352 15547 14416 15581
rect 12580 15511 14416 15547
rect 12580 15477 12660 15511
rect 12694 15477 12730 15511
rect 12764 15477 12800 15511
rect 12834 15477 12869 15511
rect 12903 15477 12938 15511
rect 12972 15477 13007 15511
rect 13041 15477 13076 15511
rect 13110 15477 13145 15511
rect 13179 15477 13214 15511
rect 13248 15477 13283 15511
rect 13317 15477 13352 15511
rect 13386 15477 13421 15511
rect 13455 15477 13490 15511
rect 13524 15477 13559 15511
rect 13593 15477 13628 15511
rect 13662 15477 13697 15511
rect 13731 15477 13766 15511
rect 13800 15477 13835 15511
rect 13869 15477 13904 15511
rect 13938 15477 13973 15511
rect 14007 15477 14042 15511
rect 14076 15477 14111 15511
rect 14145 15477 14180 15511
rect 14214 15477 14249 15511
rect 14283 15477 14318 15511
rect 14352 15477 14416 15511
rect 12580 15441 14416 15477
rect 12580 15407 12660 15441
rect 12694 15407 12730 15441
rect 12764 15407 12800 15441
rect 12834 15407 12869 15441
rect 12903 15407 12938 15441
rect 12972 15407 13007 15441
rect 13041 15407 13076 15441
rect 13110 15407 13145 15441
rect 13179 15407 13214 15441
rect 13248 15407 13283 15441
rect 13317 15407 13352 15441
rect 13386 15407 13421 15441
rect 13455 15407 13490 15441
rect 13524 15407 13559 15441
rect 13593 15407 13628 15441
rect 13662 15407 13697 15441
rect 13731 15407 13766 15441
rect 13800 15407 13835 15441
rect 13869 15407 13904 15441
rect 13938 15407 13973 15441
rect 14007 15407 14042 15441
rect 14076 15407 14111 15441
rect 14145 15407 14180 15441
rect 14214 15407 14249 15441
rect 14283 15407 14318 15441
rect 14352 15407 14416 15441
rect 12580 15371 14416 15407
rect 12580 15337 12660 15371
rect 12694 15337 12730 15371
rect 12764 15337 12800 15371
rect 12834 15337 12869 15371
rect 12903 15337 12938 15371
rect 12972 15337 13007 15371
rect 13041 15337 13076 15371
rect 13110 15337 13145 15371
rect 13179 15337 13214 15371
rect 13248 15337 13283 15371
rect 13317 15337 13352 15371
rect 13386 15337 13421 15371
rect 13455 15337 13490 15371
rect 13524 15337 13559 15371
rect 13593 15337 13628 15371
rect 13662 15337 13697 15371
rect 13731 15337 13766 15371
rect 13800 15337 13835 15371
rect 13869 15337 13904 15371
rect 13938 15337 13973 15371
rect 14007 15337 14042 15371
rect 14076 15337 14111 15371
rect 14145 15337 14180 15371
rect 14214 15337 14249 15371
rect 14283 15337 14318 15371
rect 14352 15337 14416 15371
rect 12580 15301 14416 15337
rect 12580 15267 12660 15301
rect 12694 15267 12730 15301
rect 12764 15267 12800 15301
rect 12834 15267 12869 15301
rect 12903 15267 12938 15301
rect 12972 15267 13007 15301
rect 13041 15267 13076 15301
rect 13110 15267 13145 15301
rect 13179 15267 13214 15301
rect 13248 15267 13283 15301
rect 13317 15267 13352 15301
rect 13386 15267 13421 15301
rect 13455 15267 13490 15301
rect 13524 15267 13559 15301
rect 13593 15267 13628 15301
rect 13662 15267 13697 15301
rect 13731 15267 13766 15301
rect 13800 15267 13835 15301
rect 13869 15267 13904 15301
rect 13938 15267 13973 15301
rect 14007 15267 14042 15301
rect 14076 15267 14111 15301
rect 14145 15267 14180 15301
rect 14214 15267 14249 15301
rect 14283 15267 14318 15301
rect 14352 15267 14416 15301
rect 12580 15231 14416 15267
rect 12580 15197 12660 15231
rect 12694 15197 12730 15231
rect 12764 15197 12800 15231
rect 12834 15197 12869 15231
rect 12903 15197 12938 15231
rect 12972 15197 13007 15231
rect 13041 15197 13076 15231
rect 13110 15197 13145 15231
rect 13179 15197 13214 15231
rect 13248 15197 13283 15231
rect 13317 15197 13352 15231
rect 13386 15197 13421 15231
rect 13455 15197 13490 15231
rect 13524 15197 13559 15231
rect 13593 15197 13628 15231
rect 13662 15197 13697 15231
rect 13731 15197 13766 15231
rect 13800 15197 13835 15231
rect 13869 15197 13904 15231
rect 13938 15197 13973 15231
rect 14007 15197 14042 15231
rect 14076 15197 14111 15231
rect 14145 15197 14180 15231
rect 14214 15197 14249 15231
rect 14283 15197 14318 15231
rect 14352 15197 14416 15231
rect 12580 15161 14416 15197
rect 12580 15127 12660 15161
rect 12694 15127 12730 15161
rect 12764 15127 12800 15161
rect 12834 15127 12869 15161
rect 12903 15127 12938 15161
rect 12972 15127 13007 15161
rect 13041 15127 13076 15161
rect 13110 15127 13145 15161
rect 13179 15127 13214 15161
rect 13248 15127 13283 15161
rect 13317 15127 13352 15161
rect 13386 15127 13421 15161
rect 13455 15127 13490 15161
rect 13524 15127 13559 15161
rect 13593 15127 13628 15161
rect 13662 15127 13697 15161
rect 13731 15127 13766 15161
rect 13800 15127 13835 15161
rect 13869 15127 13904 15161
rect 13938 15127 13973 15161
rect 14007 15127 14042 15161
rect 14076 15127 14111 15161
rect 14145 15127 14180 15161
rect 14214 15127 14249 15161
rect 14283 15127 14318 15161
rect 14352 15127 14416 15161
rect 12580 15091 14416 15127
rect 12580 15057 12660 15091
rect 12694 15057 12730 15091
rect 12764 15057 12800 15091
rect 12834 15057 12869 15091
rect 12903 15057 12938 15091
rect 12972 15057 13007 15091
rect 13041 15057 13076 15091
rect 13110 15057 13145 15091
rect 13179 15057 13214 15091
rect 13248 15057 13283 15091
rect 13317 15057 13352 15091
rect 13386 15057 13421 15091
rect 13455 15057 13490 15091
rect 13524 15057 13559 15091
rect 13593 15057 13628 15091
rect 13662 15057 13697 15091
rect 13731 15057 13766 15091
rect 13800 15057 13835 15091
rect 13869 15057 13904 15091
rect 13938 15057 13973 15091
rect 14007 15057 14042 15091
rect 14076 15057 14111 15091
rect 14145 15057 14180 15091
rect 14214 15057 14249 15091
rect 14283 15057 14318 15091
rect 14352 15057 14416 15091
rect 12580 15021 14416 15057
rect 12580 14987 12660 15021
rect 12694 14987 12730 15021
rect 12764 14987 12800 15021
rect 12834 14987 12869 15021
rect 12903 14987 12938 15021
rect 12972 14987 13007 15021
rect 13041 14987 13076 15021
rect 13110 14987 13145 15021
rect 13179 14987 13214 15021
rect 13248 14987 13283 15021
rect 13317 14987 13352 15021
rect 13386 14987 13421 15021
rect 13455 14987 13490 15021
rect 13524 14987 13559 15021
rect 13593 14987 13628 15021
rect 13662 14987 13697 15021
rect 13731 14987 13766 15021
rect 13800 14987 13835 15021
rect 13869 14987 13904 15021
rect 13938 14987 13973 15021
rect 14007 14987 14042 15021
rect 14076 14987 14111 15021
rect 14145 14987 14180 15021
rect 14214 14987 14249 15021
rect 14283 14987 14318 15021
rect 14352 14987 14416 15021
rect 12580 14951 14416 14987
rect 12580 14917 12660 14951
rect 12694 14917 12730 14951
rect 12764 14917 12800 14951
rect 12834 14917 12869 14951
rect 12903 14917 12938 14951
rect 12972 14917 13007 14951
rect 13041 14917 13076 14951
rect 13110 14917 13145 14951
rect 13179 14917 13214 14951
rect 13248 14917 13283 14951
rect 13317 14917 13352 14951
rect 13386 14917 13421 14951
rect 13455 14917 13490 14951
rect 13524 14917 13559 14951
rect 13593 14917 13628 14951
rect 13662 14917 13697 14951
rect 13731 14917 13766 14951
rect 13800 14917 13835 14951
rect 13869 14917 13904 14951
rect 13938 14917 13973 14951
rect 14007 14917 14042 14951
rect 14076 14917 14111 14951
rect 14145 14917 14180 14951
rect 14214 14917 14249 14951
rect 14283 14917 14318 14951
rect 14352 14917 14416 14951
rect 12580 14881 14416 14917
rect 12580 14847 12660 14881
rect 12694 14847 12730 14881
rect 12764 14847 12800 14881
rect 12834 14847 12869 14881
rect 12903 14847 12938 14881
rect 12972 14847 13007 14881
rect 13041 14847 13076 14881
rect 13110 14847 13145 14881
rect 13179 14847 13214 14881
rect 13248 14847 13283 14881
rect 13317 14847 13352 14881
rect 13386 14847 13421 14881
rect 13455 14847 13490 14881
rect 13524 14847 13559 14881
rect 13593 14847 13628 14881
rect 13662 14847 13697 14881
rect 13731 14847 13766 14881
rect 13800 14847 13835 14881
rect 13869 14847 13904 14881
rect 13938 14847 13973 14881
rect 14007 14847 14042 14881
rect 14076 14847 14111 14881
rect 14145 14847 14180 14881
rect 14214 14847 14249 14881
rect 14283 14847 14318 14881
rect 14352 14847 14416 14881
rect 12580 14777 14416 14847
rect 8359 8808 15102 8809
rect 34 8774 15102 8808
rect 34 8740 68 8774
rect 102 8740 138 8774
rect 172 8740 208 8774
rect 242 8740 278 8774
rect 312 8740 348 8774
rect 382 8740 418 8774
rect 452 8740 488 8774
rect 522 8740 558 8774
rect 592 8740 628 8774
rect 662 8740 698 8774
rect 732 8740 768 8774
rect 802 8740 838 8774
rect 872 8740 908 8774
rect 942 8740 978 8774
rect 1012 8740 1048 8774
rect 1082 8740 1118 8774
rect 1152 8740 1188 8774
rect 1222 8740 1258 8774
rect 1292 8740 1328 8774
rect 1362 8740 1398 8774
rect 1432 8740 1467 8774
rect 1501 8740 1536 8774
rect 1570 8740 1605 8774
rect 1639 8740 1674 8774
rect 1708 8740 1743 8774
rect 1777 8740 1812 8774
rect 1846 8740 1881 8774
rect 1915 8740 1950 8774
rect 1984 8740 2019 8774
rect 2053 8740 2088 8774
rect 2122 8740 2157 8774
rect 2191 8740 2226 8774
rect 2260 8740 2295 8774
rect 2329 8740 2364 8774
rect 2398 8740 2433 8774
rect 2467 8740 2502 8774
rect 2536 8740 2571 8774
rect 2605 8740 2640 8774
rect 2674 8740 2709 8774
rect 2743 8740 2778 8774
rect 2812 8740 2847 8774
rect 2881 8773 15102 8774
rect 2881 8770 8393 8773
rect 2881 8740 2933 8770
rect 34 8736 2933 8740
rect 2967 8736 3002 8770
rect 3036 8736 3071 8770
rect 3105 8736 3139 8770
rect 3173 8736 3207 8770
rect 3241 8736 3275 8770
rect 3309 8736 3343 8770
rect 3377 8736 3411 8770
rect 3445 8736 3479 8770
rect 3513 8736 3547 8770
rect 3581 8736 3615 8770
rect 3649 8736 3683 8770
rect 3717 8736 3751 8770
rect 3785 8736 3819 8770
rect 3853 8736 3887 8770
rect 3921 8736 3955 8770
rect 3989 8736 4023 8770
rect 4057 8736 4091 8770
rect 4125 8736 4159 8770
rect 4193 8736 4227 8770
rect 4261 8736 4295 8770
rect 4329 8736 4363 8770
rect 4397 8736 4431 8770
rect 4465 8736 4499 8770
rect 4533 8736 4567 8770
rect 4601 8736 4635 8770
rect 4669 8736 4703 8770
rect 4737 8736 4771 8770
rect 4805 8736 4839 8770
rect 4873 8736 4907 8770
rect 4941 8736 4975 8770
rect 5009 8736 5043 8770
rect 5077 8736 5111 8770
rect 5145 8736 5179 8770
rect 5213 8736 5247 8770
rect 5281 8736 5315 8770
rect 5349 8736 5383 8770
rect 5417 8736 5451 8770
rect 5485 8736 5519 8770
rect 5553 8736 5587 8770
rect 5621 8736 5655 8770
rect 5689 8736 5723 8770
rect 5757 8736 5791 8770
rect 5825 8736 5859 8770
rect 5893 8736 5927 8770
rect 5961 8736 5995 8770
rect 6029 8736 6063 8770
rect 6097 8736 6131 8770
rect 6165 8736 6199 8770
rect 6233 8736 6267 8770
rect 6301 8736 6335 8770
rect 6369 8736 6403 8770
rect 6437 8736 6471 8770
rect 6505 8736 6539 8770
rect 6573 8736 6607 8770
rect 6641 8736 6675 8770
rect 6709 8736 6743 8770
rect 6777 8736 6811 8770
rect 6845 8736 6879 8770
rect 6913 8736 6947 8770
rect 6981 8736 7015 8770
rect 7049 8736 7083 8770
rect 7117 8736 7151 8770
rect 7185 8736 7219 8770
rect 7253 8736 7287 8770
rect 7321 8736 7355 8770
rect 7389 8736 7423 8770
rect 7457 8736 7491 8770
rect 7525 8736 7559 8770
rect 7593 8736 7627 8770
rect 7661 8736 7695 8770
rect 7729 8736 7763 8770
rect 7797 8736 7831 8770
rect 7865 8736 7899 8770
rect 7933 8736 7967 8770
rect 8001 8736 8035 8770
rect 8069 8736 8103 8770
rect 8137 8736 8171 8770
rect 8205 8736 8239 8770
rect 8273 8736 8307 8770
rect 8341 8739 8393 8770
rect 8427 8739 8462 8773
rect 8496 8739 8531 8773
rect 8565 8739 8600 8773
rect 8634 8739 8669 8773
rect 8703 8739 8738 8773
rect 8772 8739 8807 8773
rect 8841 8739 8876 8773
rect 8910 8739 8945 8773
rect 8979 8739 9014 8773
rect 9048 8739 9083 8773
rect 9117 8739 9152 8773
rect 9186 8739 9220 8773
rect 9254 8739 9288 8773
rect 9322 8739 9356 8773
rect 9390 8739 9424 8773
rect 9458 8739 9492 8773
rect 9526 8739 9560 8773
rect 9594 8739 9628 8773
rect 9662 8739 9696 8773
rect 9730 8739 9764 8773
rect 9798 8739 9832 8773
rect 9866 8739 9900 8773
rect 9934 8739 9968 8773
rect 10002 8739 10036 8773
rect 10070 8739 10104 8773
rect 10138 8739 10172 8773
rect 10206 8739 10240 8773
rect 10274 8739 10308 8773
rect 10342 8739 10376 8773
rect 10410 8739 10444 8773
rect 10478 8739 10512 8773
rect 10546 8739 10580 8773
rect 10614 8739 10648 8773
rect 10682 8739 10716 8773
rect 10750 8739 10784 8773
rect 10818 8739 10852 8773
rect 10886 8739 10920 8773
rect 10954 8739 10988 8773
rect 11022 8739 11056 8773
rect 11090 8739 11124 8773
rect 11158 8739 11192 8773
rect 11226 8739 11260 8773
rect 11294 8739 11328 8773
rect 11362 8739 11396 8773
rect 11430 8739 11464 8773
rect 11498 8739 11532 8773
rect 11566 8739 11600 8773
rect 11634 8739 11668 8773
rect 11702 8739 11736 8773
rect 11770 8739 11804 8773
rect 11838 8739 11872 8773
rect 11906 8739 11940 8773
rect 11974 8739 12008 8773
rect 12042 8739 12076 8773
rect 12110 8739 12144 8773
rect 12178 8739 12212 8773
rect 12246 8739 12280 8773
rect 12314 8739 12348 8773
rect 12382 8739 12416 8773
rect 12450 8739 12484 8773
rect 12518 8739 12552 8773
rect 12586 8739 12620 8773
rect 12654 8739 12688 8773
rect 12722 8739 12756 8773
rect 12790 8739 12824 8773
rect 12858 8739 12892 8773
rect 12926 8739 12960 8773
rect 12994 8739 13028 8773
rect 13062 8739 13096 8773
rect 13130 8739 13164 8773
rect 13198 8739 13232 8773
rect 13266 8739 13300 8773
rect 13334 8739 13368 8773
rect 13402 8739 13436 8773
rect 13470 8739 13504 8773
rect 13538 8739 13572 8773
rect 13606 8739 13640 8773
rect 13674 8739 13708 8773
rect 13742 8739 13776 8773
rect 13810 8739 13844 8773
rect 13878 8739 13912 8773
rect 13946 8739 13980 8773
rect 14014 8739 14048 8773
rect 14082 8739 14116 8773
rect 14150 8739 14184 8773
rect 14218 8739 14252 8773
rect 14286 8739 14320 8773
rect 14354 8739 14388 8773
rect 14422 8739 14456 8773
rect 14490 8739 14524 8773
rect 14558 8739 14592 8773
rect 14626 8739 14660 8773
rect 14694 8739 14728 8773
rect 14762 8739 14796 8773
rect 14830 8739 14864 8773
rect 14898 8739 15102 8773
rect 8341 8736 15102 8739
rect 34 8721 15102 8736
rect 34 8700 14932 8721
rect 34 8666 68 8700
rect 102 8666 138 8700
rect 172 8666 208 8700
rect 242 8666 278 8700
rect 312 8666 348 8700
rect 382 8666 418 8700
rect 452 8666 488 8700
rect 522 8666 558 8700
rect 592 8666 628 8700
rect 662 8666 698 8700
rect 732 8666 768 8700
rect 802 8666 838 8700
rect 872 8666 908 8700
rect 942 8666 978 8700
rect 1012 8666 1048 8700
rect 1082 8666 1118 8700
rect 1152 8666 1188 8700
rect 1222 8666 1258 8700
rect 1292 8666 1328 8700
rect 1362 8666 1398 8700
rect 1432 8666 1467 8700
rect 1501 8666 1536 8700
rect 1570 8666 1605 8700
rect 1639 8666 1674 8700
rect 1708 8666 1743 8700
rect 1777 8666 1812 8700
rect 1846 8666 1881 8700
rect 1915 8666 1950 8700
rect 1984 8666 2019 8700
rect 2053 8666 2088 8700
rect 2122 8666 2157 8700
rect 2191 8666 2226 8700
rect 2260 8666 2295 8700
rect 2329 8666 2364 8700
rect 2398 8666 2433 8700
rect 2467 8666 2502 8700
rect 2536 8666 2571 8700
rect 2605 8666 2640 8700
rect 2674 8666 2709 8700
rect 2743 8666 2778 8700
rect 2812 8666 2847 8700
rect 2881 8666 2933 8700
rect 2967 8666 3002 8700
rect 3036 8666 3071 8700
rect 3105 8666 3139 8700
rect 3173 8666 3207 8700
rect 3241 8666 3275 8700
rect 3309 8666 3343 8700
rect 3377 8666 3411 8700
rect 3445 8666 3479 8700
rect 3513 8666 3547 8700
rect 3581 8666 3615 8700
rect 3649 8666 3683 8700
rect 3717 8666 3751 8700
rect 3785 8666 3819 8700
rect 3853 8666 3887 8700
rect 3921 8666 3955 8700
rect 3989 8666 4023 8700
rect 4057 8666 4091 8700
rect 4125 8666 4159 8700
rect 4193 8666 4227 8700
rect 4261 8666 4295 8700
rect 4329 8666 4363 8700
rect 4397 8666 4431 8700
rect 4465 8666 4499 8700
rect 4533 8666 4567 8700
rect 4601 8666 4635 8700
rect 4669 8666 4703 8700
rect 4737 8666 4771 8700
rect 4805 8666 4839 8700
rect 4873 8666 4907 8700
rect 4941 8666 4975 8700
rect 5009 8666 5043 8700
rect 5077 8666 5111 8700
rect 5145 8666 5179 8700
rect 5213 8666 5247 8700
rect 5281 8666 5315 8700
rect 5349 8666 5383 8700
rect 5417 8666 5451 8700
rect 5485 8666 5519 8700
rect 5553 8666 5587 8700
rect 5621 8666 5655 8700
rect 5689 8666 5723 8700
rect 5757 8666 5791 8700
rect 5825 8666 5859 8700
rect 5893 8666 5927 8700
rect 5961 8666 5995 8700
rect 6029 8666 6063 8700
rect 6097 8666 6131 8700
rect 6165 8666 6199 8700
rect 6233 8666 6267 8700
rect 6301 8666 6335 8700
rect 6369 8666 6403 8700
rect 6437 8666 6471 8700
rect 6505 8666 6539 8700
rect 6573 8666 6607 8700
rect 6641 8666 6675 8700
rect 6709 8666 6743 8700
rect 6777 8666 6811 8700
rect 6845 8666 6879 8700
rect 6913 8666 6947 8700
rect 6981 8666 7015 8700
rect 7049 8666 7083 8700
rect 7117 8666 7151 8700
rect 7185 8666 7219 8700
rect 7253 8666 7287 8700
rect 7321 8666 7355 8700
rect 7389 8666 7423 8700
rect 7457 8666 7491 8700
rect 7525 8666 7559 8700
rect 7593 8666 7627 8700
rect 7661 8666 7695 8700
rect 7729 8666 7763 8700
rect 7797 8666 7831 8700
rect 7865 8666 7899 8700
rect 7933 8666 7967 8700
rect 8001 8666 8035 8700
rect 8069 8666 8103 8700
rect 8137 8666 8171 8700
rect 8205 8666 8239 8700
rect 8273 8666 8307 8700
rect 8341 8693 14932 8700
rect 8341 8666 8393 8693
rect 34 8659 8393 8666
rect 8427 8659 8462 8693
rect 8496 8659 8531 8693
rect 8565 8659 8600 8693
rect 8634 8659 8669 8693
rect 8703 8659 8738 8693
rect 8772 8659 8807 8693
rect 8841 8659 8876 8693
rect 8910 8659 8945 8693
rect 8979 8659 9014 8693
rect 9048 8659 9083 8693
rect 9117 8659 9152 8693
rect 9186 8659 9220 8693
rect 9254 8659 9288 8693
rect 9322 8659 9356 8693
rect 9390 8659 9424 8693
rect 9458 8659 9492 8693
rect 9526 8659 9560 8693
rect 9594 8659 9628 8693
rect 9662 8659 9696 8693
rect 9730 8659 9764 8693
rect 9798 8659 9832 8693
rect 9866 8659 9900 8693
rect 9934 8659 9968 8693
rect 10002 8659 10036 8693
rect 10070 8659 10104 8693
rect 10138 8659 10172 8693
rect 10206 8659 10240 8693
rect 10274 8659 10308 8693
rect 10342 8659 10376 8693
rect 10410 8659 10444 8693
rect 10478 8659 10512 8693
rect 10546 8659 10580 8693
rect 10614 8659 10648 8693
rect 10682 8659 10716 8693
rect 10750 8659 10784 8693
rect 10818 8659 10852 8693
rect 10886 8659 10920 8693
rect 10954 8659 10988 8693
rect 11022 8659 11056 8693
rect 11090 8659 11124 8693
rect 11158 8659 11192 8693
rect 11226 8659 11260 8693
rect 11294 8659 11328 8693
rect 11362 8659 11396 8693
rect 11430 8659 11464 8693
rect 11498 8659 11532 8693
rect 11566 8659 11600 8693
rect 11634 8659 11668 8693
rect 11702 8659 11736 8693
rect 11770 8659 11804 8693
rect 11838 8659 11872 8693
rect 11906 8659 11940 8693
rect 11974 8659 12008 8693
rect 12042 8659 12076 8693
rect 12110 8659 12144 8693
rect 12178 8659 12212 8693
rect 12246 8659 12280 8693
rect 12314 8659 12348 8693
rect 12382 8659 12416 8693
rect 12450 8659 12484 8693
rect 12518 8659 12552 8693
rect 12586 8659 12620 8693
rect 12654 8659 12688 8693
rect 12722 8659 12756 8693
rect 12790 8659 12824 8693
rect 12858 8659 12892 8693
rect 12926 8659 12960 8693
rect 12994 8659 13028 8693
rect 13062 8659 13096 8693
rect 13130 8659 13164 8693
rect 13198 8659 13232 8693
rect 13266 8659 13300 8693
rect 13334 8659 13368 8693
rect 13402 8659 13436 8693
rect 13470 8659 13504 8693
rect 13538 8659 13572 8693
rect 13606 8659 13640 8693
rect 13674 8659 13708 8693
rect 13742 8659 13776 8693
rect 13810 8659 13844 8693
rect 13878 8659 13912 8693
rect 13946 8659 13980 8693
rect 14014 8659 14048 8693
rect 14082 8659 14116 8693
rect 14150 8659 14184 8693
rect 14218 8659 14252 8693
rect 14286 8659 14320 8693
rect 14354 8659 14388 8693
rect 14422 8659 14456 8693
rect 14490 8659 14524 8693
rect 14558 8659 14592 8693
rect 14626 8659 14660 8693
rect 14694 8659 14728 8693
rect 14762 8659 14796 8693
rect 14830 8659 14864 8693
rect 14898 8687 14932 8693
rect 14966 8687 15000 8721
rect 15034 8687 15068 8721
rect 14898 8659 15102 8687
rect 34 8649 15102 8659
rect 34 8630 14932 8649
rect 34 8626 2933 8630
rect 34 8592 68 8626
rect 102 8592 138 8626
rect 172 8592 208 8626
rect 242 8592 278 8626
rect 312 8592 348 8626
rect 382 8592 418 8626
rect 452 8592 488 8626
rect 522 8592 558 8626
rect 592 8592 628 8626
rect 662 8592 698 8626
rect 732 8592 768 8626
rect 802 8592 838 8626
rect 872 8592 908 8626
rect 942 8592 978 8626
rect 1012 8592 1048 8626
rect 1082 8592 1118 8626
rect 1152 8592 1188 8626
rect 1222 8592 1258 8626
rect 1292 8592 1328 8626
rect 1362 8592 1398 8626
rect 1432 8592 1467 8626
rect 1501 8592 1536 8626
rect 1570 8592 1605 8626
rect 1639 8592 1674 8626
rect 1708 8592 1743 8626
rect 1777 8592 1812 8626
rect 1846 8592 1881 8626
rect 1915 8592 1950 8626
rect 1984 8592 2019 8626
rect 2053 8592 2088 8626
rect 2122 8592 2157 8626
rect 2191 8592 2226 8626
rect 2260 8592 2295 8626
rect 2329 8592 2364 8626
rect 2398 8592 2433 8626
rect 2467 8592 2502 8626
rect 2536 8592 2571 8626
rect 2605 8592 2640 8626
rect 2674 8592 2709 8626
rect 2743 8592 2778 8626
rect 2812 8592 2847 8626
rect 2881 8596 2933 8626
rect 2967 8596 3002 8630
rect 3036 8596 3071 8630
rect 3105 8596 3139 8630
rect 3173 8596 3207 8630
rect 3241 8596 3275 8630
rect 3309 8596 3343 8630
rect 3377 8596 3411 8630
rect 3445 8596 3479 8630
rect 3513 8596 3547 8630
rect 3581 8596 3615 8630
rect 3649 8596 3683 8630
rect 3717 8596 3751 8630
rect 3785 8596 3819 8630
rect 3853 8596 3887 8630
rect 3921 8596 3955 8630
rect 3989 8596 4023 8630
rect 4057 8596 4091 8630
rect 4125 8596 4159 8630
rect 4193 8596 4227 8630
rect 4261 8596 4295 8630
rect 4329 8596 4363 8630
rect 4397 8596 4431 8630
rect 4465 8596 4499 8630
rect 4533 8596 4567 8630
rect 4601 8596 4635 8630
rect 4669 8596 4703 8630
rect 4737 8596 4771 8630
rect 4805 8596 4839 8630
rect 4873 8596 4907 8630
rect 4941 8596 4975 8630
rect 5009 8596 5043 8630
rect 5077 8596 5111 8630
rect 5145 8596 5179 8630
rect 5213 8596 5247 8630
rect 5281 8596 5315 8630
rect 5349 8596 5383 8630
rect 5417 8596 5451 8630
rect 5485 8596 5519 8630
rect 5553 8596 5587 8630
rect 5621 8596 5655 8630
rect 5689 8596 5723 8630
rect 5757 8596 5791 8630
rect 5825 8596 5859 8630
rect 5893 8596 5927 8630
rect 5961 8596 5995 8630
rect 6029 8596 6063 8630
rect 6097 8596 6131 8630
rect 6165 8596 6199 8630
rect 6233 8596 6267 8630
rect 6301 8596 6335 8630
rect 6369 8596 6403 8630
rect 6437 8596 6471 8630
rect 6505 8596 6539 8630
rect 6573 8596 6607 8630
rect 6641 8596 6675 8630
rect 6709 8596 6743 8630
rect 6777 8596 6811 8630
rect 6845 8596 6879 8630
rect 6913 8596 6947 8630
rect 6981 8596 7015 8630
rect 7049 8596 7083 8630
rect 7117 8596 7151 8630
rect 7185 8596 7219 8630
rect 7253 8596 7287 8630
rect 7321 8596 7355 8630
rect 7389 8596 7423 8630
rect 7457 8596 7491 8630
rect 7525 8596 7559 8630
rect 7593 8596 7627 8630
rect 7661 8596 7695 8630
rect 7729 8596 7763 8630
rect 7797 8596 7831 8630
rect 7865 8596 7899 8630
rect 7933 8596 7967 8630
rect 8001 8596 8035 8630
rect 8069 8596 8103 8630
rect 8137 8596 8171 8630
rect 8205 8596 8239 8630
rect 8273 8596 8307 8630
rect 8341 8615 14932 8630
rect 14966 8615 15000 8649
rect 15034 8615 15068 8649
rect 8341 8613 15102 8615
rect 8341 8596 8393 8613
rect 2881 8592 8393 8596
rect 34 8579 8393 8592
rect 8427 8579 8462 8613
rect 8496 8579 8531 8613
rect 8565 8579 8600 8613
rect 8634 8579 8669 8613
rect 8703 8579 8738 8613
rect 8772 8579 8807 8613
rect 8841 8579 8876 8613
rect 8910 8579 8945 8613
rect 8979 8579 9014 8613
rect 9048 8579 9083 8613
rect 9117 8579 9152 8613
rect 9186 8579 9220 8613
rect 9254 8579 9288 8613
rect 9322 8579 9356 8613
rect 9390 8579 9424 8613
rect 9458 8579 9492 8613
rect 9526 8579 9560 8613
rect 9594 8579 9628 8613
rect 9662 8579 9696 8613
rect 9730 8579 9764 8613
rect 9798 8579 9832 8613
rect 9866 8579 9900 8613
rect 9934 8579 9968 8613
rect 10002 8579 10036 8613
rect 10070 8579 10104 8613
rect 10138 8579 10172 8613
rect 10206 8579 10240 8613
rect 10274 8579 10308 8613
rect 10342 8579 10376 8613
rect 10410 8579 10444 8613
rect 10478 8579 10512 8613
rect 10546 8579 10580 8613
rect 10614 8579 10648 8613
rect 10682 8579 10716 8613
rect 10750 8579 10784 8613
rect 10818 8579 10852 8613
rect 10886 8579 10920 8613
rect 10954 8579 10988 8613
rect 11022 8579 11056 8613
rect 11090 8579 11124 8613
rect 11158 8579 11192 8613
rect 11226 8579 11260 8613
rect 11294 8579 11328 8613
rect 11362 8579 11396 8613
rect 11430 8579 11464 8613
rect 11498 8579 11532 8613
rect 11566 8579 11600 8613
rect 11634 8579 11668 8613
rect 11702 8579 11736 8613
rect 11770 8579 11804 8613
rect 11838 8579 11872 8613
rect 11906 8579 11940 8613
rect 11974 8579 12008 8613
rect 12042 8579 12076 8613
rect 12110 8579 12144 8613
rect 12178 8579 12212 8613
rect 12246 8579 12280 8613
rect 12314 8579 12348 8613
rect 12382 8579 12416 8613
rect 12450 8579 12484 8613
rect 12518 8579 12552 8613
rect 12586 8579 12620 8613
rect 12654 8579 12688 8613
rect 12722 8579 12756 8613
rect 12790 8579 12824 8613
rect 12858 8579 12892 8613
rect 12926 8579 12960 8613
rect 12994 8579 13028 8613
rect 13062 8579 13096 8613
rect 13130 8579 13164 8613
rect 13198 8579 13232 8613
rect 13266 8579 13300 8613
rect 13334 8579 13368 8613
rect 13402 8579 13436 8613
rect 13470 8579 13504 8613
rect 13538 8579 13572 8613
rect 13606 8579 13640 8613
rect 13674 8579 13708 8613
rect 13742 8579 13776 8613
rect 13810 8579 13844 8613
rect 13878 8579 13912 8613
rect 13946 8579 13980 8613
rect 14014 8579 14048 8613
rect 14082 8579 14116 8613
rect 14150 8579 14184 8613
rect 14218 8579 14252 8613
rect 14286 8579 14320 8613
rect 14354 8579 14388 8613
rect 14422 8579 14456 8613
rect 14490 8579 14524 8613
rect 14558 8579 14592 8613
rect 14626 8579 14660 8613
rect 14694 8579 14728 8613
rect 14762 8579 14796 8613
rect 14830 8579 14864 8613
rect 14898 8579 15102 8613
rect 34 8577 15102 8579
rect 34 8560 14932 8577
rect 34 8552 2933 8560
rect 34 8518 68 8552
rect 102 8518 138 8552
rect 172 8518 208 8552
rect 242 8518 278 8552
rect 312 8518 348 8552
rect 382 8518 418 8552
rect 452 8518 488 8552
rect 522 8518 558 8552
rect 592 8518 628 8552
rect 662 8518 698 8552
rect 732 8518 768 8552
rect 802 8518 838 8552
rect 872 8518 908 8552
rect 942 8518 978 8552
rect 1012 8518 1048 8552
rect 1082 8518 1118 8552
rect 1152 8518 1188 8552
rect 1222 8518 1258 8552
rect 1292 8518 1328 8552
rect 1362 8518 1398 8552
rect 1432 8518 1467 8552
rect 1501 8518 1536 8552
rect 1570 8518 1605 8552
rect 1639 8518 1674 8552
rect 1708 8518 1743 8552
rect 1777 8518 1812 8552
rect 1846 8518 1881 8552
rect 1915 8518 1950 8552
rect 1984 8518 2019 8552
rect 2053 8518 2088 8552
rect 2122 8518 2157 8552
rect 2191 8518 2226 8552
rect 2260 8518 2295 8552
rect 2329 8518 2364 8552
rect 2398 8518 2433 8552
rect 2467 8518 2502 8552
rect 2536 8518 2571 8552
rect 2605 8518 2640 8552
rect 2674 8518 2709 8552
rect 2743 8518 2778 8552
rect 2812 8518 2847 8552
rect 2881 8526 2933 8552
rect 2967 8526 3002 8560
rect 3036 8526 3071 8560
rect 3105 8526 3139 8560
rect 3173 8526 3207 8560
rect 3241 8526 3275 8560
rect 3309 8526 3343 8560
rect 3377 8526 3411 8560
rect 3445 8526 3479 8560
rect 3513 8526 3547 8560
rect 3581 8526 3615 8560
rect 3649 8526 3683 8560
rect 3717 8526 3751 8560
rect 3785 8526 3819 8560
rect 3853 8526 3887 8560
rect 3921 8526 3955 8560
rect 3989 8526 4023 8560
rect 4057 8526 4091 8560
rect 4125 8526 4159 8560
rect 4193 8526 4227 8560
rect 4261 8526 4295 8560
rect 4329 8526 4363 8560
rect 4397 8526 4431 8560
rect 4465 8526 4499 8560
rect 4533 8526 4567 8560
rect 4601 8526 4635 8560
rect 4669 8526 4703 8560
rect 4737 8526 4771 8560
rect 4805 8526 4839 8560
rect 4873 8526 4907 8560
rect 4941 8526 4975 8560
rect 5009 8526 5043 8560
rect 5077 8526 5111 8560
rect 5145 8526 5179 8560
rect 5213 8526 5247 8560
rect 5281 8526 5315 8560
rect 5349 8526 5383 8560
rect 5417 8526 5451 8560
rect 5485 8526 5519 8560
rect 5553 8526 5587 8560
rect 5621 8526 5655 8560
rect 5689 8526 5723 8560
rect 5757 8526 5791 8560
rect 5825 8526 5859 8560
rect 5893 8526 5927 8560
rect 5961 8526 5995 8560
rect 6029 8526 6063 8560
rect 6097 8526 6131 8560
rect 6165 8526 6199 8560
rect 6233 8526 6267 8560
rect 6301 8526 6335 8560
rect 6369 8526 6403 8560
rect 6437 8526 6471 8560
rect 6505 8526 6539 8560
rect 6573 8526 6607 8560
rect 6641 8526 6675 8560
rect 6709 8526 6743 8560
rect 6777 8526 6811 8560
rect 6845 8526 6879 8560
rect 6913 8526 6947 8560
rect 6981 8526 7015 8560
rect 7049 8526 7083 8560
rect 7117 8526 7151 8560
rect 7185 8526 7219 8560
rect 7253 8526 7287 8560
rect 7321 8526 7355 8560
rect 7389 8526 7423 8560
rect 7457 8526 7491 8560
rect 7525 8526 7559 8560
rect 7593 8526 7627 8560
rect 7661 8526 7695 8560
rect 7729 8526 7763 8560
rect 7797 8526 7831 8560
rect 7865 8526 7899 8560
rect 7933 8526 7967 8560
rect 8001 8526 8035 8560
rect 8069 8526 8103 8560
rect 8137 8526 8171 8560
rect 8205 8526 8239 8560
rect 8273 8526 8307 8560
rect 8341 8543 14932 8560
rect 14966 8543 15000 8577
rect 15034 8543 15068 8577
rect 8341 8533 15102 8543
rect 8341 8526 8393 8533
rect 2881 8518 8393 8526
rect 34 8499 8393 8518
rect 8427 8499 8462 8533
rect 8496 8499 8531 8533
rect 8565 8499 8600 8533
rect 8634 8499 8669 8533
rect 8703 8499 8738 8533
rect 8772 8499 8807 8533
rect 8841 8499 8876 8533
rect 8910 8499 8945 8533
rect 8979 8499 9014 8533
rect 9048 8499 9083 8533
rect 9117 8499 9152 8533
rect 9186 8499 9220 8533
rect 9254 8499 9288 8533
rect 9322 8499 9356 8533
rect 9390 8499 9424 8533
rect 9458 8499 9492 8533
rect 9526 8499 9560 8533
rect 9594 8499 9628 8533
rect 9662 8499 9696 8533
rect 9730 8499 9764 8533
rect 9798 8499 9832 8533
rect 9866 8499 9900 8533
rect 9934 8499 9968 8533
rect 10002 8499 10036 8533
rect 10070 8499 10104 8533
rect 10138 8499 10172 8533
rect 10206 8499 10240 8533
rect 10274 8499 10308 8533
rect 10342 8499 10376 8533
rect 10410 8499 10444 8533
rect 10478 8499 10512 8533
rect 10546 8499 10580 8533
rect 10614 8499 10648 8533
rect 10682 8499 10716 8533
rect 10750 8499 10784 8533
rect 10818 8499 10852 8533
rect 10886 8499 10920 8533
rect 10954 8499 10988 8533
rect 11022 8499 11056 8533
rect 11090 8499 11124 8533
rect 11158 8499 11192 8533
rect 11226 8499 11260 8533
rect 11294 8499 11328 8533
rect 11362 8499 11396 8533
rect 11430 8499 11464 8533
rect 11498 8499 11532 8533
rect 11566 8499 11600 8533
rect 11634 8499 11668 8533
rect 11702 8499 11736 8533
rect 11770 8499 11804 8533
rect 11838 8499 11872 8533
rect 11906 8499 11940 8533
rect 11974 8499 12008 8533
rect 12042 8499 12076 8533
rect 12110 8499 12144 8533
rect 12178 8499 12212 8533
rect 12246 8499 12280 8533
rect 12314 8499 12348 8533
rect 12382 8499 12416 8533
rect 12450 8499 12484 8533
rect 12518 8499 12552 8533
rect 12586 8499 12620 8533
rect 12654 8499 12688 8533
rect 12722 8499 12756 8533
rect 12790 8499 12824 8533
rect 12858 8499 12892 8533
rect 12926 8499 12960 8533
rect 12994 8499 13028 8533
rect 13062 8499 13096 8533
rect 13130 8499 13164 8533
rect 13198 8499 13232 8533
rect 13266 8499 13300 8533
rect 13334 8499 13368 8533
rect 13402 8499 13436 8533
rect 13470 8499 13504 8533
rect 13538 8499 13572 8533
rect 13606 8499 13640 8533
rect 13674 8499 13708 8533
rect 13742 8499 13776 8533
rect 13810 8499 13844 8533
rect 13878 8499 13912 8533
rect 13946 8499 13980 8533
rect 14014 8499 14048 8533
rect 14082 8499 14116 8533
rect 14150 8499 14184 8533
rect 14218 8499 14252 8533
rect 14286 8499 14320 8533
rect 14354 8499 14388 8533
rect 14422 8499 14456 8533
rect 14490 8499 14524 8533
rect 14558 8499 14592 8533
rect 14626 8499 14660 8533
rect 14694 8499 14728 8533
rect 14762 8499 14796 8533
rect 14830 8499 14864 8533
rect 14898 8505 15102 8533
rect 14898 8499 14932 8505
rect 34 8490 14932 8499
rect 34 8484 2933 8490
rect 34 8460 136 8484
rect 34 8426 68 8460
rect 102 8426 136 8460
rect 34 8392 136 8426
rect 34 8358 68 8392
rect 102 8358 136 8392
rect 34 8324 136 8358
rect 34 8290 68 8324
rect 102 8290 136 8324
rect 34 8256 136 8290
rect 34 8222 68 8256
rect 102 8222 136 8256
rect 34 8192 136 8222
rect 2899 8456 2933 8484
rect 2967 8456 3002 8490
rect 3036 8456 3071 8490
rect 3105 8456 3139 8490
rect 3173 8456 3207 8490
rect 3241 8456 3275 8490
rect 3309 8456 3343 8490
rect 3377 8456 3411 8490
rect 3445 8456 3479 8490
rect 3513 8456 3547 8490
rect 3581 8456 3615 8490
rect 3649 8456 3683 8490
rect 3717 8456 3751 8490
rect 3785 8456 3819 8490
rect 3853 8456 3887 8490
rect 3921 8456 3955 8490
rect 3989 8456 4023 8490
rect 4057 8456 4091 8490
rect 4125 8456 4159 8490
rect 4193 8456 4227 8490
rect 4261 8456 4295 8490
rect 4329 8456 4363 8490
rect 4397 8456 4431 8490
rect 4465 8456 4499 8490
rect 4533 8456 4567 8490
rect 4601 8456 4635 8490
rect 4669 8456 4703 8490
rect 4737 8456 4771 8490
rect 4805 8456 4839 8490
rect 4873 8456 4907 8490
rect 4941 8456 4975 8490
rect 5009 8456 5043 8490
rect 5077 8456 5111 8490
rect 5145 8456 5179 8490
rect 5213 8456 5247 8490
rect 5281 8456 5315 8490
rect 5349 8456 5383 8490
rect 5417 8456 5451 8490
rect 5485 8456 5519 8490
rect 5553 8456 5587 8490
rect 5621 8456 5655 8490
rect 5689 8456 5723 8490
rect 5757 8456 5791 8490
rect 5825 8456 5859 8490
rect 5893 8456 5927 8490
rect 5961 8456 5995 8490
rect 6029 8456 6063 8490
rect 6097 8456 6131 8490
rect 6165 8456 6199 8490
rect 6233 8456 6267 8490
rect 6301 8456 6335 8490
rect 6369 8456 6403 8490
rect 6437 8456 6471 8490
rect 6505 8456 6539 8490
rect 6573 8456 6607 8490
rect 6641 8456 6675 8490
rect 6709 8456 6743 8490
rect 6777 8456 6811 8490
rect 6845 8456 6879 8490
rect 6913 8456 6947 8490
rect 6981 8456 7015 8490
rect 7049 8456 7083 8490
rect 7117 8456 7151 8490
rect 7185 8456 7219 8490
rect 7253 8456 7287 8490
rect 7321 8456 7355 8490
rect 7389 8456 7423 8490
rect 7457 8456 7491 8490
rect 7525 8456 7559 8490
rect 7593 8456 7627 8490
rect 7661 8456 7695 8490
rect 7729 8456 7763 8490
rect 7797 8456 7831 8490
rect 7865 8456 7899 8490
rect 7933 8456 7967 8490
rect 8001 8456 8035 8490
rect 8069 8456 8103 8490
rect 8137 8456 8171 8490
rect 8205 8456 8239 8490
rect 8273 8456 8307 8490
rect 8341 8471 14932 8490
rect 14966 8471 15000 8505
rect 15034 8471 15068 8505
rect 8341 8456 15102 8471
rect 2899 8453 15102 8456
rect 2899 8420 8393 8453
rect 2899 8386 2933 8420
rect 2967 8386 3002 8420
rect 3036 8386 3071 8420
rect 3105 8386 3139 8420
rect 3173 8386 3207 8420
rect 3241 8386 3275 8420
rect 3309 8386 3343 8420
rect 3377 8386 3411 8420
rect 3445 8386 3479 8420
rect 3513 8386 3547 8420
rect 3581 8386 3615 8420
rect 3649 8386 3683 8420
rect 3717 8386 3751 8420
rect 3785 8386 3819 8420
rect 3853 8386 3887 8420
rect 3921 8386 3955 8420
rect 3989 8386 4023 8420
rect 4057 8386 4091 8420
rect 4125 8386 4159 8420
rect 4193 8386 4227 8420
rect 4261 8386 4295 8420
rect 4329 8386 4363 8420
rect 4397 8386 4431 8420
rect 4465 8386 4499 8420
rect 4533 8386 4567 8420
rect 4601 8386 4635 8420
rect 4669 8386 4703 8420
rect 4737 8386 4771 8420
rect 4805 8386 4839 8420
rect 4873 8386 4907 8420
rect 4941 8386 4975 8420
rect 5009 8386 5043 8420
rect 5077 8386 5111 8420
rect 5145 8386 5179 8420
rect 5213 8386 5247 8420
rect 5281 8386 5315 8420
rect 5349 8386 5383 8420
rect 5417 8386 5451 8420
rect 5485 8386 5519 8420
rect 5553 8386 5587 8420
rect 5621 8386 5655 8420
rect 5689 8386 5723 8420
rect 5757 8386 5791 8420
rect 5825 8386 5859 8420
rect 5893 8386 5927 8420
rect 5961 8386 5995 8420
rect 6029 8386 6063 8420
rect 6097 8386 6131 8420
rect 6165 8386 6199 8420
rect 6233 8386 6267 8420
rect 6301 8386 6335 8420
rect 6369 8386 6403 8420
rect 6437 8386 6471 8420
rect 6505 8386 6539 8420
rect 6573 8386 6607 8420
rect 6641 8386 6675 8420
rect 6709 8386 6743 8420
rect 6777 8386 6811 8420
rect 6845 8386 6879 8420
rect 6913 8386 6947 8420
rect 6981 8386 7015 8420
rect 7049 8386 7083 8420
rect 7117 8386 7151 8420
rect 7185 8386 7219 8420
rect 7253 8386 7287 8420
rect 7321 8386 7355 8420
rect 7389 8386 7423 8420
rect 7457 8386 7491 8420
rect 7525 8386 7559 8420
rect 7593 8386 7627 8420
rect 7661 8386 7695 8420
rect 7729 8386 7763 8420
rect 7797 8386 7831 8420
rect 7865 8386 7899 8420
rect 7933 8386 7967 8420
rect 8001 8386 8035 8420
rect 8069 8386 8103 8420
rect 8137 8386 8171 8420
rect 8205 8386 8239 8420
rect 8273 8386 8307 8420
rect 8341 8419 8393 8420
rect 8427 8419 8462 8453
rect 8496 8419 8531 8453
rect 8565 8419 8600 8453
rect 8634 8419 8669 8453
rect 8703 8419 8738 8453
rect 8772 8419 8807 8453
rect 8841 8419 8876 8453
rect 8910 8419 8945 8453
rect 8979 8419 9014 8453
rect 9048 8419 9083 8453
rect 9117 8419 9152 8453
rect 9186 8419 9220 8453
rect 9254 8419 9288 8453
rect 9322 8419 9356 8453
rect 9390 8419 9424 8453
rect 9458 8419 9492 8453
rect 9526 8419 9560 8453
rect 9594 8419 9628 8453
rect 9662 8419 9696 8453
rect 9730 8419 9764 8453
rect 9798 8419 9832 8453
rect 9866 8419 9900 8453
rect 9934 8419 9968 8453
rect 10002 8419 10036 8453
rect 10070 8419 10104 8453
rect 10138 8419 10172 8453
rect 10206 8419 10240 8453
rect 10274 8419 10308 8453
rect 10342 8419 10376 8453
rect 10410 8419 10444 8453
rect 10478 8419 10512 8453
rect 10546 8419 10580 8453
rect 10614 8419 10648 8453
rect 10682 8419 10716 8453
rect 10750 8419 10784 8453
rect 10818 8419 10852 8453
rect 10886 8419 10920 8453
rect 10954 8419 10988 8453
rect 11022 8419 11056 8453
rect 11090 8419 11124 8453
rect 11158 8419 11192 8453
rect 11226 8419 11260 8453
rect 11294 8419 11328 8453
rect 11362 8419 11396 8453
rect 11430 8419 11464 8453
rect 11498 8419 11532 8453
rect 11566 8419 11600 8453
rect 11634 8419 11668 8453
rect 11702 8419 11736 8453
rect 11770 8419 11804 8453
rect 11838 8419 11872 8453
rect 11906 8419 11940 8453
rect 11974 8419 12008 8453
rect 12042 8419 12076 8453
rect 12110 8419 12144 8453
rect 12178 8419 12212 8453
rect 12246 8419 12280 8453
rect 12314 8419 12348 8453
rect 12382 8419 12416 8453
rect 12450 8419 12484 8453
rect 12518 8419 12552 8453
rect 12586 8419 12620 8453
rect 12654 8419 12688 8453
rect 12722 8419 12756 8453
rect 12790 8419 12824 8453
rect 12858 8419 12892 8453
rect 12926 8419 12960 8453
rect 12994 8419 13028 8453
rect 13062 8419 13096 8453
rect 13130 8419 13164 8453
rect 13198 8419 13232 8453
rect 13266 8419 13300 8453
rect 13334 8419 13368 8453
rect 13402 8419 13436 8453
rect 13470 8419 13504 8453
rect 13538 8419 13572 8453
rect 13606 8419 13640 8453
rect 13674 8419 13708 8453
rect 13742 8419 13776 8453
rect 13810 8419 13844 8453
rect 13878 8419 13912 8453
rect 13946 8419 13980 8453
rect 14014 8419 14048 8453
rect 14082 8419 14116 8453
rect 14150 8419 14184 8453
rect 14218 8419 14252 8453
rect 14286 8419 14320 8453
rect 14354 8419 14388 8453
rect 14422 8419 14456 8453
rect 14490 8419 14524 8453
rect 14558 8419 14592 8453
rect 14626 8419 14660 8453
rect 14694 8419 14728 8453
rect 14762 8419 14796 8453
rect 14830 8419 14864 8453
rect 14898 8433 15102 8453
rect 14898 8419 14932 8433
rect 8341 8399 14932 8419
rect 14966 8399 15000 8433
rect 15034 8399 15068 8433
rect 8341 8386 15102 8399
rect 2899 8383 15102 8386
rect 2899 8350 8375 8383
rect 2899 8316 2933 8350
rect 2967 8316 3002 8350
rect 3036 8316 3071 8350
rect 3105 8316 3139 8350
rect 3173 8316 3207 8350
rect 3241 8316 3275 8350
rect 3309 8316 3343 8350
rect 3377 8316 3411 8350
rect 3445 8316 3479 8350
rect 3513 8316 3547 8350
rect 3581 8316 3615 8350
rect 3649 8316 3683 8350
rect 3717 8316 3751 8350
rect 3785 8316 3819 8350
rect 3853 8316 3887 8350
rect 3921 8316 3955 8350
rect 3989 8316 4023 8350
rect 4057 8316 4091 8350
rect 4125 8316 4159 8350
rect 4193 8316 4227 8350
rect 4261 8316 4295 8350
rect 4329 8316 4363 8350
rect 4397 8316 4431 8350
rect 4465 8316 4499 8350
rect 4533 8316 4567 8350
rect 4601 8316 4635 8350
rect 4669 8316 4703 8350
rect 4737 8316 4771 8350
rect 4805 8316 4839 8350
rect 4873 8316 4907 8350
rect 4941 8316 4975 8350
rect 5009 8316 5043 8350
rect 5077 8316 5111 8350
rect 5145 8316 5179 8350
rect 5213 8316 5247 8350
rect 5281 8316 5315 8350
rect 5349 8316 5383 8350
rect 5417 8316 5451 8350
rect 5485 8316 5519 8350
rect 5553 8316 5587 8350
rect 5621 8316 5655 8350
rect 5689 8316 5723 8350
rect 5757 8316 5791 8350
rect 5825 8316 5859 8350
rect 5893 8316 5927 8350
rect 5961 8316 5995 8350
rect 6029 8316 6063 8350
rect 6097 8316 6131 8350
rect 6165 8316 6199 8350
rect 6233 8316 6267 8350
rect 6301 8316 6335 8350
rect 6369 8316 6403 8350
rect 6437 8316 6471 8350
rect 6505 8316 6539 8350
rect 6573 8316 6607 8350
rect 6641 8316 6675 8350
rect 6709 8316 6743 8350
rect 6777 8316 6811 8350
rect 6845 8316 6879 8350
rect 6913 8316 6947 8350
rect 6981 8316 7015 8350
rect 7049 8316 7083 8350
rect 7117 8316 7151 8350
rect 7185 8316 7219 8350
rect 7253 8316 7287 8350
rect 7321 8316 7355 8350
rect 7389 8316 7423 8350
rect 7457 8316 7491 8350
rect 7525 8316 7559 8350
rect 7593 8316 7627 8350
rect 7661 8316 7695 8350
rect 7729 8316 7763 8350
rect 7797 8316 7831 8350
rect 7865 8316 7899 8350
rect 7933 8316 7967 8350
rect 8001 8316 8035 8350
rect 8069 8316 8103 8350
rect 8137 8316 8171 8350
rect 8205 8316 8239 8350
rect 8273 8316 8307 8350
rect 8341 8316 8375 8350
rect 2899 8280 8375 8316
rect 13498 8361 15102 8383
rect 13498 8357 14932 8361
rect 13498 8323 13532 8357
rect 13566 8323 13603 8357
rect 13637 8323 13674 8357
rect 13708 8323 13744 8357
rect 13778 8323 13814 8357
rect 13848 8323 13884 8357
rect 13918 8323 13954 8357
rect 13988 8323 14024 8357
rect 14058 8323 14094 8357
rect 14128 8323 14164 8357
rect 14198 8323 14234 8357
rect 14268 8323 14304 8357
rect 14338 8323 14374 8357
rect 14408 8323 14444 8357
rect 14478 8323 14514 8357
rect 14548 8323 14584 8357
rect 14618 8323 14654 8357
rect 14688 8323 14724 8357
rect 14758 8323 14794 8357
rect 14828 8323 14864 8357
rect 14898 8327 14932 8357
rect 14966 8327 15000 8361
rect 15034 8327 15068 8361
rect 14898 8323 15102 8327
rect 13498 8289 15102 8323
rect 2899 8246 2933 8280
rect 2967 8246 3002 8280
rect 3036 8246 3071 8280
rect 3105 8246 3139 8280
rect 3173 8246 3207 8280
rect 3241 8246 3275 8280
rect 3309 8246 3343 8280
rect 3377 8246 3411 8280
rect 3445 8246 3479 8280
rect 3513 8246 3547 8280
rect 3581 8246 3615 8280
rect 3649 8246 3683 8280
rect 3717 8246 3751 8280
rect 3785 8246 3819 8280
rect 3853 8246 3887 8280
rect 3921 8246 3955 8280
rect 3989 8246 4023 8280
rect 4057 8246 4091 8280
rect 4125 8246 4159 8280
rect 4193 8246 4227 8280
rect 4261 8246 4295 8280
rect 4329 8246 4363 8280
rect 4397 8246 4431 8280
rect 4465 8246 4499 8280
rect 4533 8246 4567 8280
rect 4601 8246 4635 8280
rect 4669 8246 4703 8280
rect 4737 8246 4771 8280
rect 4805 8246 4839 8280
rect 4873 8246 4907 8280
rect 4941 8246 4975 8280
rect 5009 8246 5043 8280
rect 5077 8246 5111 8280
rect 5145 8246 5179 8280
rect 5213 8246 5247 8280
rect 5281 8246 5315 8280
rect 5349 8246 5383 8280
rect 5417 8246 5451 8280
rect 5485 8246 5519 8280
rect 5553 8246 5587 8280
rect 5621 8246 5655 8280
rect 5689 8246 5723 8280
rect 5757 8246 5791 8280
rect 5825 8246 5859 8280
rect 5893 8246 5927 8280
rect 5961 8246 5995 8280
rect 6029 8246 6063 8280
rect 6097 8246 6131 8280
rect 6165 8246 6199 8280
rect 6233 8246 6267 8280
rect 6301 8246 6335 8280
rect 6369 8246 6403 8280
rect 6437 8246 6471 8280
rect 6505 8246 6539 8280
rect 6573 8246 6607 8280
rect 6641 8246 6675 8280
rect 6709 8246 6743 8280
rect 6777 8246 6811 8280
rect 6845 8246 6879 8280
rect 6913 8246 6947 8280
rect 6981 8246 7015 8280
rect 7049 8246 7083 8280
rect 7117 8246 7151 8280
rect 7185 8246 7219 8280
rect 7253 8246 7287 8280
rect 7321 8246 7355 8280
rect 7389 8246 7423 8280
rect 7457 8246 7491 8280
rect 7525 8246 7559 8280
rect 7593 8246 7627 8280
rect 7661 8246 7695 8280
rect 7729 8246 7763 8280
rect 7797 8246 7831 8280
rect 7865 8246 7899 8280
rect 7933 8246 7967 8280
rect 8001 8246 8035 8280
rect 8069 8246 8103 8280
rect 8137 8246 8171 8280
rect 8205 8246 8239 8280
rect 8273 8246 8307 8280
rect 8341 8246 8375 8280
rect 2899 8210 8375 8246
rect 2899 8192 2933 8210
rect 34 8176 2933 8192
rect 2967 8176 3002 8210
rect 3036 8176 3071 8210
rect 3105 8176 3139 8210
rect 3173 8176 3207 8210
rect 3241 8176 3275 8210
rect 3309 8176 3343 8210
rect 3377 8176 3411 8210
rect 3445 8176 3479 8210
rect 3513 8176 3547 8210
rect 3581 8176 3615 8210
rect 3649 8176 3683 8210
rect 3717 8176 3751 8210
rect 3785 8176 3819 8210
rect 3853 8176 3887 8210
rect 3921 8176 3955 8210
rect 3989 8176 4023 8210
rect 4057 8176 4091 8210
rect 4125 8176 4159 8210
rect 4193 8176 4227 8210
rect 4261 8176 4295 8210
rect 4329 8176 4363 8210
rect 4397 8176 4431 8210
rect 4465 8176 4499 8210
rect 4533 8176 4567 8210
rect 4601 8176 4635 8210
rect 4669 8176 4703 8210
rect 4737 8176 4771 8210
rect 4805 8176 4839 8210
rect 4873 8176 4907 8210
rect 4941 8176 4975 8210
rect 5009 8176 5043 8210
rect 5077 8176 5111 8210
rect 5145 8176 5179 8210
rect 5213 8176 5247 8210
rect 5281 8176 5315 8210
rect 5349 8176 5383 8210
rect 5417 8176 5451 8210
rect 5485 8176 5519 8210
rect 5553 8176 5587 8210
rect 5621 8176 5655 8210
rect 5689 8176 5723 8210
rect 5757 8176 5791 8210
rect 5825 8176 5859 8210
rect 5893 8176 5927 8210
rect 5961 8176 5995 8210
rect 6029 8176 6063 8210
rect 6097 8176 6131 8210
rect 6165 8176 6199 8210
rect 6233 8176 6267 8210
rect 6301 8176 6335 8210
rect 6369 8176 6403 8210
rect 6437 8176 6471 8210
rect 6505 8176 6539 8210
rect 6573 8176 6607 8210
rect 6641 8176 6675 8210
rect 6709 8176 6743 8210
rect 6777 8176 6811 8210
rect 6845 8176 6879 8210
rect 6913 8176 6947 8210
rect 6981 8176 7015 8210
rect 7049 8176 7083 8210
rect 7117 8176 7151 8210
rect 7185 8176 7219 8210
rect 7253 8176 7287 8210
rect 7321 8176 7355 8210
rect 7389 8176 7423 8210
rect 7457 8176 7491 8210
rect 7525 8176 7559 8210
rect 7593 8176 7627 8210
rect 7661 8176 7695 8210
rect 7729 8176 7763 8210
rect 7797 8176 7831 8210
rect 7865 8176 7899 8210
rect 7933 8176 7967 8210
rect 8001 8176 8035 8210
rect 8069 8176 8103 8210
rect 8137 8176 8171 8210
rect 8205 8176 8239 8210
rect 8273 8176 8307 8210
rect 8341 8176 8375 8210
rect 34 8157 8375 8176
rect 34 8123 68 8157
rect 102 8123 138 8157
rect 172 8123 208 8157
rect 242 8123 278 8157
rect 312 8123 348 8157
rect 382 8123 418 8157
rect 452 8123 488 8157
rect 522 8123 558 8157
rect 592 8123 628 8157
rect 662 8123 698 8157
rect 732 8123 768 8157
rect 802 8123 838 8157
rect 872 8123 908 8157
rect 942 8123 978 8157
rect 1012 8123 1048 8157
rect 1082 8123 1118 8157
rect 1152 8123 1188 8157
rect 1222 8123 1258 8157
rect 1292 8123 1328 8157
rect 1362 8123 1398 8157
rect 1432 8123 1467 8157
rect 1501 8123 1536 8157
rect 1570 8123 1605 8157
rect 1639 8123 1674 8157
rect 1708 8123 1743 8157
rect 1777 8123 1812 8157
rect 1846 8123 1881 8157
rect 1915 8123 1950 8157
rect 1984 8123 2019 8157
rect 2053 8123 2088 8157
rect 2122 8123 2157 8157
rect 2191 8123 2226 8157
rect 2260 8123 2295 8157
rect 2329 8123 2364 8157
rect 2398 8123 2433 8157
rect 2467 8123 2502 8157
rect 2536 8123 2571 8157
rect 2605 8123 2640 8157
rect 2674 8123 2709 8157
rect 2743 8123 2778 8157
rect 2812 8123 2847 8157
rect 2881 8140 8375 8157
rect 2881 8123 2933 8140
rect 34 8106 2933 8123
rect 2967 8106 3002 8140
rect 3036 8106 3071 8140
rect 3105 8106 3139 8140
rect 3173 8106 3207 8140
rect 3241 8106 3275 8140
rect 3309 8106 3343 8140
rect 3377 8106 3411 8140
rect 3445 8106 3479 8140
rect 3513 8106 3547 8140
rect 3581 8106 3615 8140
rect 3649 8106 3683 8140
rect 3717 8106 3751 8140
rect 3785 8106 3819 8140
rect 3853 8106 3887 8140
rect 3921 8106 3955 8140
rect 3989 8106 4023 8140
rect 4057 8106 4091 8140
rect 4125 8106 4159 8140
rect 4193 8106 4227 8140
rect 4261 8106 4295 8140
rect 4329 8106 4363 8140
rect 4397 8106 4431 8140
rect 4465 8106 4499 8140
rect 4533 8106 4567 8140
rect 4601 8106 4635 8140
rect 4669 8106 4703 8140
rect 4737 8106 4771 8140
rect 4805 8106 4839 8140
rect 4873 8106 4907 8140
rect 4941 8106 4975 8140
rect 5009 8106 5043 8140
rect 5077 8106 5111 8140
rect 5145 8106 5179 8140
rect 5213 8106 5247 8140
rect 5281 8106 5315 8140
rect 5349 8106 5383 8140
rect 5417 8106 5451 8140
rect 5485 8106 5519 8140
rect 5553 8106 5587 8140
rect 5621 8106 5655 8140
rect 5689 8106 5723 8140
rect 5757 8106 5791 8140
rect 5825 8106 5859 8140
rect 5893 8106 5927 8140
rect 5961 8106 5995 8140
rect 6029 8106 6063 8140
rect 6097 8106 6131 8140
rect 6165 8106 6199 8140
rect 6233 8106 6267 8140
rect 6301 8106 6335 8140
rect 6369 8106 6403 8140
rect 6437 8106 6471 8140
rect 6505 8106 6539 8140
rect 6573 8106 6607 8140
rect 6641 8106 6675 8140
rect 6709 8106 6743 8140
rect 6777 8106 6811 8140
rect 6845 8106 6879 8140
rect 6913 8106 6947 8140
rect 6981 8106 7015 8140
rect 7049 8106 7083 8140
rect 7117 8106 7151 8140
rect 7185 8106 7219 8140
rect 7253 8106 7287 8140
rect 7321 8106 7355 8140
rect 7389 8106 7423 8140
rect 7457 8106 7491 8140
rect 7525 8106 7559 8140
rect 7593 8106 7627 8140
rect 7661 8106 7695 8140
rect 7729 8106 7763 8140
rect 7797 8106 7831 8140
rect 7865 8106 7899 8140
rect 7933 8106 7967 8140
rect 8001 8106 8035 8140
rect 8069 8106 8103 8140
rect 8137 8106 8171 8140
rect 8205 8106 8239 8140
rect 8273 8106 8307 8140
rect 8341 8106 8375 8140
rect 34 8082 8375 8106
rect 34 8048 68 8082
rect 102 8048 138 8082
rect 172 8048 208 8082
rect 242 8048 278 8082
rect 312 8048 348 8082
rect 382 8048 418 8082
rect 452 8048 488 8082
rect 522 8048 558 8082
rect 592 8048 628 8082
rect 662 8048 698 8082
rect 732 8048 768 8082
rect 802 8048 838 8082
rect 872 8048 908 8082
rect 942 8048 978 8082
rect 1012 8048 1048 8082
rect 1082 8048 1118 8082
rect 1152 8048 1188 8082
rect 1222 8048 1258 8082
rect 1292 8048 1328 8082
rect 1362 8048 1398 8082
rect 1432 8048 1467 8082
rect 1501 8048 1536 8082
rect 1570 8048 1605 8082
rect 1639 8048 1674 8082
rect 1708 8048 1743 8082
rect 1777 8048 1812 8082
rect 1846 8048 1881 8082
rect 1915 8048 1950 8082
rect 1984 8048 2019 8082
rect 2053 8048 2088 8082
rect 2122 8048 2157 8082
rect 2191 8048 2226 8082
rect 2260 8048 2295 8082
rect 2329 8048 2364 8082
rect 2398 8048 2433 8082
rect 2467 8048 2502 8082
rect 2536 8048 2571 8082
rect 2605 8048 2640 8082
rect 2674 8048 2709 8082
rect 2743 8048 2778 8082
rect 2812 8048 2847 8082
rect 2881 8070 8375 8082
rect 2881 8048 2933 8070
rect 34 8036 2933 8048
rect 2967 8036 3002 8070
rect 3036 8036 3071 8070
rect 3105 8036 3139 8070
rect 3173 8036 3207 8070
rect 3241 8036 3275 8070
rect 3309 8036 3343 8070
rect 3377 8036 3411 8070
rect 3445 8036 3479 8070
rect 3513 8036 3547 8070
rect 3581 8036 3615 8070
rect 3649 8036 3683 8070
rect 3717 8036 3751 8070
rect 3785 8036 3819 8070
rect 3853 8036 3887 8070
rect 3921 8036 3955 8070
rect 3989 8036 4023 8070
rect 4057 8036 4091 8070
rect 4125 8036 4159 8070
rect 4193 8036 4227 8070
rect 4261 8036 4295 8070
rect 4329 8036 4363 8070
rect 4397 8036 4431 8070
rect 4465 8036 4499 8070
rect 4533 8036 4567 8070
rect 4601 8036 4635 8070
rect 4669 8036 4703 8070
rect 4737 8036 4771 8070
rect 4805 8036 4839 8070
rect 4873 8036 4907 8070
rect 4941 8036 4975 8070
rect 5009 8036 5043 8070
rect 5077 8036 5111 8070
rect 5145 8036 5179 8070
rect 5213 8036 5247 8070
rect 5281 8036 5315 8070
rect 5349 8036 5383 8070
rect 5417 8036 5451 8070
rect 5485 8036 5519 8070
rect 5553 8036 5587 8070
rect 5621 8036 5655 8070
rect 5689 8036 5723 8070
rect 5757 8036 5791 8070
rect 5825 8036 5859 8070
rect 5893 8036 5927 8070
rect 5961 8036 5995 8070
rect 6029 8036 6063 8070
rect 6097 8036 6131 8070
rect 6165 8036 6199 8070
rect 6233 8036 6267 8070
rect 6301 8036 6335 8070
rect 6369 8036 6403 8070
rect 6437 8036 6471 8070
rect 6505 8036 6539 8070
rect 6573 8036 6607 8070
rect 6641 8036 6675 8070
rect 6709 8036 6743 8070
rect 6777 8036 6811 8070
rect 6845 8036 6879 8070
rect 6913 8036 6947 8070
rect 6981 8036 7015 8070
rect 7049 8036 7083 8070
rect 7117 8036 7151 8070
rect 7185 8036 7219 8070
rect 7253 8036 7287 8070
rect 7321 8036 7355 8070
rect 7389 8036 7423 8070
rect 7457 8036 7491 8070
rect 7525 8036 7559 8070
rect 7593 8036 7627 8070
rect 7661 8036 7695 8070
rect 7729 8036 7763 8070
rect 7797 8036 7831 8070
rect 7865 8036 7899 8070
rect 7933 8036 7967 8070
rect 8001 8036 8035 8070
rect 8069 8036 8103 8070
rect 8137 8036 8171 8070
rect 8205 8036 8239 8070
rect 8273 8036 8307 8070
rect 8341 8036 8375 8070
rect 34 8007 8375 8036
rect 34 7973 68 8007
rect 102 7973 138 8007
rect 172 7973 208 8007
rect 242 7973 278 8007
rect 312 7973 348 8007
rect 382 7973 418 8007
rect 452 7973 488 8007
rect 522 7973 558 8007
rect 592 7973 628 8007
rect 662 7973 698 8007
rect 732 7973 768 8007
rect 802 7973 838 8007
rect 872 7973 908 8007
rect 942 7973 978 8007
rect 1012 7973 1048 8007
rect 1082 7973 1118 8007
rect 1152 7973 1188 8007
rect 1222 7973 1258 8007
rect 1292 7973 1328 8007
rect 1362 7973 1398 8007
rect 1432 7973 1467 8007
rect 1501 7973 1536 8007
rect 1570 7973 1605 8007
rect 1639 7973 1674 8007
rect 1708 7973 1743 8007
rect 1777 7973 1812 8007
rect 1846 7973 1881 8007
rect 1915 7973 1950 8007
rect 1984 7973 2019 8007
rect 2053 7973 2088 8007
rect 2122 7973 2157 8007
rect 2191 7973 2226 8007
rect 2260 7973 2295 8007
rect 2329 7973 2364 8007
rect 2398 7973 2433 8007
rect 2467 7973 2502 8007
rect 2536 7973 2571 8007
rect 2605 7973 2640 8007
rect 2674 7973 2709 8007
rect 2743 7973 2778 8007
rect 2812 7973 2847 8007
rect 2881 8000 8375 8007
rect 2881 7973 2933 8000
rect 34 7966 2933 7973
rect 2967 7966 3002 8000
rect 3036 7966 3071 8000
rect 3105 7966 3139 8000
rect 3173 7966 3207 8000
rect 3241 7966 3275 8000
rect 3309 7966 3343 8000
rect 3377 7966 3411 8000
rect 3445 7966 3479 8000
rect 3513 7966 3547 8000
rect 3581 7966 3615 8000
rect 3649 7966 3683 8000
rect 3717 7966 3751 8000
rect 3785 7966 3819 8000
rect 3853 7966 3887 8000
rect 3921 7966 3955 8000
rect 3989 7966 4023 8000
rect 4057 7966 4091 8000
rect 4125 7966 4159 8000
rect 4193 7966 4227 8000
rect 4261 7966 4295 8000
rect 4329 7966 4363 8000
rect 4397 7966 4431 8000
rect 4465 7966 4499 8000
rect 4533 7966 4567 8000
rect 4601 7966 4635 8000
rect 4669 7966 4703 8000
rect 4737 7966 4771 8000
rect 4805 7966 4839 8000
rect 4873 7966 4907 8000
rect 4941 7966 4975 8000
rect 5009 7966 5043 8000
rect 5077 7966 5111 8000
rect 5145 7966 5179 8000
rect 5213 7966 5247 8000
rect 5281 7966 5315 8000
rect 5349 7966 5383 8000
rect 5417 7966 5451 8000
rect 5485 7966 5519 8000
rect 5553 7966 5587 8000
rect 5621 7966 5655 8000
rect 5689 7966 5723 8000
rect 5757 7966 5791 8000
rect 5825 7966 5859 8000
rect 5893 7966 5927 8000
rect 5961 7966 5995 8000
rect 6029 7966 6063 8000
rect 6097 7966 6131 8000
rect 6165 7966 6199 8000
rect 6233 7966 6267 8000
rect 6301 7966 6335 8000
rect 6369 7966 6403 8000
rect 6437 7966 6471 8000
rect 6505 7966 6539 8000
rect 6573 7966 6607 8000
rect 6641 7966 6675 8000
rect 6709 7966 6743 8000
rect 6777 7966 6811 8000
rect 6845 7966 6879 8000
rect 6913 7966 6947 8000
rect 6981 7966 7015 8000
rect 7049 7966 7083 8000
rect 7117 7966 7151 8000
rect 7185 7966 7219 8000
rect 7253 7966 7287 8000
rect 7321 7966 7355 8000
rect 7389 7966 7423 8000
rect 7457 7966 7491 8000
rect 7525 7966 7559 8000
rect 7593 7966 7627 8000
rect 7661 7966 7695 8000
rect 7729 7966 7763 8000
rect 7797 7966 7831 8000
rect 7865 7966 7899 8000
rect 7933 7966 7967 8000
rect 8001 7966 8035 8000
rect 8069 7966 8103 8000
rect 8137 7966 8171 8000
rect 8205 7966 8239 8000
rect 8273 7966 8307 8000
rect 8341 7966 8375 8000
rect 34 7932 8375 7966
rect 34 7898 68 7932
rect 102 7898 138 7932
rect 172 7898 208 7932
rect 242 7898 278 7932
rect 312 7898 348 7932
rect 382 7898 418 7932
rect 452 7898 488 7932
rect 522 7898 558 7932
rect 592 7898 628 7932
rect 662 7898 698 7932
rect 732 7898 768 7932
rect 802 7898 838 7932
rect 872 7898 908 7932
rect 942 7898 978 7932
rect 1012 7898 1048 7932
rect 1082 7898 1118 7932
rect 1152 7898 1188 7932
rect 1222 7898 1258 7932
rect 1292 7898 1328 7932
rect 1362 7898 1398 7932
rect 1432 7898 1467 7932
rect 1501 7898 1536 7932
rect 1570 7898 1605 7932
rect 1639 7898 1674 7932
rect 1708 7898 1743 7932
rect 1777 7898 1812 7932
rect 1846 7898 1881 7932
rect 1915 7898 1950 7932
rect 1984 7898 2019 7932
rect 2053 7898 2088 7932
rect 2122 7898 2157 7932
rect 2191 7898 2226 7932
rect 2260 7898 2295 7932
rect 2329 7898 2364 7932
rect 2398 7898 2433 7932
rect 2467 7898 2502 7932
rect 2536 7898 2571 7932
rect 2605 7898 2640 7932
rect 2674 7898 2709 7932
rect 2743 7898 2778 7932
rect 2812 7898 2847 7932
rect 2881 7930 8375 7932
rect 2881 7898 2933 7930
rect 34 7896 2933 7898
rect 2967 7896 3002 7930
rect 3036 7896 3071 7930
rect 3105 7896 3139 7930
rect 3173 7896 3207 7930
rect 3241 7896 3275 7930
rect 3309 7896 3343 7930
rect 3377 7896 3411 7930
rect 3445 7896 3479 7930
rect 3513 7896 3547 7930
rect 3581 7896 3615 7930
rect 3649 7896 3683 7930
rect 3717 7896 3751 7930
rect 3785 7896 3819 7930
rect 3853 7896 3887 7930
rect 3921 7896 3955 7930
rect 3989 7896 4023 7930
rect 4057 7896 4091 7930
rect 4125 7896 4159 7930
rect 4193 7896 4227 7930
rect 4261 7896 4295 7930
rect 4329 7896 4363 7930
rect 4397 7896 4431 7930
rect 4465 7896 4499 7930
rect 4533 7896 4567 7930
rect 4601 7896 4635 7930
rect 4669 7896 4703 7930
rect 4737 7896 4771 7930
rect 4805 7896 4839 7930
rect 4873 7896 4907 7930
rect 4941 7896 4975 7930
rect 5009 7896 5043 7930
rect 5077 7896 5111 7930
rect 5145 7896 5179 7930
rect 5213 7896 5247 7930
rect 5281 7896 5315 7930
rect 5349 7896 5383 7930
rect 5417 7896 5451 7930
rect 5485 7896 5519 7930
rect 5553 7896 5587 7930
rect 5621 7896 5655 7930
rect 5689 7896 5723 7930
rect 5757 7896 5791 7930
rect 5825 7896 5859 7930
rect 5893 7896 5927 7930
rect 5961 7896 5995 7930
rect 6029 7896 6063 7930
rect 6097 7896 6131 7930
rect 6165 7896 6199 7930
rect 6233 7896 6267 7930
rect 6301 7896 6335 7930
rect 6369 7896 6403 7930
rect 6437 7896 6471 7930
rect 6505 7896 6539 7930
rect 6573 7896 6607 7930
rect 6641 7896 6675 7930
rect 6709 7896 6743 7930
rect 6777 7896 6811 7930
rect 6845 7896 6879 7930
rect 6913 7896 6947 7930
rect 6981 7896 7015 7930
rect 7049 7896 7083 7930
rect 7117 7896 7151 7930
rect 7185 7896 7219 7930
rect 7253 7896 7287 7930
rect 7321 7896 7355 7930
rect 7389 7896 7423 7930
rect 7457 7896 7491 7930
rect 7525 7896 7559 7930
rect 7593 7896 7627 7930
rect 7661 7896 7695 7930
rect 7729 7896 7763 7930
rect 7797 7896 7831 7930
rect 7865 7896 7899 7930
rect 7933 7896 7967 7930
rect 8001 7896 8035 7930
rect 8069 7896 8103 7930
rect 8137 7896 8171 7930
rect 8205 7896 8239 7930
rect 8273 7896 8307 7930
rect 8341 7896 8375 7930
rect 34 7860 8375 7896
rect 13498 8283 14932 8289
rect 13498 8249 13532 8283
rect 13566 8249 13603 8283
rect 13637 8249 13674 8283
rect 13708 8249 13744 8283
rect 13778 8249 13814 8283
rect 13848 8249 13884 8283
rect 13918 8249 13954 8283
rect 13988 8249 14024 8283
rect 14058 8249 14094 8283
rect 14128 8249 14164 8283
rect 14198 8249 14234 8283
rect 14268 8249 14304 8283
rect 14338 8249 14374 8283
rect 14408 8249 14444 8283
rect 14478 8249 14514 8283
rect 14548 8249 14584 8283
rect 14618 8249 14654 8283
rect 14688 8249 14724 8283
rect 14758 8249 14794 8283
rect 14828 8249 14864 8283
rect 14898 8255 14932 8283
rect 14966 8255 15000 8289
rect 15034 8255 15068 8289
rect 14898 8249 15102 8255
rect 13498 8217 15102 8249
rect 13498 8209 14932 8217
rect 13498 8175 13532 8209
rect 13566 8175 13603 8209
rect 13637 8175 13674 8209
rect 13708 8175 13744 8209
rect 13778 8175 13814 8209
rect 13848 8175 13884 8209
rect 13918 8175 13954 8209
rect 13988 8175 14024 8209
rect 14058 8175 14094 8209
rect 14128 8175 14164 8209
rect 14198 8175 14234 8209
rect 14268 8175 14304 8209
rect 14338 8175 14374 8209
rect 14408 8175 14444 8209
rect 14478 8175 14514 8209
rect 14548 8175 14584 8209
rect 14618 8175 14654 8209
rect 14688 8175 14724 8209
rect 14758 8175 14794 8209
rect 14828 8175 14864 8209
rect 14898 8183 14932 8209
rect 14966 8183 15000 8217
rect 15034 8183 15068 8217
rect 14898 8175 15102 8183
rect 13498 8145 15102 8175
rect 13498 8135 14932 8145
rect 13498 8101 13532 8135
rect 13566 8101 13603 8135
rect 13637 8101 13674 8135
rect 13708 8101 13744 8135
rect 13778 8101 13814 8135
rect 13848 8101 13884 8135
rect 13918 8101 13954 8135
rect 13988 8101 14024 8135
rect 14058 8101 14094 8135
rect 14128 8101 14164 8135
rect 14198 8101 14234 8135
rect 14268 8101 14304 8135
rect 14338 8101 14374 8135
rect 14408 8101 14444 8135
rect 14478 8101 14514 8135
rect 14548 8101 14584 8135
rect 14618 8101 14654 8135
rect 14688 8101 14724 8135
rect 14758 8101 14794 8135
rect 14828 8101 14864 8135
rect 14898 8111 14932 8135
rect 14966 8111 15000 8145
rect 15034 8111 15068 8145
rect 14898 8101 15102 8111
rect 13498 8073 15102 8101
rect 13498 8061 14932 8073
rect 13498 8027 13532 8061
rect 13566 8027 13603 8061
rect 13637 8027 13674 8061
rect 13708 8027 13744 8061
rect 13778 8027 13814 8061
rect 13848 8027 13884 8061
rect 13918 8027 13954 8061
rect 13988 8027 14024 8061
rect 14058 8027 14094 8061
rect 14128 8027 14164 8061
rect 14198 8027 14234 8061
rect 14268 8027 14304 8061
rect 14338 8027 14374 8061
rect 14408 8027 14444 8061
rect 14478 8027 14514 8061
rect 14548 8027 14584 8061
rect 14618 8027 14654 8061
rect 14688 8027 14724 8061
rect 14758 8027 14794 8061
rect 14828 8027 14864 8061
rect 14898 8039 14932 8061
rect 14966 8039 15000 8073
rect 15034 8039 15068 8073
rect 14898 8027 15102 8039
rect 13498 8001 15102 8027
rect 13498 7987 14932 8001
rect 13498 7953 13532 7987
rect 13566 7953 13603 7987
rect 13637 7953 13674 7987
rect 13708 7953 13744 7987
rect 13778 7953 13814 7987
rect 13848 7953 13884 7987
rect 13918 7953 13954 7987
rect 13988 7953 14024 7987
rect 14058 7953 14094 7987
rect 14128 7953 14164 7987
rect 14198 7953 14234 7987
rect 14268 7953 14304 7987
rect 14338 7953 14374 7987
rect 14408 7953 14444 7987
rect 14478 7953 14514 7987
rect 14548 7953 14584 7987
rect 14618 7953 14654 7987
rect 14688 7953 14724 7987
rect 14758 7953 14794 7987
rect 14828 7953 14864 7987
rect 14898 7967 14932 7987
rect 14966 7967 15000 8001
rect 15034 7967 15068 8001
rect 14898 7953 15102 7967
rect 13498 7929 15102 7953
rect 13498 7913 14932 7929
rect 34 7857 2933 7860
rect 34 7823 68 7857
rect 102 7823 138 7857
rect 172 7823 208 7857
rect 242 7823 278 7857
rect 312 7823 348 7857
rect 382 7823 418 7857
rect 452 7823 488 7857
rect 522 7823 558 7857
rect 592 7823 628 7857
rect 662 7823 698 7857
rect 732 7823 768 7857
rect 802 7823 838 7857
rect 872 7823 908 7857
rect 942 7823 978 7857
rect 1012 7823 1048 7857
rect 1082 7823 1118 7857
rect 1152 7823 1188 7857
rect 1222 7823 1258 7857
rect 1292 7823 1328 7857
rect 1362 7823 1398 7857
rect 1432 7823 1467 7857
rect 1501 7823 1536 7857
rect 1570 7823 1605 7857
rect 1639 7823 1674 7857
rect 1708 7823 1743 7857
rect 1777 7823 1812 7857
rect 1846 7823 1881 7857
rect 1915 7823 1950 7857
rect 1984 7823 2019 7857
rect 2053 7823 2088 7857
rect 2122 7823 2157 7857
rect 2191 7823 2226 7857
rect 2260 7823 2295 7857
rect 2329 7823 2364 7857
rect 2398 7823 2433 7857
rect 2467 7823 2502 7857
rect 2536 7823 2571 7857
rect 2605 7823 2640 7857
rect 2674 7823 2709 7857
rect 2743 7823 2778 7857
rect 2812 7823 2847 7857
rect 2881 7826 2933 7857
rect 2967 7826 3002 7860
rect 3036 7826 3071 7860
rect 3105 7826 3139 7860
rect 3173 7826 3207 7860
rect 3241 7826 3275 7860
rect 3309 7826 3343 7860
rect 3377 7826 3411 7860
rect 3445 7826 3479 7860
rect 3513 7826 3547 7860
rect 3581 7826 3615 7860
rect 3649 7826 3683 7860
rect 3717 7826 3751 7860
rect 3785 7826 3819 7860
rect 3853 7826 3887 7860
rect 3921 7826 3955 7860
rect 3989 7826 4023 7860
rect 4057 7826 4091 7860
rect 4125 7826 4159 7860
rect 4193 7826 4227 7860
rect 4261 7826 4295 7860
rect 4329 7826 4363 7860
rect 4397 7826 4431 7860
rect 4465 7826 4499 7860
rect 4533 7826 4567 7860
rect 4601 7826 4635 7860
rect 4669 7826 4703 7860
rect 4737 7826 4771 7860
rect 4805 7826 4839 7860
rect 4873 7826 4907 7860
rect 4941 7826 4975 7860
rect 5009 7826 5043 7860
rect 5077 7826 5111 7860
rect 5145 7826 5179 7860
rect 5213 7826 5247 7860
rect 5281 7826 5315 7860
rect 5349 7826 5383 7860
rect 5417 7826 5451 7860
rect 5485 7826 5519 7860
rect 5553 7826 5587 7860
rect 5621 7826 5655 7860
rect 5689 7826 5723 7860
rect 5757 7826 5791 7860
rect 5825 7826 5859 7860
rect 5893 7826 5927 7860
rect 5961 7826 5995 7860
rect 6029 7826 6063 7860
rect 6097 7826 6131 7860
rect 6165 7826 6199 7860
rect 6233 7826 6267 7860
rect 6301 7826 6335 7860
rect 6369 7826 6403 7860
rect 6437 7826 6471 7860
rect 6505 7826 6539 7860
rect 6573 7826 6607 7860
rect 6641 7826 6675 7860
rect 6709 7826 6743 7860
rect 6777 7826 6811 7860
rect 6845 7826 6879 7860
rect 6913 7826 6947 7860
rect 6981 7826 7015 7860
rect 7049 7826 7083 7860
rect 7117 7826 7151 7860
rect 7185 7826 7219 7860
rect 7253 7826 7287 7860
rect 7321 7826 7355 7860
rect 7389 7826 7423 7860
rect 7457 7826 7491 7860
rect 7525 7826 7559 7860
rect 7593 7826 7627 7860
rect 7661 7826 7695 7860
rect 7729 7826 7763 7860
rect 7797 7826 7831 7860
rect 7865 7826 7899 7860
rect 7933 7826 7967 7860
rect 8001 7826 8035 7860
rect 8069 7826 8103 7860
rect 8137 7826 8171 7860
rect 8205 7826 8239 7860
rect 8273 7826 8307 7860
rect 8341 7826 8375 7860
rect 2881 7823 8375 7826
rect 34 7788 8375 7823
rect 13498 7879 13532 7913
rect 13566 7879 13603 7913
rect 13637 7879 13674 7913
rect 13708 7879 13744 7913
rect 13778 7879 13814 7913
rect 13848 7879 13884 7913
rect 13918 7879 13954 7913
rect 13988 7879 14024 7913
rect 14058 7879 14094 7913
rect 14128 7879 14164 7913
rect 14198 7879 14234 7913
rect 14268 7879 14304 7913
rect 14338 7879 14374 7913
rect 14408 7879 14444 7913
rect 14478 7879 14514 7913
rect 14548 7879 14584 7913
rect 14618 7879 14654 7913
rect 14688 7879 14724 7913
rect 14758 7879 14794 7913
rect 14828 7879 14864 7913
rect 14898 7895 14932 7913
rect 14966 7895 15000 7929
rect 15034 7895 15068 7929
rect 14898 7879 15102 7895
rect 13498 7857 15102 7879
rect 13498 7839 14932 7857
rect 13498 7805 13532 7839
rect 13566 7805 13603 7839
rect 13637 7805 13674 7839
rect 13708 7805 13744 7839
rect 13778 7805 13814 7839
rect 13848 7805 13884 7839
rect 13918 7805 13954 7839
rect 13988 7805 14024 7839
rect 14058 7805 14094 7839
rect 14128 7805 14164 7839
rect 14198 7805 14234 7839
rect 14268 7805 14304 7839
rect 14338 7805 14374 7839
rect 14408 7805 14444 7839
rect 14478 7805 14514 7839
rect 14548 7805 14584 7839
rect 14618 7805 14654 7839
rect 14688 7805 14724 7839
rect 14758 7805 14794 7839
rect 14828 7805 14864 7839
rect 14898 7823 14932 7839
rect 14966 7823 15000 7857
rect 15034 7823 15068 7857
rect 14898 7805 15102 7823
rect 13498 7788 15102 7805
rect 34 7785 15102 7788
rect 34 7751 14932 7785
rect 14966 7751 15000 7785
rect 15034 7751 15068 7785
rect 34 7749 15102 7751
rect 34 7715 68 7749
rect 102 7715 137 7749
rect 171 7715 206 7749
rect 240 7715 275 7749
rect 309 7715 344 7749
rect 378 7715 413 7749
rect 447 7715 482 7749
rect 516 7715 551 7749
rect 585 7715 620 7749
rect 654 7715 689 7749
rect 723 7715 758 7749
rect 792 7715 827 7749
rect 861 7715 896 7749
rect 930 7715 965 7749
rect 999 7715 1034 7749
rect 1068 7715 1103 7749
rect 1137 7715 1172 7749
rect 1206 7715 1241 7749
rect 1275 7715 1310 7749
rect 1344 7715 1379 7749
rect 1413 7715 1448 7749
rect 1482 7715 1517 7749
rect 1551 7715 1586 7749
rect 1620 7715 1655 7749
rect 1689 7715 1724 7749
rect 1758 7715 1793 7749
rect 1827 7715 1862 7749
rect 1896 7715 1931 7749
rect 1965 7715 2000 7749
rect 2034 7715 2069 7749
rect 2103 7715 2138 7749
rect 2172 7715 2207 7749
rect 2241 7715 2276 7749
rect 2310 7715 2345 7749
rect 2379 7715 2414 7749
rect 2448 7715 2483 7749
rect 2517 7715 2552 7749
rect 2586 7715 2621 7749
rect 2655 7715 2690 7749
rect 2724 7715 2759 7749
rect 2793 7715 2828 7749
rect 2862 7715 2896 7749
rect 2930 7715 2964 7749
rect 2998 7715 3032 7749
rect 3066 7715 3100 7749
rect 3134 7715 3168 7749
rect 3202 7715 3236 7749
rect 3270 7715 3304 7749
rect 3338 7715 3372 7749
rect 3406 7715 3440 7749
rect 3474 7715 3508 7749
rect 3542 7715 3576 7749
rect 3610 7715 3644 7749
rect 3678 7715 3712 7749
rect 3746 7715 3780 7749
rect 3814 7715 3848 7749
rect 3882 7715 3916 7749
rect 3950 7715 3984 7749
rect 4018 7715 4052 7749
rect 4086 7715 4120 7749
rect 4154 7715 4188 7749
rect 4222 7715 4256 7749
rect 4290 7715 4324 7749
rect 4358 7715 4392 7749
rect 4426 7715 4460 7749
rect 4494 7715 4528 7749
rect 4562 7715 4596 7749
rect 4630 7715 4664 7749
rect 4698 7715 4732 7749
rect 4766 7715 4800 7749
rect 4834 7715 4868 7749
rect 4902 7715 4936 7749
rect 4970 7715 5004 7749
rect 5038 7715 5072 7749
rect 5106 7715 5140 7749
rect 5174 7715 5208 7749
rect 5242 7715 5276 7749
rect 5310 7715 5344 7749
rect 5378 7715 5412 7749
rect 5446 7715 5480 7749
rect 5514 7715 5548 7749
rect 5582 7715 5616 7749
rect 5650 7715 5684 7749
rect 5718 7715 5752 7749
rect 5786 7715 5820 7749
rect 5854 7715 5888 7749
rect 5922 7715 5956 7749
rect 5990 7715 6024 7749
rect 6058 7715 6092 7749
rect 6126 7715 6160 7749
rect 6194 7715 6228 7749
rect 6262 7715 6296 7749
rect 6330 7715 6364 7749
rect 6398 7715 6432 7749
rect 6466 7715 6500 7749
rect 6534 7715 6568 7749
rect 6602 7715 6636 7749
rect 6670 7715 6704 7749
rect 6738 7715 6772 7749
rect 6806 7715 6840 7749
rect 6874 7715 6908 7749
rect 6942 7715 6976 7749
rect 7010 7715 7044 7749
rect 7078 7715 7112 7749
rect 7146 7715 7180 7749
rect 7214 7715 7248 7749
rect 7282 7715 7316 7749
rect 7350 7715 7384 7749
rect 7418 7715 7452 7749
rect 7486 7715 7520 7749
rect 7554 7715 7588 7749
rect 7622 7715 7656 7749
rect 7690 7715 7724 7749
rect 7758 7715 7792 7749
rect 7826 7715 7860 7749
rect 7894 7715 7928 7749
rect 7962 7715 7996 7749
rect 8030 7715 8064 7749
rect 8098 7715 8132 7749
rect 8166 7715 8200 7749
rect 8234 7715 8268 7749
rect 8302 7715 8336 7749
rect 8370 7715 8404 7749
rect 8438 7715 8472 7749
rect 8506 7715 8540 7749
rect 8574 7715 8608 7749
rect 8642 7715 8676 7749
rect 8710 7715 8744 7749
rect 8778 7715 8812 7749
rect 8846 7715 8880 7749
rect 8914 7715 8948 7749
rect 8982 7715 9016 7749
rect 9050 7715 9084 7749
rect 9118 7715 9152 7749
rect 9186 7715 9220 7749
rect 9254 7715 9288 7749
rect 9322 7715 9356 7749
rect 9390 7715 9424 7749
rect 9458 7715 9492 7749
rect 9526 7715 9560 7749
rect 9594 7715 9628 7749
rect 9662 7715 9696 7749
rect 9730 7715 9764 7749
rect 9798 7715 9832 7749
rect 9866 7715 9900 7749
rect 9934 7715 9968 7749
rect 10002 7715 10036 7749
rect 10070 7715 10104 7749
rect 10138 7715 10172 7749
rect 10206 7715 10240 7749
rect 10274 7715 10308 7749
rect 10342 7715 10376 7749
rect 10410 7715 10444 7749
rect 10478 7715 10512 7749
rect 10546 7715 10580 7749
rect 10614 7715 10648 7749
rect 10682 7715 10716 7749
rect 10750 7715 10784 7749
rect 10818 7715 10852 7749
rect 10886 7715 10920 7749
rect 10954 7715 10988 7749
rect 11022 7715 11056 7749
rect 11090 7715 11124 7749
rect 11158 7715 11192 7749
rect 11226 7715 11260 7749
rect 11294 7715 11328 7749
rect 11362 7715 11396 7749
rect 11430 7715 11464 7749
rect 11498 7715 11532 7749
rect 11566 7715 11600 7749
rect 11634 7715 11668 7749
rect 11702 7715 11736 7749
rect 11770 7715 11804 7749
rect 11838 7715 11872 7749
rect 11906 7715 11940 7749
rect 11974 7715 12008 7749
rect 12042 7715 12076 7749
rect 12110 7715 12144 7749
rect 12178 7715 12212 7749
rect 12246 7715 12280 7749
rect 12314 7715 12348 7749
rect 12382 7715 12416 7749
rect 12450 7715 12484 7749
rect 12518 7715 12552 7749
rect 12586 7715 12620 7749
rect 12654 7715 12688 7749
rect 12722 7715 12756 7749
rect 12790 7715 12824 7749
rect 12858 7715 12892 7749
rect 12926 7715 12960 7749
rect 12994 7715 13028 7749
rect 13062 7715 13096 7749
rect 13130 7715 13164 7749
rect 13198 7715 13232 7749
rect 13266 7715 13300 7749
rect 13334 7715 13368 7749
rect 13402 7715 13436 7749
rect 13470 7715 13504 7749
rect 13538 7715 13572 7749
rect 13606 7715 13640 7749
rect 13674 7715 13708 7749
rect 13742 7715 13776 7749
rect 13810 7715 13844 7749
rect 13878 7715 13912 7749
rect 13946 7715 13980 7749
rect 14014 7715 14048 7749
rect 14082 7715 14116 7749
rect 14150 7715 14184 7749
rect 14218 7715 14252 7749
rect 14286 7715 14320 7749
rect 14354 7715 14388 7749
rect 14422 7715 14456 7749
rect 14490 7715 14524 7749
rect 14558 7715 14592 7749
rect 14626 7715 14660 7749
rect 14694 7715 14728 7749
rect 14762 7715 14796 7749
rect 14830 7715 14864 7749
rect 14898 7715 15102 7749
rect 34 7713 15102 7715
rect 34 7679 14932 7713
rect 14966 7679 15000 7713
rect 15034 7679 15068 7713
rect 34 7676 15102 7679
rect 34 7642 2733 7676
rect 34 7608 68 7642
rect 102 7608 137 7642
rect 171 7608 206 7642
rect 240 7608 275 7642
rect 309 7608 344 7642
rect 378 7608 413 7642
rect 447 7608 482 7642
rect 516 7608 551 7642
rect 585 7608 620 7642
rect 654 7608 689 7642
rect 723 7608 758 7642
rect 792 7608 827 7642
rect 861 7608 896 7642
rect 930 7608 965 7642
rect 999 7608 1033 7642
rect 1067 7608 1101 7642
rect 1135 7608 1169 7642
rect 1203 7608 1237 7642
rect 1271 7608 1305 7642
rect 1339 7608 1373 7642
rect 1407 7608 1441 7642
rect 1475 7608 1509 7642
rect 1543 7608 1577 7642
rect 1611 7608 1645 7642
rect 1679 7608 1713 7642
rect 1747 7608 1781 7642
rect 1815 7608 1849 7642
rect 1883 7608 1917 7642
rect 1951 7608 1985 7642
rect 2019 7608 2053 7642
rect 2087 7608 2121 7642
rect 2155 7608 2189 7642
rect 2223 7608 2257 7642
rect 2291 7608 2325 7642
rect 2359 7608 2393 7642
rect 2427 7608 2461 7642
rect 2495 7608 2529 7642
rect 2563 7608 2597 7642
rect 2631 7608 2665 7642
rect 2699 7608 2733 7642
rect 34 7570 2733 7608
rect 34 7536 68 7570
rect 102 7536 137 7570
rect 171 7536 206 7570
rect 240 7536 275 7570
rect 309 7536 344 7570
rect 378 7536 413 7570
rect 447 7536 482 7570
rect 516 7536 551 7570
rect 585 7536 620 7570
rect 654 7536 689 7570
rect 723 7536 758 7570
rect 792 7536 827 7570
rect 861 7536 896 7570
rect 930 7536 965 7570
rect 999 7536 1033 7570
rect 1067 7536 1101 7570
rect 1135 7536 1169 7570
rect 1203 7536 1237 7570
rect 1271 7536 1305 7570
rect 1339 7536 1373 7570
rect 1407 7536 1441 7570
rect 1475 7536 1509 7570
rect 1543 7536 1577 7570
rect 1611 7536 1645 7570
rect 1679 7536 1713 7570
rect 1747 7536 1781 7570
rect 1815 7536 1849 7570
rect 1883 7536 1917 7570
rect 1951 7536 1985 7570
rect 2019 7536 2053 7570
rect 2087 7536 2121 7570
rect 2155 7536 2189 7570
rect 2223 7536 2257 7570
rect 2291 7536 2325 7570
rect 2359 7536 2393 7570
rect 2427 7536 2461 7570
rect 2495 7536 2529 7570
rect 2563 7536 2597 7570
rect 2631 7536 2665 7570
rect 2699 7536 2733 7570
rect 34 7498 2733 7536
rect 34 7464 68 7498
rect 102 7464 137 7498
rect 171 7464 206 7498
rect 240 7464 275 7498
rect 309 7464 344 7498
rect 378 7464 413 7498
rect 447 7464 482 7498
rect 516 7464 551 7498
rect 585 7464 620 7498
rect 654 7464 689 7498
rect 723 7464 758 7498
rect 792 7464 827 7498
rect 861 7464 896 7498
rect 930 7464 965 7498
rect 999 7464 1033 7498
rect 1067 7464 1101 7498
rect 1135 7464 1169 7498
rect 1203 7464 1237 7498
rect 1271 7464 1305 7498
rect 1339 7464 1373 7498
rect 1407 7464 1441 7498
rect 1475 7464 1509 7498
rect 1543 7464 1577 7498
rect 1611 7464 1645 7498
rect 1679 7464 1713 7498
rect 1747 7464 1781 7498
rect 1815 7464 1849 7498
rect 1883 7464 1917 7498
rect 1951 7464 1985 7498
rect 2019 7464 2053 7498
rect 2087 7464 2121 7498
rect 2155 7464 2189 7498
rect 2223 7464 2257 7498
rect 2291 7464 2325 7498
rect 2359 7464 2393 7498
rect 2427 7464 2461 7498
rect 2495 7464 2529 7498
rect 2563 7464 2597 7498
rect 2631 7464 2665 7498
rect 2699 7464 2733 7498
rect 34 7426 2733 7464
rect 34 7392 68 7426
rect 102 7392 137 7426
rect 171 7392 206 7426
rect 240 7392 275 7426
rect 309 7392 344 7426
rect 378 7392 413 7426
rect 447 7392 482 7426
rect 516 7392 551 7426
rect 585 7392 620 7426
rect 654 7392 689 7426
rect 723 7392 758 7426
rect 792 7392 827 7426
rect 861 7392 896 7426
rect 930 7392 965 7426
rect 999 7392 1033 7426
rect 1067 7392 1101 7426
rect 1135 7392 1169 7426
rect 1203 7392 1237 7426
rect 1271 7392 1305 7426
rect 1339 7392 1373 7426
rect 1407 7392 1441 7426
rect 1475 7392 1509 7426
rect 1543 7392 1577 7426
rect 1611 7392 1645 7426
rect 1679 7392 1713 7426
rect 1747 7392 1781 7426
rect 1815 7392 1849 7426
rect 1883 7392 1917 7426
rect 1951 7392 1985 7426
rect 2019 7392 2053 7426
rect 2087 7392 2121 7426
rect 2155 7392 2189 7426
rect 2223 7392 2257 7426
rect 2291 7392 2325 7426
rect 2359 7392 2393 7426
rect 2427 7392 2461 7426
rect 2495 7392 2529 7426
rect 2563 7392 2597 7426
rect 2631 7392 2665 7426
rect 2699 7392 2733 7426
rect 34 7354 2733 7392
rect 34 7320 68 7354
rect 102 7320 137 7354
rect 171 7320 206 7354
rect 240 7320 275 7354
rect 309 7320 344 7354
rect 378 7320 413 7354
rect 447 7320 482 7354
rect 516 7320 551 7354
rect 585 7320 620 7354
rect 654 7320 689 7354
rect 723 7320 758 7354
rect 792 7320 827 7354
rect 861 7320 896 7354
rect 930 7320 965 7354
rect 999 7320 1033 7354
rect 1067 7320 1101 7354
rect 1135 7320 1169 7354
rect 1203 7320 1237 7354
rect 1271 7320 1305 7354
rect 1339 7320 1373 7354
rect 1407 7320 1441 7354
rect 1475 7320 1509 7354
rect 1543 7320 1577 7354
rect 1611 7320 1645 7354
rect 1679 7320 1713 7354
rect 1747 7320 1781 7354
rect 1815 7320 1849 7354
rect 1883 7320 1917 7354
rect 1951 7320 1985 7354
rect 2019 7320 2053 7354
rect 2087 7320 2121 7354
rect 2155 7320 2189 7354
rect 2223 7320 2257 7354
rect 2291 7320 2325 7354
rect 2359 7320 2393 7354
rect 2427 7320 2461 7354
rect 2495 7320 2529 7354
rect 2563 7320 2597 7354
rect 2631 7320 2665 7354
rect 2699 7320 2733 7354
rect 34 7282 2733 7320
rect 12490 7641 15102 7676
rect 12490 7640 14932 7641
rect 12490 7606 12524 7640
rect 12558 7606 12593 7640
rect 12627 7606 12662 7640
rect 12696 7606 12731 7640
rect 12765 7606 12800 7640
rect 12834 7606 12869 7640
rect 12903 7606 12938 7640
rect 12972 7606 13007 7640
rect 13041 7606 13076 7640
rect 13110 7606 13145 7640
rect 13179 7606 13214 7640
rect 13248 7606 13283 7640
rect 13317 7606 13352 7640
rect 13386 7606 13421 7640
rect 13455 7606 13490 7640
rect 13524 7606 13559 7640
rect 13593 7606 13628 7640
rect 13662 7606 13697 7640
rect 13731 7606 13766 7640
rect 13800 7606 13835 7640
rect 13869 7606 13904 7640
rect 13938 7606 13973 7640
rect 14007 7606 14042 7640
rect 14076 7606 14111 7640
rect 14145 7606 14180 7640
rect 14214 7606 14249 7640
rect 14283 7606 14318 7640
rect 14352 7606 14387 7640
rect 14421 7606 14456 7640
rect 14490 7606 14524 7640
rect 14558 7606 14592 7640
rect 14626 7606 14660 7640
rect 14694 7606 14728 7640
rect 14762 7606 14796 7640
rect 14830 7606 14864 7640
rect 14898 7607 14932 7640
rect 14966 7607 15000 7641
rect 15034 7607 15068 7641
rect 14898 7606 15102 7607
rect 12490 7569 15102 7606
rect 12490 7556 14932 7569
rect 12490 7522 12524 7556
rect 12558 7522 12593 7556
rect 12627 7522 12662 7556
rect 12696 7522 12731 7556
rect 12765 7522 12800 7556
rect 12834 7522 12869 7556
rect 12903 7522 12938 7556
rect 12972 7522 13007 7556
rect 13041 7522 13076 7556
rect 13110 7522 13145 7556
rect 13179 7522 13214 7556
rect 13248 7522 13283 7556
rect 13317 7522 13352 7556
rect 13386 7522 13421 7556
rect 13455 7522 13490 7556
rect 13524 7522 13559 7556
rect 13593 7522 13628 7556
rect 13662 7522 13697 7556
rect 13731 7522 13766 7556
rect 13800 7522 13835 7556
rect 13869 7522 13904 7556
rect 13938 7522 13973 7556
rect 14007 7522 14042 7556
rect 14076 7522 14111 7556
rect 14145 7522 14180 7556
rect 14214 7522 14249 7556
rect 14283 7522 14318 7556
rect 14352 7522 14387 7556
rect 14421 7522 14456 7556
rect 14490 7522 14524 7556
rect 14558 7522 14592 7556
rect 14626 7522 14660 7556
rect 14694 7522 14728 7556
rect 14762 7522 14796 7556
rect 14830 7522 14864 7556
rect 14898 7535 14932 7556
rect 14966 7535 15000 7569
rect 15034 7535 15068 7569
rect 14898 7522 15102 7535
rect 12490 7497 15102 7522
rect 12490 7472 14932 7497
rect 12490 7438 12524 7472
rect 12558 7438 12593 7472
rect 12627 7438 12662 7472
rect 12696 7438 12731 7472
rect 12765 7438 12800 7472
rect 12834 7438 12869 7472
rect 12903 7438 12938 7472
rect 12972 7438 13007 7472
rect 13041 7438 13076 7472
rect 13110 7438 13145 7472
rect 13179 7438 13214 7472
rect 13248 7438 13283 7472
rect 13317 7438 13352 7472
rect 13386 7438 13421 7472
rect 13455 7438 13490 7472
rect 13524 7438 13559 7472
rect 13593 7438 13628 7472
rect 13662 7438 13697 7472
rect 13731 7438 13766 7472
rect 13800 7438 13835 7472
rect 13869 7438 13904 7472
rect 13938 7438 13973 7472
rect 14007 7438 14042 7472
rect 14076 7438 14111 7472
rect 14145 7438 14180 7472
rect 14214 7438 14249 7472
rect 14283 7438 14318 7472
rect 14352 7438 14387 7472
rect 14421 7438 14456 7472
rect 14490 7438 14524 7472
rect 14558 7438 14592 7472
rect 14626 7438 14660 7472
rect 14694 7438 14728 7472
rect 14762 7438 14796 7472
rect 14830 7438 14864 7472
rect 14898 7463 14932 7472
rect 14966 7463 15000 7497
rect 15034 7463 15068 7497
rect 14898 7438 15102 7463
rect 12490 7425 15102 7438
rect 12490 7391 14932 7425
rect 14966 7391 15000 7425
rect 15034 7391 15068 7425
rect 12490 7388 15102 7391
rect 12490 7354 12524 7388
rect 12558 7354 12593 7388
rect 12627 7354 12662 7388
rect 12696 7354 12731 7388
rect 12765 7354 12800 7388
rect 12834 7354 12869 7388
rect 12903 7354 12938 7388
rect 12972 7354 13007 7388
rect 13041 7354 13076 7388
rect 13110 7354 13145 7388
rect 13179 7354 13214 7388
rect 13248 7354 13283 7388
rect 13317 7354 13352 7388
rect 13386 7354 13421 7388
rect 13455 7354 13490 7388
rect 13524 7354 13559 7388
rect 13593 7354 13628 7388
rect 13662 7354 13697 7388
rect 13731 7354 13766 7388
rect 13800 7354 13835 7388
rect 13869 7354 13904 7388
rect 13938 7354 13973 7388
rect 14007 7354 14042 7388
rect 14076 7354 14111 7388
rect 14145 7354 14180 7388
rect 14214 7354 14249 7388
rect 14283 7354 14318 7388
rect 14352 7354 14387 7388
rect 14421 7354 14456 7388
rect 14490 7354 14524 7388
rect 14558 7354 14592 7388
rect 14626 7354 14660 7388
rect 14694 7354 14728 7388
rect 14762 7354 14796 7388
rect 14830 7354 14864 7388
rect 14898 7354 15102 7388
rect 12490 7353 15102 7354
rect 12490 7319 14932 7353
rect 14966 7319 15000 7353
rect 15034 7319 15068 7353
rect 12490 7317 15102 7319
rect 34 7248 68 7282
rect 102 7248 137 7282
rect 171 7248 206 7282
rect 240 7248 275 7282
rect 309 7248 344 7282
rect 378 7248 413 7282
rect 447 7248 482 7282
rect 516 7248 551 7282
rect 585 7248 620 7282
rect 654 7248 689 7282
rect 723 7248 758 7282
rect 792 7248 827 7282
rect 861 7248 896 7282
rect 930 7248 965 7282
rect 999 7248 1033 7282
rect 1067 7248 1101 7282
rect 1135 7248 1169 7282
rect 1203 7248 1237 7282
rect 1271 7248 1305 7282
rect 1339 7248 1373 7282
rect 1407 7248 1441 7282
rect 1475 7248 1509 7282
rect 1543 7248 1577 7282
rect 1611 7248 1645 7282
rect 1679 7248 1713 7282
rect 1747 7248 1781 7282
rect 1815 7248 1849 7282
rect 1883 7248 1917 7282
rect 1951 7248 1985 7282
rect 2019 7248 2053 7282
rect 2087 7248 2121 7282
rect 2155 7248 2189 7282
rect 2223 7248 2257 7282
rect 2291 7248 2325 7282
rect 2359 7248 2393 7282
rect 2427 7248 2461 7282
rect 2495 7248 2529 7282
rect 2563 7248 2597 7282
rect 2631 7248 2665 7282
rect 2699 7248 2733 7282
rect 34 7210 2733 7248
rect 34 7176 68 7210
rect 102 7176 137 7210
rect 171 7176 206 7210
rect 240 7176 275 7210
rect 309 7176 344 7210
rect 378 7176 413 7210
rect 447 7176 482 7210
rect 516 7176 551 7210
rect 585 7176 620 7210
rect 654 7176 689 7210
rect 723 7176 758 7210
rect 792 7176 827 7210
rect 861 7176 896 7210
rect 930 7176 965 7210
rect 999 7176 1033 7210
rect 1067 7176 1101 7210
rect 1135 7176 1169 7210
rect 1203 7176 1237 7210
rect 1271 7176 1305 7210
rect 1339 7176 1373 7210
rect 1407 7176 1441 7210
rect 1475 7176 1509 7210
rect 1543 7176 1577 7210
rect 1611 7176 1645 7210
rect 1679 7176 1713 7210
rect 1747 7176 1781 7210
rect 1815 7176 1849 7210
rect 1883 7176 1917 7210
rect 1951 7176 1985 7210
rect 2019 7176 2053 7210
rect 2087 7176 2121 7210
rect 2155 7176 2189 7210
rect 2223 7176 2257 7210
rect 2291 7176 2325 7210
rect 2359 7176 2393 7210
rect 2427 7176 2461 7210
rect 2495 7176 2529 7210
rect 2563 7176 2597 7210
rect 2631 7176 2665 7210
rect 2699 7176 2733 7210
rect 34 7138 2733 7176
rect 34 7104 68 7138
rect 102 7104 137 7138
rect 171 7104 206 7138
rect 240 7104 275 7138
rect 309 7104 344 7138
rect 378 7104 413 7138
rect 447 7104 482 7138
rect 516 7104 551 7138
rect 585 7104 620 7138
rect 654 7104 689 7138
rect 723 7104 758 7138
rect 792 7104 827 7138
rect 861 7104 896 7138
rect 930 7104 965 7138
rect 999 7104 1033 7138
rect 1067 7104 1101 7138
rect 1135 7104 1169 7138
rect 1203 7104 1237 7138
rect 1271 7104 1305 7138
rect 1339 7104 1373 7138
rect 1407 7104 1441 7138
rect 1475 7104 1509 7138
rect 1543 7104 1577 7138
rect 1611 7104 1645 7138
rect 1679 7104 1713 7138
rect 1747 7104 1781 7138
rect 1815 7104 1849 7138
rect 1883 7104 1917 7138
rect 1951 7104 1985 7138
rect 2019 7104 2053 7138
rect 2087 7104 2121 7138
rect 2155 7104 2189 7138
rect 2223 7104 2257 7138
rect 2291 7104 2325 7138
rect 2359 7104 2393 7138
rect 2427 7104 2461 7138
rect 2495 7104 2529 7138
rect 2563 7104 2597 7138
rect 2631 7104 2665 7138
rect 2699 7104 2733 7138
rect 34 7066 2733 7104
rect 34 7032 68 7066
rect 102 7032 137 7066
rect 171 7032 206 7066
rect 240 7032 275 7066
rect 309 7032 344 7066
rect 378 7032 413 7066
rect 447 7032 482 7066
rect 516 7032 551 7066
rect 585 7032 620 7066
rect 654 7032 689 7066
rect 723 7032 758 7066
rect 792 7032 827 7066
rect 861 7032 896 7066
rect 930 7032 965 7066
rect 999 7032 1033 7066
rect 1067 7032 1101 7066
rect 1135 7032 1169 7066
rect 1203 7032 1237 7066
rect 1271 7032 1305 7066
rect 1339 7032 1373 7066
rect 1407 7032 1441 7066
rect 1475 7032 1509 7066
rect 1543 7032 1577 7066
rect 1611 7032 1645 7066
rect 1679 7032 1713 7066
rect 1747 7032 1781 7066
rect 1815 7032 1849 7066
rect 1883 7032 1917 7066
rect 1951 7032 1985 7066
rect 2019 7032 2053 7066
rect 2087 7032 2121 7066
rect 2155 7032 2189 7066
rect 2223 7032 2257 7066
rect 2291 7032 2325 7066
rect 2359 7032 2393 7066
rect 2427 7032 2461 7066
rect 2495 7032 2529 7066
rect 2563 7032 2597 7066
rect 2631 7032 2665 7066
rect 2699 7063 2733 7066
rect 8176 7282 15102 7317
rect 8176 7248 8210 7282
rect 8244 7248 8279 7282
rect 8313 7248 8348 7282
rect 8382 7248 8417 7282
rect 8451 7248 8486 7282
rect 8520 7248 8555 7282
rect 8589 7248 8624 7282
rect 8658 7248 8693 7282
rect 8727 7248 8762 7282
rect 8796 7248 8831 7282
rect 8865 7248 8900 7282
rect 8934 7248 8969 7282
rect 9003 7248 9038 7282
rect 9072 7248 9107 7282
rect 9141 7248 9176 7282
rect 9210 7248 9245 7282
rect 9279 7248 9314 7282
rect 9348 7248 9383 7282
rect 9417 7248 9452 7282
rect 9486 7248 9521 7282
rect 9555 7248 9590 7282
rect 9624 7248 9659 7282
rect 9693 7248 9728 7282
rect 9762 7248 9797 7282
rect 9831 7248 9866 7282
rect 9900 7248 9935 7282
rect 9969 7248 10004 7282
rect 10038 7248 10073 7282
rect 10107 7248 10142 7282
rect 10176 7248 10211 7282
rect 10245 7248 10280 7282
rect 10314 7248 10349 7282
rect 10383 7248 10418 7282
rect 10452 7248 10487 7282
rect 10521 7248 10556 7282
rect 10590 7248 10625 7282
rect 10659 7248 10694 7282
rect 10728 7248 10763 7282
rect 10797 7248 10832 7282
rect 10866 7248 10901 7282
rect 10935 7248 10970 7282
rect 11004 7248 11039 7282
rect 11073 7248 11108 7282
rect 11142 7248 11177 7282
rect 11211 7248 11246 7282
rect 11280 7248 11315 7282
rect 11349 7248 11384 7282
rect 11418 7248 11453 7282
rect 11487 7248 11522 7282
rect 11556 7248 11591 7282
rect 11625 7248 11660 7282
rect 11694 7248 11729 7282
rect 11763 7248 11798 7282
rect 11832 7248 11867 7282
rect 11901 7248 11936 7282
rect 11970 7248 12005 7282
rect 12039 7248 12074 7282
rect 12108 7248 12143 7282
rect 12177 7248 12212 7282
rect 12246 7248 12280 7282
rect 12314 7248 12348 7282
rect 12382 7248 12416 7282
rect 12450 7248 12484 7282
rect 12518 7248 12552 7282
rect 12586 7248 12620 7282
rect 12654 7248 12688 7282
rect 12722 7248 12756 7282
rect 12790 7248 12824 7282
rect 12858 7248 12892 7282
rect 12926 7248 12960 7282
rect 12994 7248 13028 7282
rect 13062 7248 13096 7282
rect 13130 7248 13164 7282
rect 13198 7248 13232 7282
rect 13266 7248 13300 7282
rect 13334 7248 13368 7282
rect 13402 7248 13436 7282
rect 13470 7248 13504 7282
rect 13538 7248 13572 7282
rect 13606 7248 13640 7282
rect 13674 7248 13708 7282
rect 13742 7248 13776 7282
rect 13810 7248 13844 7282
rect 13878 7248 13912 7282
rect 13946 7248 13980 7282
rect 14014 7248 14048 7282
rect 14082 7248 14116 7282
rect 14150 7248 14184 7282
rect 14218 7248 14252 7282
rect 14286 7248 14320 7282
rect 14354 7248 14388 7282
rect 14422 7248 14456 7282
rect 14490 7248 14524 7282
rect 14558 7248 14592 7282
rect 14626 7248 14660 7282
rect 14694 7248 14728 7282
rect 14762 7248 14796 7282
rect 14830 7248 14864 7282
rect 14898 7281 15102 7282
rect 14898 7248 14932 7281
rect 8176 7247 14932 7248
rect 14966 7247 15000 7281
rect 15034 7247 15068 7281
rect 8176 7210 15102 7247
rect 8176 7176 8210 7210
rect 8244 7176 8279 7210
rect 8313 7176 8348 7210
rect 8382 7176 8417 7210
rect 8451 7176 8486 7210
rect 8520 7176 8555 7210
rect 8589 7176 8624 7210
rect 8658 7176 8693 7210
rect 8727 7176 8762 7210
rect 8796 7176 8831 7210
rect 8865 7176 8900 7210
rect 8934 7176 8969 7210
rect 9003 7176 9038 7210
rect 9072 7176 9107 7210
rect 9141 7176 9176 7210
rect 9210 7176 9245 7210
rect 9279 7176 9314 7210
rect 9348 7176 9383 7210
rect 9417 7176 9452 7210
rect 9486 7176 9521 7210
rect 9555 7176 9590 7210
rect 9624 7176 9659 7210
rect 9693 7176 9728 7210
rect 9762 7176 9797 7210
rect 9831 7176 9866 7210
rect 9900 7176 9935 7210
rect 9969 7176 10004 7210
rect 10038 7176 10073 7210
rect 10107 7176 10142 7210
rect 10176 7176 10211 7210
rect 10245 7176 10280 7210
rect 10314 7176 10349 7210
rect 10383 7176 10418 7210
rect 10452 7176 10487 7210
rect 10521 7176 10556 7210
rect 10590 7176 10625 7210
rect 10659 7176 10694 7210
rect 10728 7176 10763 7210
rect 10797 7176 10832 7210
rect 10866 7176 10901 7210
rect 10935 7176 10970 7210
rect 11004 7176 11039 7210
rect 11073 7176 11108 7210
rect 11142 7176 11177 7210
rect 11211 7176 11246 7210
rect 11280 7176 11315 7210
rect 11349 7176 11384 7210
rect 11418 7176 11453 7210
rect 11487 7176 11522 7210
rect 11556 7176 11591 7210
rect 11625 7176 11660 7210
rect 11694 7176 11729 7210
rect 11763 7176 11798 7210
rect 11832 7176 11867 7210
rect 11901 7176 11936 7210
rect 11970 7176 12005 7210
rect 12039 7176 12074 7210
rect 12108 7176 12143 7210
rect 12177 7176 12212 7210
rect 12246 7176 12280 7210
rect 12314 7176 12348 7210
rect 12382 7176 12416 7210
rect 12450 7176 12484 7210
rect 12518 7176 12552 7210
rect 12586 7176 12620 7210
rect 12654 7176 12688 7210
rect 12722 7176 12756 7210
rect 12790 7176 12824 7210
rect 12858 7176 12892 7210
rect 12926 7176 12960 7210
rect 12994 7176 13028 7210
rect 13062 7176 13096 7210
rect 13130 7176 13164 7210
rect 13198 7176 13232 7210
rect 13266 7176 13300 7210
rect 13334 7176 13368 7210
rect 13402 7176 13436 7210
rect 13470 7176 13504 7210
rect 13538 7176 13572 7210
rect 13606 7176 13640 7210
rect 13674 7176 13708 7210
rect 13742 7176 13776 7210
rect 13810 7176 13844 7210
rect 13878 7176 13912 7210
rect 13946 7176 13980 7210
rect 14014 7176 14048 7210
rect 14082 7176 14116 7210
rect 14150 7176 14184 7210
rect 14218 7176 14252 7210
rect 14286 7176 14320 7210
rect 14354 7176 14388 7210
rect 14422 7176 14456 7210
rect 14490 7176 14524 7210
rect 14558 7176 14592 7210
rect 14626 7176 14660 7210
rect 14694 7176 14728 7210
rect 14762 7176 14796 7210
rect 14830 7176 14864 7210
rect 14898 7209 15102 7210
rect 14898 7176 14932 7209
rect 8176 7175 14932 7176
rect 14966 7175 15000 7209
rect 15034 7175 15068 7209
rect 8176 7138 15102 7175
rect 8176 7104 8210 7138
rect 8244 7104 8279 7138
rect 8313 7104 8348 7138
rect 8382 7104 8417 7138
rect 8451 7104 8486 7138
rect 8520 7104 8555 7138
rect 8589 7104 8624 7138
rect 8658 7104 8693 7138
rect 8727 7104 8762 7138
rect 8796 7104 8831 7138
rect 8865 7104 8900 7138
rect 8934 7104 8969 7138
rect 9003 7104 9038 7138
rect 9072 7104 9107 7138
rect 9141 7104 9176 7138
rect 9210 7104 9245 7138
rect 9279 7104 9314 7138
rect 9348 7104 9383 7138
rect 9417 7104 9452 7138
rect 9486 7104 9521 7138
rect 9555 7104 9590 7138
rect 9624 7104 9659 7138
rect 9693 7104 9728 7138
rect 9762 7104 9797 7138
rect 9831 7104 9866 7138
rect 9900 7104 9935 7138
rect 9969 7104 10004 7138
rect 10038 7104 10073 7138
rect 10107 7104 10142 7138
rect 10176 7104 10211 7138
rect 10245 7104 10280 7138
rect 10314 7104 10349 7138
rect 10383 7104 10418 7138
rect 10452 7104 10487 7138
rect 10521 7104 10556 7138
rect 10590 7104 10625 7138
rect 10659 7104 10694 7138
rect 10728 7104 10763 7138
rect 10797 7104 10832 7138
rect 10866 7104 10901 7138
rect 10935 7104 10970 7138
rect 11004 7104 11039 7138
rect 11073 7104 11108 7138
rect 11142 7104 11177 7138
rect 11211 7104 11246 7138
rect 11280 7104 11315 7138
rect 11349 7104 11384 7138
rect 11418 7104 11453 7138
rect 11487 7104 11522 7138
rect 11556 7104 11591 7138
rect 11625 7104 11660 7138
rect 11694 7104 11729 7138
rect 11763 7104 11798 7138
rect 11832 7104 11867 7138
rect 11901 7104 11936 7138
rect 11970 7104 12005 7138
rect 12039 7104 12074 7138
rect 12108 7104 12143 7138
rect 12177 7104 12212 7138
rect 12246 7104 12280 7138
rect 12314 7104 12348 7138
rect 12382 7104 12416 7138
rect 12450 7104 12484 7138
rect 12518 7104 12552 7138
rect 12586 7104 12620 7138
rect 12654 7104 12688 7138
rect 12722 7104 12756 7138
rect 12790 7104 12824 7138
rect 12858 7104 12892 7138
rect 12926 7104 12960 7138
rect 12994 7104 13028 7138
rect 13062 7104 13096 7138
rect 13130 7104 13164 7138
rect 13198 7104 13232 7138
rect 13266 7104 13300 7138
rect 13334 7104 13368 7138
rect 13402 7104 13436 7138
rect 13470 7104 13504 7138
rect 13538 7104 13572 7138
rect 13606 7104 13640 7138
rect 13674 7104 13708 7138
rect 13742 7104 13776 7138
rect 13810 7104 13844 7138
rect 13878 7104 13912 7138
rect 13946 7104 13980 7138
rect 14014 7104 14048 7138
rect 14082 7104 14116 7138
rect 14150 7104 14184 7138
rect 14218 7104 14252 7138
rect 14286 7104 14320 7138
rect 14354 7104 14388 7138
rect 14422 7104 14456 7138
rect 14490 7104 14524 7138
rect 14558 7104 14592 7138
rect 14626 7104 14660 7138
rect 14694 7104 14728 7138
rect 14762 7104 14796 7138
rect 14830 7104 14864 7138
rect 14898 7137 15102 7138
rect 14898 7104 14932 7137
rect 8176 7103 14932 7104
rect 14966 7103 15000 7137
rect 15034 7103 15068 7137
rect 8176 7066 15102 7103
rect 2699 7047 7756 7063
rect 2699 7032 2757 7047
rect 34 7013 2757 7032
rect 2791 7013 2825 7047
rect 2859 7013 2893 7047
rect 2927 7013 2961 7047
rect 2995 7013 3029 7047
rect 3063 7013 3097 7047
rect 3131 7013 3165 7047
rect 3199 7013 3233 7047
rect 3267 7013 3301 7047
rect 3335 7013 3369 7047
rect 3403 7013 3437 7047
rect 3471 7013 3505 7047
rect 3539 7013 3573 7047
rect 3607 7013 3641 7047
rect 3675 7013 3709 7047
rect 3743 7013 3777 7047
rect 3811 7013 3845 7047
rect 3879 7013 3913 7047
rect 3947 7013 3981 7047
rect 4015 7013 4049 7047
rect 4083 7013 4117 7047
rect 4151 7013 4185 7047
rect 4219 7013 4253 7047
rect 4287 7013 4321 7047
rect 4355 7013 4389 7047
rect 4423 7013 4457 7047
rect 4491 7013 4525 7047
rect 4559 7013 4593 7047
rect 4627 7013 4661 7047
rect 4695 7013 4729 7047
rect 4763 7013 4797 7047
rect 4831 7013 4865 7047
rect 4899 7013 4933 7047
rect 4967 7013 5001 7047
rect 5035 7013 5069 7047
rect 5103 7013 5137 7047
rect 5171 7013 5205 7047
rect 5239 7013 5273 7047
rect 5307 7013 5341 7047
rect 5375 7013 5409 7047
rect 5443 7013 5477 7047
rect 5511 7013 5545 7047
rect 5579 7013 5613 7047
rect 5647 7013 5681 7047
rect 5715 7013 5749 7047
rect 5783 7013 5817 7047
rect 5851 7013 5885 7047
rect 5919 7013 5953 7047
rect 5987 7013 6021 7047
rect 6055 7013 6089 7047
rect 6123 7013 6157 7047
rect 6191 7013 6225 7047
rect 6259 7013 6293 7047
rect 6327 7013 6361 7047
rect 6395 7013 6429 7047
rect 6463 7013 6497 7047
rect 6531 7013 6565 7047
rect 6599 7013 6633 7047
rect 6667 7013 6701 7047
rect 6735 7013 6769 7047
rect 6803 7013 6837 7047
rect 6871 7013 6905 7047
rect 6939 7013 6973 7047
rect 7007 7013 7041 7047
rect 7075 7013 7109 7047
rect 7143 7013 7177 7047
rect 7211 7013 7245 7047
rect 7279 7013 7313 7047
rect 7347 7013 7381 7047
rect 7415 7013 7449 7047
rect 7483 7013 7517 7047
rect 7551 7013 7585 7047
rect 7619 7013 7653 7047
rect 7687 7013 7756 7047
rect 34 6997 7756 7013
rect 8176 7032 8210 7066
rect 8244 7032 8279 7066
rect 8313 7032 8348 7066
rect 8382 7032 8417 7066
rect 8451 7032 8486 7066
rect 8520 7032 8555 7066
rect 8589 7032 8624 7066
rect 8658 7032 8693 7066
rect 8727 7032 8762 7066
rect 8796 7032 8831 7066
rect 8865 7032 8900 7066
rect 8934 7032 8969 7066
rect 9003 7032 9038 7066
rect 9072 7032 9107 7066
rect 9141 7032 9176 7066
rect 9210 7032 9245 7066
rect 9279 7032 9314 7066
rect 9348 7032 9383 7066
rect 9417 7032 9452 7066
rect 9486 7032 9521 7066
rect 9555 7032 9590 7066
rect 9624 7032 9659 7066
rect 9693 7032 9728 7066
rect 9762 7032 9797 7066
rect 9831 7032 9866 7066
rect 9900 7032 9935 7066
rect 9969 7032 10004 7066
rect 10038 7032 10073 7066
rect 10107 7032 10142 7066
rect 10176 7032 10211 7066
rect 10245 7032 10280 7066
rect 10314 7032 10349 7066
rect 10383 7032 10418 7066
rect 10452 7032 10487 7066
rect 10521 7032 10556 7066
rect 10590 7032 10625 7066
rect 10659 7032 10694 7066
rect 10728 7032 10763 7066
rect 10797 7032 10832 7066
rect 10866 7032 10901 7066
rect 10935 7032 10970 7066
rect 11004 7032 11039 7066
rect 11073 7032 11108 7066
rect 11142 7032 11177 7066
rect 11211 7032 11246 7066
rect 11280 7032 11315 7066
rect 11349 7032 11384 7066
rect 11418 7032 11453 7066
rect 11487 7032 11522 7066
rect 11556 7032 11591 7066
rect 11625 7032 11660 7066
rect 11694 7032 11729 7066
rect 11763 7032 11798 7066
rect 11832 7032 11867 7066
rect 11901 7032 11936 7066
rect 11970 7032 12005 7066
rect 12039 7032 12074 7066
rect 12108 7032 12143 7066
rect 12177 7032 12212 7066
rect 12246 7032 12280 7066
rect 12314 7032 12348 7066
rect 12382 7032 12416 7066
rect 12450 7032 12484 7066
rect 12518 7032 12552 7066
rect 12586 7032 12620 7066
rect 12654 7032 12688 7066
rect 12722 7032 12756 7066
rect 12790 7032 12824 7066
rect 12858 7032 12892 7066
rect 12926 7032 12960 7066
rect 12994 7032 13028 7066
rect 13062 7032 13096 7066
rect 13130 7032 13164 7066
rect 13198 7032 13232 7066
rect 13266 7032 13300 7066
rect 13334 7032 13368 7066
rect 13402 7032 13436 7066
rect 13470 7032 13504 7066
rect 13538 7032 13572 7066
rect 13606 7032 13640 7066
rect 13674 7032 13708 7066
rect 13742 7032 13776 7066
rect 13810 7032 13844 7066
rect 13878 7032 13912 7066
rect 13946 7032 13980 7066
rect 14014 7032 14048 7066
rect 14082 7032 14116 7066
rect 14150 7032 14184 7066
rect 14218 7032 14252 7066
rect 14286 7032 14320 7066
rect 14354 7032 14388 7066
rect 14422 7032 14456 7066
rect 14490 7032 14524 7066
rect 14558 7032 14592 7066
rect 14626 7032 14660 7066
rect 14694 7032 14728 7066
rect 14762 7032 14796 7066
rect 14830 7032 14864 7066
rect 14898 7065 15102 7066
rect 14898 7032 14932 7065
rect 8176 7031 14932 7032
rect 14966 7031 15000 7065
rect 15034 7031 15068 7065
rect 8176 6997 15102 7031
<< mvpsubdiffcont >>
rect -932 9613 -898 9647
rect -864 9613 -830 9647
rect -796 9613 -762 9647
rect -723 9646 -689 9680
rect -654 9646 -620 9680
rect -585 9646 -551 9680
rect -516 9646 -482 9680
rect -447 9646 -413 9680
rect -378 9646 -344 9680
rect -309 9646 -275 9680
rect -240 9646 -206 9680
rect -171 9646 -137 9680
rect -102 9646 -68 9680
rect -723 9578 -689 9612
rect -654 9578 -620 9612
rect -585 9578 -551 9612
rect -516 9578 -482 9612
rect -447 9578 -413 9612
rect -378 9578 -344 9612
rect -309 9578 -275 9612
rect -240 9578 -206 9612
rect -171 9578 -137 9612
rect -102 9578 -68 9612
rect -932 9537 -898 9571
rect -864 9537 -830 9571
rect -796 9537 -762 9571
rect -723 9510 -689 9544
rect -654 9510 -620 9544
rect -585 9510 -551 9544
rect -516 9510 -482 9544
rect -447 9510 -413 9544
rect -378 9510 -344 9544
rect -309 9510 -275 9544
rect -240 9510 -206 9544
rect -171 9510 -137 9544
rect -102 9510 -68 9544
rect -932 9461 -898 9495
rect -864 9461 -830 9495
rect -796 9461 -762 9495
rect -723 9442 -689 9476
rect -654 9442 -620 9476
rect -585 9442 -551 9476
rect -516 9442 -482 9476
rect -447 9442 -413 9476
rect -378 9442 -344 9476
rect -309 9442 -275 9476
rect -240 9442 -206 9476
rect -171 9442 -137 9476
rect -102 9442 -68 9476
rect -932 9384 -898 9418
rect -864 9384 -830 9418
rect -796 9384 -762 9418
rect -723 9374 -689 9408
rect -654 9374 -620 9408
rect -585 9374 -551 9408
rect -516 9374 -482 9408
rect -447 9374 -413 9408
rect -378 9374 -344 9408
rect -309 9374 -275 9408
rect -240 9374 -206 9408
rect -171 9374 -137 9408
rect -102 9374 -68 9408
rect -932 9307 -898 9341
rect -864 9307 -830 9341
rect -796 9307 -762 9341
rect -723 9306 -689 9340
rect -654 9306 -620 9340
rect -585 9306 -551 9340
rect -516 9306 -482 9340
rect -447 9306 -413 9340
rect -378 9306 -344 9340
rect -309 9306 -275 9340
rect -240 9306 -206 9340
rect -171 9306 -137 9340
rect -102 9306 -68 9340
rect -932 9230 -898 9264
rect -864 9230 -830 9264
rect -796 9230 -762 9264
rect -723 9238 -689 9272
rect -654 9238 -620 9272
rect -585 9238 -551 9272
rect -516 9238 -482 9272
rect -447 9238 -413 9272
rect -378 9238 -344 9272
rect -309 9238 -275 9272
rect -240 9238 -206 9272
rect -171 9238 -137 9272
rect -102 9238 -68 9272
rect -932 9153 -898 9187
rect -864 9153 -830 9187
rect -796 9153 -762 9187
rect -723 9170 -689 9204
rect -654 9170 -620 9204
rect -585 9170 -551 9204
rect -516 9170 -482 9204
rect -447 9170 -413 9204
rect -378 9170 -344 9204
rect -309 9170 -275 9204
rect -240 9170 -206 9204
rect -171 9170 -137 9204
rect -102 9170 -68 9204
rect -932 9076 -898 9110
rect -864 9076 -830 9110
rect -796 9076 -762 9110
rect -723 9102 -689 9136
rect -654 9102 -620 9136
rect -585 9102 -551 9136
rect -516 9102 -482 9136
rect -447 9102 -413 9136
rect -378 9102 -344 9136
rect -309 9102 -275 9136
rect -240 9102 -206 9136
rect -171 9102 -137 9136
rect -102 9102 -68 9136
rect -723 9034 -689 9068
rect -654 9034 -620 9068
rect -585 9034 -551 9068
rect -516 9034 -482 9068
rect -447 9034 -413 9068
rect -378 9034 -344 9068
rect -309 9034 -275 9068
rect -240 9034 -206 9068
rect -171 9034 -137 9068
rect -102 9034 -68 9068
rect -932 8999 -898 9033
rect -864 8999 -830 9033
rect -796 8999 -762 9033
rect -723 8966 -689 9000
rect -654 8966 -620 9000
rect -585 8966 -551 9000
rect -516 8966 -482 9000
rect -447 8966 -413 9000
rect -378 8966 -344 9000
rect -309 8966 -275 9000
rect -240 8966 -206 9000
rect -171 8966 -137 9000
rect -102 8966 -68 9000
rect -33 8966 14893 9680
rect 14932 9613 14966 9647
rect 15000 9613 15034 9647
rect 15068 9613 15102 9647
rect 14932 9537 14966 9571
rect 15000 9537 15034 9571
rect 15068 9537 15102 9571
rect 14932 9461 14966 9495
rect 15000 9461 15034 9495
rect 15068 9461 15102 9495
rect 14932 9384 14966 9418
rect 15000 9384 15034 9418
rect 15068 9384 15102 9418
rect 14932 9307 14966 9341
rect 15000 9307 15034 9341
rect 15068 9307 15102 9341
rect 14932 9230 14966 9264
rect 15000 9230 15034 9264
rect 15068 9230 15102 9264
rect 14932 9153 14966 9187
rect 15000 9153 15034 9187
rect 15068 9153 15102 9187
rect 14932 9076 14966 9110
rect 15000 9076 15034 9110
rect 15068 9076 15102 9110
rect 14932 8999 14966 9033
rect 15000 8999 15034 9033
rect 15068 8999 15102 9033
rect 68 6809 102 6843
rect 137 6809 171 6843
rect 206 6809 240 6843
rect 275 6809 309 6843
rect 344 6809 378 6843
rect 413 6809 447 6843
rect 482 6809 516 6843
rect 551 6809 585 6843
rect 620 6809 654 6843
rect 689 6809 723 6843
rect 758 6809 792 6843
rect 827 6809 861 6843
rect 896 6809 930 6843
rect 965 6809 999 6843
rect 1034 6809 1068 6843
rect 1103 6809 1137 6843
rect 1172 6809 1206 6843
rect 1241 6809 1275 6843
rect 1310 6809 1344 6843
rect 1379 6809 1413 6843
rect 1448 6809 1482 6843
rect 1517 6809 1551 6843
rect 1586 6809 1620 6843
rect 1655 6809 1689 6843
rect 1724 6809 1758 6843
rect 1793 6809 1827 6843
rect 1862 6809 1896 6843
rect 1931 6809 1965 6843
rect 2000 6809 2034 6843
rect 2069 6809 2103 6843
rect 2138 6809 2172 6843
rect 2207 6809 2241 6843
rect 2276 6809 2310 6843
rect 2345 6809 2379 6843
rect 2414 6809 2448 6843
rect 2483 6809 2517 6843
rect 2552 6809 2586 6843
rect 2621 6809 2655 6843
rect 2690 6809 2724 6843
rect 2759 6809 2793 6843
rect 2828 6809 2862 6843
rect 2897 6809 2931 6843
rect 2966 6809 3000 6843
rect 3035 6809 3069 6843
rect 3104 6809 3138 6843
rect 3173 6809 3207 6843
rect 3242 6809 3276 6843
rect 3310 6809 3344 6843
rect 3378 6809 3412 6843
rect 3446 6809 3480 6843
rect 3514 6809 3548 6843
rect 3582 6809 3616 6843
rect 3650 6809 3684 6843
rect 3718 6809 3752 6843
rect 3786 6809 3820 6843
rect 3854 6809 3888 6843
rect 3922 6809 3956 6843
rect 3990 6809 4024 6843
rect 4058 6809 4092 6843
rect 4126 6809 4160 6843
rect 4194 6809 4228 6843
rect 4262 6809 4296 6843
rect 4330 6809 4364 6843
rect 4398 6809 4432 6843
rect 4466 6809 4500 6843
rect 4534 6809 4568 6843
rect 4602 6809 4636 6843
rect 4670 6809 4704 6843
rect 4738 6809 4772 6843
rect 4806 6809 4840 6843
rect 4874 6809 4908 6843
rect 4942 6809 4976 6843
rect 5010 6809 5044 6843
rect 5078 6809 5112 6843
rect 5146 6809 5180 6843
rect 5214 6809 5248 6843
rect 5282 6809 5316 6843
rect 5350 6809 5384 6843
rect 5418 6809 5452 6843
rect 5486 6809 5520 6843
rect 5554 6809 5588 6843
rect 5622 6809 5656 6843
rect 5690 6809 5724 6843
rect 5758 6809 5792 6843
rect 5826 6809 5860 6843
rect 5894 6809 5928 6843
rect 5962 6809 5996 6843
rect 6030 6809 6064 6843
rect 6098 6809 6132 6843
rect 6166 6809 6200 6843
rect 6234 6809 6268 6843
rect 6302 6809 6336 6843
rect 6370 6809 6404 6843
rect 6438 6809 6472 6843
rect 6506 6809 6540 6843
rect 6574 6809 6608 6843
rect 6642 6809 6676 6843
rect 6710 6809 6744 6843
rect 6778 6809 6812 6843
rect 6846 6809 6880 6843
rect 6914 6809 6948 6843
rect 6982 6809 7016 6843
rect 7050 6809 7084 6843
rect 68 6722 102 6756
rect 137 6722 171 6756
rect 206 6722 240 6756
rect 275 6722 309 6756
rect 344 6722 378 6756
rect 413 6722 447 6756
rect 482 6722 516 6756
rect 551 6722 585 6756
rect 620 6722 654 6756
rect 689 6722 723 6756
rect 758 6722 792 6756
rect 827 6722 861 6756
rect 896 6722 930 6756
rect 965 6722 999 6756
rect 1034 6722 1068 6756
rect 1103 6722 1137 6756
rect 1172 6722 1206 6756
rect 1241 6722 1275 6756
rect 1310 6722 1344 6756
rect 1379 6722 1413 6756
rect 1448 6722 1482 6756
rect 1517 6722 1551 6756
rect 1586 6722 1620 6756
rect 1655 6722 1689 6756
rect 1724 6722 1758 6756
rect 1793 6722 1827 6756
rect 1862 6722 1896 6756
rect 1931 6722 1965 6756
rect 2000 6722 2034 6756
rect 2069 6722 2103 6756
rect 2138 6722 2172 6756
rect 2207 6722 2241 6756
rect 2276 6722 2310 6756
rect 2345 6722 2379 6756
rect 2414 6722 2448 6756
rect 2483 6722 2517 6756
rect 2552 6722 2586 6756
rect 2621 6722 2655 6756
rect 2690 6722 2724 6756
rect 2759 6722 2793 6756
rect 2828 6722 2862 6756
rect 2897 6722 2931 6756
rect 2966 6722 3000 6756
rect 3035 6722 3069 6756
rect 3104 6722 3138 6756
rect 3173 6722 3207 6756
rect 3242 6722 3276 6756
rect 3310 6722 3344 6756
rect 3378 6722 3412 6756
rect 3446 6722 3480 6756
rect 3514 6722 3548 6756
rect 3582 6722 3616 6756
rect 3650 6722 3684 6756
rect 3718 6722 3752 6756
rect 3786 6722 3820 6756
rect 3854 6722 3888 6756
rect 3922 6722 3956 6756
rect 3990 6722 4024 6756
rect 4058 6722 4092 6756
rect 4126 6722 4160 6756
rect 4194 6722 4228 6756
rect 4262 6722 4296 6756
rect 4330 6722 4364 6756
rect 4398 6722 4432 6756
rect 4466 6722 4500 6756
rect 4534 6722 4568 6756
rect 4602 6722 4636 6756
rect 4670 6722 4704 6756
rect 4738 6722 4772 6756
rect 4806 6722 4840 6756
rect 4874 6722 4908 6756
rect 4942 6722 4976 6756
rect 5010 6722 5044 6756
rect 5078 6722 5112 6756
rect 5146 6722 5180 6756
rect 5214 6722 5248 6756
rect 5282 6722 5316 6756
rect 5350 6722 5384 6756
rect 5418 6722 5452 6756
rect 5486 6722 5520 6756
rect 5554 6722 5588 6756
rect 5622 6722 5656 6756
rect 5690 6722 5724 6756
rect 5758 6722 5792 6756
rect 5826 6722 5860 6756
rect 5894 6722 5928 6756
rect 5962 6722 5996 6756
rect 6030 6722 6064 6756
rect 6098 6722 6132 6756
rect 6166 6722 6200 6756
rect 6234 6722 6268 6756
rect 6302 6722 6336 6756
rect 6370 6722 6404 6756
rect 6438 6722 6472 6756
rect 6506 6722 6540 6756
rect 6574 6722 6608 6756
rect 6642 6722 6676 6756
rect 6710 6722 6744 6756
rect 6778 6722 6812 6756
rect 6846 6722 6880 6756
rect 6914 6722 6948 6756
rect 6982 6722 7016 6756
rect 7050 6722 7084 6756
rect 68 6635 102 6669
rect 137 6635 171 6669
rect 206 6635 240 6669
rect 275 6635 309 6669
rect 344 6635 378 6669
rect 413 6635 447 6669
rect 482 6635 516 6669
rect 551 6635 585 6669
rect 620 6635 654 6669
rect 689 6635 723 6669
rect 758 6635 792 6669
rect 827 6635 861 6669
rect 896 6635 930 6669
rect 965 6635 999 6669
rect 1034 6635 1068 6669
rect 1103 6635 1137 6669
rect 1172 6635 1206 6669
rect 1241 6635 1275 6669
rect 1310 6635 1344 6669
rect 1379 6635 1413 6669
rect 1448 6635 1482 6669
rect 1517 6635 1551 6669
rect 1586 6635 1620 6669
rect 1655 6635 1689 6669
rect 1724 6635 1758 6669
rect 1793 6635 1827 6669
rect 1862 6635 1896 6669
rect 1931 6635 1965 6669
rect 2000 6635 2034 6669
rect 2069 6635 2103 6669
rect 2138 6635 2172 6669
rect 2207 6635 2241 6669
rect 2276 6635 2310 6669
rect 2345 6635 2379 6669
rect 2414 6635 2448 6669
rect 2483 6635 2517 6669
rect 2552 6635 2586 6669
rect 2621 6635 2655 6669
rect 2690 6635 2724 6669
rect 2759 6635 2793 6669
rect 2828 6635 2862 6669
rect 2897 6635 2931 6669
rect 2966 6635 3000 6669
rect 3035 6635 3069 6669
rect 3104 6635 3138 6669
rect 3173 6635 3207 6669
rect 3242 6635 3276 6669
rect 3310 6635 3344 6669
rect 3378 6635 3412 6669
rect 3446 6635 3480 6669
rect 3514 6635 3548 6669
rect 3582 6635 3616 6669
rect 3650 6635 3684 6669
rect 3718 6635 3752 6669
rect 3786 6635 3820 6669
rect 3854 6635 3888 6669
rect 3922 6635 3956 6669
rect 3990 6635 4024 6669
rect 4058 6635 4092 6669
rect 4126 6635 4160 6669
rect 4194 6635 4228 6669
rect 4262 6635 4296 6669
rect 4330 6635 4364 6669
rect 4398 6635 4432 6669
rect 4466 6635 4500 6669
rect 4534 6635 4568 6669
rect 4602 6635 4636 6669
rect 4670 6635 4704 6669
rect 4738 6635 4772 6669
rect 4806 6635 4840 6669
rect 4874 6635 4908 6669
rect 4942 6635 4976 6669
rect 5010 6635 5044 6669
rect 5078 6635 5112 6669
rect 5146 6635 5180 6669
rect 5214 6635 5248 6669
rect 5282 6635 5316 6669
rect 5350 6635 5384 6669
rect 5418 6635 5452 6669
rect 5486 6635 5520 6669
rect 5554 6635 5588 6669
rect 5622 6635 5656 6669
rect 5690 6635 5724 6669
rect 5758 6635 5792 6669
rect 5826 6635 5860 6669
rect 5894 6635 5928 6669
rect 5962 6635 5996 6669
rect 6030 6635 6064 6669
rect 6098 6635 6132 6669
rect 6166 6635 6200 6669
rect 6234 6635 6268 6669
rect 6302 6635 6336 6669
rect 6370 6635 6404 6669
rect 6438 6635 6472 6669
rect 6506 6635 6540 6669
rect 6574 6635 6608 6669
rect 6642 6635 6676 6669
rect 6710 6635 6744 6669
rect 6778 6635 6812 6669
rect 6846 6635 6880 6669
rect 6914 6635 6948 6669
rect 6982 6635 7016 6669
rect 7050 6635 7084 6669
rect 12517 6809 12551 6843
rect 12586 6809 12620 6843
rect 12655 6809 12689 6843
rect 12724 6809 12758 6843
rect 12793 6809 12827 6843
rect 12862 6809 12896 6843
rect 12931 6809 12965 6843
rect 13000 6809 13034 6843
rect 13069 6809 13103 6843
rect 13138 6809 13172 6843
rect 13207 6809 13241 6843
rect 13276 6809 13310 6843
rect 13345 6809 13379 6843
rect 13414 6809 13448 6843
rect 13483 6809 13517 6843
rect 13552 6809 13586 6843
rect 13621 6809 13655 6843
rect 13690 6809 13724 6843
rect 13759 6809 13793 6843
rect 13828 6809 13862 6843
rect 13897 6809 13931 6843
rect 13966 6809 14000 6843
rect 14035 6809 14069 6843
rect 14104 6809 14138 6843
rect 14173 6809 14207 6843
rect 14242 6809 14276 6843
rect 14311 6809 14345 6843
rect 14380 6809 14414 6843
rect 14449 6809 14483 6843
rect 14518 6809 14552 6843
rect 14587 6809 14621 6843
rect 14655 6809 14689 6843
rect 14723 6809 14757 6843
rect 14791 6809 14825 6843
rect 14859 6809 14893 6843
rect 14932 6771 14966 6805
rect 15000 6771 15034 6805
rect 15068 6771 15102 6805
rect 12517 6722 12551 6756
rect 12586 6722 12620 6756
rect 12655 6722 12689 6756
rect 12724 6722 12758 6756
rect 12793 6722 12827 6756
rect 12862 6722 12896 6756
rect 12931 6722 12965 6756
rect 13000 6722 13034 6756
rect 13069 6722 13103 6756
rect 13138 6722 13172 6756
rect 13207 6722 13241 6756
rect 13276 6722 13310 6756
rect 13345 6722 13379 6756
rect 13414 6722 13448 6756
rect 13483 6722 13517 6756
rect 13552 6722 13586 6756
rect 13621 6722 13655 6756
rect 13690 6722 13724 6756
rect 13759 6722 13793 6756
rect 13828 6722 13862 6756
rect 13897 6722 13931 6756
rect 13966 6722 14000 6756
rect 14035 6722 14069 6756
rect 14104 6722 14138 6756
rect 14173 6722 14207 6756
rect 14242 6722 14276 6756
rect 14311 6722 14345 6756
rect 14380 6722 14414 6756
rect 14449 6722 14483 6756
rect 14518 6722 14552 6756
rect 14587 6722 14621 6756
rect 14655 6722 14689 6756
rect 14723 6722 14757 6756
rect 14791 6722 14825 6756
rect 14859 6722 14893 6756
rect 14932 6697 14966 6731
rect 15000 6697 15034 6731
rect 15068 6697 15102 6731
rect 12517 6635 12551 6669
rect 12586 6635 12620 6669
rect 12655 6635 12689 6669
rect 12724 6635 12758 6669
rect 12793 6635 12827 6669
rect 12862 6635 12896 6669
rect 12931 6635 12965 6669
rect 13000 6635 13034 6669
rect 13069 6635 13103 6669
rect 13138 6635 13172 6669
rect 13207 6635 13241 6669
rect 13276 6635 13310 6669
rect 13345 6635 13379 6669
rect 13414 6635 13448 6669
rect 13483 6635 13517 6669
rect 13552 6635 13586 6669
rect 13621 6635 13655 6669
rect 13690 6635 13724 6669
rect 13759 6635 13793 6669
rect 13828 6635 13862 6669
rect 13897 6635 13931 6669
rect 13966 6635 14000 6669
rect 14035 6635 14069 6669
rect 14104 6635 14138 6669
rect 14173 6635 14207 6669
rect 14242 6635 14276 6669
rect 14311 6635 14345 6669
rect 14380 6635 14414 6669
rect 14449 6635 14483 6669
rect 14518 6635 14552 6669
rect 14587 6635 14621 6669
rect 14655 6635 14689 6669
rect 14723 6635 14757 6669
rect 14791 6635 14825 6669
rect 14859 6635 14893 6669
rect 14932 6623 14966 6657
rect 15000 6623 15034 6657
rect 15068 6623 15102 6657
rect 68 6548 102 6582
rect 137 6548 171 6582
rect 206 6548 240 6582
rect 275 6548 309 6582
rect 344 6548 378 6582
rect 413 6548 447 6582
rect 482 6548 516 6582
rect 551 6548 585 6582
rect 620 6548 654 6582
rect 689 6548 723 6582
rect 758 6548 792 6582
rect 827 6548 861 6582
rect 896 6548 930 6582
rect 965 6548 999 6582
rect 1034 6548 1068 6582
rect 1103 6548 1137 6582
rect 1172 6548 1206 6582
rect 1241 6548 1275 6582
rect 1310 6548 1344 6582
rect 1379 6548 1413 6582
rect 1448 6548 1482 6582
rect 1517 6548 1551 6582
rect 1586 6548 1620 6582
rect 1655 6548 1689 6582
rect 1724 6548 1758 6582
rect 1793 6548 1827 6582
rect 1862 6548 1896 6582
rect 1931 6548 1965 6582
rect 2000 6548 2034 6582
rect 2069 6548 2103 6582
rect 2138 6548 2172 6582
rect 2207 6548 2241 6582
rect 2276 6548 2310 6582
rect 2345 6548 2379 6582
rect 2414 6548 2448 6582
rect 2483 6548 2517 6582
rect 2551 6548 2585 6582
rect 2619 6548 2653 6582
rect 2687 6548 2721 6582
rect 2755 6548 2789 6582
rect 2823 6548 2857 6582
rect 2891 6548 2925 6582
rect 2959 6548 2993 6582
rect 3027 6548 3061 6582
rect 3095 6548 3129 6582
rect 3163 6548 3197 6582
rect 3231 6548 3265 6582
rect 3299 6548 3333 6582
rect 3367 6548 3401 6582
rect 3435 6548 3469 6582
rect 3503 6548 3537 6582
rect 3571 6548 3605 6582
rect 3639 6548 3673 6582
rect 3707 6548 3741 6582
rect 3775 6548 3809 6582
rect 3843 6548 3877 6582
rect 3911 6548 3945 6582
rect 3979 6548 4013 6582
rect 4047 6548 4081 6582
rect 4115 6548 4149 6582
rect 4183 6548 4217 6582
rect 4251 6548 4285 6582
rect 4319 6548 4353 6582
rect 4387 6548 4421 6582
rect 4455 6548 4489 6582
rect 4523 6548 4557 6582
rect 4591 6548 4625 6582
rect 4659 6548 4693 6582
rect 4727 6548 4761 6582
rect 4795 6548 4829 6582
rect 4863 6548 4897 6582
rect 4931 6548 4965 6582
rect 4999 6548 5033 6582
rect 5067 6548 5101 6582
rect 5135 6548 5169 6582
rect 5203 6548 5237 6582
rect 5271 6548 5305 6582
rect 5339 6548 5373 6582
rect 5407 6548 5441 6582
rect 5475 6548 5509 6582
rect 5543 6548 5577 6582
rect 5611 6548 5645 6582
rect 5679 6548 5713 6582
rect 5747 6548 5781 6582
rect 5815 6548 5849 6582
rect 5883 6548 5917 6582
rect 5951 6548 5985 6582
rect 6019 6548 6053 6582
rect 6087 6548 6121 6582
rect 6155 6548 6189 6582
rect 6223 6548 6257 6582
rect 6291 6548 6325 6582
rect 6359 6548 6393 6582
rect 6427 6548 6461 6582
rect 6495 6548 6529 6582
rect 6563 6548 6597 6582
rect 6631 6548 6665 6582
rect 6699 6548 6733 6582
rect 6767 6548 6801 6582
rect 6835 6548 6869 6582
rect 6903 6548 6937 6582
rect 6971 6548 7005 6582
rect 7039 6548 7073 6582
rect 7107 6548 7141 6582
rect 7175 6548 7209 6582
rect 7243 6548 7277 6582
rect 7311 6548 7345 6582
rect 7379 6548 7413 6582
rect 7447 6548 7481 6582
rect 7515 6548 7549 6582
rect 7583 6548 7617 6582
rect 7651 6548 7685 6582
rect 7719 6548 7753 6582
rect 7787 6548 7821 6582
rect 7855 6548 7889 6582
rect 7923 6548 7957 6582
rect 7991 6548 8025 6582
rect 8059 6548 8093 6582
rect 8127 6548 8161 6582
rect 8195 6548 8229 6582
rect 8263 6548 8297 6582
rect 8331 6548 8365 6582
rect 8399 6548 8433 6582
rect 8467 6548 8501 6582
rect 8535 6548 8569 6582
rect 8603 6548 8637 6582
rect 8671 6548 8705 6582
rect 8739 6548 8773 6582
rect 8807 6548 8841 6582
rect 8875 6548 8909 6582
rect 8943 6548 8977 6582
rect 9011 6548 9045 6582
rect 9079 6548 9113 6582
rect 9147 6548 9181 6582
rect 9215 6548 9249 6582
rect 9283 6548 9317 6582
rect 9351 6548 9385 6582
rect 9419 6548 9453 6582
rect 9487 6548 9521 6582
rect 9555 6548 9589 6582
rect 9623 6548 9657 6582
rect 9691 6548 9725 6582
rect 9759 6548 9793 6582
rect 9827 6548 9861 6582
rect 9895 6548 9929 6582
rect 9963 6548 9997 6582
rect 10031 6548 10065 6582
rect 10099 6548 10133 6582
rect 10167 6548 10201 6582
rect 10235 6548 10269 6582
rect 10303 6548 10337 6582
rect 10371 6548 10405 6582
rect 10439 6548 10473 6582
rect 10507 6548 10541 6582
rect 10575 6548 10609 6582
rect 10643 6548 10677 6582
rect 10711 6548 10745 6582
rect 10779 6548 10813 6582
rect 10847 6548 10881 6582
rect 10915 6548 10949 6582
rect 10983 6548 11017 6582
rect 11051 6548 11085 6582
rect 11119 6548 11153 6582
rect 11187 6548 11221 6582
rect 11255 6548 11289 6582
rect 11323 6548 11357 6582
rect 11391 6548 11425 6582
rect 11459 6548 11493 6582
rect 11527 6548 11561 6582
rect 11595 6548 11629 6582
rect 11663 6548 11697 6582
rect 11731 6548 11765 6582
rect 11799 6548 11833 6582
rect 11867 6548 11901 6582
rect 11935 6548 11969 6582
rect 12003 6548 12037 6582
rect 12071 6548 12105 6582
rect 12139 6548 12173 6582
rect 12207 6548 12241 6582
rect 12275 6548 12309 6582
rect 12343 6548 12377 6582
rect 12411 6548 12445 6582
rect 12479 6548 12513 6582
rect 12547 6548 12581 6582
rect 12615 6548 12649 6582
rect 12683 6548 12717 6582
rect 12751 6548 12785 6582
rect 12819 6548 12853 6582
rect 12887 6548 12921 6582
rect 12955 6548 12989 6582
rect 13023 6548 13057 6582
rect 13091 6548 13125 6582
rect 13159 6548 13193 6582
rect 13227 6548 13261 6582
rect 13295 6548 13329 6582
rect 13363 6548 13397 6582
rect 13431 6548 13465 6582
rect 13499 6548 13533 6582
rect 13567 6548 13601 6582
rect 13635 6548 13669 6582
rect 13703 6548 13737 6582
rect 13771 6548 13805 6582
rect 13839 6548 13873 6582
rect 13907 6548 13941 6582
rect 13975 6548 14009 6582
rect 14043 6548 14077 6582
rect 14111 6548 14145 6582
rect 14179 6548 14213 6582
rect 14247 6548 14281 6582
rect 14315 6548 14349 6582
rect 14383 6548 14417 6582
rect 14451 6548 14485 6582
rect 14519 6548 14553 6582
rect 14587 6548 14621 6582
rect 14655 6548 14689 6582
rect 14723 6548 14757 6582
rect 14791 6548 14825 6582
rect 14859 6548 14893 6582
rect 14932 6549 14966 6583
rect 15000 6549 15034 6583
rect 15068 6549 15102 6583
rect 68 6474 102 6508
rect 137 6474 171 6508
rect 206 6474 240 6508
rect 275 6474 309 6508
rect 344 6474 378 6508
rect 413 6474 447 6508
rect 482 6474 516 6508
rect 551 6474 585 6508
rect 620 6474 654 6508
rect 689 6474 723 6508
rect 758 6474 792 6508
rect 827 6474 861 6508
rect 896 6474 930 6508
rect 965 6474 999 6508
rect 1034 6474 1068 6508
rect 1103 6474 1137 6508
rect 1172 6474 1206 6508
rect 1241 6474 1275 6508
rect 1310 6474 1344 6508
rect 1379 6474 1413 6508
rect 1448 6474 1482 6508
rect 1517 6474 1551 6508
rect 1586 6474 1620 6508
rect 1655 6474 1689 6508
rect 1724 6474 1758 6508
rect 1793 6474 1827 6508
rect 1862 6474 1896 6508
rect 1931 6474 1965 6508
rect 2000 6474 2034 6508
rect 2069 6474 2103 6508
rect 2138 6474 2172 6508
rect 2207 6474 2241 6508
rect 2276 6474 2310 6508
rect 2345 6474 2379 6508
rect 2414 6474 2448 6508
rect 2483 6474 2517 6508
rect 2551 6474 2585 6508
rect 2619 6474 2653 6508
rect 2687 6474 2721 6508
rect 2755 6474 2789 6508
rect 2823 6474 2857 6508
rect 2891 6474 2925 6508
rect 2959 6474 2993 6508
rect 3027 6474 3061 6508
rect 3095 6474 3129 6508
rect 3163 6474 3197 6508
rect 3231 6474 3265 6508
rect 3299 6474 3333 6508
rect 3367 6474 3401 6508
rect 3435 6474 3469 6508
rect 3503 6474 3537 6508
rect 3571 6474 3605 6508
rect 3639 6474 3673 6508
rect 3707 6474 3741 6508
rect 3775 6474 3809 6508
rect 3843 6474 3877 6508
rect 3911 6474 3945 6508
rect 3979 6474 4013 6508
rect 4047 6474 4081 6508
rect 4115 6474 4149 6508
rect 4183 6474 4217 6508
rect 4251 6474 4285 6508
rect 4319 6474 4353 6508
rect 4387 6474 4421 6508
rect 4455 6474 4489 6508
rect 4523 6474 4557 6508
rect 4591 6474 4625 6508
rect 4659 6474 4693 6508
rect 4727 6474 4761 6508
rect 4795 6474 4829 6508
rect 4863 6474 4897 6508
rect 4931 6474 4965 6508
rect 4999 6474 5033 6508
rect 5067 6474 5101 6508
rect 5135 6474 5169 6508
rect 5203 6474 5237 6508
rect 5271 6474 5305 6508
rect 5339 6474 5373 6508
rect 5407 6474 5441 6508
rect 5475 6474 5509 6508
rect 5543 6474 5577 6508
rect 5611 6474 5645 6508
rect 5679 6474 5713 6508
rect 5747 6474 5781 6508
rect 5815 6474 5849 6508
rect 5883 6474 5917 6508
rect 5951 6474 5985 6508
rect 6019 6474 6053 6508
rect 6087 6474 6121 6508
rect 6155 6474 6189 6508
rect 6223 6474 6257 6508
rect 6291 6474 6325 6508
rect 6359 6474 6393 6508
rect 6427 6474 6461 6508
rect 6495 6474 6529 6508
rect 6563 6474 6597 6508
rect 6631 6474 6665 6508
rect 6699 6474 6733 6508
rect 6767 6474 6801 6508
rect 6835 6474 6869 6508
rect 6903 6474 6937 6508
rect 6971 6474 7005 6508
rect 7039 6474 7073 6508
rect 7107 6474 7141 6508
rect 7175 6474 7209 6508
rect 7243 6474 7277 6508
rect 7311 6474 7345 6508
rect 7379 6474 7413 6508
rect 7447 6474 7481 6508
rect 7515 6474 7549 6508
rect 7583 6474 7617 6508
rect 7651 6474 7685 6508
rect 7719 6474 7753 6508
rect 7787 6474 7821 6508
rect 7855 6474 7889 6508
rect 7923 6474 7957 6508
rect 7991 6474 8025 6508
rect 8059 6474 8093 6508
rect 8127 6474 8161 6508
rect 8195 6474 8229 6508
rect 8263 6474 8297 6508
rect 8331 6474 8365 6508
rect 8399 6474 8433 6508
rect 8467 6474 8501 6508
rect 8535 6474 8569 6508
rect 8603 6474 8637 6508
rect 8671 6474 8705 6508
rect 8739 6474 8773 6508
rect 8807 6474 8841 6508
rect 8875 6474 8909 6508
rect 8943 6474 8977 6508
rect 9011 6474 9045 6508
rect 9079 6474 9113 6508
rect 9147 6474 9181 6508
rect 9215 6474 9249 6508
rect 9283 6474 9317 6508
rect 9351 6474 9385 6508
rect 9419 6474 9453 6508
rect 9487 6474 9521 6508
rect 9555 6474 9589 6508
rect 9623 6474 9657 6508
rect 9691 6474 9725 6508
rect 9759 6474 9793 6508
rect 9827 6474 9861 6508
rect 9895 6474 9929 6508
rect 9963 6474 9997 6508
rect 10031 6474 10065 6508
rect 10099 6474 10133 6508
rect 10167 6474 10201 6508
rect 10235 6474 10269 6508
rect 10303 6474 10337 6508
rect 10371 6474 10405 6508
rect 10439 6474 10473 6508
rect 10507 6474 10541 6508
rect 10575 6474 10609 6508
rect 10643 6474 10677 6508
rect 10711 6474 10745 6508
rect 10779 6474 10813 6508
rect 10847 6474 10881 6508
rect 10915 6474 10949 6508
rect 10983 6474 11017 6508
rect 11051 6474 11085 6508
rect 11119 6474 11153 6508
rect 11187 6474 11221 6508
rect 11255 6474 11289 6508
rect 11323 6474 11357 6508
rect 11391 6474 11425 6508
rect 11459 6474 11493 6508
rect 11527 6474 11561 6508
rect 11595 6474 11629 6508
rect 11663 6474 11697 6508
rect 11731 6474 11765 6508
rect 11799 6474 11833 6508
rect 11867 6474 11901 6508
rect 11935 6474 11969 6508
rect 12003 6474 12037 6508
rect 12071 6474 12105 6508
rect 12139 6474 12173 6508
rect 12207 6474 12241 6508
rect 12275 6474 12309 6508
rect 12343 6474 12377 6508
rect 12411 6474 12445 6508
rect 12479 6474 12513 6508
rect 12547 6474 12581 6508
rect 12615 6474 12649 6508
rect 12683 6474 12717 6508
rect 12751 6474 12785 6508
rect 12819 6474 12853 6508
rect 12887 6474 12921 6508
rect 12955 6474 12989 6508
rect 13023 6474 13057 6508
rect 13091 6474 13125 6508
rect 13159 6474 13193 6508
rect 13227 6474 13261 6508
rect 13295 6474 13329 6508
rect 13363 6474 13397 6508
rect 13431 6474 13465 6508
rect 13499 6474 13533 6508
rect 13567 6474 13601 6508
rect 13635 6474 13669 6508
rect 13703 6474 13737 6508
rect 13771 6474 13805 6508
rect 13839 6474 13873 6508
rect 13907 6474 13941 6508
rect 13975 6474 14009 6508
rect 14043 6474 14077 6508
rect 14111 6474 14145 6508
rect 14179 6474 14213 6508
rect 14247 6474 14281 6508
rect 14315 6474 14349 6508
rect 14383 6474 14417 6508
rect 14451 6474 14485 6508
rect 14519 6474 14553 6508
rect 14587 6474 14621 6508
rect 14655 6474 14689 6508
rect 14723 6474 14757 6508
rect 14791 6474 14825 6508
rect 14859 6474 14893 6508
rect 14932 6475 14966 6509
rect 15000 6475 15034 6509
rect 15068 6475 15102 6509
rect 68 6400 102 6434
rect 137 6400 171 6434
rect 206 6400 240 6434
rect 275 6400 309 6434
rect 344 6400 378 6434
rect 413 6400 447 6434
rect 482 6400 516 6434
rect 551 6400 585 6434
rect 620 6400 654 6434
rect 689 6400 723 6434
rect 758 6400 792 6434
rect 827 6400 861 6434
rect 896 6400 930 6434
rect 965 6400 999 6434
rect 1034 6400 1068 6434
rect 1103 6400 1137 6434
rect 1172 6400 1206 6434
rect 1241 6400 1275 6434
rect 1310 6400 1344 6434
rect 1379 6400 1413 6434
rect 1448 6400 1482 6434
rect 1517 6400 1551 6434
rect 1586 6400 1620 6434
rect 1655 6400 1689 6434
rect 1724 6400 1758 6434
rect 1793 6400 1827 6434
rect 1862 6400 1896 6434
rect 1931 6400 1965 6434
rect 2000 6400 2034 6434
rect 2069 6400 2103 6434
rect 2138 6400 2172 6434
rect 2207 6400 2241 6434
rect 2276 6400 2310 6434
rect 2345 6400 2379 6434
rect 2414 6400 2448 6434
rect 2483 6400 2517 6434
rect 2551 6400 2585 6434
rect 2619 6400 2653 6434
rect 2687 6400 2721 6434
rect 2755 6400 2789 6434
rect 2823 6400 2857 6434
rect 2891 6400 2925 6434
rect 2959 6400 2993 6434
rect 3027 6400 3061 6434
rect 3095 6400 3129 6434
rect 3163 6400 3197 6434
rect 3231 6400 3265 6434
rect 3299 6400 3333 6434
rect 3367 6400 3401 6434
rect 3435 6400 3469 6434
rect 3503 6400 3537 6434
rect 3571 6400 3605 6434
rect 3639 6400 3673 6434
rect 3707 6400 3741 6434
rect 3775 6400 3809 6434
rect 3843 6400 3877 6434
rect 3911 6400 3945 6434
rect 3979 6400 4013 6434
rect 4047 6400 4081 6434
rect 4115 6400 4149 6434
rect 4183 6400 4217 6434
rect 4251 6400 4285 6434
rect 4319 6400 4353 6434
rect 4387 6400 4421 6434
rect 4455 6400 4489 6434
rect 4523 6400 4557 6434
rect 4591 6400 4625 6434
rect 4659 6400 4693 6434
rect 4727 6400 4761 6434
rect 4795 6400 4829 6434
rect 4863 6400 4897 6434
rect 4931 6400 4965 6434
rect 4999 6400 5033 6434
rect 5067 6400 5101 6434
rect 5135 6400 5169 6434
rect 5203 6400 5237 6434
rect 5271 6400 5305 6434
rect 5339 6400 5373 6434
rect 5407 6400 5441 6434
rect 5475 6400 5509 6434
rect 5543 6400 5577 6434
rect 5611 6400 5645 6434
rect 5679 6400 5713 6434
rect 5747 6400 5781 6434
rect 5815 6400 5849 6434
rect 5883 6400 5917 6434
rect 5951 6400 5985 6434
rect 6019 6400 6053 6434
rect 6087 6400 6121 6434
rect 6155 6400 6189 6434
rect 6223 6400 6257 6434
rect 6291 6400 6325 6434
rect 6359 6400 6393 6434
rect 6427 6400 6461 6434
rect 6495 6400 6529 6434
rect 6563 6400 6597 6434
rect 6631 6400 6665 6434
rect 6699 6400 6733 6434
rect 6767 6400 6801 6434
rect 6835 6400 6869 6434
rect 6903 6400 6937 6434
rect 6971 6400 7005 6434
rect 7039 6400 7073 6434
rect 7107 6400 7141 6434
rect 7175 6400 7209 6434
rect 7243 6400 7277 6434
rect 7311 6400 7345 6434
rect 7379 6400 7413 6434
rect 7447 6400 7481 6434
rect 7515 6400 7549 6434
rect 7583 6400 7617 6434
rect 7651 6400 7685 6434
rect 7719 6400 7753 6434
rect 7787 6400 7821 6434
rect 7855 6400 7889 6434
rect 7923 6400 7957 6434
rect 7991 6400 8025 6434
rect 8059 6400 8093 6434
rect 8127 6400 8161 6434
rect 8195 6400 8229 6434
rect 8263 6400 8297 6434
rect 8331 6400 8365 6434
rect 8399 6400 8433 6434
rect 8467 6400 8501 6434
rect 8535 6400 8569 6434
rect 8603 6400 8637 6434
rect 8671 6400 8705 6434
rect 8739 6400 8773 6434
rect 8807 6400 8841 6434
rect 8875 6400 8909 6434
rect 8943 6400 8977 6434
rect 9011 6400 9045 6434
rect 9079 6400 9113 6434
rect 9147 6400 9181 6434
rect 9215 6400 9249 6434
rect 9283 6400 9317 6434
rect 9351 6400 9385 6434
rect 9419 6400 9453 6434
rect 9487 6400 9521 6434
rect 9555 6400 9589 6434
rect 9623 6400 9657 6434
rect 9691 6400 9725 6434
rect 9759 6400 9793 6434
rect 9827 6400 9861 6434
rect 9895 6400 9929 6434
rect 9963 6400 9997 6434
rect 10031 6400 10065 6434
rect 10099 6400 10133 6434
rect 10167 6400 10201 6434
rect 10235 6400 10269 6434
rect 10303 6400 10337 6434
rect 10371 6400 10405 6434
rect 10439 6400 10473 6434
rect 10507 6400 10541 6434
rect 10575 6400 10609 6434
rect 10643 6400 10677 6434
rect 10711 6400 10745 6434
rect 10779 6400 10813 6434
rect 10847 6400 10881 6434
rect 10915 6400 10949 6434
rect 10983 6400 11017 6434
rect 11051 6400 11085 6434
rect 11119 6400 11153 6434
rect 11187 6400 11221 6434
rect 11255 6400 11289 6434
rect 11323 6400 11357 6434
rect 11391 6400 11425 6434
rect 11459 6400 11493 6434
rect 11527 6400 11561 6434
rect 11595 6400 11629 6434
rect 11663 6400 11697 6434
rect 11731 6400 11765 6434
rect 11799 6400 11833 6434
rect 11867 6400 11901 6434
rect 11935 6400 11969 6434
rect 12003 6400 12037 6434
rect 12071 6400 12105 6434
rect 12139 6400 12173 6434
rect 12207 6400 12241 6434
rect 12275 6400 12309 6434
rect 12343 6400 12377 6434
rect 12411 6400 12445 6434
rect 12479 6400 12513 6434
rect 12547 6400 12581 6434
rect 12615 6400 12649 6434
rect 12683 6400 12717 6434
rect 12751 6400 12785 6434
rect 12819 6400 12853 6434
rect 12887 6400 12921 6434
rect 12955 6400 12989 6434
rect 13023 6400 13057 6434
rect 13091 6400 13125 6434
rect 13159 6400 13193 6434
rect 13227 6400 13261 6434
rect 13295 6400 13329 6434
rect 13363 6400 13397 6434
rect 13431 6400 13465 6434
rect 13499 6400 13533 6434
rect 13567 6400 13601 6434
rect 13635 6400 13669 6434
rect 13703 6400 13737 6434
rect 13771 6400 13805 6434
rect 13839 6400 13873 6434
rect 13907 6400 13941 6434
rect 13975 6400 14009 6434
rect 14043 6400 14077 6434
rect 14111 6400 14145 6434
rect 14179 6400 14213 6434
rect 14247 6400 14281 6434
rect 14315 6400 14349 6434
rect 14383 6400 14417 6434
rect 14451 6400 14485 6434
rect 14519 6400 14553 6434
rect 14587 6400 14621 6434
rect 14655 6400 14689 6434
rect 14723 6400 14757 6434
rect 14791 6400 14825 6434
rect 14859 6400 14893 6434
rect 14932 6401 14966 6435
rect 15000 6401 15034 6435
rect 15068 6401 15102 6435
rect 68 6326 102 6360
rect 137 6326 171 6360
rect 206 6326 240 6360
rect 275 6326 309 6360
rect 344 6326 378 6360
rect 413 6326 447 6360
rect 482 6326 516 6360
rect 551 6326 585 6360
rect 620 6326 654 6360
rect 689 6326 723 6360
rect 758 6326 792 6360
rect 827 6326 861 6360
rect 896 6326 930 6360
rect 965 6326 999 6360
rect 1034 6326 1068 6360
rect 1103 6326 1137 6360
rect 1172 6326 1206 6360
rect 1241 6326 1275 6360
rect 1310 6326 1344 6360
rect 1379 6326 1413 6360
rect 1448 6326 1482 6360
rect 1517 6326 1551 6360
rect 1586 6326 1620 6360
rect 1655 6326 1689 6360
rect 1724 6326 1758 6360
rect 1793 6326 1827 6360
rect 1862 6326 1896 6360
rect 1931 6326 1965 6360
rect 2000 6326 2034 6360
rect 2069 6326 2103 6360
rect 2138 6326 2172 6360
rect 2207 6326 2241 6360
rect 2276 6326 2310 6360
rect 2345 6326 2379 6360
rect 2414 6326 2448 6360
rect 2483 6326 2517 6360
rect 2551 6326 2585 6360
rect 2619 6326 2653 6360
rect 2687 6326 2721 6360
rect 2755 6326 2789 6360
rect 2823 6326 2857 6360
rect 2891 6326 2925 6360
rect 2959 6326 2993 6360
rect 3027 6326 3061 6360
rect 3095 6326 3129 6360
rect 3163 6326 3197 6360
rect 3231 6326 3265 6360
rect 3299 6326 3333 6360
rect 3367 6326 3401 6360
rect 3435 6326 3469 6360
rect 3503 6326 3537 6360
rect 3571 6326 3605 6360
rect 3639 6326 3673 6360
rect 3707 6326 3741 6360
rect 3775 6326 3809 6360
rect 3843 6326 3877 6360
rect 3911 6326 3945 6360
rect 3979 6326 4013 6360
rect 4047 6326 4081 6360
rect 4115 6326 4149 6360
rect 4183 6326 4217 6360
rect 4251 6326 4285 6360
rect 4319 6326 4353 6360
rect 4387 6326 4421 6360
rect 4455 6326 4489 6360
rect 4523 6326 4557 6360
rect 4591 6326 4625 6360
rect 4659 6326 4693 6360
rect 4727 6326 4761 6360
rect 4795 6326 4829 6360
rect 4863 6326 4897 6360
rect 4931 6326 4965 6360
rect 4999 6326 5033 6360
rect 5067 6326 5101 6360
rect 5135 6326 5169 6360
rect 5203 6326 5237 6360
rect 5271 6326 5305 6360
rect 5339 6326 5373 6360
rect 5407 6326 5441 6360
rect 5475 6326 5509 6360
rect 5543 6326 5577 6360
rect 5611 6326 5645 6360
rect 5679 6326 5713 6360
rect 5747 6326 5781 6360
rect 5815 6326 5849 6360
rect 5883 6326 5917 6360
rect 5951 6326 5985 6360
rect 6019 6326 6053 6360
rect 6087 6326 6121 6360
rect 6155 6326 6189 6360
rect 6223 6326 6257 6360
rect 6291 6326 6325 6360
rect 6359 6326 6393 6360
rect 6427 6326 6461 6360
rect 6495 6326 6529 6360
rect 6563 6326 6597 6360
rect 6631 6326 6665 6360
rect 6699 6326 6733 6360
rect 6767 6326 6801 6360
rect 6835 6326 6869 6360
rect 6903 6326 6937 6360
rect 6971 6326 7005 6360
rect 7039 6326 7073 6360
rect 7107 6326 7141 6360
rect 7175 6326 7209 6360
rect 7243 6326 7277 6360
rect 7311 6326 7345 6360
rect 7379 6326 7413 6360
rect 7447 6326 7481 6360
rect 7515 6326 7549 6360
rect 7583 6326 7617 6360
rect 7651 6326 7685 6360
rect 7719 6326 7753 6360
rect 7787 6326 7821 6360
rect 7855 6326 7889 6360
rect 7923 6326 7957 6360
rect 7991 6326 8025 6360
rect 8059 6326 8093 6360
rect 8127 6326 8161 6360
rect 8195 6326 8229 6360
rect 8263 6326 8297 6360
rect 8331 6326 8365 6360
rect 8399 6326 8433 6360
rect 8467 6326 8501 6360
rect 8535 6326 8569 6360
rect 8603 6326 8637 6360
rect 8671 6326 8705 6360
rect 8739 6326 8773 6360
rect 8807 6326 8841 6360
rect 8875 6326 8909 6360
rect 8943 6326 8977 6360
rect 9011 6326 9045 6360
rect 9079 6326 9113 6360
rect 9147 6326 9181 6360
rect 9215 6326 9249 6360
rect 9283 6326 9317 6360
rect 9351 6326 9385 6360
rect 9419 6326 9453 6360
rect 9487 6326 9521 6360
rect 9555 6326 9589 6360
rect 9623 6326 9657 6360
rect 9691 6326 9725 6360
rect 9759 6326 9793 6360
rect 9827 6326 9861 6360
rect 9895 6326 9929 6360
rect 9963 6326 9997 6360
rect 10031 6326 10065 6360
rect 10099 6326 10133 6360
rect 10167 6326 10201 6360
rect 10235 6326 10269 6360
rect 10303 6326 10337 6360
rect 10371 6326 10405 6360
rect 10439 6326 10473 6360
rect 10507 6326 10541 6360
rect 10575 6326 10609 6360
rect 10643 6326 10677 6360
rect 10711 6326 10745 6360
rect 10779 6326 10813 6360
rect 10847 6326 10881 6360
rect 10915 6326 10949 6360
rect 10983 6326 11017 6360
rect 11051 6326 11085 6360
rect 11119 6326 11153 6360
rect 11187 6326 11221 6360
rect 11255 6326 11289 6360
rect 11323 6326 11357 6360
rect 11391 6326 11425 6360
rect 11459 6326 11493 6360
rect 11527 6326 11561 6360
rect 11595 6326 11629 6360
rect 11663 6326 11697 6360
rect 11731 6326 11765 6360
rect 11799 6326 11833 6360
rect 11867 6326 11901 6360
rect 11935 6326 11969 6360
rect 12003 6326 12037 6360
rect 12071 6326 12105 6360
rect 12139 6326 12173 6360
rect 12207 6326 12241 6360
rect 12275 6326 12309 6360
rect 12343 6326 12377 6360
rect 12411 6326 12445 6360
rect 12479 6326 12513 6360
rect 12547 6326 12581 6360
rect 12615 6326 12649 6360
rect 12683 6326 12717 6360
rect 12751 6326 12785 6360
rect 12819 6326 12853 6360
rect 12887 6326 12921 6360
rect 12955 6326 12989 6360
rect 13023 6326 13057 6360
rect 13091 6326 13125 6360
rect 13159 6326 13193 6360
rect 13227 6326 13261 6360
rect 13295 6326 13329 6360
rect 13363 6326 13397 6360
rect 13431 6326 13465 6360
rect 13499 6326 13533 6360
rect 13567 6326 13601 6360
rect 13635 6326 13669 6360
rect 13703 6326 13737 6360
rect 13771 6326 13805 6360
rect 13839 6326 13873 6360
rect 13907 6326 13941 6360
rect 13975 6326 14009 6360
rect 14043 6326 14077 6360
rect 14111 6326 14145 6360
rect 14179 6326 14213 6360
rect 14247 6326 14281 6360
rect 14315 6326 14349 6360
rect 14383 6326 14417 6360
rect 14451 6326 14485 6360
rect 14519 6326 14553 6360
rect 14587 6326 14621 6360
rect 14655 6326 14689 6360
rect 14723 6326 14757 6360
rect 14791 6326 14825 6360
rect 14859 6326 14893 6360
rect 14932 6326 14966 6360
rect 15000 6326 15034 6360
rect 15068 6326 15102 6360
rect 68 6252 102 6286
rect 137 6252 171 6286
rect 206 6252 240 6286
rect 275 6252 309 6286
rect 344 6252 378 6286
rect 413 6252 447 6286
rect 482 6252 516 6286
rect 551 6252 585 6286
rect 620 6252 654 6286
rect 689 6252 723 6286
rect 758 6252 792 6286
rect 827 6252 861 6286
rect 896 6252 930 6286
rect 965 6252 999 6286
rect 1034 6252 1068 6286
rect 1103 6252 1137 6286
rect 1172 6252 1206 6286
rect 1241 6252 1275 6286
rect 1310 6252 1344 6286
rect 1379 6252 1413 6286
rect 1448 6252 1482 6286
rect 1517 6252 1551 6286
rect 1586 6252 1620 6286
rect 1655 6252 1689 6286
rect 1724 6252 1758 6286
rect 1793 6252 1827 6286
rect 1862 6252 1896 6286
rect 1931 6252 1965 6286
rect 2000 6252 2034 6286
rect 2069 6252 2103 6286
rect 2138 6252 2172 6286
rect 2207 6252 2241 6286
rect 2276 6252 2310 6286
rect 2345 6252 2379 6286
rect 2414 6252 2448 6286
rect 2483 6252 2517 6286
rect 2551 6252 2585 6286
rect 2619 6252 2653 6286
rect 2687 6252 2721 6286
rect 2755 6252 2789 6286
rect 2823 6252 2857 6286
rect 2891 6252 2925 6286
rect 2959 6252 2993 6286
rect 3027 6252 3061 6286
rect 3095 6252 3129 6286
rect 3163 6252 3197 6286
rect 3231 6252 3265 6286
rect 3299 6252 3333 6286
rect 3367 6252 3401 6286
rect 3435 6252 3469 6286
rect 3503 6252 3537 6286
rect 3571 6252 3605 6286
rect 3639 6252 3673 6286
rect 3707 6252 3741 6286
rect 3775 6252 3809 6286
rect 3843 6252 3877 6286
rect 3911 6252 3945 6286
rect 3979 6252 4013 6286
rect 4047 6252 4081 6286
rect 4115 6252 4149 6286
rect 4183 6252 4217 6286
rect 4251 6252 4285 6286
rect 4319 6252 4353 6286
rect 4387 6252 4421 6286
rect 4455 6252 4489 6286
rect 4523 6252 4557 6286
rect 4591 6252 4625 6286
rect 4659 6252 4693 6286
rect 4727 6252 4761 6286
rect 4795 6252 4829 6286
rect 4863 6252 4897 6286
rect 4931 6252 4965 6286
rect 4999 6252 5033 6286
rect 5067 6252 5101 6286
rect 5135 6252 5169 6286
rect 5203 6252 5237 6286
rect 5271 6252 5305 6286
rect 5339 6252 5373 6286
rect 5407 6252 5441 6286
rect 5475 6252 5509 6286
rect 5543 6252 5577 6286
rect 5611 6252 5645 6286
rect 5679 6252 5713 6286
rect 5747 6252 5781 6286
rect 5815 6252 5849 6286
rect 5883 6252 5917 6286
rect 5951 6252 5985 6286
rect 6019 6252 6053 6286
rect 6087 6252 6121 6286
rect 6155 6252 6189 6286
rect 6223 6252 6257 6286
rect 6291 6252 6325 6286
rect 6359 6252 6393 6286
rect 6427 6252 6461 6286
rect 6495 6252 6529 6286
rect 6563 6252 6597 6286
rect 6631 6252 6665 6286
rect 6699 6252 6733 6286
rect 6767 6252 6801 6286
rect 6835 6252 6869 6286
rect 6903 6252 6937 6286
rect 6971 6252 7005 6286
rect 7039 6252 7073 6286
rect 7107 6252 7141 6286
rect 7175 6252 7209 6286
rect 7243 6252 7277 6286
rect 7311 6252 7345 6286
rect 7379 6252 7413 6286
rect 7447 6252 7481 6286
rect 7515 6252 7549 6286
rect 7583 6252 7617 6286
rect 7651 6252 7685 6286
rect 7719 6252 7753 6286
rect 7787 6252 7821 6286
rect 7855 6252 7889 6286
rect 7923 6252 7957 6286
rect 7991 6252 8025 6286
rect 8059 6252 8093 6286
rect 8127 6252 8161 6286
rect 8195 6252 8229 6286
rect 8263 6252 8297 6286
rect 8331 6252 8365 6286
rect 8399 6252 8433 6286
rect 8467 6252 8501 6286
rect 8535 6252 8569 6286
rect 8603 6252 8637 6286
rect 8671 6252 8705 6286
rect 8739 6252 8773 6286
rect 8807 6252 8841 6286
rect 8875 6252 8909 6286
rect 8943 6252 8977 6286
rect 9011 6252 9045 6286
rect 9079 6252 9113 6286
rect 9147 6252 9181 6286
rect 9215 6252 9249 6286
rect 9283 6252 9317 6286
rect 9351 6252 9385 6286
rect 9419 6252 9453 6286
rect 9487 6252 9521 6286
rect 9555 6252 9589 6286
rect 9623 6252 9657 6286
rect 9691 6252 9725 6286
rect 9759 6252 9793 6286
rect 9827 6252 9861 6286
rect 9895 6252 9929 6286
rect 9963 6252 9997 6286
rect 10031 6252 10065 6286
rect 10099 6252 10133 6286
rect 10167 6252 10201 6286
rect 10235 6252 10269 6286
rect 10303 6252 10337 6286
rect 10371 6252 10405 6286
rect 10439 6252 10473 6286
rect 10507 6252 10541 6286
rect 10575 6252 10609 6286
rect 10643 6252 10677 6286
rect 10711 6252 10745 6286
rect 10779 6252 10813 6286
rect 10847 6252 10881 6286
rect 10915 6252 10949 6286
rect 10983 6252 11017 6286
rect 11051 6252 11085 6286
rect 11119 6252 11153 6286
rect 11187 6252 11221 6286
rect 11255 6252 11289 6286
rect 11323 6252 11357 6286
rect 11391 6252 11425 6286
rect 11459 6252 11493 6286
rect 11527 6252 11561 6286
rect 11595 6252 11629 6286
rect 11663 6252 11697 6286
rect 11731 6252 11765 6286
rect 11799 6252 11833 6286
rect 11867 6252 11901 6286
rect 11935 6252 11969 6286
rect 12003 6252 12037 6286
rect 12071 6252 12105 6286
rect 12139 6252 12173 6286
rect 12207 6252 12241 6286
rect 12275 6252 12309 6286
rect 12343 6252 12377 6286
rect 12411 6252 12445 6286
rect 12479 6252 12513 6286
rect 12547 6252 12581 6286
rect 12615 6252 12649 6286
rect 12683 6252 12717 6286
rect 12751 6252 12785 6286
rect 12819 6252 12853 6286
rect 12887 6252 12921 6286
rect 12955 6252 12989 6286
rect 13023 6252 13057 6286
rect 13091 6252 13125 6286
rect 13159 6252 13193 6286
rect 13227 6252 13261 6286
rect 13295 6252 13329 6286
rect 13363 6252 13397 6286
rect 13431 6252 13465 6286
rect 13499 6252 13533 6286
rect 13567 6252 13601 6286
rect 13635 6252 13669 6286
rect 13703 6252 13737 6286
rect 13771 6252 13805 6286
rect 13839 6252 13873 6286
rect 13907 6252 13941 6286
rect 13975 6252 14009 6286
rect 14043 6252 14077 6286
rect 14111 6252 14145 6286
rect 14179 6252 14213 6286
rect 14247 6252 14281 6286
rect 14315 6252 14349 6286
rect 14383 6252 14417 6286
rect 14451 6252 14485 6286
rect 14519 6252 14553 6286
rect 14587 6252 14621 6286
rect 14655 6252 14689 6286
rect 14723 6252 14757 6286
rect 14791 6252 14825 6286
rect 14859 6252 14893 6286
rect 14932 6251 14966 6285
rect 15000 6251 15034 6285
rect 15068 6251 15102 6285
rect 68 6178 102 6212
rect 137 6178 171 6212
rect 206 6178 240 6212
rect 275 6178 309 6212
rect 344 6178 378 6212
rect 413 6178 447 6212
rect 482 6178 516 6212
rect 551 6178 585 6212
rect 620 6178 654 6212
rect 689 6178 723 6212
rect 758 6178 792 6212
rect 827 6178 861 6212
rect 896 6178 930 6212
rect 965 6178 999 6212
rect 1034 6178 1068 6212
rect 1103 6178 1137 6212
rect 1172 6178 1206 6212
rect 1241 6178 1275 6212
rect 1310 6178 1344 6212
rect 1379 6178 1413 6212
rect 1448 6178 1482 6212
rect 1517 6178 1551 6212
rect 1586 6178 1620 6212
rect 1655 6178 1689 6212
rect 1724 6178 1758 6212
rect 1793 6178 1827 6212
rect 1862 6178 1896 6212
rect 1931 6178 1965 6212
rect 2000 6178 2034 6212
rect 2069 6178 2103 6212
rect 2138 6178 2172 6212
rect 2207 6178 2241 6212
rect 2276 6178 2310 6212
rect 2345 6178 2379 6212
rect 2414 6178 2448 6212
rect 2483 6178 2517 6212
rect 2551 6178 2585 6212
rect 2619 6178 2653 6212
rect 2687 6178 2721 6212
rect 2755 6178 2789 6212
rect 2823 6178 2857 6212
rect 2891 6178 2925 6212
rect 2959 6178 2993 6212
rect 3027 6178 3061 6212
rect 3095 6178 3129 6212
rect 3163 6178 3197 6212
rect 3231 6178 3265 6212
rect 3299 6178 3333 6212
rect 3367 6178 3401 6212
rect 3435 6178 3469 6212
rect 3503 6178 3537 6212
rect 3571 6178 3605 6212
rect 3639 6178 3673 6212
rect 3707 6178 3741 6212
rect 3775 6178 3809 6212
rect 3843 6178 3877 6212
rect 3911 6178 3945 6212
rect 3979 6178 4013 6212
rect 4047 6178 4081 6212
rect 4115 6178 4149 6212
rect 4183 6178 4217 6212
rect 4251 6178 4285 6212
rect 4319 6178 4353 6212
rect 4387 6178 4421 6212
rect 4455 6178 4489 6212
rect 4523 6178 4557 6212
rect 4591 6178 4625 6212
rect 4659 6178 4693 6212
rect 4727 6178 4761 6212
rect 4795 6178 4829 6212
rect 4863 6178 4897 6212
rect 4931 6178 4965 6212
rect 4999 6178 5033 6212
rect 5067 6178 5101 6212
rect 5135 6178 5169 6212
rect 5203 6178 5237 6212
rect 5271 6178 5305 6212
rect 5339 6178 5373 6212
rect 5407 6178 5441 6212
rect 5475 6178 5509 6212
rect 5543 6178 5577 6212
rect 5611 6178 5645 6212
rect 5679 6178 5713 6212
rect 5747 6178 5781 6212
rect 5815 6178 5849 6212
rect 5883 6178 5917 6212
rect 5951 6178 5985 6212
rect 6019 6178 6053 6212
rect 6087 6178 6121 6212
rect 6155 6178 6189 6212
rect 6223 6178 6257 6212
rect 6291 6178 6325 6212
rect 6359 6178 6393 6212
rect 6427 6178 6461 6212
rect 6495 6178 6529 6212
rect 6563 6178 6597 6212
rect 6631 6178 6665 6212
rect 6699 6178 6733 6212
rect 6767 6178 6801 6212
rect 6835 6178 6869 6212
rect 6903 6178 6937 6212
rect 6971 6178 7005 6212
rect 7039 6178 7073 6212
rect 7107 6178 7141 6212
rect 7175 6178 7209 6212
rect 7243 6178 7277 6212
rect 7311 6178 7345 6212
rect 7379 6178 7413 6212
rect 7447 6178 7481 6212
rect 7515 6178 7549 6212
rect 7583 6178 7617 6212
rect 7651 6178 7685 6212
rect 7719 6178 7753 6212
rect 7787 6178 7821 6212
rect 7855 6178 7889 6212
rect 7923 6178 7957 6212
rect 7991 6178 8025 6212
rect 8059 6178 8093 6212
rect 8127 6178 8161 6212
rect 8195 6178 8229 6212
rect 8263 6178 8297 6212
rect 8331 6178 8365 6212
rect 8399 6178 8433 6212
rect 8467 6178 8501 6212
rect 8535 6178 8569 6212
rect 8603 6178 8637 6212
rect 8671 6178 8705 6212
rect 8739 6178 8773 6212
rect 8807 6178 8841 6212
rect 8875 6178 8909 6212
rect 8943 6178 8977 6212
rect 9011 6178 9045 6212
rect 9079 6178 9113 6212
rect 9147 6178 9181 6212
rect 9215 6178 9249 6212
rect 9283 6178 9317 6212
rect 9351 6178 9385 6212
rect 9419 6178 9453 6212
rect 9487 6178 9521 6212
rect 9555 6178 9589 6212
rect 9623 6178 9657 6212
rect 9691 6178 9725 6212
rect 9759 6178 9793 6212
rect 9827 6178 9861 6212
rect 9895 6178 9929 6212
rect 9963 6178 9997 6212
rect 10031 6178 10065 6212
rect 10099 6178 10133 6212
rect 10167 6178 10201 6212
rect 10235 6178 10269 6212
rect 10303 6178 10337 6212
rect 10371 6178 10405 6212
rect 10439 6178 10473 6212
rect 10507 6178 10541 6212
rect 10575 6178 10609 6212
rect 10643 6178 10677 6212
rect 10711 6178 10745 6212
rect 10779 6178 10813 6212
rect 10847 6178 10881 6212
rect 10915 6178 10949 6212
rect 10983 6178 11017 6212
rect 11051 6178 11085 6212
rect 11119 6178 11153 6212
rect 11187 6178 11221 6212
rect 11255 6178 11289 6212
rect 11323 6178 11357 6212
rect 11391 6178 11425 6212
rect 11459 6178 11493 6212
rect 11527 6178 11561 6212
rect 11595 6178 11629 6212
rect 11663 6178 11697 6212
rect 11731 6178 11765 6212
rect 11799 6178 11833 6212
rect 11867 6178 11901 6212
rect 11935 6178 11969 6212
rect 12003 6178 12037 6212
rect 12071 6178 12105 6212
rect 12139 6178 12173 6212
rect 12207 6178 12241 6212
rect 12275 6178 12309 6212
rect 12343 6178 12377 6212
rect 12411 6178 12445 6212
rect 12479 6178 12513 6212
rect 12547 6178 12581 6212
rect 12615 6178 12649 6212
rect 12683 6178 12717 6212
rect 12751 6178 12785 6212
rect 12819 6178 12853 6212
rect 12887 6178 12921 6212
rect 12955 6178 12989 6212
rect 13023 6178 13057 6212
rect 13091 6178 13125 6212
rect 13159 6178 13193 6212
rect 13227 6178 13261 6212
rect 13295 6178 13329 6212
rect 13363 6178 13397 6212
rect 13431 6178 13465 6212
rect 13499 6178 13533 6212
rect 13567 6178 13601 6212
rect 13635 6178 13669 6212
rect 13703 6178 13737 6212
rect 13771 6178 13805 6212
rect 13839 6178 13873 6212
rect 13907 6178 13941 6212
rect 13975 6178 14009 6212
rect 14043 6178 14077 6212
rect 14111 6178 14145 6212
rect 14179 6178 14213 6212
rect 14247 6178 14281 6212
rect 14315 6178 14349 6212
rect 14383 6178 14417 6212
rect 14451 6178 14485 6212
rect 14519 6178 14553 6212
rect 14587 6178 14621 6212
rect 14655 6178 14689 6212
rect 14723 6178 14757 6212
rect 14791 6178 14825 6212
rect 14859 6178 14893 6212
rect 14932 6176 14966 6210
rect 15000 6176 15034 6210
rect 15068 6176 15102 6210
rect 68 6104 102 6138
rect 137 6104 171 6138
rect 206 6104 240 6138
rect 275 6104 309 6138
rect 344 6104 378 6138
rect 413 6104 447 6138
rect 482 6104 516 6138
rect 551 6104 585 6138
rect 620 6104 654 6138
rect 689 6104 723 6138
rect 758 6104 792 6138
rect 827 6104 861 6138
rect 896 6104 930 6138
rect 965 6104 999 6138
rect 1034 6104 1068 6138
rect 1103 6104 1137 6138
rect 1172 6104 1206 6138
rect 1241 6104 1275 6138
rect 1310 6104 1344 6138
rect 1379 6104 1413 6138
rect 1448 6104 1482 6138
rect 1517 6104 1551 6138
rect 1586 6104 1620 6138
rect 1655 6104 1689 6138
rect 1724 6104 1758 6138
rect 1793 6104 1827 6138
rect 1862 6104 1896 6138
rect 1931 6104 1965 6138
rect 2000 6104 2034 6138
rect 2069 6104 2103 6138
rect 2138 6104 2172 6138
rect 2207 6104 2241 6138
rect 2276 6104 2310 6138
rect 2345 6104 2379 6138
rect 2414 6104 2448 6138
rect 2483 6104 2517 6138
rect 2551 6104 2585 6138
rect 2619 6104 2653 6138
rect 2687 6104 2721 6138
rect 2755 6104 2789 6138
rect 2823 6104 2857 6138
rect 2891 6104 2925 6138
rect 2959 6104 2993 6138
rect 3027 6104 3061 6138
rect 3095 6104 3129 6138
rect 3163 6104 3197 6138
rect 3231 6104 3265 6138
rect 3299 6104 3333 6138
rect 3367 6104 3401 6138
rect 3435 6104 3469 6138
rect 3503 6104 3537 6138
rect 3571 6104 3605 6138
rect 3639 6104 3673 6138
rect 3707 6104 3741 6138
rect 3775 6104 3809 6138
rect 3843 6104 3877 6138
rect 3911 6104 3945 6138
rect 3979 6104 4013 6138
rect 4047 6104 4081 6138
rect 4115 6104 4149 6138
rect 4183 6104 4217 6138
rect 4251 6104 4285 6138
rect 4319 6104 4353 6138
rect 4387 6104 4421 6138
rect 4455 6104 4489 6138
rect 4523 6104 4557 6138
rect 4591 6104 4625 6138
rect 4659 6104 4693 6138
rect 4727 6104 4761 6138
rect 4795 6104 4829 6138
rect 4863 6104 4897 6138
rect 4931 6104 4965 6138
rect 4999 6104 5033 6138
rect 5067 6104 5101 6138
rect 5135 6104 5169 6138
rect 5203 6104 5237 6138
rect 5271 6104 5305 6138
rect 5339 6104 5373 6138
rect 5407 6104 5441 6138
rect 5475 6104 5509 6138
rect 5543 6104 5577 6138
rect 5611 6104 5645 6138
rect 5679 6104 5713 6138
rect 5747 6104 5781 6138
rect 5815 6104 5849 6138
rect 5883 6104 5917 6138
rect 5951 6104 5985 6138
rect 6019 6104 6053 6138
rect 6087 6104 6121 6138
rect 6155 6104 6189 6138
rect 6223 6104 6257 6138
rect 6291 6104 6325 6138
rect 6359 6104 6393 6138
rect 6427 6104 6461 6138
rect 6495 6104 6529 6138
rect 6563 6104 6597 6138
rect 6631 6104 6665 6138
rect 6699 6104 6733 6138
rect 6767 6104 6801 6138
rect 6835 6104 6869 6138
rect 6903 6104 6937 6138
rect 6971 6104 7005 6138
rect 7039 6104 7073 6138
rect 7107 6104 7141 6138
rect 7175 6104 7209 6138
rect 7243 6104 7277 6138
rect 7311 6104 7345 6138
rect 7379 6104 7413 6138
rect 7447 6104 7481 6138
rect 7515 6104 7549 6138
rect 7583 6104 7617 6138
rect 7651 6104 7685 6138
rect 7719 6104 7753 6138
rect 7787 6104 7821 6138
rect 7855 6104 7889 6138
rect 7923 6104 7957 6138
rect 7991 6104 8025 6138
rect 8059 6104 8093 6138
rect 8127 6104 8161 6138
rect 8195 6104 8229 6138
rect 8263 6104 8297 6138
rect 8331 6104 8365 6138
rect 8399 6104 8433 6138
rect 8467 6104 8501 6138
rect 8535 6104 8569 6138
rect 8603 6104 8637 6138
rect 8671 6104 8705 6138
rect 8739 6104 8773 6138
rect 8807 6104 8841 6138
rect 8875 6104 8909 6138
rect 8943 6104 8977 6138
rect 9011 6104 9045 6138
rect 9079 6104 9113 6138
rect 9147 6104 9181 6138
rect 9215 6104 9249 6138
rect 9283 6104 9317 6138
rect 9351 6104 9385 6138
rect 9419 6104 9453 6138
rect 9487 6104 9521 6138
rect 9555 6104 9589 6138
rect 9623 6104 9657 6138
rect 9691 6104 9725 6138
rect 9759 6104 9793 6138
rect 9827 6104 9861 6138
rect 9895 6104 9929 6138
rect 9963 6104 9997 6138
rect 10031 6104 10065 6138
rect 10099 6104 10133 6138
rect 10167 6104 10201 6138
rect 10235 6104 10269 6138
rect 10303 6104 10337 6138
rect 10371 6104 10405 6138
rect 10439 6104 10473 6138
rect 10507 6104 10541 6138
rect 10575 6104 10609 6138
rect 10643 6104 10677 6138
rect 10711 6104 10745 6138
rect 10779 6104 10813 6138
rect 10847 6104 10881 6138
rect 10915 6104 10949 6138
rect 10983 6104 11017 6138
rect 11051 6104 11085 6138
rect 11119 6104 11153 6138
rect 11187 6104 11221 6138
rect 11255 6104 11289 6138
rect 11323 6104 11357 6138
rect 11391 6104 11425 6138
rect 11459 6104 11493 6138
rect 11527 6104 11561 6138
rect 11595 6104 11629 6138
rect 11663 6104 11697 6138
rect 11731 6104 11765 6138
rect 11799 6104 11833 6138
rect 11867 6104 11901 6138
rect 11935 6104 11969 6138
rect 12003 6104 12037 6138
rect 12071 6104 12105 6138
rect 12139 6104 12173 6138
rect 12207 6104 12241 6138
rect 12275 6104 12309 6138
rect 12343 6104 12377 6138
rect 12411 6104 12445 6138
rect 12479 6104 12513 6138
rect 12547 6104 12581 6138
rect 12615 6104 12649 6138
rect 12683 6104 12717 6138
rect 12751 6104 12785 6138
rect 12819 6104 12853 6138
rect 12887 6104 12921 6138
rect 12955 6104 12989 6138
rect 13023 6104 13057 6138
rect 13091 6104 13125 6138
rect 13159 6104 13193 6138
rect 13227 6104 13261 6138
rect 13295 6104 13329 6138
rect 13363 6104 13397 6138
rect 13431 6104 13465 6138
rect 13499 6104 13533 6138
rect 13567 6104 13601 6138
rect 13635 6104 13669 6138
rect 13703 6104 13737 6138
rect 13771 6104 13805 6138
rect 13839 6104 13873 6138
rect 13907 6104 13941 6138
rect 13975 6104 14009 6138
rect 14043 6104 14077 6138
rect 14111 6104 14145 6138
rect 14179 6104 14213 6138
rect 14247 6104 14281 6138
rect 14315 6104 14349 6138
rect 14383 6104 14417 6138
rect 14451 6104 14485 6138
rect 14519 6104 14553 6138
rect 14587 6104 14621 6138
rect 14655 6104 14689 6138
rect 14723 6104 14757 6138
rect 14791 6104 14825 6138
rect 14859 6104 14893 6138
rect 14932 6101 14966 6135
rect 15000 6101 15034 6135
rect 15068 6101 15102 6135
rect 14932 6026 14966 6060
rect 15000 6026 15034 6060
rect 15068 6026 15102 6060
rect 15000 4628 15102 5954
rect 15000 4559 15034 4593
rect 15068 4559 15102 4593
rect 15000 4490 15034 4524
rect 15068 4490 15102 4524
rect 15000 4421 15034 4455
rect 15068 4421 15102 4455
rect 15000 4352 15034 4386
rect 15068 4352 15102 4386
rect 15000 4283 15034 4317
rect 15068 4283 15102 4317
rect 15000 4214 15034 4248
rect 15068 4214 15102 4248
rect 15000 4145 15034 4179
rect 15068 4145 15102 4179
rect 15000 4076 15034 4110
rect 15068 4076 15102 4110
rect 15000 4007 15034 4041
rect 15068 4007 15102 4041
rect 15000 3938 15034 3972
rect 15068 3938 15102 3972
rect 15000 3869 15034 3903
rect 15068 3869 15102 3903
rect 15000 3800 15034 3834
rect 15068 3800 15102 3834
rect 15000 3731 15034 3765
rect 15068 3731 15102 3765
rect 15000 3662 15034 3696
rect 15068 3662 15102 3696
rect 15000 3593 15034 3627
rect 15068 3593 15102 3627
rect 15000 3524 15034 3558
rect 15068 3524 15102 3558
rect 15000 3455 15034 3489
rect 15068 3455 15102 3489
rect 15000 3386 15034 3420
rect 15068 3386 15102 3420
rect 15000 3317 15034 3351
rect 15068 3317 15102 3351
rect 15000 3248 15034 3282
rect 15068 3248 15102 3282
rect 15000 3179 15034 3213
rect 15068 3179 15102 3213
rect 15000 3110 15034 3144
rect 15068 3110 15102 3144
rect 15000 3041 15034 3075
rect 15068 3041 15102 3075
rect 15000 2972 15034 3006
rect 15068 2972 15102 3006
rect 15000 2903 15034 2937
rect 15068 2903 15102 2937
rect 15000 2834 15034 2868
rect 15068 2834 15102 2868
rect 15000 2765 15034 2799
rect 15068 2765 15102 2799
rect 15000 2696 15034 2730
rect 15068 2696 15102 2730
rect 15000 2627 15034 2661
rect 15068 2627 15102 2661
rect 15000 2558 15034 2592
rect 15068 2558 15102 2592
rect 15000 2489 15034 2523
rect 15068 2489 15102 2523
rect 15000 2420 15034 2454
rect 15068 2420 15102 2454
rect 15000 2351 15034 2385
rect 15068 2351 15102 2385
rect 15000 2282 15034 2316
rect 15068 2282 15102 2316
rect 15000 2213 15034 2247
rect 15068 2213 15102 2247
rect 15000 2144 15034 2178
rect 15068 2144 15102 2178
rect 15000 2075 15034 2109
rect 15068 2075 15102 2109
rect 15000 2006 15034 2040
rect 15068 2006 15102 2040
rect 15000 1937 15034 1971
rect 15068 1937 15102 1971
rect 15000 1868 15034 1902
rect 15068 1868 15102 1902
rect 15000 1799 15034 1833
rect 15068 1799 15102 1833
rect 15000 1730 15034 1764
rect 15068 1730 15102 1764
rect 15000 1661 15034 1695
rect 15068 1661 15102 1695
rect 15000 1592 15034 1626
rect 15068 1592 15102 1626
rect 15000 1523 15034 1557
rect 15068 1523 15102 1557
rect 15000 1454 15034 1488
rect 15068 1454 15102 1488
rect 15000 1385 15034 1419
rect 15068 1385 15102 1419
rect 15000 1316 15034 1350
rect 15068 1316 15102 1350
rect 7068 1223 7102 1257
rect 7137 1223 7171 1257
rect 7206 1223 7240 1257
rect 7275 1223 7309 1257
rect 7344 1223 7378 1257
rect 7413 1223 7447 1257
rect 7482 1223 7516 1257
rect 7551 1223 7585 1257
rect 7620 1223 7654 1257
rect 7689 1223 7723 1257
rect 7758 1223 7792 1257
rect 7827 1223 7861 1257
rect 7896 1223 7930 1257
rect 7965 1223 7999 1257
rect 8034 1223 8068 1257
rect 8103 1223 8137 1257
rect 8172 1223 8206 1257
rect 8241 1223 8275 1257
rect 8310 1223 8344 1257
rect 8379 1223 8413 1257
rect 8448 1223 8482 1257
rect 8517 1223 8551 1257
rect 8586 1223 8620 1257
rect 8655 1223 8689 1257
rect 8724 1223 8758 1257
rect 8793 1223 8827 1257
rect 8862 1223 8896 1257
rect 8931 1223 8965 1257
rect 9000 1223 9034 1257
rect 9069 1223 9103 1257
rect 9138 1223 9172 1257
rect 9207 1223 9241 1257
rect 9276 1223 9310 1257
rect 9345 1223 9379 1257
rect 9414 1223 9448 1257
rect 9483 1223 9517 1257
rect 9552 1223 9586 1257
rect 9621 1223 9655 1257
rect 9690 1223 9724 1257
rect 7068 1155 7102 1189
rect 7137 1155 7171 1189
rect 7206 1155 7240 1189
rect 7275 1155 7309 1189
rect 7344 1155 7378 1189
rect 7413 1155 7447 1189
rect 7482 1155 7516 1189
rect 7551 1155 7585 1189
rect 7620 1155 7654 1189
rect 7689 1155 7723 1189
rect 7758 1155 7792 1189
rect 7827 1155 7861 1189
rect 7896 1155 7930 1189
rect 7965 1155 7999 1189
rect 8034 1155 8068 1189
rect 8103 1155 8137 1189
rect 8172 1155 8206 1189
rect 8241 1155 8275 1189
rect 8310 1155 8344 1189
rect 8379 1155 8413 1189
rect 8448 1155 8482 1189
rect 8517 1155 8551 1189
rect 8586 1155 8620 1189
rect 8655 1155 8689 1189
rect 8724 1155 8758 1189
rect 8793 1155 8827 1189
rect 8862 1155 8896 1189
rect 8931 1155 8965 1189
rect 9000 1155 9034 1189
rect 9069 1155 9103 1189
rect 9138 1155 9172 1189
rect 9207 1155 9241 1189
rect 9276 1155 9310 1189
rect 9345 1155 9379 1189
rect 9414 1155 9448 1189
rect 9483 1155 9517 1189
rect 9552 1155 9586 1189
rect 9621 1155 9655 1189
rect 9690 1155 9724 1189
rect 7068 1087 7102 1121
rect 7137 1087 7171 1121
rect 7206 1087 7240 1121
rect 7275 1087 7309 1121
rect 7344 1087 7378 1121
rect 7413 1087 7447 1121
rect 7482 1087 7516 1121
rect 7551 1087 7585 1121
rect 7620 1087 7654 1121
rect 7689 1087 7723 1121
rect 7758 1087 7792 1121
rect 7827 1087 7861 1121
rect 7896 1087 7930 1121
rect 7965 1087 7999 1121
rect 8034 1087 8068 1121
rect 8103 1087 8137 1121
rect 8172 1087 8206 1121
rect 8241 1087 8275 1121
rect 8310 1087 8344 1121
rect 8379 1087 8413 1121
rect 8448 1087 8482 1121
rect 8517 1087 8551 1121
rect 8586 1087 8620 1121
rect 8655 1087 8689 1121
rect 8724 1087 8758 1121
rect 8793 1087 8827 1121
rect 8862 1087 8896 1121
rect 8931 1087 8965 1121
rect 9000 1087 9034 1121
rect 9069 1087 9103 1121
rect 9138 1087 9172 1121
rect 9207 1087 9241 1121
rect 9276 1087 9310 1121
rect 9345 1087 9379 1121
rect 9414 1087 9448 1121
rect 9483 1087 9517 1121
rect 9552 1087 9586 1121
rect 9621 1087 9655 1121
rect 9690 1087 9724 1121
rect 7068 1019 7102 1053
rect 7137 1019 7171 1053
rect 7206 1019 7240 1053
rect 7275 1019 7309 1053
rect 7344 1019 7378 1053
rect 7413 1019 7447 1053
rect 7482 1019 7516 1053
rect 7551 1019 7585 1053
rect 7620 1019 7654 1053
rect 7689 1019 7723 1053
rect 7758 1019 7792 1053
rect 7827 1019 7861 1053
rect 7896 1019 7930 1053
rect 7965 1019 7999 1053
rect 8034 1019 8068 1053
rect 8103 1019 8137 1053
rect 8172 1019 8206 1053
rect 8241 1019 8275 1053
rect 8310 1019 8344 1053
rect 8379 1019 8413 1053
rect 8448 1019 8482 1053
rect 8517 1019 8551 1053
rect 8586 1019 8620 1053
rect 8655 1019 8689 1053
rect 8724 1019 8758 1053
rect 8793 1019 8827 1053
rect 8862 1019 8896 1053
rect 8931 1019 8965 1053
rect 9000 1019 9034 1053
rect 9069 1019 9103 1053
rect 9138 1019 9172 1053
rect 9207 1019 9241 1053
rect 9276 1019 9310 1053
rect 9345 1019 9379 1053
rect 9414 1019 9448 1053
rect 9483 1019 9517 1053
rect 9552 1019 9586 1053
rect 9621 1019 9655 1053
rect 9690 1019 9724 1053
rect 9759 1019 14893 1257
rect 14932 1210 14966 1244
rect 15000 1210 15034 1244
rect 15068 1210 15102 1244
rect 14932 1138 14966 1172
rect 15000 1138 15034 1172
rect 15068 1138 15102 1172
rect 14932 1066 14966 1100
rect 15000 1066 15034 1100
rect 15068 1066 15102 1100
rect 14932 994 14966 1028
rect 15000 994 15034 1028
rect 15068 994 15102 1028
rect 7067 913 7101 947
rect 7137 913 7171 947
rect 7207 913 7241 947
rect 7277 913 7311 947
rect 7347 913 7381 947
rect 7417 913 7451 947
rect 7487 913 7521 947
rect 7557 913 7591 947
rect 7627 913 7661 947
rect 7696 913 7730 947
rect 7067 841 7101 875
rect 7137 841 7171 875
rect 7207 841 7241 875
rect 7277 841 7311 875
rect 7347 841 7381 875
rect 7417 841 7451 875
rect 7487 841 7521 875
rect 7557 841 7591 875
rect 7627 841 7661 875
rect 7696 841 7730 875
rect 7067 769 7101 803
rect 7137 769 7171 803
rect 7207 769 7241 803
rect 7277 769 7311 803
rect 7347 769 7381 803
rect 7417 769 7451 803
rect 7487 769 7521 803
rect 7557 769 7591 803
rect 7627 769 7661 803
rect 7696 769 7730 803
rect 7067 697 7101 731
rect 7137 697 7171 731
rect 7207 697 7241 731
rect 7277 697 7311 731
rect 7347 697 7381 731
rect 7417 697 7451 731
rect 7487 697 7521 731
rect 7557 697 7591 731
rect 7627 697 7661 731
rect 7696 697 7730 731
rect 7067 625 7101 659
rect 7137 625 7171 659
rect 7207 625 7241 659
rect 7277 625 7311 659
rect 7347 625 7381 659
rect 7417 625 7451 659
rect 7487 625 7521 659
rect 7557 625 7591 659
rect 7627 625 7661 659
rect 7696 625 7730 659
rect 7067 553 7101 587
rect 7137 553 7171 587
rect 7207 553 7241 587
rect 7277 553 7311 587
rect 7347 553 7381 587
rect 7417 553 7451 587
rect 7487 553 7521 587
rect 7557 553 7591 587
rect 7627 553 7661 587
rect 7696 553 7730 587
rect 7067 481 7101 515
rect 7137 481 7171 515
rect 7207 481 7241 515
rect 7277 481 7311 515
rect 7347 481 7381 515
rect 7417 481 7451 515
rect 7487 481 7521 515
rect 7557 481 7591 515
rect 7627 481 7661 515
rect 7696 481 7730 515
rect 7067 409 7101 443
rect 7137 409 7171 443
rect 7207 409 7241 443
rect 7277 409 7311 443
rect 7347 409 7381 443
rect 7417 409 7451 443
rect 7487 409 7521 443
rect 7557 409 7591 443
rect 7627 409 7661 443
rect 7696 409 7730 443
rect 9711 913 9745 947
rect 9781 913 9815 947
rect 9851 913 9885 947
rect 9921 913 9955 947
rect 9991 913 10025 947
rect 10061 913 10095 947
rect 10131 913 10165 947
rect 10201 913 10235 947
rect 10271 913 10305 947
rect 10341 913 10375 947
rect 10411 913 10445 947
rect 10481 913 10515 947
rect 10551 913 10585 947
rect 10621 913 10655 947
rect 10691 913 10725 947
rect 10761 913 10795 947
rect 10831 913 10865 947
rect 10901 913 10935 947
rect 10971 913 11005 947
rect 11041 913 11075 947
rect 11111 913 11145 947
rect 11181 913 11215 947
rect 11251 913 11285 947
rect 11321 913 11355 947
rect 11391 913 11425 947
rect 11460 913 11494 947
rect 11529 913 11563 947
rect 11598 913 11632 947
rect 11680 921 11714 955
rect 11750 921 11784 955
rect 11820 921 11854 955
rect 11890 921 11924 955
rect 11960 921 11994 955
rect 12030 921 12064 955
rect 12099 921 12133 955
rect 12168 921 12202 955
rect 12237 921 12271 955
rect 12306 921 12340 955
rect 12375 921 12409 955
rect 12444 921 12478 955
rect 12513 921 12547 955
rect 12582 921 12616 955
rect 12651 921 12685 955
rect 12720 921 12754 955
rect 12789 921 12823 955
rect 12858 921 12892 955
rect 12927 921 12961 955
rect 12996 921 13030 955
rect 13065 921 13099 955
rect 13134 921 13168 955
rect 13203 921 13237 955
rect 13272 921 13306 955
rect 13341 921 13375 955
rect 13410 921 13444 955
rect 13479 921 13513 955
rect 13548 921 13582 955
rect 13617 921 13651 955
rect 13686 921 13720 955
rect 13755 921 13789 955
rect 13824 921 13858 955
rect 13893 921 13927 955
rect 13962 921 13996 955
rect 14031 921 14065 955
rect 14100 921 14134 955
rect 14169 921 14203 955
rect 14238 921 14272 955
rect 14307 921 14341 955
rect 14376 921 14410 955
rect 14445 921 14479 955
rect 14514 921 14548 955
rect 14583 921 14617 955
rect 14652 921 14686 955
rect 14721 921 14755 955
rect 14790 921 14824 955
rect 14859 921 14893 955
rect 14932 922 14966 956
rect 15000 922 15034 956
rect 15068 922 15102 956
rect 9711 841 9745 875
rect 9781 841 9815 875
rect 9851 841 9885 875
rect 9921 841 9955 875
rect 9991 841 10025 875
rect 10061 841 10095 875
rect 10131 841 10165 875
rect 10201 841 10235 875
rect 10271 841 10305 875
rect 10341 841 10375 875
rect 10411 841 10445 875
rect 10481 841 10515 875
rect 10551 841 10585 875
rect 10621 841 10655 875
rect 10691 841 10725 875
rect 10761 841 10795 875
rect 10831 841 10865 875
rect 10901 841 10935 875
rect 10971 841 11005 875
rect 11041 841 11075 875
rect 11111 841 11145 875
rect 11181 841 11215 875
rect 11251 841 11285 875
rect 11321 841 11355 875
rect 11391 841 11425 875
rect 11460 841 11494 875
rect 11529 841 11563 875
rect 11598 841 11632 875
rect 11680 841 11714 875
rect 11750 841 11784 875
rect 11820 841 11854 875
rect 11890 841 11924 875
rect 11960 841 11994 875
rect 12030 841 12064 875
rect 12099 841 12133 875
rect 12168 841 12202 875
rect 12237 841 12271 875
rect 12306 841 12340 875
rect 12375 841 12409 875
rect 12444 841 12478 875
rect 12513 841 12547 875
rect 12582 841 12616 875
rect 12651 841 12685 875
rect 12720 841 12754 875
rect 12789 841 12823 875
rect 12858 841 12892 875
rect 12927 841 12961 875
rect 12996 841 13030 875
rect 13065 841 13099 875
rect 13134 841 13168 875
rect 13203 841 13237 875
rect 13272 841 13306 875
rect 13341 841 13375 875
rect 13410 841 13444 875
rect 13479 841 13513 875
rect 13548 841 13582 875
rect 13617 841 13651 875
rect 13686 841 13720 875
rect 13755 841 13789 875
rect 13824 841 13858 875
rect 13893 841 13927 875
rect 13962 841 13996 875
rect 14031 841 14065 875
rect 14100 841 14134 875
rect 14169 841 14203 875
rect 14238 841 14272 875
rect 14307 841 14341 875
rect 14376 841 14410 875
rect 14445 841 14479 875
rect 14514 841 14548 875
rect 14583 841 14617 875
rect 14652 841 14686 875
rect 14721 841 14755 875
rect 14790 841 14824 875
rect 14859 841 14893 875
rect 14932 850 14966 884
rect 15000 850 15034 884
rect 15068 850 15102 884
rect 9711 769 9745 803
rect 9781 769 9815 803
rect 9851 769 9885 803
rect 9921 769 9955 803
rect 9991 769 10025 803
rect 10061 769 10095 803
rect 10131 769 10165 803
rect 10201 769 10235 803
rect 10271 769 10305 803
rect 10341 769 10375 803
rect 10411 769 10445 803
rect 10481 769 10515 803
rect 10551 769 10585 803
rect 10621 769 10655 803
rect 10691 769 10725 803
rect 10761 769 10795 803
rect 10831 769 10865 803
rect 10901 769 10935 803
rect 10971 769 11005 803
rect 11041 769 11075 803
rect 11111 769 11145 803
rect 11181 769 11215 803
rect 11251 769 11285 803
rect 11321 769 11355 803
rect 11391 769 11425 803
rect 11460 769 11494 803
rect 11529 769 11563 803
rect 11598 769 11632 803
rect 11680 761 11714 795
rect 11750 761 11784 795
rect 11820 761 11854 795
rect 11890 761 11924 795
rect 11960 761 11994 795
rect 12030 761 12064 795
rect 12099 761 12133 795
rect 12168 761 12202 795
rect 12237 761 12271 795
rect 12306 761 12340 795
rect 12375 761 12409 795
rect 12444 761 12478 795
rect 12513 761 12547 795
rect 12582 761 12616 795
rect 12651 761 12685 795
rect 12720 761 12754 795
rect 12789 761 12823 795
rect 12858 761 12892 795
rect 12927 761 12961 795
rect 12996 761 13030 795
rect 13065 761 13099 795
rect 13134 761 13168 795
rect 13203 761 13237 795
rect 13272 761 13306 795
rect 13341 761 13375 795
rect 13410 761 13444 795
rect 13479 761 13513 795
rect 13548 761 13582 795
rect 13617 761 13651 795
rect 13686 761 13720 795
rect 13755 761 13789 795
rect 13824 761 13858 795
rect 13893 761 13927 795
rect 13962 761 13996 795
rect 14031 761 14065 795
rect 14100 761 14134 795
rect 14169 761 14203 795
rect 14238 761 14272 795
rect 14307 761 14341 795
rect 14376 761 14410 795
rect 14445 761 14479 795
rect 14514 761 14548 795
rect 14583 761 14617 795
rect 14652 761 14686 795
rect 14721 761 14755 795
rect 14790 761 14824 795
rect 14859 761 14893 795
rect 14932 778 14966 812
rect 15000 778 15034 812
rect 15068 778 15102 812
rect 9711 697 9745 731
rect 9781 697 9815 731
rect 9851 697 9885 731
rect 9921 697 9955 731
rect 9991 697 10025 731
rect 10061 697 10095 731
rect 10131 697 10165 731
rect 10201 697 10235 731
rect 10271 697 10305 731
rect 10341 697 10375 731
rect 10411 697 10445 731
rect 10481 697 10515 731
rect 10551 697 10585 731
rect 10621 697 10655 731
rect 10691 697 10725 731
rect 10761 697 10795 731
rect 10831 697 10865 731
rect 10901 697 10935 731
rect 10971 697 11005 731
rect 11041 697 11075 731
rect 11111 697 11145 731
rect 11181 697 11215 731
rect 11251 697 11285 731
rect 11321 697 11355 731
rect 11391 697 11425 731
rect 11460 697 11494 731
rect 11529 697 11563 731
rect 11598 697 11632 731
rect 9711 625 9745 659
rect 9781 625 9815 659
rect 9851 625 9885 659
rect 9921 625 9955 659
rect 9991 625 10025 659
rect 10061 625 10095 659
rect 10131 625 10165 659
rect 10201 625 10235 659
rect 10271 625 10305 659
rect 10341 625 10375 659
rect 10411 625 10445 659
rect 10481 625 10515 659
rect 10551 625 10585 659
rect 10621 625 10655 659
rect 10691 625 10725 659
rect 10761 625 10795 659
rect 10831 625 10865 659
rect 10901 625 10935 659
rect 10971 625 11005 659
rect 11041 625 11075 659
rect 11111 625 11145 659
rect 11181 625 11215 659
rect 11251 625 11285 659
rect 11321 625 11355 659
rect 11391 625 11425 659
rect 11460 625 11494 659
rect 11529 625 11563 659
rect 11598 625 11632 659
rect 9711 553 9745 587
rect 9781 553 9815 587
rect 9851 553 9885 587
rect 9921 553 9955 587
rect 9991 553 10025 587
rect 10061 553 10095 587
rect 10131 553 10165 587
rect 10201 553 10235 587
rect 10271 553 10305 587
rect 10341 553 10375 587
rect 10411 553 10445 587
rect 10481 553 10515 587
rect 10551 553 10585 587
rect 10621 553 10655 587
rect 10691 553 10725 587
rect 10761 553 10795 587
rect 10831 553 10865 587
rect 10901 553 10935 587
rect 10971 553 11005 587
rect 11041 553 11075 587
rect 11111 553 11145 587
rect 11181 553 11215 587
rect 11251 553 11285 587
rect 11321 553 11355 587
rect 11391 553 11425 587
rect 11460 553 11494 587
rect 11529 553 11563 587
rect 11598 553 11632 587
rect 9711 481 9745 515
rect 9781 481 9815 515
rect 9851 481 9885 515
rect 9921 481 9955 515
rect 9991 481 10025 515
rect 10061 481 10095 515
rect 10131 481 10165 515
rect 10201 481 10235 515
rect 10271 481 10305 515
rect 10341 481 10375 515
rect 10411 481 10445 515
rect 10481 481 10515 515
rect 10551 481 10585 515
rect 10621 481 10655 515
rect 10691 481 10725 515
rect 10761 481 10795 515
rect 10831 481 10865 515
rect 10901 481 10935 515
rect 10971 481 11005 515
rect 11041 481 11075 515
rect 11111 481 11145 515
rect 11181 481 11215 515
rect 11251 481 11285 515
rect 11321 481 11355 515
rect 11391 481 11425 515
rect 11460 481 11494 515
rect 11529 481 11563 515
rect 11598 481 11632 515
rect 9711 409 9745 443
rect 9781 409 9815 443
rect 9851 409 9885 443
rect 9921 409 9955 443
rect 9991 409 10025 443
rect 10061 409 10095 443
rect 10131 409 10165 443
rect 10201 409 10235 443
rect 10271 409 10305 443
rect 10341 409 10375 443
rect 10411 409 10445 443
rect 10481 409 10515 443
rect 10551 409 10585 443
rect 10621 409 10655 443
rect 10691 409 10725 443
rect 10761 409 10795 443
rect 10831 409 10865 443
rect 10901 409 10935 443
rect 10971 409 11005 443
rect 11041 409 11075 443
rect 11111 409 11145 443
rect 11181 409 11215 443
rect 11251 409 11285 443
rect 11321 409 11355 443
rect 11391 409 11425 443
rect 11460 409 11494 443
rect 11529 409 11563 443
rect 11598 409 11632 443
rect 14932 706 14966 740
rect 15000 706 15034 740
rect 15068 706 15102 740
rect 14465 661 14499 695
rect 14543 661 14577 695
rect 14621 661 14655 695
rect 14698 661 14732 695
rect 14775 661 14809 695
rect 14852 661 14886 695
rect 14932 634 14966 668
rect 15000 634 15034 668
rect 15068 634 15102 668
rect 14465 575 14499 609
rect 14543 575 14577 609
rect 14621 575 14655 609
rect 14698 575 14732 609
rect 14775 575 14809 609
rect 14852 575 14886 609
rect 14932 562 14966 596
rect 15000 562 15034 596
rect 15068 562 15102 596
rect 14465 489 14499 523
rect 14543 489 14577 523
rect 14621 489 14655 523
rect 14698 489 14732 523
rect 14775 489 14809 523
rect 14852 489 14886 523
rect 14932 490 14966 524
rect 15000 490 15034 524
rect 15068 490 15102 524
rect 14465 403 14499 437
rect 14543 403 14577 437
rect 14621 403 14655 437
rect 14698 403 14732 437
rect 14775 403 14809 437
rect 14852 403 14886 437
rect 14932 418 14966 452
rect 15000 418 15034 452
rect 15068 418 15102 452
rect 7056 333 7090 367
rect 7125 333 7159 367
rect 7194 333 7228 367
rect 7263 333 7297 367
rect 7332 333 7366 367
rect 7401 333 7435 367
rect 7470 333 7504 367
rect 7539 333 7573 367
rect 7608 333 7642 367
rect 7677 333 7711 367
rect 7746 333 7780 367
rect 7815 333 7849 367
rect 7884 333 7918 367
rect 7953 333 7987 367
rect 8022 333 8056 367
rect 8091 333 8125 367
rect 8160 333 8194 367
rect 8229 333 8263 367
rect 8298 333 8332 367
rect 8367 333 8401 367
rect 8436 333 8470 367
rect 8505 333 8539 367
rect 8574 333 8608 367
rect 8643 333 8677 367
rect 8712 333 8746 367
rect 8781 333 8815 367
rect 8850 333 8884 367
rect 8919 333 8953 367
rect 8988 333 9022 367
rect 9057 333 9091 367
rect 9126 333 9160 367
rect 9195 333 9229 367
rect 9264 333 9298 367
rect 9333 333 9367 367
rect 9402 333 9436 367
rect 9471 333 9505 367
rect 9540 333 9574 367
rect 9609 333 9643 367
rect 9678 333 9712 367
rect 9747 333 9781 367
rect 9816 333 9850 367
rect 9885 333 9919 367
rect 9954 333 9988 367
rect 10023 333 10057 367
rect 10092 333 10126 367
rect 10161 333 10195 367
rect 10230 333 10264 367
rect 10299 333 10333 367
rect 10368 333 10402 367
rect 10437 333 10471 367
rect 10506 333 10540 367
rect 10575 333 10609 367
rect 10643 333 10677 367
rect 10711 333 10745 367
rect 10779 333 10813 367
rect 10847 333 10881 367
rect 10915 333 10949 367
rect 10983 333 11017 367
rect 11051 333 11085 367
rect 11119 333 11153 367
rect 11187 333 11221 367
rect 11255 333 11289 367
rect 11323 333 11357 367
rect 11391 333 11425 367
rect 11459 333 11493 367
rect 11527 333 11561 367
rect 11595 333 11629 367
rect 11663 333 11697 367
rect 11731 333 11765 367
rect 11799 333 11833 367
rect 11867 333 11901 367
rect 11935 333 11969 367
rect 12003 333 12037 367
rect 12071 333 12105 367
rect 12139 333 12173 367
rect 12207 333 12241 367
rect 12275 333 12309 367
rect 12343 333 12377 367
rect 12411 333 12445 367
rect 12479 333 12513 367
rect 12547 333 12581 367
rect 12615 333 12649 367
rect 12683 333 12717 367
rect 12751 333 12785 367
rect 12819 333 12853 367
rect 12887 333 12921 367
rect 12955 333 12989 367
rect 13023 333 13057 367
rect 13091 333 13125 367
rect 13159 333 13193 367
rect 13227 333 13261 367
rect 13295 333 13329 367
rect 13363 333 13397 367
rect 13431 333 13465 367
rect 13499 333 13533 367
rect 13567 333 13601 367
rect 13635 333 13669 367
rect 13703 333 13737 367
rect 13771 333 13805 367
rect 13839 333 13873 367
rect 13907 333 13941 367
rect 13975 333 14009 367
rect 14043 333 14077 367
rect 14111 333 14145 367
rect 14179 333 14213 367
rect 14247 333 14281 367
rect 14315 333 14349 367
rect 14383 333 14417 367
rect 14451 333 14485 367
rect 14519 333 14553 367
rect 14587 333 14621 367
rect 14655 333 14689 367
rect 14723 333 14757 367
rect 14791 333 14825 367
rect 14859 333 14893 367
rect 14932 346 14966 380
rect 15000 346 15034 380
rect 15068 346 15102 380
rect 7056 255 7090 289
rect 7125 255 7159 289
rect 7194 255 7228 289
rect 7263 255 7297 289
rect 7332 255 7366 289
rect 7401 255 7435 289
rect 7470 255 7504 289
rect 7539 255 7573 289
rect 7608 255 7642 289
rect 7677 255 7711 289
rect 7746 255 7780 289
rect 7815 255 7849 289
rect 7884 255 7918 289
rect 7953 255 7987 289
rect 8022 255 8056 289
rect 8091 255 8125 289
rect 8160 255 8194 289
rect 8229 255 8263 289
rect 8298 255 8332 289
rect 8367 255 8401 289
rect 8436 255 8470 289
rect 8505 255 8539 289
rect 8574 255 8608 289
rect 8643 255 8677 289
rect 8712 255 8746 289
rect 8781 255 8815 289
rect 8850 255 8884 289
rect 8919 255 8953 289
rect 8988 255 9022 289
rect 9057 255 9091 289
rect 9126 255 9160 289
rect 9195 255 9229 289
rect 9264 255 9298 289
rect 9333 255 9367 289
rect 9402 255 9436 289
rect 9471 255 9505 289
rect 9540 255 9574 289
rect 9609 255 9643 289
rect 9678 255 9712 289
rect 9747 255 9781 289
rect 9816 255 9850 289
rect 9885 255 9919 289
rect 9954 255 9988 289
rect 10023 255 10057 289
rect 10092 255 10126 289
rect 10161 255 10195 289
rect 10230 255 10264 289
rect 10299 255 10333 289
rect 10368 255 10402 289
rect 10437 255 10471 289
rect 10506 255 10540 289
rect 10575 255 10609 289
rect 10643 255 10677 289
rect 10711 255 10745 289
rect 10779 255 10813 289
rect 10847 255 10881 289
rect 10915 255 10949 289
rect 10983 255 11017 289
rect 11051 255 11085 289
rect 11119 255 11153 289
rect 11187 255 11221 289
rect 11255 255 11289 289
rect 11323 255 11357 289
rect 11391 255 11425 289
rect 11459 255 11493 289
rect 11527 255 11561 289
rect 11595 255 11629 289
rect 11663 255 11697 289
rect 11731 255 11765 289
rect 11799 255 11833 289
rect 11867 255 11901 289
rect 11935 255 11969 289
rect 12003 255 12037 289
rect 12071 255 12105 289
rect 12139 255 12173 289
rect 12207 255 12241 289
rect 12275 255 12309 289
rect 12343 255 12377 289
rect 12411 255 12445 289
rect 12479 255 12513 289
rect 12547 255 12581 289
rect 12615 255 12649 289
rect 12683 255 12717 289
rect 12751 255 12785 289
rect 12819 255 12853 289
rect 12887 255 12921 289
rect 12955 255 12989 289
rect 13023 255 13057 289
rect 13091 255 13125 289
rect 13159 255 13193 289
rect 13227 255 13261 289
rect 13295 255 13329 289
rect 13363 255 13397 289
rect 13431 255 13465 289
rect 13499 255 13533 289
rect 13567 255 13601 289
rect 13635 255 13669 289
rect 13703 255 13737 289
rect 13771 255 13805 289
rect 13839 255 13873 289
rect 13907 255 13941 289
rect 13975 255 14009 289
rect 14043 255 14077 289
rect 14111 255 14145 289
rect 14179 255 14213 289
rect 14247 255 14281 289
rect 14315 255 14349 289
rect 14383 255 14417 289
rect 14451 255 14485 289
rect 14519 255 14553 289
rect 14587 255 14621 289
rect 14655 255 14689 289
rect 14723 255 14757 289
rect 14791 255 14825 289
rect 14859 255 14893 289
rect 14932 274 14966 308
rect 15000 274 15034 308
rect 15068 274 15102 308
rect 7056 177 7090 211
rect 7125 177 7159 211
rect 7194 177 7228 211
rect 7263 177 7297 211
rect 7332 177 7366 211
rect 7401 177 7435 211
rect 7470 177 7504 211
rect 7539 177 7573 211
rect 7608 177 7642 211
rect 7677 177 7711 211
rect 7746 177 7780 211
rect 7815 177 7849 211
rect 7884 177 7918 211
rect 7953 177 7987 211
rect 8022 177 8056 211
rect 8091 177 8125 211
rect 8160 177 8194 211
rect 8229 177 8263 211
rect 8298 177 8332 211
rect 8367 177 8401 211
rect 8436 177 8470 211
rect 8505 177 8539 211
rect 8574 177 8608 211
rect 8643 177 8677 211
rect 8712 177 8746 211
rect 8781 177 8815 211
rect 8850 177 8884 211
rect 8919 177 8953 211
rect 8988 177 9022 211
rect 9057 177 9091 211
rect 9126 177 9160 211
rect 9195 177 9229 211
rect 9264 177 9298 211
rect 9333 177 9367 211
rect 9402 177 9436 211
rect 9471 177 9505 211
rect 9540 177 9574 211
rect 9609 177 9643 211
rect 9678 177 9712 211
rect 9747 177 9781 211
rect 9816 177 9850 211
rect 9885 177 9919 211
rect 9954 177 9988 211
rect 10023 177 10057 211
rect 10092 177 10126 211
rect 10161 177 10195 211
rect 10230 177 10264 211
rect 10299 177 10333 211
rect 10368 177 10402 211
rect 10437 177 10471 211
rect 10506 177 10540 211
rect 10575 177 10609 211
rect 10643 177 10677 211
rect 10711 177 10745 211
rect 10779 177 10813 211
rect 10847 177 10881 211
rect 10915 177 10949 211
rect 10983 177 11017 211
rect 11051 177 11085 211
rect 11119 177 11153 211
rect 11187 177 11221 211
rect 11255 177 11289 211
rect 11323 177 11357 211
rect 11391 177 11425 211
rect 11459 177 11493 211
rect 11527 177 11561 211
rect 11595 177 11629 211
rect 11663 177 11697 211
rect 11731 177 11765 211
rect 11799 177 11833 211
rect 11867 177 11901 211
rect 11935 177 11969 211
rect 12003 177 12037 211
rect 12071 177 12105 211
rect 12139 177 12173 211
rect 12207 177 12241 211
rect 12275 177 12309 211
rect 12343 177 12377 211
rect 12411 177 12445 211
rect 12479 177 12513 211
rect 12547 177 12581 211
rect 12615 177 12649 211
rect 12683 177 12717 211
rect 12751 177 12785 211
rect 12819 177 12853 211
rect 12887 177 12921 211
rect 12955 177 12989 211
rect 13023 177 13057 211
rect 13091 177 13125 211
rect 13159 177 13193 211
rect 13227 177 13261 211
rect 13295 177 13329 211
rect 13363 177 13397 211
rect 13431 177 13465 211
rect 13499 177 13533 211
rect 13567 177 13601 211
rect 13635 177 13669 211
rect 13703 177 13737 211
rect 13771 177 13805 211
rect 13839 177 13873 211
rect 13907 177 13941 211
rect 13975 177 14009 211
rect 14043 177 14077 211
rect 14111 177 14145 211
rect 14179 177 14213 211
rect 14247 177 14281 211
rect 14315 177 14349 211
rect 14383 177 14417 211
rect 14451 177 14485 211
rect 14519 177 14553 211
rect 14587 177 14621 211
rect 14655 177 14689 211
rect 14723 177 14757 211
rect 14791 177 14825 211
rect 14859 177 14893 211
rect 14932 202 14966 236
rect 15000 202 15034 236
rect 15068 202 15102 236
rect 7056 99 7090 133
rect 7125 99 7159 133
rect 7194 99 7228 133
rect 7263 99 7297 133
rect 7332 99 7366 133
rect 7401 99 7435 133
rect 7470 99 7504 133
rect 7539 99 7573 133
rect 7608 99 7642 133
rect 7677 99 7711 133
rect 7746 99 7780 133
rect 7815 99 7849 133
rect 7884 99 7918 133
rect 7953 99 7987 133
rect 8022 99 8056 133
rect 8091 99 8125 133
rect 8160 99 8194 133
rect 8229 99 8263 133
rect 8298 99 8332 133
rect 8367 99 8401 133
rect 8436 99 8470 133
rect 8505 99 8539 133
rect 8574 99 8608 133
rect 8643 99 8677 133
rect 8712 99 8746 133
rect 8781 99 8815 133
rect 8850 99 8884 133
rect 8919 99 8953 133
rect 8988 99 9022 133
rect 9057 99 9091 133
rect 9126 99 9160 133
rect 9195 99 9229 133
rect 9264 99 9298 133
rect 9333 99 9367 133
rect 9402 99 9436 133
rect 9471 99 9505 133
rect 9540 99 9574 133
rect 9609 99 9643 133
rect 9678 99 9712 133
rect 9747 99 9781 133
rect 9816 99 9850 133
rect 9885 99 9919 133
rect 9954 99 9988 133
rect 10023 99 10057 133
rect 10092 99 10126 133
rect 10161 99 10195 133
rect 10230 99 10264 133
rect 10299 99 10333 133
rect 10368 99 10402 133
rect 10437 99 10471 133
rect 10506 99 10540 133
rect 10575 99 10609 133
rect 10643 99 10677 133
rect 10711 99 10745 133
rect 10779 99 10813 133
rect 10847 99 10881 133
rect 10915 99 10949 133
rect 10983 99 11017 133
rect 11051 99 11085 133
rect 11119 99 11153 133
rect 11187 99 11221 133
rect 11255 99 11289 133
rect 11323 99 11357 133
rect 11391 99 11425 133
rect 11459 99 11493 133
rect 11527 99 11561 133
rect 11595 99 11629 133
rect 11663 99 11697 133
rect 11731 99 11765 133
rect 11799 99 11833 133
rect 11867 99 11901 133
rect 11935 99 11969 133
rect 12003 99 12037 133
rect 12071 99 12105 133
rect 12139 99 12173 133
rect 12207 99 12241 133
rect 12275 99 12309 133
rect 12343 99 12377 133
rect 12411 99 12445 133
rect 12479 99 12513 133
rect 12547 99 12581 133
rect 12615 99 12649 133
rect 12683 99 12717 133
rect 12751 99 12785 133
rect 12819 99 12853 133
rect 12887 99 12921 133
rect 12955 99 12989 133
rect 13023 99 13057 133
rect 13091 99 13125 133
rect 13159 99 13193 133
rect 13227 99 13261 133
rect 13295 99 13329 133
rect 13363 99 13397 133
rect 13431 99 13465 133
rect 13499 99 13533 133
rect 13567 99 13601 133
rect 13635 99 13669 133
rect 13703 99 13737 133
rect 13771 99 13805 133
rect 13839 99 13873 133
rect 13907 99 13941 133
rect 13975 99 14009 133
rect 14043 99 14077 133
rect 14111 99 14145 133
rect 14179 99 14213 133
rect 14247 99 14281 133
rect 14315 99 14349 133
rect 14383 99 14417 133
rect 14451 99 14485 133
rect 14519 99 14553 133
rect 14587 99 14621 133
rect 14655 99 14689 133
rect 14723 99 14757 133
rect 14791 99 14825 133
rect 14859 99 14893 133
rect 14932 130 14966 164
rect 15000 130 15034 164
rect 15068 130 15102 164
rect 14932 57 14966 91
rect 15000 57 15034 91
rect 15068 57 15102 91
rect 7056 21 7090 55
rect 7125 21 7159 55
rect 7194 21 7228 55
rect 7263 21 7297 55
rect 7332 21 7366 55
rect 7401 21 7435 55
rect 7470 21 7504 55
rect 7539 21 7573 55
rect 7608 21 7642 55
rect 7677 21 7711 55
rect 7746 21 7780 55
rect 7815 21 7849 55
rect 7884 21 7918 55
rect 7953 21 7987 55
rect 8022 21 8056 55
rect 8091 21 8125 55
rect 8160 21 8194 55
rect 8229 21 8263 55
rect 8298 21 8332 55
rect 8367 21 8401 55
rect 8436 21 8470 55
rect 8505 21 8539 55
rect 8574 21 8608 55
rect 8643 21 8677 55
rect 8712 21 8746 55
rect 8781 21 8815 55
rect 8850 21 8884 55
rect 8919 21 8953 55
rect 8988 21 9022 55
rect 9057 21 9091 55
rect 9126 21 9160 55
rect 9195 21 9229 55
rect 9264 21 9298 55
rect 9333 21 9367 55
rect 9402 21 9436 55
rect 9471 21 9505 55
rect 9540 21 9574 55
rect 9609 21 9643 55
rect 9678 21 9712 55
rect 9747 21 9781 55
rect 9816 21 9850 55
rect 9885 21 9919 55
rect 9954 21 9988 55
rect 10023 21 10057 55
rect 10092 21 10126 55
rect 10161 21 10195 55
rect 10230 21 10264 55
rect 10299 21 10333 55
rect 10368 21 10402 55
rect 10437 21 10471 55
rect 10506 21 10540 55
rect 10575 21 10609 55
rect 10643 21 10677 55
rect 10711 21 10745 55
rect 10779 21 10813 55
rect 10847 21 10881 55
rect 10915 21 10949 55
rect 10983 21 11017 55
rect 11051 21 11085 55
rect 11119 21 11153 55
rect 11187 21 11221 55
rect 11255 21 11289 55
rect 11323 21 11357 55
rect 11391 21 11425 55
rect 11459 21 11493 55
rect 11527 21 11561 55
rect 11595 21 11629 55
rect 11663 21 11697 55
rect 11731 21 11765 55
rect 11799 21 11833 55
rect 11867 21 11901 55
rect 11935 21 11969 55
rect 12003 21 12037 55
rect 12071 21 12105 55
rect 12139 21 12173 55
rect 12207 21 12241 55
rect 12275 21 12309 55
rect 12343 21 12377 55
rect 12411 21 12445 55
rect 12479 21 12513 55
rect 12547 21 12581 55
rect 12615 21 12649 55
rect 12683 21 12717 55
rect 12751 21 12785 55
rect 12819 21 12853 55
rect 12887 21 12921 55
rect 12955 21 12989 55
rect 13023 21 13057 55
rect 13091 21 13125 55
rect 13159 21 13193 55
rect 13227 21 13261 55
rect 13295 21 13329 55
rect 13363 21 13397 55
rect 13431 21 13465 55
rect 13499 21 13533 55
rect 13567 21 13601 55
rect 13635 21 13669 55
rect 13703 21 13737 55
rect 13771 21 13805 55
rect 13839 21 13873 55
rect 13907 21 13941 55
rect 13975 21 14009 55
rect 14043 21 14077 55
rect 14111 21 14145 55
rect 14179 21 14213 55
rect 14247 21 14281 55
rect 14315 21 14349 55
rect 14383 21 14417 55
rect 14451 21 14485 55
rect 14519 21 14553 55
rect 14587 21 14621 55
rect 14655 21 14689 55
rect 14723 21 14757 55
rect 14791 21 14825 55
rect 14859 21 14893 55
<< mvnsubdiffcont >>
rect 12660 15617 12694 15651
rect 12730 15617 12764 15651
rect 12800 15617 12834 15651
rect 12869 15617 12903 15651
rect 12938 15617 12972 15651
rect 13007 15617 13041 15651
rect 13076 15617 13110 15651
rect 13145 15617 13179 15651
rect 13214 15617 13248 15651
rect 13283 15617 13317 15651
rect 13352 15617 13386 15651
rect 13421 15617 13455 15651
rect 13490 15617 13524 15651
rect 13559 15617 13593 15651
rect 13628 15617 13662 15651
rect 13697 15617 13731 15651
rect 13766 15617 13800 15651
rect 13835 15617 13869 15651
rect 13904 15617 13938 15651
rect 13973 15617 14007 15651
rect 14042 15617 14076 15651
rect 14111 15617 14145 15651
rect 14180 15617 14214 15651
rect 14249 15617 14283 15651
rect 14318 15617 14352 15651
rect 12660 15547 12694 15581
rect 12730 15547 12764 15581
rect 12800 15547 12834 15581
rect 12869 15547 12903 15581
rect 12938 15547 12972 15581
rect 13007 15547 13041 15581
rect 13076 15547 13110 15581
rect 13145 15547 13179 15581
rect 13214 15547 13248 15581
rect 13283 15547 13317 15581
rect 13352 15547 13386 15581
rect 13421 15547 13455 15581
rect 13490 15547 13524 15581
rect 13559 15547 13593 15581
rect 13628 15547 13662 15581
rect 13697 15547 13731 15581
rect 13766 15547 13800 15581
rect 13835 15547 13869 15581
rect 13904 15547 13938 15581
rect 13973 15547 14007 15581
rect 14042 15547 14076 15581
rect 14111 15547 14145 15581
rect 14180 15547 14214 15581
rect 14249 15547 14283 15581
rect 14318 15547 14352 15581
rect 12660 15477 12694 15511
rect 12730 15477 12764 15511
rect 12800 15477 12834 15511
rect 12869 15477 12903 15511
rect 12938 15477 12972 15511
rect 13007 15477 13041 15511
rect 13076 15477 13110 15511
rect 13145 15477 13179 15511
rect 13214 15477 13248 15511
rect 13283 15477 13317 15511
rect 13352 15477 13386 15511
rect 13421 15477 13455 15511
rect 13490 15477 13524 15511
rect 13559 15477 13593 15511
rect 13628 15477 13662 15511
rect 13697 15477 13731 15511
rect 13766 15477 13800 15511
rect 13835 15477 13869 15511
rect 13904 15477 13938 15511
rect 13973 15477 14007 15511
rect 14042 15477 14076 15511
rect 14111 15477 14145 15511
rect 14180 15477 14214 15511
rect 14249 15477 14283 15511
rect 14318 15477 14352 15511
rect 12660 15407 12694 15441
rect 12730 15407 12764 15441
rect 12800 15407 12834 15441
rect 12869 15407 12903 15441
rect 12938 15407 12972 15441
rect 13007 15407 13041 15441
rect 13076 15407 13110 15441
rect 13145 15407 13179 15441
rect 13214 15407 13248 15441
rect 13283 15407 13317 15441
rect 13352 15407 13386 15441
rect 13421 15407 13455 15441
rect 13490 15407 13524 15441
rect 13559 15407 13593 15441
rect 13628 15407 13662 15441
rect 13697 15407 13731 15441
rect 13766 15407 13800 15441
rect 13835 15407 13869 15441
rect 13904 15407 13938 15441
rect 13973 15407 14007 15441
rect 14042 15407 14076 15441
rect 14111 15407 14145 15441
rect 14180 15407 14214 15441
rect 14249 15407 14283 15441
rect 14318 15407 14352 15441
rect 12660 15337 12694 15371
rect 12730 15337 12764 15371
rect 12800 15337 12834 15371
rect 12869 15337 12903 15371
rect 12938 15337 12972 15371
rect 13007 15337 13041 15371
rect 13076 15337 13110 15371
rect 13145 15337 13179 15371
rect 13214 15337 13248 15371
rect 13283 15337 13317 15371
rect 13352 15337 13386 15371
rect 13421 15337 13455 15371
rect 13490 15337 13524 15371
rect 13559 15337 13593 15371
rect 13628 15337 13662 15371
rect 13697 15337 13731 15371
rect 13766 15337 13800 15371
rect 13835 15337 13869 15371
rect 13904 15337 13938 15371
rect 13973 15337 14007 15371
rect 14042 15337 14076 15371
rect 14111 15337 14145 15371
rect 14180 15337 14214 15371
rect 14249 15337 14283 15371
rect 14318 15337 14352 15371
rect 12660 15267 12694 15301
rect 12730 15267 12764 15301
rect 12800 15267 12834 15301
rect 12869 15267 12903 15301
rect 12938 15267 12972 15301
rect 13007 15267 13041 15301
rect 13076 15267 13110 15301
rect 13145 15267 13179 15301
rect 13214 15267 13248 15301
rect 13283 15267 13317 15301
rect 13352 15267 13386 15301
rect 13421 15267 13455 15301
rect 13490 15267 13524 15301
rect 13559 15267 13593 15301
rect 13628 15267 13662 15301
rect 13697 15267 13731 15301
rect 13766 15267 13800 15301
rect 13835 15267 13869 15301
rect 13904 15267 13938 15301
rect 13973 15267 14007 15301
rect 14042 15267 14076 15301
rect 14111 15267 14145 15301
rect 14180 15267 14214 15301
rect 14249 15267 14283 15301
rect 14318 15267 14352 15301
rect 12660 15197 12694 15231
rect 12730 15197 12764 15231
rect 12800 15197 12834 15231
rect 12869 15197 12903 15231
rect 12938 15197 12972 15231
rect 13007 15197 13041 15231
rect 13076 15197 13110 15231
rect 13145 15197 13179 15231
rect 13214 15197 13248 15231
rect 13283 15197 13317 15231
rect 13352 15197 13386 15231
rect 13421 15197 13455 15231
rect 13490 15197 13524 15231
rect 13559 15197 13593 15231
rect 13628 15197 13662 15231
rect 13697 15197 13731 15231
rect 13766 15197 13800 15231
rect 13835 15197 13869 15231
rect 13904 15197 13938 15231
rect 13973 15197 14007 15231
rect 14042 15197 14076 15231
rect 14111 15197 14145 15231
rect 14180 15197 14214 15231
rect 14249 15197 14283 15231
rect 14318 15197 14352 15231
rect 12660 15127 12694 15161
rect 12730 15127 12764 15161
rect 12800 15127 12834 15161
rect 12869 15127 12903 15161
rect 12938 15127 12972 15161
rect 13007 15127 13041 15161
rect 13076 15127 13110 15161
rect 13145 15127 13179 15161
rect 13214 15127 13248 15161
rect 13283 15127 13317 15161
rect 13352 15127 13386 15161
rect 13421 15127 13455 15161
rect 13490 15127 13524 15161
rect 13559 15127 13593 15161
rect 13628 15127 13662 15161
rect 13697 15127 13731 15161
rect 13766 15127 13800 15161
rect 13835 15127 13869 15161
rect 13904 15127 13938 15161
rect 13973 15127 14007 15161
rect 14042 15127 14076 15161
rect 14111 15127 14145 15161
rect 14180 15127 14214 15161
rect 14249 15127 14283 15161
rect 14318 15127 14352 15161
rect 12660 15057 12694 15091
rect 12730 15057 12764 15091
rect 12800 15057 12834 15091
rect 12869 15057 12903 15091
rect 12938 15057 12972 15091
rect 13007 15057 13041 15091
rect 13076 15057 13110 15091
rect 13145 15057 13179 15091
rect 13214 15057 13248 15091
rect 13283 15057 13317 15091
rect 13352 15057 13386 15091
rect 13421 15057 13455 15091
rect 13490 15057 13524 15091
rect 13559 15057 13593 15091
rect 13628 15057 13662 15091
rect 13697 15057 13731 15091
rect 13766 15057 13800 15091
rect 13835 15057 13869 15091
rect 13904 15057 13938 15091
rect 13973 15057 14007 15091
rect 14042 15057 14076 15091
rect 14111 15057 14145 15091
rect 14180 15057 14214 15091
rect 14249 15057 14283 15091
rect 14318 15057 14352 15091
rect 12660 14987 12694 15021
rect 12730 14987 12764 15021
rect 12800 14987 12834 15021
rect 12869 14987 12903 15021
rect 12938 14987 12972 15021
rect 13007 14987 13041 15021
rect 13076 14987 13110 15021
rect 13145 14987 13179 15021
rect 13214 14987 13248 15021
rect 13283 14987 13317 15021
rect 13352 14987 13386 15021
rect 13421 14987 13455 15021
rect 13490 14987 13524 15021
rect 13559 14987 13593 15021
rect 13628 14987 13662 15021
rect 13697 14987 13731 15021
rect 13766 14987 13800 15021
rect 13835 14987 13869 15021
rect 13904 14987 13938 15021
rect 13973 14987 14007 15021
rect 14042 14987 14076 15021
rect 14111 14987 14145 15021
rect 14180 14987 14214 15021
rect 14249 14987 14283 15021
rect 14318 14987 14352 15021
rect 12660 14917 12694 14951
rect 12730 14917 12764 14951
rect 12800 14917 12834 14951
rect 12869 14917 12903 14951
rect 12938 14917 12972 14951
rect 13007 14917 13041 14951
rect 13076 14917 13110 14951
rect 13145 14917 13179 14951
rect 13214 14917 13248 14951
rect 13283 14917 13317 14951
rect 13352 14917 13386 14951
rect 13421 14917 13455 14951
rect 13490 14917 13524 14951
rect 13559 14917 13593 14951
rect 13628 14917 13662 14951
rect 13697 14917 13731 14951
rect 13766 14917 13800 14951
rect 13835 14917 13869 14951
rect 13904 14917 13938 14951
rect 13973 14917 14007 14951
rect 14042 14917 14076 14951
rect 14111 14917 14145 14951
rect 14180 14917 14214 14951
rect 14249 14917 14283 14951
rect 14318 14917 14352 14951
rect 12660 14847 12694 14881
rect 12730 14847 12764 14881
rect 12800 14847 12834 14881
rect 12869 14847 12903 14881
rect 12938 14847 12972 14881
rect 13007 14847 13041 14881
rect 13076 14847 13110 14881
rect 13145 14847 13179 14881
rect 13214 14847 13248 14881
rect 13283 14847 13317 14881
rect 13352 14847 13386 14881
rect 13421 14847 13455 14881
rect 13490 14847 13524 14881
rect 13559 14847 13593 14881
rect 13628 14847 13662 14881
rect 13697 14847 13731 14881
rect 13766 14847 13800 14881
rect 13835 14847 13869 14881
rect 13904 14847 13938 14881
rect 13973 14847 14007 14881
rect 14042 14847 14076 14881
rect 14111 14847 14145 14881
rect 14180 14847 14214 14881
rect 14249 14847 14283 14881
rect 14318 14847 14352 14881
rect 68 8740 102 8774
rect 138 8740 172 8774
rect 208 8740 242 8774
rect 278 8740 312 8774
rect 348 8740 382 8774
rect 418 8740 452 8774
rect 488 8740 522 8774
rect 558 8740 592 8774
rect 628 8740 662 8774
rect 698 8740 732 8774
rect 768 8740 802 8774
rect 838 8740 872 8774
rect 908 8740 942 8774
rect 978 8740 1012 8774
rect 1048 8740 1082 8774
rect 1118 8740 1152 8774
rect 1188 8740 1222 8774
rect 1258 8740 1292 8774
rect 1328 8740 1362 8774
rect 1398 8740 1432 8774
rect 1467 8740 1501 8774
rect 1536 8740 1570 8774
rect 1605 8740 1639 8774
rect 1674 8740 1708 8774
rect 1743 8740 1777 8774
rect 1812 8740 1846 8774
rect 1881 8740 1915 8774
rect 1950 8740 1984 8774
rect 2019 8740 2053 8774
rect 2088 8740 2122 8774
rect 2157 8740 2191 8774
rect 2226 8740 2260 8774
rect 2295 8740 2329 8774
rect 2364 8740 2398 8774
rect 2433 8740 2467 8774
rect 2502 8740 2536 8774
rect 2571 8740 2605 8774
rect 2640 8740 2674 8774
rect 2709 8740 2743 8774
rect 2778 8740 2812 8774
rect 2847 8740 2881 8774
rect 2933 8736 2967 8770
rect 3002 8736 3036 8770
rect 3071 8736 3105 8770
rect 3139 8736 3173 8770
rect 3207 8736 3241 8770
rect 3275 8736 3309 8770
rect 3343 8736 3377 8770
rect 3411 8736 3445 8770
rect 3479 8736 3513 8770
rect 3547 8736 3581 8770
rect 3615 8736 3649 8770
rect 3683 8736 3717 8770
rect 3751 8736 3785 8770
rect 3819 8736 3853 8770
rect 3887 8736 3921 8770
rect 3955 8736 3989 8770
rect 4023 8736 4057 8770
rect 4091 8736 4125 8770
rect 4159 8736 4193 8770
rect 4227 8736 4261 8770
rect 4295 8736 4329 8770
rect 4363 8736 4397 8770
rect 4431 8736 4465 8770
rect 4499 8736 4533 8770
rect 4567 8736 4601 8770
rect 4635 8736 4669 8770
rect 4703 8736 4737 8770
rect 4771 8736 4805 8770
rect 4839 8736 4873 8770
rect 4907 8736 4941 8770
rect 4975 8736 5009 8770
rect 5043 8736 5077 8770
rect 5111 8736 5145 8770
rect 5179 8736 5213 8770
rect 5247 8736 5281 8770
rect 5315 8736 5349 8770
rect 5383 8736 5417 8770
rect 5451 8736 5485 8770
rect 5519 8736 5553 8770
rect 5587 8736 5621 8770
rect 5655 8736 5689 8770
rect 5723 8736 5757 8770
rect 5791 8736 5825 8770
rect 5859 8736 5893 8770
rect 5927 8736 5961 8770
rect 5995 8736 6029 8770
rect 6063 8736 6097 8770
rect 6131 8736 6165 8770
rect 6199 8736 6233 8770
rect 6267 8736 6301 8770
rect 6335 8736 6369 8770
rect 6403 8736 6437 8770
rect 6471 8736 6505 8770
rect 6539 8736 6573 8770
rect 6607 8736 6641 8770
rect 6675 8736 6709 8770
rect 6743 8736 6777 8770
rect 6811 8736 6845 8770
rect 6879 8736 6913 8770
rect 6947 8736 6981 8770
rect 7015 8736 7049 8770
rect 7083 8736 7117 8770
rect 7151 8736 7185 8770
rect 7219 8736 7253 8770
rect 7287 8736 7321 8770
rect 7355 8736 7389 8770
rect 7423 8736 7457 8770
rect 7491 8736 7525 8770
rect 7559 8736 7593 8770
rect 7627 8736 7661 8770
rect 7695 8736 7729 8770
rect 7763 8736 7797 8770
rect 7831 8736 7865 8770
rect 7899 8736 7933 8770
rect 7967 8736 8001 8770
rect 8035 8736 8069 8770
rect 8103 8736 8137 8770
rect 8171 8736 8205 8770
rect 8239 8736 8273 8770
rect 8307 8736 8341 8770
rect 8393 8739 8427 8773
rect 8462 8739 8496 8773
rect 8531 8739 8565 8773
rect 8600 8739 8634 8773
rect 8669 8739 8703 8773
rect 8738 8739 8772 8773
rect 8807 8739 8841 8773
rect 8876 8739 8910 8773
rect 8945 8739 8979 8773
rect 9014 8739 9048 8773
rect 9083 8739 9117 8773
rect 9152 8739 9186 8773
rect 9220 8739 9254 8773
rect 9288 8739 9322 8773
rect 9356 8739 9390 8773
rect 9424 8739 9458 8773
rect 9492 8739 9526 8773
rect 9560 8739 9594 8773
rect 9628 8739 9662 8773
rect 9696 8739 9730 8773
rect 9764 8739 9798 8773
rect 9832 8739 9866 8773
rect 9900 8739 9934 8773
rect 9968 8739 10002 8773
rect 10036 8739 10070 8773
rect 10104 8739 10138 8773
rect 10172 8739 10206 8773
rect 10240 8739 10274 8773
rect 10308 8739 10342 8773
rect 10376 8739 10410 8773
rect 10444 8739 10478 8773
rect 10512 8739 10546 8773
rect 10580 8739 10614 8773
rect 10648 8739 10682 8773
rect 10716 8739 10750 8773
rect 10784 8739 10818 8773
rect 10852 8739 10886 8773
rect 10920 8739 10954 8773
rect 10988 8739 11022 8773
rect 11056 8739 11090 8773
rect 11124 8739 11158 8773
rect 11192 8739 11226 8773
rect 11260 8739 11294 8773
rect 11328 8739 11362 8773
rect 11396 8739 11430 8773
rect 11464 8739 11498 8773
rect 11532 8739 11566 8773
rect 11600 8739 11634 8773
rect 11668 8739 11702 8773
rect 11736 8739 11770 8773
rect 11804 8739 11838 8773
rect 11872 8739 11906 8773
rect 11940 8739 11974 8773
rect 12008 8739 12042 8773
rect 12076 8739 12110 8773
rect 12144 8739 12178 8773
rect 12212 8739 12246 8773
rect 12280 8739 12314 8773
rect 12348 8739 12382 8773
rect 12416 8739 12450 8773
rect 12484 8739 12518 8773
rect 12552 8739 12586 8773
rect 12620 8739 12654 8773
rect 12688 8739 12722 8773
rect 12756 8739 12790 8773
rect 12824 8739 12858 8773
rect 12892 8739 12926 8773
rect 12960 8739 12994 8773
rect 13028 8739 13062 8773
rect 13096 8739 13130 8773
rect 13164 8739 13198 8773
rect 13232 8739 13266 8773
rect 13300 8739 13334 8773
rect 13368 8739 13402 8773
rect 13436 8739 13470 8773
rect 13504 8739 13538 8773
rect 13572 8739 13606 8773
rect 13640 8739 13674 8773
rect 13708 8739 13742 8773
rect 13776 8739 13810 8773
rect 13844 8739 13878 8773
rect 13912 8739 13946 8773
rect 13980 8739 14014 8773
rect 14048 8739 14082 8773
rect 14116 8739 14150 8773
rect 14184 8739 14218 8773
rect 14252 8739 14286 8773
rect 14320 8739 14354 8773
rect 14388 8739 14422 8773
rect 14456 8739 14490 8773
rect 14524 8739 14558 8773
rect 14592 8739 14626 8773
rect 14660 8739 14694 8773
rect 14728 8739 14762 8773
rect 14796 8739 14830 8773
rect 14864 8739 14898 8773
rect 68 8666 102 8700
rect 138 8666 172 8700
rect 208 8666 242 8700
rect 278 8666 312 8700
rect 348 8666 382 8700
rect 418 8666 452 8700
rect 488 8666 522 8700
rect 558 8666 592 8700
rect 628 8666 662 8700
rect 698 8666 732 8700
rect 768 8666 802 8700
rect 838 8666 872 8700
rect 908 8666 942 8700
rect 978 8666 1012 8700
rect 1048 8666 1082 8700
rect 1118 8666 1152 8700
rect 1188 8666 1222 8700
rect 1258 8666 1292 8700
rect 1328 8666 1362 8700
rect 1398 8666 1432 8700
rect 1467 8666 1501 8700
rect 1536 8666 1570 8700
rect 1605 8666 1639 8700
rect 1674 8666 1708 8700
rect 1743 8666 1777 8700
rect 1812 8666 1846 8700
rect 1881 8666 1915 8700
rect 1950 8666 1984 8700
rect 2019 8666 2053 8700
rect 2088 8666 2122 8700
rect 2157 8666 2191 8700
rect 2226 8666 2260 8700
rect 2295 8666 2329 8700
rect 2364 8666 2398 8700
rect 2433 8666 2467 8700
rect 2502 8666 2536 8700
rect 2571 8666 2605 8700
rect 2640 8666 2674 8700
rect 2709 8666 2743 8700
rect 2778 8666 2812 8700
rect 2847 8666 2881 8700
rect 2933 8666 2967 8700
rect 3002 8666 3036 8700
rect 3071 8666 3105 8700
rect 3139 8666 3173 8700
rect 3207 8666 3241 8700
rect 3275 8666 3309 8700
rect 3343 8666 3377 8700
rect 3411 8666 3445 8700
rect 3479 8666 3513 8700
rect 3547 8666 3581 8700
rect 3615 8666 3649 8700
rect 3683 8666 3717 8700
rect 3751 8666 3785 8700
rect 3819 8666 3853 8700
rect 3887 8666 3921 8700
rect 3955 8666 3989 8700
rect 4023 8666 4057 8700
rect 4091 8666 4125 8700
rect 4159 8666 4193 8700
rect 4227 8666 4261 8700
rect 4295 8666 4329 8700
rect 4363 8666 4397 8700
rect 4431 8666 4465 8700
rect 4499 8666 4533 8700
rect 4567 8666 4601 8700
rect 4635 8666 4669 8700
rect 4703 8666 4737 8700
rect 4771 8666 4805 8700
rect 4839 8666 4873 8700
rect 4907 8666 4941 8700
rect 4975 8666 5009 8700
rect 5043 8666 5077 8700
rect 5111 8666 5145 8700
rect 5179 8666 5213 8700
rect 5247 8666 5281 8700
rect 5315 8666 5349 8700
rect 5383 8666 5417 8700
rect 5451 8666 5485 8700
rect 5519 8666 5553 8700
rect 5587 8666 5621 8700
rect 5655 8666 5689 8700
rect 5723 8666 5757 8700
rect 5791 8666 5825 8700
rect 5859 8666 5893 8700
rect 5927 8666 5961 8700
rect 5995 8666 6029 8700
rect 6063 8666 6097 8700
rect 6131 8666 6165 8700
rect 6199 8666 6233 8700
rect 6267 8666 6301 8700
rect 6335 8666 6369 8700
rect 6403 8666 6437 8700
rect 6471 8666 6505 8700
rect 6539 8666 6573 8700
rect 6607 8666 6641 8700
rect 6675 8666 6709 8700
rect 6743 8666 6777 8700
rect 6811 8666 6845 8700
rect 6879 8666 6913 8700
rect 6947 8666 6981 8700
rect 7015 8666 7049 8700
rect 7083 8666 7117 8700
rect 7151 8666 7185 8700
rect 7219 8666 7253 8700
rect 7287 8666 7321 8700
rect 7355 8666 7389 8700
rect 7423 8666 7457 8700
rect 7491 8666 7525 8700
rect 7559 8666 7593 8700
rect 7627 8666 7661 8700
rect 7695 8666 7729 8700
rect 7763 8666 7797 8700
rect 7831 8666 7865 8700
rect 7899 8666 7933 8700
rect 7967 8666 8001 8700
rect 8035 8666 8069 8700
rect 8103 8666 8137 8700
rect 8171 8666 8205 8700
rect 8239 8666 8273 8700
rect 8307 8666 8341 8700
rect 8393 8659 8427 8693
rect 8462 8659 8496 8693
rect 8531 8659 8565 8693
rect 8600 8659 8634 8693
rect 8669 8659 8703 8693
rect 8738 8659 8772 8693
rect 8807 8659 8841 8693
rect 8876 8659 8910 8693
rect 8945 8659 8979 8693
rect 9014 8659 9048 8693
rect 9083 8659 9117 8693
rect 9152 8659 9186 8693
rect 9220 8659 9254 8693
rect 9288 8659 9322 8693
rect 9356 8659 9390 8693
rect 9424 8659 9458 8693
rect 9492 8659 9526 8693
rect 9560 8659 9594 8693
rect 9628 8659 9662 8693
rect 9696 8659 9730 8693
rect 9764 8659 9798 8693
rect 9832 8659 9866 8693
rect 9900 8659 9934 8693
rect 9968 8659 10002 8693
rect 10036 8659 10070 8693
rect 10104 8659 10138 8693
rect 10172 8659 10206 8693
rect 10240 8659 10274 8693
rect 10308 8659 10342 8693
rect 10376 8659 10410 8693
rect 10444 8659 10478 8693
rect 10512 8659 10546 8693
rect 10580 8659 10614 8693
rect 10648 8659 10682 8693
rect 10716 8659 10750 8693
rect 10784 8659 10818 8693
rect 10852 8659 10886 8693
rect 10920 8659 10954 8693
rect 10988 8659 11022 8693
rect 11056 8659 11090 8693
rect 11124 8659 11158 8693
rect 11192 8659 11226 8693
rect 11260 8659 11294 8693
rect 11328 8659 11362 8693
rect 11396 8659 11430 8693
rect 11464 8659 11498 8693
rect 11532 8659 11566 8693
rect 11600 8659 11634 8693
rect 11668 8659 11702 8693
rect 11736 8659 11770 8693
rect 11804 8659 11838 8693
rect 11872 8659 11906 8693
rect 11940 8659 11974 8693
rect 12008 8659 12042 8693
rect 12076 8659 12110 8693
rect 12144 8659 12178 8693
rect 12212 8659 12246 8693
rect 12280 8659 12314 8693
rect 12348 8659 12382 8693
rect 12416 8659 12450 8693
rect 12484 8659 12518 8693
rect 12552 8659 12586 8693
rect 12620 8659 12654 8693
rect 12688 8659 12722 8693
rect 12756 8659 12790 8693
rect 12824 8659 12858 8693
rect 12892 8659 12926 8693
rect 12960 8659 12994 8693
rect 13028 8659 13062 8693
rect 13096 8659 13130 8693
rect 13164 8659 13198 8693
rect 13232 8659 13266 8693
rect 13300 8659 13334 8693
rect 13368 8659 13402 8693
rect 13436 8659 13470 8693
rect 13504 8659 13538 8693
rect 13572 8659 13606 8693
rect 13640 8659 13674 8693
rect 13708 8659 13742 8693
rect 13776 8659 13810 8693
rect 13844 8659 13878 8693
rect 13912 8659 13946 8693
rect 13980 8659 14014 8693
rect 14048 8659 14082 8693
rect 14116 8659 14150 8693
rect 14184 8659 14218 8693
rect 14252 8659 14286 8693
rect 14320 8659 14354 8693
rect 14388 8659 14422 8693
rect 14456 8659 14490 8693
rect 14524 8659 14558 8693
rect 14592 8659 14626 8693
rect 14660 8659 14694 8693
rect 14728 8659 14762 8693
rect 14796 8659 14830 8693
rect 14864 8659 14898 8693
rect 14932 8687 14966 8721
rect 15000 8687 15034 8721
rect 15068 8687 15102 8721
rect 68 8592 102 8626
rect 138 8592 172 8626
rect 208 8592 242 8626
rect 278 8592 312 8626
rect 348 8592 382 8626
rect 418 8592 452 8626
rect 488 8592 522 8626
rect 558 8592 592 8626
rect 628 8592 662 8626
rect 698 8592 732 8626
rect 768 8592 802 8626
rect 838 8592 872 8626
rect 908 8592 942 8626
rect 978 8592 1012 8626
rect 1048 8592 1082 8626
rect 1118 8592 1152 8626
rect 1188 8592 1222 8626
rect 1258 8592 1292 8626
rect 1328 8592 1362 8626
rect 1398 8592 1432 8626
rect 1467 8592 1501 8626
rect 1536 8592 1570 8626
rect 1605 8592 1639 8626
rect 1674 8592 1708 8626
rect 1743 8592 1777 8626
rect 1812 8592 1846 8626
rect 1881 8592 1915 8626
rect 1950 8592 1984 8626
rect 2019 8592 2053 8626
rect 2088 8592 2122 8626
rect 2157 8592 2191 8626
rect 2226 8592 2260 8626
rect 2295 8592 2329 8626
rect 2364 8592 2398 8626
rect 2433 8592 2467 8626
rect 2502 8592 2536 8626
rect 2571 8592 2605 8626
rect 2640 8592 2674 8626
rect 2709 8592 2743 8626
rect 2778 8592 2812 8626
rect 2847 8592 2881 8626
rect 2933 8596 2967 8630
rect 3002 8596 3036 8630
rect 3071 8596 3105 8630
rect 3139 8596 3173 8630
rect 3207 8596 3241 8630
rect 3275 8596 3309 8630
rect 3343 8596 3377 8630
rect 3411 8596 3445 8630
rect 3479 8596 3513 8630
rect 3547 8596 3581 8630
rect 3615 8596 3649 8630
rect 3683 8596 3717 8630
rect 3751 8596 3785 8630
rect 3819 8596 3853 8630
rect 3887 8596 3921 8630
rect 3955 8596 3989 8630
rect 4023 8596 4057 8630
rect 4091 8596 4125 8630
rect 4159 8596 4193 8630
rect 4227 8596 4261 8630
rect 4295 8596 4329 8630
rect 4363 8596 4397 8630
rect 4431 8596 4465 8630
rect 4499 8596 4533 8630
rect 4567 8596 4601 8630
rect 4635 8596 4669 8630
rect 4703 8596 4737 8630
rect 4771 8596 4805 8630
rect 4839 8596 4873 8630
rect 4907 8596 4941 8630
rect 4975 8596 5009 8630
rect 5043 8596 5077 8630
rect 5111 8596 5145 8630
rect 5179 8596 5213 8630
rect 5247 8596 5281 8630
rect 5315 8596 5349 8630
rect 5383 8596 5417 8630
rect 5451 8596 5485 8630
rect 5519 8596 5553 8630
rect 5587 8596 5621 8630
rect 5655 8596 5689 8630
rect 5723 8596 5757 8630
rect 5791 8596 5825 8630
rect 5859 8596 5893 8630
rect 5927 8596 5961 8630
rect 5995 8596 6029 8630
rect 6063 8596 6097 8630
rect 6131 8596 6165 8630
rect 6199 8596 6233 8630
rect 6267 8596 6301 8630
rect 6335 8596 6369 8630
rect 6403 8596 6437 8630
rect 6471 8596 6505 8630
rect 6539 8596 6573 8630
rect 6607 8596 6641 8630
rect 6675 8596 6709 8630
rect 6743 8596 6777 8630
rect 6811 8596 6845 8630
rect 6879 8596 6913 8630
rect 6947 8596 6981 8630
rect 7015 8596 7049 8630
rect 7083 8596 7117 8630
rect 7151 8596 7185 8630
rect 7219 8596 7253 8630
rect 7287 8596 7321 8630
rect 7355 8596 7389 8630
rect 7423 8596 7457 8630
rect 7491 8596 7525 8630
rect 7559 8596 7593 8630
rect 7627 8596 7661 8630
rect 7695 8596 7729 8630
rect 7763 8596 7797 8630
rect 7831 8596 7865 8630
rect 7899 8596 7933 8630
rect 7967 8596 8001 8630
rect 8035 8596 8069 8630
rect 8103 8596 8137 8630
rect 8171 8596 8205 8630
rect 8239 8596 8273 8630
rect 8307 8596 8341 8630
rect 14932 8615 14966 8649
rect 15000 8615 15034 8649
rect 15068 8615 15102 8649
rect 8393 8579 8427 8613
rect 8462 8579 8496 8613
rect 8531 8579 8565 8613
rect 8600 8579 8634 8613
rect 8669 8579 8703 8613
rect 8738 8579 8772 8613
rect 8807 8579 8841 8613
rect 8876 8579 8910 8613
rect 8945 8579 8979 8613
rect 9014 8579 9048 8613
rect 9083 8579 9117 8613
rect 9152 8579 9186 8613
rect 9220 8579 9254 8613
rect 9288 8579 9322 8613
rect 9356 8579 9390 8613
rect 9424 8579 9458 8613
rect 9492 8579 9526 8613
rect 9560 8579 9594 8613
rect 9628 8579 9662 8613
rect 9696 8579 9730 8613
rect 9764 8579 9798 8613
rect 9832 8579 9866 8613
rect 9900 8579 9934 8613
rect 9968 8579 10002 8613
rect 10036 8579 10070 8613
rect 10104 8579 10138 8613
rect 10172 8579 10206 8613
rect 10240 8579 10274 8613
rect 10308 8579 10342 8613
rect 10376 8579 10410 8613
rect 10444 8579 10478 8613
rect 10512 8579 10546 8613
rect 10580 8579 10614 8613
rect 10648 8579 10682 8613
rect 10716 8579 10750 8613
rect 10784 8579 10818 8613
rect 10852 8579 10886 8613
rect 10920 8579 10954 8613
rect 10988 8579 11022 8613
rect 11056 8579 11090 8613
rect 11124 8579 11158 8613
rect 11192 8579 11226 8613
rect 11260 8579 11294 8613
rect 11328 8579 11362 8613
rect 11396 8579 11430 8613
rect 11464 8579 11498 8613
rect 11532 8579 11566 8613
rect 11600 8579 11634 8613
rect 11668 8579 11702 8613
rect 11736 8579 11770 8613
rect 11804 8579 11838 8613
rect 11872 8579 11906 8613
rect 11940 8579 11974 8613
rect 12008 8579 12042 8613
rect 12076 8579 12110 8613
rect 12144 8579 12178 8613
rect 12212 8579 12246 8613
rect 12280 8579 12314 8613
rect 12348 8579 12382 8613
rect 12416 8579 12450 8613
rect 12484 8579 12518 8613
rect 12552 8579 12586 8613
rect 12620 8579 12654 8613
rect 12688 8579 12722 8613
rect 12756 8579 12790 8613
rect 12824 8579 12858 8613
rect 12892 8579 12926 8613
rect 12960 8579 12994 8613
rect 13028 8579 13062 8613
rect 13096 8579 13130 8613
rect 13164 8579 13198 8613
rect 13232 8579 13266 8613
rect 13300 8579 13334 8613
rect 13368 8579 13402 8613
rect 13436 8579 13470 8613
rect 13504 8579 13538 8613
rect 13572 8579 13606 8613
rect 13640 8579 13674 8613
rect 13708 8579 13742 8613
rect 13776 8579 13810 8613
rect 13844 8579 13878 8613
rect 13912 8579 13946 8613
rect 13980 8579 14014 8613
rect 14048 8579 14082 8613
rect 14116 8579 14150 8613
rect 14184 8579 14218 8613
rect 14252 8579 14286 8613
rect 14320 8579 14354 8613
rect 14388 8579 14422 8613
rect 14456 8579 14490 8613
rect 14524 8579 14558 8613
rect 14592 8579 14626 8613
rect 14660 8579 14694 8613
rect 14728 8579 14762 8613
rect 14796 8579 14830 8613
rect 14864 8579 14898 8613
rect 68 8518 102 8552
rect 138 8518 172 8552
rect 208 8518 242 8552
rect 278 8518 312 8552
rect 348 8518 382 8552
rect 418 8518 452 8552
rect 488 8518 522 8552
rect 558 8518 592 8552
rect 628 8518 662 8552
rect 698 8518 732 8552
rect 768 8518 802 8552
rect 838 8518 872 8552
rect 908 8518 942 8552
rect 978 8518 1012 8552
rect 1048 8518 1082 8552
rect 1118 8518 1152 8552
rect 1188 8518 1222 8552
rect 1258 8518 1292 8552
rect 1328 8518 1362 8552
rect 1398 8518 1432 8552
rect 1467 8518 1501 8552
rect 1536 8518 1570 8552
rect 1605 8518 1639 8552
rect 1674 8518 1708 8552
rect 1743 8518 1777 8552
rect 1812 8518 1846 8552
rect 1881 8518 1915 8552
rect 1950 8518 1984 8552
rect 2019 8518 2053 8552
rect 2088 8518 2122 8552
rect 2157 8518 2191 8552
rect 2226 8518 2260 8552
rect 2295 8518 2329 8552
rect 2364 8518 2398 8552
rect 2433 8518 2467 8552
rect 2502 8518 2536 8552
rect 2571 8518 2605 8552
rect 2640 8518 2674 8552
rect 2709 8518 2743 8552
rect 2778 8518 2812 8552
rect 2847 8518 2881 8552
rect 2933 8526 2967 8560
rect 3002 8526 3036 8560
rect 3071 8526 3105 8560
rect 3139 8526 3173 8560
rect 3207 8526 3241 8560
rect 3275 8526 3309 8560
rect 3343 8526 3377 8560
rect 3411 8526 3445 8560
rect 3479 8526 3513 8560
rect 3547 8526 3581 8560
rect 3615 8526 3649 8560
rect 3683 8526 3717 8560
rect 3751 8526 3785 8560
rect 3819 8526 3853 8560
rect 3887 8526 3921 8560
rect 3955 8526 3989 8560
rect 4023 8526 4057 8560
rect 4091 8526 4125 8560
rect 4159 8526 4193 8560
rect 4227 8526 4261 8560
rect 4295 8526 4329 8560
rect 4363 8526 4397 8560
rect 4431 8526 4465 8560
rect 4499 8526 4533 8560
rect 4567 8526 4601 8560
rect 4635 8526 4669 8560
rect 4703 8526 4737 8560
rect 4771 8526 4805 8560
rect 4839 8526 4873 8560
rect 4907 8526 4941 8560
rect 4975 8526 5009 8560
rect 5043 8526 5077 8560
rect 5111 8526 5145 8560
rect 5179 8526 5213 8560
rect 5247 8526 5281 8560
rect 5315 8526 5349 8560
rect 5383 8526 5417 8560
rect 5451 8526 5485 8560
rect 5519 8526 5553 8560
rect 5587 8526 5621 8560
rect 5655 8526 5689 8560
rect 5723 8526 5757 8560
rect 5791 8526 5825 8560
rect 5859 8526 5893 8560
rect 5927 8526 5961 8560
rect 5995 8526 6029 8560
rect 6063 8526 6097 8560
rect 6131 8526 6165 8560
rect 6199 8526 6233 8560
rect 6267 8526 6301 8560
rect 6335 8526 6369 8560
rect 6403 8526 6437 8560
rect 6471 8526 6505 8560
rect 6539 8526 6573 8560
rect 6607 8526 6641 8560
rect 6675 8526 6709 8560
rect 6743 8526 6777 8560
rect 6811 8526 6845 8560
rect 6879 8526 6913 8560
rect 6947 8526 6981 8560
rect 7015 8526 7049 8560
rect 7083 8526 7117 8560
rect 7151 8526 7185 8560
rect 7219 8526 7253 8560
rect 7287 8526 7321 8560
rect 7355 8526 7389 8560
rect 7423 8526 7457 8560
rect 7491 8526 7525 8560
rect 7559 8526 7593 8560
rect 7627 8526 7661 8560
rect 7695 8526 7729 8560
rect 7763 8526 7797 8560
rect 7831 8526 7865 8560
rect 7899 8526 7933 8560
rect 7967 8526 8001 8560
rect 8035 8526 8069 8560
rect 8103 8526 8137 8560
rect 8171 8526 8205 8560
rect 8239 8526 8273 8560
rect 8307 8526 8341 8560
rect 14932 8543 14966 8577
rect 15000 8543 15034 8577
rect 15068 8543 15102 8577
rect 8393 8499 8427 8533
rect 8462 8499 8496 8533
rect 8531 8499 8565 8533
rect 8600 8499 8634 8533
rect 8669 8499 8703 8533
rect 8738 8499 8772 8533
rect 8807 8499 8841 8533
rect 8876 8499 8910 8533
rect 8945 8499 8979 8533
rect 9014 8499 9048 8533
rect 9083 8499 9117 8533
rect 9152 8499 9186 8533
rect 9220 8499 9254 8533
rect 9288 8499 9322 8533
rect 9356 8499 9390 8533
rect 9424 8499 9458 8533
rect 9492 8499 9526 8533
rect 9560 8499 9594 8533
rect 9628 8499 9662 8533
rect 9696 8499 9730 8533
rect 9764 8499 9798 8533
rect 9832 8499 9866 8533
rect 9900 8499 9934 8533
rect 9968 8499 10002 8533
rect 10036 8499 10070 8533
rect 10104 8499 10138 8533
rect 10172 8499 10206 8533
rect 10240 8499 10274 8533
rect 10308 8499 10342 8533
rect 10376 8499 10410 8533
rect 10444 8499 10478 8533
rect 10512 8499 10546 8533
rect 10580 8499 10614 8533
rect 10648 8499 10682 8533
rect 10716 8499 10750 8533
rect 10784 8499 10818 8533
rect 10852 8499 10886 8533
rect 10920 8499 10954 8533
rect 10988 8499 11022 8533
rect 11056 8499 11090 8533
rect 11124 8499 11158 8533
rect 11192 8499 11226 8533
rect 11260 8499 11294 8533
rect 11328 8499 11362 8533
rect 11396 8499 11430 8533
rect 11464 8499 11498 8533
rect 11532 8499 11566 8533
rect 11600 8499 11634 8533
rect 11668 8499 11702 8533
rect 11736 8499 11770 8533
rect 11804 8499 11838 8533
rect 11872 8499 11906 8533
rect 11940 8499 11974 8533
rect 12008 8499 12042 8533
rect 12076 8499 12110 8533
rect 12144 8499 12178 8533
rect 12212 8499 12246 8533
rect 12280 8499 12314 8533
rect 12348 8499 12382 8533
rect 12416 8499 12450 8533
rect 12484 8499 12518 8533
rect 12552 8499 12586 8533
rect 12620 8499 12654 8533
rect 12688 8499 12722 8533
rect 12756 8499 12790 8533
rect 12824 8499 12858 8533
rect 12892 8499 12926 8533
rect 12960 8499 12994 8533
rect 13028 8499 13062 8533
rect 13096 8499 13130 8533
rect 13164 8499 13198 8533
rect 13232 8499 13266 8533
rect 13300 8499 13334 8533
rect 13368 8499 13402 8533
rect 13436 8499 13470 8533
rect 13504 8499 13538 8533
rect 13572 8499 13606 8533
rect 13640 8499 13674 8533
rect 13708 8499 13742 8533
rect 13776 8499 13810 8533
rect 13844 8499 13878 8533
rect 13912 8499 13946 8533
rect 13980 8499 14014 8533
rect 14048 8499 14082 8533
rect 14116 8499 14150 8533
rect 14184 8499 14218 8533
rect 14252 8499 14286 8533
rect 14320 8499 14354 8533
rect 14388 8499 14422 8533
rect 14456 8499 14490 8533
rect 14524 8499 14558 8533
rect 14592 8499 14626 8533
rect 14660 8499 14694 8533
rect 14728 8499 14762 8533
rect 14796 8499 14830 8533
rect 14864 8499 14898 8533
rect 68 8426 102 8460
rect 68 8358 102 8392
rect 68 8290 102 8324
rect 68 8222 102 8256
rect 2933 8456 2967 8490
rect 3002 8456 3036 8490
rect 3071 8456 3105 8490
rect 3139 8456 3173 8490
rect 3207 8456 3241 8490
rect 3275 8456 3309 8490
rect 3343 8456 3377 8490
rect 3411 8456 3445 8490
rect 3479 8456 3513 8490
rect 3547 8456 3581 8490
rect 3615 8456 3649 8490
rect 3683 8456 3717 8490
rect 3751 8456 3785 8490
rect 3819 8456 3853 8490
rect 3887 8456 3921 8490
rect 3955 8456 3989 8490
rect 4023 8456 4057 8490
rect 4091 8456 4125 8490
rect 4159 8456 4193 8490
rect 4227 8456 4261 8490
rect 4295 8456 4329 8490
rect 4363 8456 4397 8490
rect 4431 8456 4465 8490
rect 4499 8456 4533 8490
rect 4567 8456 4601 8490
rect 4635 8456 4669 8490
rect 4703 8456 4737 8490
rect 4771 8456 4805 8490
rect 4839 8456 4873 8490
rect 4907 8456 4941 8490
rect 4975 8456 5009 8490
rect 5043 8456 5077 8490
rect 5111 8456 5145 8490
rect 5179 8456 5213 8490
rect 5247 8456 5281 8490
rect 5315 8456 5349 8490
rect 5383 8456 5417 8490
rect 5451 8456 5485 8490
rect 5519 8456 5553 8490
rect 5587 8456 5621 8490
rect 5655 8456 5689 8490
rect 5723 8456 5757 8490
rect 5791 8456 5825 8490
rect 5859 8456 5893 8490
rect 5927 8456 5961 8490
rect 5995 8456 6029 8490
rect 6063 8456 6097 8490
rect 6131 8456 6165 8490
rect 6199 8456 6233 8490
rect 6267 8456 6301 8490
rect 6335 8456 6369 8490
rect 6403 8456 6437 8490
rect 6471 8456 6505 8490
rect 6539 8456 6573 8490
rect 6607 8456 6641 8490
rect 6675 8456 6709 8490
rect 6743 8456 6777 8490
rect 6811 8456 6845 8490
rect 6879 8456 6913 8490
rect 6947 8456 6981 8490
rect 7015 8456 7049 8490
rect 7083 8456 7117 8490
rect 7151 8456 7185 8490
rect 7219 8456 7253 8490
rect 7287 8456 7321 8490
rect 7355 8456 7389 8490
rect 7423 8456 7457 8490
rect 7491 8456 7525 8490
rect 7559 8456 7593 8490
rect 7627 8456 7661 8490
rect 7695 8456 7729 8490
rect 7763 8456 7797 8490
rect 7831 8456 7865 8490
rect 7899 8456 7933 8490
rect 7967 8456 8001 8490
rect 8035 8456 8069 8490
rect 8103 8456 8137 8490
rect 8171 8456 8205 8490
rect 8239 8456 8273 8490
rect 8307 8456 8341 8490
rect 14932 8471 14966 8505
rect 15000 8471 15034 8505
rect 15068 8471 15102 8505
rect 2933 8386 2967 8420
rect 3002 8386 3036 8420
rect 3071 8386 3105 8420
rect 3139 8386 3173 8420
rect 3207 8386 3241 8420
rect 3275 8386 3309 8420
rect 3343 8386 3377 8420
rect 3411 8386 3445 8420
rect 3479 8386 3513 8420
rect 3547 8386 3581 8420
rect 3615 8386 3649 8420
rect 3683 8386 3717 8420
rect 3751 8386 3785 8420
rect 3819 8386 3853 8420
rect 3887 8386 3921 8420
rect 3955 8386 3989 8420
rect 4023 8386 4057 8420
rect 4091 8386 4125 8420
rect 4159 8386 4193 8420
rect 4227 8386 4261 8420
rect 4295 8386 4329 8420
rect 4363 8386 4397 8420
rect 4431 8386 4465 8420
rect 4499 8386 4533 8420
rect 4567 8386 4601 8420
rect 4635 8386 4669 8420
rect 4703 8386 4737 8420
rect 4771 8386 4805 8420
rect 4839 8386 4873 8420
rect 4907 8386 4941 8420
rect 4975 8386 5009 8420
rect 5043 8386 5077 8420
rect 5111 8386 5145 8420
rect 5179 8386 5213 8420
rect 5247 8386 5281 8420
rect 5315 8386 5349 8420
rect 5383 8386 5417 8420
rect 5451 8386 5485 8420
rect 5519 8386 5553 8420
rect 5587 8386 5621 8420
rect 5655 8386 5689 8420
rect 5723 8386 5757 8420
rect 5791 8386 5825 8420
rect 5859 8386 5893 8420
rect 5927 8386 5961 8420
rect 5995 8386 6029 8420
rect 6063 8386 6097 8420
rect 6131 8386 6165 8420
rect 6199 8386 6233 8420
rect 6267 8386 6301 8420
rect 6335 8386 6369 8420
rect 6403 8386 6437 8420
rect 6471 8386 6505 8420
rect 6539 8386 6573 8420
rect 6607 8386 6641 8420
rect 6675 8386 6709 8420
rect 6743 8386 6777 8420
rect 6811 8386 6845 8420
rect 6879 8386 6913 8420
rect 6947 8386 6981 8420
rect 7015 8386 7049 8420
rect 7083 8386 7117 8420
rect 7151 8386 7185 8420
rect 7219 8386 7253 8420
rect 7287 8386 7321 8420
rect 7355 8386 7389 8420
rect 7423 8386 7457 8420
rect 7491 8386 7525 8420
rect 7559 8386 7593 8420
rect 7627 8386 7661 8420
rect 7695 8386 7729 8420
rect 7763 8386 7797 8420
rect 7831 8386 7865 8420
rect 7899 8386 7933 8420
rect 7967 8386 8001 8420
rect 8035 8386 8069 8420
rect 8103 8386 8137 8420
rect 8171 8386 8205 8420
rect 8239 8386 8273 8420
rect 8307 8386 8341 8420
rect 8393 8419 8427 8453
rect 8462 8419 8496 8453
rect 8531 8419 8565 8453
rect 8600 8419 8634 8453
rect 8669 8419 8703 8453
rect 8738 8419 8772 8453
rect 8807 8419 8841 8453
rect 8876 8419 8910 8453
rect 8945 8419 8979 8453
rect 9014 8419 9048 8453
rect 9083 8419 9117 8453
rect 9152 8419 9186 8453
rect 9220 8419 9254 8453
rect 9288 8419 9322 8453
rect 9356 8419 9390 8453
rect 9424 8419 9458 8453
rect 9492 8419 9526 8453
rect 9560 8419 9594 8453
rect 9628 8419 9662 8453
rect 9696 8419 9730 8453
rect 9764 8419 9798 8453
rect 9832 8419 9866 8453
rect 9900 8419 9934 8453
rect 9968 8419 10002 8453
rect 10036 8419 10070 8453
rect 10104 8419 10138 8453
rect 10172 8419 10206 8453
rect 10240 8419 10274 8453
rect 10308 8419 10342 8453
rect 10376 8419 10410 8453
rect 10444 8419 10478 8453
rect 10512 8419 10546 8453
rect 10580 8419 10614 8453
rect 10648 8419 10682 8453
rect 10716 8419 10750 8453
rect 10784 8419 10818 8453
rect 10852 8419 10886 8453
rect 10920 8419 10954 8453
rect 10988 8419 11022 8453
rect 11056 8419 11090 8453
rect 11124 8419 11158 8453
rect 11192 8419 11226 8453
rect 11260 8419 11294 8453
rect 11328 8419 11362 8453
rect 11396 8419 11430 8453
rect 11464 8419 11498 8453
rect 11532 8419 11566 8453
rect 11600 8419 11634 8453
rect 11668 8419 11702 8453
rect 11736 8419 11770 8453
rect 11804 8419 11838 8453
rect 11872 8419 11906 8453
rect 11940 8419 11974 8453
rect 12008 8419 12042 8453
rect 12076 8419 12110 8453
rect 12144 8419 12178 8453
rect 12212 8419 12246 8453
rect 12280 8419 12314 8453
rect 12348 8419 12382 8453
rect 12416 8419 12450 8453
rect 12484 8419 12518 8453
rect 12552 8419 12586 8453
rect 12620 8419 12654 8453
rect 12688 8419 12722 8453
rect 12756 8419 12790 8453
rect 12824 8419 12858 8453
rect 12892 8419 12926 8453
rect 12960 8419 12994 8453
rect 13028 8419 13062 8453
rect 13096 8419 13130 8453
rect 13164 8419 13198 8453
rect 13232 8419 13266 8453
rect 13300 8419 13334 8453
rect 13368 8419 13402 8453
rect 13436 8419 13470 8453
rect 13504 8419 13538 8453
rect 13572 8419 13606 8453
rect 13640 8419 13674 8453
rect 13708 8419 13742 8453
rect 13776 8419 13810 8453
rect 13844 8419 13878 8453
rect 13912 8419 13946 8453
rect 13980 8419 14014 8453
rect 14048 8419 14082 8453
rect 14116 8419 14150 8453
rect 14184 8419 14218 8453
rect 14252 8419 14286 8453
rect 14320 8419 14354 8453
rect 14388 8419 14422 8453
rect 14456 8419 14490 8453
rect 14524 8419 14558 8453
rect 14592 8419 14626 8453
rect 14660 8419 14694 8453
rect 14728 8419 14762 8453
rect 14796 8419 14830 8453
rect 14864 8419 14898 8453
rect 14932 8399 14966 8433
rect 15000 8399 15034 8433
rect 15068 8399 15102 8433
rect 2933 8316 2967 8350
rect 3002 8316 3036 8350
rect 3071 8316 3105 8350
rect 3139 8316 3173 8350
rect 3207 8316 3241 8350
rect 3275 8316 3309 8350
rect 3343 8316 3377 8350
rect 3411 8316 3445 8350
rect 3479 8316 3513 8350
rect 3547 8316 3581 8350
rect 3615 8316 3649 8350
rect 3683 8316 3717 8350
rect 3751 8316 3785 8350
rect 3819 8316 3853 8350
rect 3887 8316 3921 8350
rect 3955 8316 3989 8350
rect 4023 8316 4057 8350
rect 4091 8316 4125 8350
rect 4159 8316 4193 8350
rect 4227 8316 4261 8350
rect 4295 8316 4329 8350
rect 4363 8316 4397 8350
rect 4431 8316 4465 8350
rect 4499 8316 4533 8350
rect 4567 8316 4601 8350
rect 4635 8316 4669 8350
rect 4703 8316 4737 8350
rect 4771 8316 4805 8350
rect 4839 8316 4873 8350
rect 4907 8316 4941 8350
rect 4975 8316 5009 8350
rect 5043 8316 5077 8350
rect 5111 8316 5145 8350
rect 5179 8316 5213 8350
rect 5247 8316 5281 8350
rect 5315 8316 5349 8350
rect 5383 8316 5417 8350
rect 5451 8316 5485 8350
rect 5519 8316 5553 8350
rect 5587 8316 5621 8350
rect 5655 8316 5689 8350
rect 5723 8316 5757 8350
rect 5791 8316 5825 8350
rect 5859 8316 5893 8350
rect 5927 8316 5961 8350
rect 5995 8316 6029 8350
rect 6063 8316 6097 8350
rect 6131 8316 6165 8350
rect 6199 8316 6233 8350
rect 6267 8316 6301 8350
rect 6335 8316 6369 8350
rect 6403 8316 6437 8350
rect 6471 8316 6505 8350
rect 6539 8316 6573 8350
rect 6607 8316 6641 8350
rect 6675 8316 6709 8350
rect 6743 8316 6777 8350
rect 6811 8316 6845 8350
rect 6879 8316 6913 8350
rect 6947 8316 6981 8350
rect 7015 8316 7049 8350
rect 7083 8316 7117 8350
rect 7151 8316 7185 8350
rect 7219 8316 7253 8350
rect 7287 8316 7321 8350
rect 7355 8316 7389 8350
rect 7423 8316 7457 8350
rect 7491 8316 7525 8350
rect 7559 8316 7593 8350
rect 7627 8316 7661 8350
rect 7695 8316 7729 8350
rect 7763 8316 7797 8350
rect 7831 8316 7865 8350
rect 7899 8316 7933 8350
rect 7967 8316 8001 8350
rect 8035 8316 8069 8350
rect 8103 8316 8137 8350
rect 8171 8316 8205 8350
rect 8239 8316 8273 8350
rect 8307 8316 8341 8350
rect 13532 8323 13566 8357
rect 13603 8323 13637 8357
rect 13674 8323 13708 8357
rect 13744 8323 13778 8357
rect 13814 8323 13848 8357
rect 13884 8323 13918 8357
rect 13954 8323 13988 8357
rect 14024 8323 14058 8357
rect 14094 8323 14128 8357
rect 14164 8323 14198 8357
rect 14234 8323 14268 8357
rect 14304 8323 14338 8357
rect 14374 8323 14408 8357
rect 14444 8323 14478 8357
rect 14514 8323 14548 8357
rect 14584 8323 14618 8357
rect 14654 8323 14688 8357
rect 14724 8323 14758 8357
rect 14794 8323 14828 8357
rect 14864 8323 14898 8357
rect 14932 8327 14966 8361
rect 15000 8327 15034 8361
rect 15068 8327 15102 8361
rect 2933 8246 2967 8280
rect 3002 8246 3036 8280
rect 3071 8246 3105 8280
rect 3139 8246 3173 8280
rect 3207 8246 3241 8280
rect 3275 8246 3309 8280
rect 3343 8246 3377 8280
rect 3411 8246 3445 8280
rect 3479 8246 3513 8280
rect 3547 8246 3581 8280
rect 3615 8246 3649 8280
rect 3683 8246 3717 8280
rect 3751 8246 3785 8280
rect 3819 8246 3853 8280
rect 3887 8246 3921 8280
rect 3955 8246 3989 8280
rect 4023 8246 4057 8280
rect 4091 8246 4125 8280
rect 4159 8246 4193 8280
rect 4227 8246 4261 8280
rect 4295 8246 4329 8280
rect 4363 8246 4397 8280
rect 4431 8246 4465 8280
rect 4499 8246 4533 8280
rect 4567 8246 4601 8280
rect 4635 8246 4669 8280
rect 4703 8246 4737 8280
rect 4771 8246 4805 8280
rect 4839 8246 4873 8280
rect 4907 8246 4941 8280
rect 4975 8246 5009 8280
rect 5043 8246 5077 8280
rect 5111 8246 5145 8280
rect 5179 8246 5213 8280
rect 5247 8246 5281 8280
rect 5315 8246 5349 8280
rect 5383 8246 5417 8280
rect 5451 8246 5485 8280
rect 5519 8246 5553 8280
rect 5587 8246 5621 8280
rect 5655 8246 5689 8280
rect 5723 8246 5757 8280
rect 5791 8246 5825 8280
rect 5859 8246 5893 8280
rect 5927 8246 5961 8280
rect 5995 8246 6029 8280
rect 6063 8246 6097 8280
rect 6131 8246 6165 8280
rect 6199 8246 6233 8280
rect 6267 8246 6301 8280
rect 6335 8246 6369 8280
rect 6403 8246 6437 8280
rect 6471 8246 6505 8280
rect 6539 8246 6573 8280
rect 6607 8246 6641 8280
rect 6675 8246 6709 8280
rect 6743 8246 6777 8280
rect 6811 8246 6845 8280
rect 6879 8246 6913 8280
rect 6947 8246 6981 8280
rect 7015 8246 7049 8280
rect 7083 8246 7117 8280
rect 7151 8246 7185 8280
rect 7219 8246 7253 8280
rect 7287 8246 7321 8280
rect 7355 8246 7389 8280
rect 7423 8246 7457 8280
rect 7491 8246 7525 8280
rect 7559 8246 7593 8280
rect 7627 8246 7661 8280
rect 7695 8246 7729 8280
rect 7763 8246 7797 8280
rect 7831 8246 7865 8280
rect 7899 8246 7933 8280
rect 7967 8246 8001 8280
rect 8035 8246 8069 8280
rect 8103 8246 8137 8280
rect 8171 8246 8205 8280
rect 8239 8246 8273 8280
rect 8307 8246 8341 8280
rect 2933 8176 2967 8210
rect 3002 8176 3036 8210
rect 3071 8176 3105 8210
rect 3139 8176 3173 8210
rect 3207 8176 3241 8210
rect 3275 8176 3309 8210
rect 3343 8176 3377 8210
rect 3411 8176 3445 8210
rect 3479 8176 3513 8210
rect 3547 8176 3581 8210
rect 3615 8176 3649 8210
rect 3683 8176 3717 8210
rect 3751 8176 3785 8210
rect 3819 8176 3853 8210
rect 3887 8176 3921 8210
rect 3955 8176 3989 8210
rect 4023 8176 4057 8210
rect 4091 8176 4125 8210
rect 4159 8176 4193 8210
rect 4227 8176 4261 8210
rect 4295 8176 4329 8210
rect 4363 8176 4397 8210
rect 4431 8176 4465 8210
rect 4499 8176 4533 8210
rect 4567 8176 4601 8210
rect 4635 8176 4669 8210
rect 4703 8176 4737 8210
rect 4771 8176 4805 8210
rect 4839 8176 4873 8210
rect 4907 8176 4941 8210
rect 4975 8176 5009 8210
rect 5043 8176 5077 8210
rect 5111 8176 5145 8210
rect 5179 8176 5213 8210
rect 5247 8176 5281 8210
rect 5315 8176 5349 8210
rect 5383 8176 5417 8210
rect 5451 8176 5485 8210
rect 5519 8176 5553 8210
rect 5587 8176 5621 8210
rect 5655 8176 5689 8210
rect 5723 8176 5757 8210
rect 5791 8176 5825 8210
rect 5859 8176 5893 8210
rect 5927 8176 5961 8210
rect 5995 8176 6029 8210
rect 6063 8176 6097 8210
rect 6131 8176 6165 8210
rect 6199 8176 6233 8210
rect 6267 8176 6301 8210
rect 6335 8176 6369 8210
rect 6403 8176 6437 8210
rect 6471 8176 6505 8210
rect 6539 8176 6573 8210
rect 6607 8176 6641 8210
rect 6675 8176 6709 8210
rect 6743 8176 6777 8210
rect 6811 8176 6845 8210
rect 6879 8176 6913 8210
rect 6947 8176 6981 8210
rect 7015 8176 7049 8210
rect 7083 8176 7117 8210
rect 7151 8176 7185 8210
rect 7219 8176 7253 8210
rect 7287 8176 7321 8210
rect 7355 8176 7389 8210
rect 7423 8176 7457 8210
rect 7491 8176 7525 8210
rect 7559 8176 7593 8210
rect 7627 8176 7661 8210
rect 7695 8176 7729 8210
rect 7763 8176 7797 8210
rect 7831 8176 7865 8210
rect 7899 8176 7933 8210
rect 7967 8176 8001 8210
rect 8035 8176 8069 8210
rect 8103 8176 8137 8210
rect 8171 8176 8205 8210
rect 8239 8176 8273 8210
rect 8307 8176 8341 8210
rect 68 8123 102 8157
rect 138 8123 172 8157
rect 208 8123 242 8157
rect 278 8123 312 8157
rect 348 8123 382 8157
rect 418 8123 452 8157
rect 488 8123 522 8157
rect 558 8123 592 8157
rect 628 8123 662 8157
rect 698 8123 732 8157
rect 768 8123 802 8157
rect 838 8123 872 8157
rect 908 8123 942 8157
rect 978 8123 1012 8157
rect 1048 8123 1082 8157
rect 1118 8123 1152 8157
rect 1188 8123 1222 8157
rect 1258 8123 1292 8157
rect 1328 8123 1362 8157
rect 1398 8123 1432 8157
rect 1467 8123 1501 8157
rect 1536 8123 1570 8157
rect 1605 8123 1639 8157
rect 1674 8123 1708 8157
rect 1743 8123 1777 8157
rect 1812 8123 1846 8157
rect 1881 8123 1915 8157
rect 1950 8123 1984 8157
rect 2019 8123 2053 8157
rect 2088 8123 2122 8157
rect 2157 8123 2191 8157
rect 2226 8123 2260 8157
rect 2295 8123 2329 8157
rect 2364 8123 2398 8157
rect 2433 8123 2467 8157
rect 2502 8123 2536 8157
rect 2571 8123 2605 8157
rect 2640 8123 2674 8157
rect 2709 8123 2743 8157
rect 2778 8123 2812 8157
rect 2847 8123 2881 8157
rect 2933 8106 2967 8140
rect 3002 8106 3036 8140
rect 3071 8106 3105 8140
rect 3139 8106 3173 8140
rect 3207 8106 3241 8140
rect 3275 8106 3309 8140
rect 3343 8106 3377 8140
rect 3411 8106 3445 8140
rect 3479 8106 3513 8140
rect 3547 8106 3581 8140
rect 3615 8106 3649 8140
rect 3683 8106 3717 8140
rect 3751 8106 3785 8140
rect 3819 8106 3853 8140
rect 3887 8106 3921 8140
rect 3955 8106 3989 8140
rect 4023 8106 4057 8140
rect 4091 8106 4125 8140
rect 4159 8106 4193 8140
rect 4227 8106 4261 8140
rect 4295 8106 4329 8140
rect 4363 8106 4397 8140
rect 4431 8106 4465 8140
rect 4499 8106 4533 8140
rect 4567 8106 4601 8140
rect 4635 8106 4669 8140
rect 4703 8106 4737 8140
rect 4771 8106 4805 8140
rect 4839 8106 4873 8140
rect 4907 8106 4941 8140
rect 4975 8106 5009 8140
rect 5043 8106 5077 8140
rect 5111 8106 5145 8140
rect 5179 8106 5213 8140
rect 5247 8106 5281 8140
rect 5315 8106 5349 8140
rect 5383 8106 5417 8140
rect 5451 8106 5485 8140
rect 5519 8106 5553 8140
rect 5587 8106 5621 8140
rect 5655 8106 5689 8140
rect 5723 8106 5757 8140
rect 5791 8106 5825 8140
rect 5859 8106 5893 8140
rect 5927 8106 5961 8140
rect 5995 8106 6029 8140
rect 6063 8106 6097 8140
rect 6131 8106 6165 8140
rect 6199 8106 6233 8140
rect 6267 8106 6301 8140
rect 6335 8106 6369 8140
rect 6403 8106 6437 8140
rect 6471 8106 6505 8140
rect 6539 8106 6573 8140
rect 6607 8106 6641 8140
rect 6675 8106 6709 8140
rect 6743 8106 6777 8140
rect 6811 8106 6845 8140
rect 6879 8106 6913 8140
rect 6947 8106 6981 8140
rect 7015 8106 7049 8140
rect 7083 8106 7117 8140
rect 7151 8106 7185 8140
rect 7219 8106 7253 8140
rect 7287 8106 7321 8140
rect 7355 8106 7389 8140
rect 7423 8106 7457 8140
rect 7491 8106 7525 8140
rect 7559 8106 7593 8140
rect 7627 8106 7661 8140
rect 7695 8106 7729 8140
rect 7763 8106 7797 8140
rect 7831 8106 7865 8140
rect 7899 8106 7933 8140
rect 7967 8106 8001 8140
rect 8035 8106 8069 8140
rect 8103 8106 8137 8140
rect 8171 8106 8205 8140
rect 8239 8106 8273 8140
rect 8307 8106 8341 8140
rect 68 8048 102 8082
rect 138 8048 172 8082
rect 208 8048 242 8082
rect 278 8048 312 8082
rect 348 8048 382 8082
rect 418 8048 452 8082
rect 488 8048 522 8082
rect 558 8048 592 8082
rect 628 8048 662 8082
rect 698 8048 732 8082
rect 768 8048 802 8082
rect 838 8048 872 8082
rect 908 8048 942 8082
rect 978 8048 1012 8082
rect 1048 8048 1082 8082
rect 1118 8048 1152 8082
rect 1188 8048 1222 8082
rect 1258 8048 1292 8082
rect 1328 8048 1362 8082
rect 1398 8048 1432 8082
rect 1467 8048 1501 8082
rect 1536 8048 1570 8082
rect 1605 8048 1639 8082
rect 1674 8048 1708 8082
rect 1743 8048 1777 8082
rect 1812 8048 1846 8082
rect 1881 8048 1915 8082
rect 1950 8048 1984 8082
rect 2019 8048 2053 8082
rect 2088 8048 2122 8082
rect 2157 8048 2191 8082
rect 2226 8048 2260 8082
rect 2295 8048 2329 8082
rect 2364 8048 2398 8082
rect 2433 8048 2467 8082
rect 2502 8048 2536 8082
rect 2571 8048 2605 8082
rect 2640 8048 2674 8082
rect 2709 8048 2743 8082
rect 2778 8048 2812 8082
rect 2847 8048 2881 8082
rect 2933 8036 2967 8070
rect 3002 8036 3036 8070
rect 3071 8036 3105 8070
rect 3139 8036 3173 8070
rect 3207 8036 3241 8070
rect 3275 8036 3309 8070
rect 3343 8036 3377 8070
rect 3411 8036 3445 8070
rect 3479 8036 3513 8070
rect 3547 8036 3581 8070
rect 3615 8036 3649 8070
rect 3683 8036 3717 8070
rect 3751 8036 3785 8070
rect 3819 8036 3853 8070
rect 3887 8036 3921 8070
rect 3955 8036 3989 8070
rect 4023 8036 4057 8070
rect 4091 8036 4125 8070
rect 4159 8036 4193 8070
rect 4227 8036 4261 8070
rect 4295 8036 4329 8070
rect 4363 8036 4397 8070
rect 4431 8036 4465 8070
rect 4499 8036 4533 8070
rect 4567 8036 4601 8070
rect 4635 8036 4669 8070
rect 4703 8036 4737 8070
rect 4771 8036 4805 8070
rect 4839 8036 4873 8070
rect 4907 8036 4941 8070
rect 4975 8036 5009 8070
rect 5043 8036 5077 8070
rect 5111 8036 5145 8070
rect 5179 8036 5213 8070
rect 5247 8036 5281 8070
rect 5315 8036 5349 8070
rect 5383 8036 5417 8070
rect 5451 8036 5485 8070
rect 5519 8036 5553 8070
rect 5587 8036 5621 8070
rect 5655 8036 5689 8070
rect 5723 8036 5757 8070
rect 5791 8036 5825 8070
rect 5859 8036 5893 8070
rect 5927 8036 5961 8070
rect 5995 8036 6029 8070
rect 6063 8036 6097 8070
rect 6131 8036 6165 8070
rect 6199 8036 6233 8070
rect 6267 8036 6301 8070
rect 6335 8036 6369 8070
rect 6403 8036 6437 8070
rect 6471 8036 6505 8070
rect 6539 8036 6573 8070
rect 6607 8036 6641 8070
rect 6675 8036 6709 8070
rect 6743 8036 6777 8070
rect 6811 8036 6845 8070
rect 6879 8036 6913 8070
rect 6947 8036 6981 8070
rect 7015 8036 7049 8070
rect 7083 8036 7117 8070
rect 7151 8036 7185 8070
rect 7219 8036 7253 8070
rect 7287 8036 7321 8070
rect 7355 8036 7389 8070
rect 7423 8036 7457 8070
rect 7491 8036 7525 8070
rect 7559 8036 7593 8070
rect 7627 8036 7661 8070
rect 7695 8036 7729 8070
rect 7763 8036 7797 8070
rect 7831 8036 7865 8070
rect 7899 8036 7933 8070
rect 7967 8036 8001 8070
rect 8035 8036 8069 8070
rect 8103 8036 8137 8070
rect 8171 8036 8205 8070
rect 8239 8036 8273 8070
rect 8307 8036 8341 8070
rect 68 7973 102 8007
rect 138 7973 172 8007
rect 208 7973 242 8007
rect 278 7973 312 8007
rect 348 7973 382 8007
rect 418 7973 452 8007
rect 488 7973 522 8007
rect 558 7973 592 8007
rect 628 7973 662 8007
rect 698 7973 732 8007
rect 768 7973 802 8007
rect 838 7973 872 8007
rect 908 7973 942 8007
rect 978 7973 1012 8007
rect 1048 7973 1082 8007
rect 1118 7973 1152 8007
rect 1188 7973 1222 8007
rect 1258 7973 1292 8007
rect 1328 7973 1362 8007
rect 1398 7973 1432 8007
rect 1467 7973 1501 8007
rect 1536 7973 1570 8007
rect 1605 7973 1639 8007
rect 1674 7973 1708 8007
rect 1743 7973 1777 8007
rect 1812 7973 1846 8007
rect 1881 7973 1915 8007
rect 1950 7973 1984 8007
rect 2019 7973 2053 8007
rect 2088 7973 2122 8007
rect 2157 7973 2191 8007
rect 2226 7973 2260 8007
rect 2295 7973 2329 8007
rect 2364 7973 2398 8007
rect 2433 7973 2467 8007
rect 2502 7973 2536 8007
rect 2571 7973 2605 8007
rect 2640 7973 2674 8007
rect 2709 7973 2743 8007
rect 2778 7973 2812 8007
rect 2847 7973 2881 8007
rect 2933 7966 2967 8000
rect 3002 7966 3036 8000
rect 3071 7966 3105 8000
rect 3139 7966 3173 8000
rect 3207 7966 3241 8000
rect 3275 7966 3309 8000
rect 3343 7966 3377 8000
rect 3411 7966 3445 8000
rect 3479 7966 3513 8000
rect 3547 7966 3581 8000
rect 3615 7966 3649 8000
rect 3683 7966 3717 8000
rect 3751 7966 3785 8000
rect 3819 7966 3853 8000
rect 3887 7966 3921 8000
rect 3955 7966 3989 8000
rect 4023 7966 4057 8000
rect 4091 7966 4125 8000
rect 4159 7966 4193 8000
rect 4227 7966 4261 8000
rect 4295 7966 4329 8000
rect 4363 7966 4397 8000
rect 4431 7966 4465 8000
rect 4499 7966 4533 8000
rect 4567 7966 4601 8000
rect 4635 7966 4669 8000
rect 4703 7966 4737 8000
rect 4771 7966 4805 8000
rect 4839 7966 4873 8000
rect 4907 7966 4941 8000
rect 4975 7966 5009 8000
rect 5043 7966 5077 8000
rect 5111 7966 5145 8000
rect 5179 7966 5213 8000
rect 5247 7966 5281 8000
rect 5315 7966 5349 8000
rect 5383 7966 5417 8000
rect 5451 7966 5485 8000
rect 5519 7966 5553 8000
rect 5587 7966 5621 8000
rect 5655 7966 5689 8000
rect 5723 7966 5757 8000
rect 5791 7966 5825 8000
rect 5859 7966 5893 8000
rect 5927 7966 5961 8000
rect 5995 7966 6029 8000
rect 6063 7966 6097 8000
rect 6131 7966 6165 8000
rect 6199 7966 6233 8000
rect 6267 7966 6301 8000
rect 6335 7966 6369 8000
rect 6403 7966 6437 8000
rect 6471 7966 6505 8000
rect 6539 7966 6573 8000
rect 6607 7966 6641 8000
rect 6675 7966 6709 8000
rect 6743 7966 6777 8000
rect 6811 7966 6845 8000
rect 6879 7966 6913 8000
rect 6947 7966 6981 8000
rect 7015 7966 7049 8000
rect 7083 7966 7117 8000
rect 7151 7966 7185 8000
rect 7219 7966 7253 8000
rect 7287 7966 7321 8000
rect 7355 7966 7389 8000
rect 7423 7966 7457 8000
rect 7491 7966 7525 8000
rect 7559 7966 7593 8000
rect 7627 7966 7661 8000
rect 7695 7966 7729 8000
rect 7763 7966 7797 8000
rect 7831 7966 7865 8000
rect 7899 7966 7933 8000
rect 7967 7966 8001 8000
rect 8035 7966 8069 8000
rect 8103 7966 8137 8000
rect 8171 7966 8205 8000
rect 8239 7966 8273 8000
rect 8307 7966 8341 8000
rect 68 7898 102 7932
rect 138 7898 172 7932
rect 208 7898 242 7932
rect 278 7898 312 7932
rect 348 7898 382 7932
rect 418 7898 452 7932
rect 488 7898 522 7932
rect 558 7898 592 7932
rect 628 7898 662 7932
rect 698 7898 732 7932
rect 768 7898 802 7932
rect 838 7898 872 7932
rect 908 7898 942 7932
rect 978 7898 1012 7932
rect 1048 7898 1082 7932
rect 1118 7898 1152 7932
rect 1188 7898 1222 7932
rect 1258 7898 1292 7932
rect 1328 7898 1362 7932
rect 1398 7898 1432 7932
rect 1467 7898 1501 7932
rect 1536 7898 1570 7932
rect 1605 7898 1639 7932
rect 1674 7898 1708 7932
rect 1743 7898 1777 7932
rect 1812 7898 1846 7932
rect 1881 7898 1915 7932
rect 1950 7898 1984 7932
rect 2019 7898 2053 7932
rect 2088 7898 2122 7932
rect 2157 7898 2191 7932
rect 2226 7898 2260 7932
rect 2295 7898 2329 7932
rect 2364 7898 2398 7932
rect 2433 7898 2467 7932
rect 2502 7898 2536 7932
rect 2571 7898 2605 7932
rect 2640 7898 2674 7932
rect 2709 7898 2743 7932
rect 2778 7898 2812 7932
rect 2847 7898 2881 7932
rect 2933 7896 2967 7930
rect 3002 7896 3036 7930
rect 3071 7896 3105 7930
rect 3139 7896 3173 7930
rect 3207 7896 3241 7930
rect 3275 7896 3309 7930
rect 3343 7896 3377 7930
rect 3411 7896 3445 7930
rect 3479 7896 3513 7930
rect 3547 7896 3581 7930
rect 3615 7896 3649 7930
rect 3683 7896 3717 7930
rect 3751 7896 3785 7930
rect 3819 7896 3853 7930
rect 3887 7896 3921 7930
rect 3955 7896 3989 7930
rect 4023 7896 4057 7930
rect 4091 7896 4125 7930
rect 4159 7896 4193 7930
rect 4227 7896 4261 7930
rect 4295 7896 4329 7930
rect 4363 7896 4397 7930
rect 4431 7896 4465 7930
rect 4499 7896 4533 7930
rect 4567 7896 4601 7930
rect 4635 7896 4669 7930
rect 4703 7896 4737 7930
rect 4771 7896 4805 7930
rect 4839 7896 4873 7930
rect 4907 7896 4941 7930
rect 4975 7896 5009 7930
rect 5043 7896 5077 7930
rect 5111 7896 5145 7930
rect 5179 7896 5213 7930
rect 5247 7896 5281 7930
rect 5315 7896 5349 7930
rect 5383 7896 5417 7930
rect 5451 7896 5485 7930
rect 5519 7896 5553 7930
rect 5587 7896 5621 7930
rect 5655 7896 5689 7930
rect 5723 7896 5757 7930
rect 5791 7896 5825 7930
rect 5859 7896 5893 7930
rect 5927 7896 5961 7930
rect 5995 7896 6029 7930
rect 6063 7896 6097 7930
rect 6131 7896 6165 7930
rect 6199 7896 6233 7930
rect 6267 7896 6301 7930
rect 6335 7896 6369 7930
rect 6403 7896 6437 7930
rect 6471 7896 6505 7930
rect 6539 7896 6573 7930
rect 6607 7896 6641 7930
rect 6675 7896 6709 7930
rect 6743 7896 6777 7930
rect 6811 7896 6845 7930
rect 6879 7896 6913 7930
rect 6947 7896 6981 7930
rect 7015 7896 7049 7930
rect 7083 7896 7117 7930
rect 7151 7896 7185 7930
rect 7219 7896 7253 7930
rect 7287 7896 7321 7930
rect 7355 7896 7389 7930
rect 7423 7896 7457 7930
rect 7491 7896 7525 7930
rect 7559 7896 7593 7930
rect 7627 7896 7661 7930
rect 7695 7896 7729 7930
rect 7763 7896 7797 7930
rect 7831 7896 7865 7930
rect 7899 7896 7933 7930
rect 7967 7896 8001 7930
rect 8035 7896 8069 7930
rect 8103 7896 8137 7930
rect 8171 7896 8205 7930
rect 8239 7896 8273 7930
rect 8307 7896 8341 7930
rect 13532 8249 13566 8283
rect 13603 8249 13637 8283
rect 13674 8249 13708 8283
rect 13744 8249 13778 8283
rect 13814 8249 13848 8283
rect 13884 8249 13918 8283
rect 13954 8249 13988 8283
rect 14024 8249 14058 8283
rect 14094 8249 14128 8283
rect 14164 8249 14198 8283
rect 14234 8249 14268 8283
rect 14304 8249 14338 8283
rect 14374 8249 14408 8283
rect 14444 8249 14478 8283
rect 14514 8249 14548 8283
rect 14584 8249 14618 8283
rect 14654 8249 14688 8283
rect 14724 8249 14758 8283
rect 14794 8249 14828 8283
rect 14864 8249 14898 8283
rect 14932 8255 14966 8289
rect 15000 8255 15034 8289
rect 15068 8255 15102 8289
rect 13532 8175 13566 8209
rect 13603 8175 13637 8209
rect 13674 8175 13708 8209
rect 13744 8175 13778 8209
rect 13814 8175 13848 8209
rect 13884 8175 13918 8209
rect 13954 8175 13988 8209
rect 14024 8175 14058 8209
rect 14094 8175 14128 8209
rect 14164 8175 14198 8209
rect 14234 8175 14268 8209
rect 14304 8175 14338 8209
rect 14374 8175 14408 8209
rect 14444 8175 14478 8209
rect 14514 8175 14548 8209
rect 14584 8175 14618 8209
rect 14654 8175 14688 8209
rect 14724 8175 14758 8209
rect 14794 8175 14828 8209
rect 14864 8175 14898 8209
rect 14932 8183 14966 8217
rect 15000 8183 15034 8217
rect 15068 8183 15102 8217
rect 13532 8101 13566 8135
rect 13603 8101 13637 8135
rect 13674 8101 13708 8135
rect 13744 8101 13778 8135
rect 13814 8101 13848 8135
rect 13884 8101 13918 8135
rect 13954 8101 13988 8135
rect 14024 8101 14058 8135
rect 14094 8101 14128 8135
rect 14164 8101 14198 8135
rect 14234 8101 14268 8135
rect 14304 8101 14338 8135
rect 14374 8101 14408 8135
rect 14444 8101 14478 8135
rect 14514 8101 14548 8135
rect 14584 8101 14618 8135
rect 14654 8101 14688 8135
rect 14724 8101 14758 8135
rect 14794 8101 14828 8135
rect 14864 8101 14898 8135
rect 14932 8111 14966 8145
rect 15000 8111 15034 8145
rect 15068 8111 15102 8145
rect 13532 8027 13566 8061
rect 13603 8027 13637 8061
rect 13674 8027 13708 8061
rect 13744 8027 13778 8061
rect 13814 8027 13848 8061
rect 13884 8027 13918 8061
rect 13954 8027 13988 8061
rect 14024 8027 14058 8061
rect 14094 8027 14128 8061
rect 14164 8027 14198 8061
rect 14234 8027 14268 8061
rect 14304 8027 14338 8061
rect 14374 8027 14408 8061
rect 14444 8027 14478 8061
rect 14514 8027 14548 8061
rect 14584 8027 14618 8061
rect 14654 8027 14688 8061
rect 14724 8027 14758 8061
rect 14794 8027 14828 8061
rect 14864 8027 14898 8061
rect 14932 8039 14966 8073
rect 15000 8039 15034 8073
rect 15068 8039 15102 8073
rect 13532 7953 13566 7987
rect 13603 7953 13637 7987
rect 13674 7953 13708 7987
rect 13744 7953 13778 7987
rect 13814 7953 13848 7987
rect 13884 7953 13918 7987
rect 13954 7953 13988 7987
rect 14024 7953 14058 7987
rect 14094 7953 14128 7987
rect 14164 7953 14198 7987
rect 14234 7953 14268 7987
rect 14304 7953 14338 7987
rect 14374 7953 14408 7987
rect 14444 7953 14478 7987
rect 14514 7953 14548 7987
rect 14584 7953 14618 7987
rect 14654 7953 14688 7987
rect 14724 7953 14758 7987
rect 14794 7953 14828 7987
rect 14864 7953 14898 7987
rect 14932 7967 14966 8001
rect 15000 7967 15034 8001
rect 15068 7967 15102 8001
rect 68 7823 102 7857
rect 138 7823 172 7857
rect 208 7823 242 7857
rect 278 7823 312 7857
rect 348 7823 382 7857
rect 418 7823 452 7857
rect 488 7823 522 7857
rect 558 7823 592 7857
rect 628 7823 662 7857
rect 698 7823 732 7857
rect 768 7823 802 7857
rect 838 7823 872 7857
rect 908 7823 942 7857
rect 978 7823 1012 7857
rect 1048 7823 1082 7857
rect 1118 7823 1152 7857
rect 1188 7823 1222 7857
rect 1258 7823 1292 7857
rect 1328 7823 1362 7857
rect 1398 7823 1432 7857
rect 1467 7823 1501 7857
rect 1536 7823 1570 7857
rect 1605 7823 1639 7857
rect 1674 7823 1708 7857
rect 1743 7823 1777 7857
rect 1812 7823 1846 7857
rect 1881 7823 1915 7857
rect 1950 7823 1984 7857
rect 2019 7823 2053 7857
rect 2088 7823 2122 7857
rect 2157 7823 2191 7857
rect 2226 7823 2260 7857
rect 2295 7823 2329 7857
rect 2364 7823 2398 7857
rect 2433 7823 2467 7857
rect 2502 7823 2536 7857
rect 2571 7823 2605 7857
rect 2640 7823 2674 7857
rect 2709 7823 2743 7857
rect 2778 7823 2812 7857
rect 2847 7823 2881 7857
rect 2933 7826 2967 7860
rect 3002 7826 3036 7860
rect 3071 7826 3105 7860
rect 3139 7826 3173 7860
rect 3207 7826 3241 7860
rect 3275 7826 3309 7860
rect 3343 7826 3377 7860
rect 3411 7826 3445 7860
rect 3479 7826 3513 7860
rect 3547 7826 3581 7860
rect 3615 7826 3649 7860
rect 3683 7826 3717 7860
rect 3751 7826 3785 7860
rect 3819 7826 3853 7860
rect 3887 7826 3921 7860
rect 3955 7826 3989 7860
rect 4023 7826 4057 7860
rect 4091 7826 4125 7860
rect 4159 7826 4193 7860
rect 4227 7826 4261 7860
rect 4295 7826 4329 7860
rect 4363 7826 4397 7860
rect 4431 7826 4465 7860
rect 4499 7826 4533 7860
rect 4567 7826 4601 7860
rect 4635 7826 4669 7860
rect 4703 7826 4737 7860
rect 4771 7826 4805 7860
rect 4839 7826 4873 7860
rect 4907 7826 4941 7860
rect 4975 7826 5009 7860
rect 5043 7826 5077 7860
rect 5111 7826 5145 7860
rect 5179 7826 5213 7860
rect 5247 7826 5281 7860
rect 5315 7826 5349 7860
rect 5383 7826 5417 7860
rect 5451 7826 5485 7860
rect 5519 7826 5553 7860
rect 5587 7826 5621 7860
rect 5655 7826 5689 7860
rect 5723 7826 5757 7860
rect 5791 7826 5825 7860
rect 5859 7826 5893 7860
rect 5927 7826 5961 7860
rect 5995 7826 6029 7860
rect 6063 7826 6097 7860
rect 6131 7826 6165 7860
rect 6199 7826 6233 7860
rect 6267 7826 6301 7860
rect 6335 7826 6369 7860
rect 6403 7826 6437 7860
rect 6471 7826 6505 7860
rect 6539 7826 6573 7860
rect 6607 7826 6641 7860
rect 6675 7826 6709 7860
rect 6743 7826 6777 7860
rect 6811 7826 6845 7860
rect 6879 7826 6913 7860
rect 6947 7826 6981 7860
rect 7015 7826 7049 7860
rect 7083 7826 7117 7860
rect 7151 7826 7185 7860
rect 7219 7826 7253 7860
rect 7287 7826 7321 7860
rect 7355 7826 7389 7860
rect 7423 7826 7457 7860
rect 7491 7826 7525 7860
rect 7559 7826 7593 7860
rect 7627 7826 7661 7860
rect 7695 7826 7729 7860
rect 7763 7826 7797 7860
rect 7831 7826 7865 7860
rect 7899 7826 7933 7860
rect 7967 7826 8001 7860
rect 8035 7826 8069 7860
rect 8103 7826 8137 7860
rect 8171 7826 8205 7860
rect 8239 7826 8273 7860
rect 8307 7826 8341 7860
rect 13532 7879 13566 7913
rect 13603 7879 13637 7913
rect 13674 7879 13708 7913
rect 13744 7879 13778 7913
rect 13814 7879 13848 7913
rect 13884 7879 13918 7913
rect 13954 7879 13988 7913
rect 14024 7879 14058 7913
rect 14094 7879 14128 7913
rect 14164 7879 14198 7913
rect 14234 7879 14268 7913
rect 14304 7879 14338 7913
rect 14374 7879 14408 7913
rect 14444 7879 14478 7913
rect 14514 7879 14548 7913
rect 14584 7879 14618 7913
rect 14654 7879 14688 7913
rect 14724 7879 14758 7913
rect 14794 7879 14828 7913
rect 14864 7879 14898 7913
rect 14932 7895 14966 7929
rect 15000 7895 15034 7929
rect 15068 7895 15102 7929
rect 13532 7805 13566 7839
rect 13603 7805 13637 7839
rect 13674 7805 13708 7839
rect 13744 7805 13778 7839
rect 13814 7805 13848 7839
rect 13884 7805 13918 7839
rect 13954 7805 13988 7839
rect 14024 7805 14058 7839
rect 14094 7805 14128 7839
rect 14164 7805 14198 7839
rect 14234 7805 14268 7839
rect 14304 7805 14338 7839
rect 14374 7805 14408 7839
rect 14444 7805 14478 7839
rect 14514 7805 14548 7839
rect 14584 7805 14618 7839
rect 14654 7805 14688 7839
rect 14724 7805 14758 7839
rect 14794 7805 14828 7839
rect 14864 7805 14898 7839
rect 14932 7823 14966 7857
rect 15000 7823 15034 7857
rect 15068 7823 15102 7857
rect 14932 7751 14966 7785
rect 15000 7751 15034 7785
rect 15068 7751 15102 7785
rect 68 7715 102 7749
rect 137 7715 171 7749
rect 206 7715 240 7749
rect 275 7715 309 7749
rect 344 7715 378 7749
rect 413 7715 447 7749
rect 482 7715 516 7749
rect 551 7715 585 7749
rect 620 7715 654 7749
rect 689 7715 723 7749
rect 758 7715 792 7749
rect 827 7715 861 7749
rect 896 7715 930 7749
rect 965 7715 999 7749
rect 1034 7715 1068 7749
rect 1103 7715 1137 7749
rect 1172 7715 1206 7749
rect 1241 7715 1275 7749
rect 1310 7715 1344 7749
rect 1379 7715 1413 7749
rect 1448 7715 1482 7749
rect 1517 7715 1551 7749
rect 1586 7715 1620 7749
rect 1655 7715 1689 7749
rect 1724 7715 1758 7749
rect 1793 7715 1827 7749
rect 1862 7715 1896 7749
rect 1931 7715 1965 7749
rect 2000 7715 2034 7749
rect 2069 7715 2103 7749
rect 2138 7715 2172 7749
rect 2207 7715 2241 7749
rect 2276 7715 2310 7749
rect 2345 7715 2379 7749
rect 2414 7715 2448 7749
rect 2483 7715 2517 7749
rect 2552 7715 2586 7749
rect 2621 7715 2655 7749
rect 2690 7715 2724 7749
rect 2759 7715 2793 7749
rect 2828 7715 2862 7749
rect 2896 7715 2930 7749
rect 2964 7715 2998 7749
rect 3032 7715 3066 7749
rect 3100 7715 3134 7749
rect 3168 7715 3202 7749
rect 3236 7715 3270 7749
rect 3304 7715 3338 7749
rect 3372 7715 3406 7749
rect 3440 7715 3474 7749
rect 3508 7715 3542 7749
rect 3576 7715 3610 7749
rect 3644 7715 3678 7749
rect 3712 7715 3746 7749
rect 3780 7715 3814 7749
rect 3848 7715 3882 7749
rect 3916 7715 3950 7749
rect 3984 7715 4018 7749
rect 4052 7715 4086 7749
rect 4120 7715 4154 7749
rect 4188 7715 4222 7749
rect 4256 7715 4290 7749
rect 4324 7715 4358 7749
rect 4392 7715 4426 7749
rect 4460 7715 4494 7749
rect 4528 7715 4562 7749
rect 4596 7715 4630 7749
rect 4664 7715 4698 7749
rect 4732 7715 4766 7749
rect 4800 7715 4834 7749
rect 4868 7715 4902 7749
rect 4936 7715 4970 7749
rect 5004 7715 5038 7749
rect 5072 7715 5106 7749
rect 5140 7715 5174 7749
rect 5208 7715 5242 7749
rect 5276 7715 5310 7749
rect 5344 7715 5378 7749
rect 5412 7715 5446 7749
rect 5480 7715 5514 7749
rect 5548 7715 5582 7749
rect 5616 7715 5650 7749
rect 5684 7715 5718 7749
rect 5752 7715 5786 7749
rect 5820 7715 5854 7749
rect 5888 7715 5922 7749
rect 5956 7715 5990 7749
rect 6024 7715 6058 7749
rect 6092 7715 6126 7749
rect 6160 7715 6194 7749
rect 6228 7715 6262 7749
rect 6296 7715 6330 7749
rect 6364 7715 6398 7749
rect 6432 7715 6466 7749
rect 6500 7715 6534 7749
rect 6568 7715 6602 7749
rect 6636 7715 6670 7749
rect 6704 7715 6738 7749
rect 6772 7715 6806 7749
rect 6840 7715 6874 7749
rect 6908 7715 6942 7749
rect 6976 7715 7010 7749
rect 7044 7715 7078 7749
rect 7112 7715 7146 7749
rect 7180 7715 7214 7749
rect 7248 7715 7282 7749
rect 7316 7715 7350 7749
rect 7384 7715 7418 7749
rect 7452 7715 7486 7749
rect 7520 7715 7554 7749
rect 7588 7715 7622 7749
rect 7656 7715 7690 7749
rect 7724 7715 7758 7749
rect 7792 7715 7826 7749
rect 7860 7715 7894 7749
rect 7928 7715 7962 7749
rect 7996 7715 8030 7749
rect 8064 7715 8098 7749
rect 8132 7715 8166 7749
rect 8200 7715 8234 7749
rect 8268 7715 8302 7749
rect 8336 7715 8370 7749
rect 8404 7715 8438 7749
rect 8472 7715 8506 7749
rect 8540 7715 8574 7749
rect 8608 7715 8642 7749
rect 8676 7715 8710 7749
rect 8744 7715 8778 7749
rect 8812 7715 8846 7749
rect 8880 7715 8914 7749
rect 8948 7715 8982 7749
rect 9016 7715 9050 7749
rect 9084 7715 9118 7749
rect 9152 7715 9186 7749
rect 9220 7715 9254 7749
rect 9288 7715 9322 7749
rect 9356 7715 9390 7749
rect 9424 7715 9458 7749
rect 9492 7715 9526 7749
rect 9560 7715 9594 7749
rect 9628 7715 9662 7749
rect 9696 7715 9730 7749
rect 9764 7715 9798 7749
rect 9832 7715 9866 7749
rect 9900 7715 9934 7749
rect 9968 7715 10002 7749
rect 10036 7715 10070 7749
rect 10104 7715 10138 7749
rect 10172 7715 10206 7749
rect 10240 7715 10274 7749
rect 10308 7715 10342 7749
rect 10376 7715 10410 7749
rect 10444 7715 10478 7749
rect 10512 7715 10546 7749
rect 10580 7715 10614 7749
rect 10648 7715 10682 7749
rect 10716 7715 10750 7749
rect 10784 7715 10818 7749
rect 10852 7715 10886 7749
rect 10920 7715 10954 7749
rect 10988 7715 11022 7749
rect 11056 7715 11090 7749
rect 11124 7715 11158 7749
rect 11192 7715 11226 7749
rect 11260 7715 11294 7749
rect 11328 7715 11362 7749
rect 11396 7715 11430 7749
rect 11464 7715 11498 7749
rect 11532 7715 11566 7749
rect 11600 7715 11634 7749
rect 11668 7715 11702 7749
rect 11736 7715 11770 7749
rect 11804 7715 11838 7749
rect 11872 7715 11906 7749
rect 11940 7715 11974 7749
rect 12008 7715 12042 7749
rect 12076 7715 12110 7749
rect 12144 7715 12178 7749
rect 12212 7715 12246 7749
rect 12280 7715 12314 7749
rect 12348 7715 12382 7749
rect 12416 7715 12450 7749
rect 12484 7715 12518 7749
rect 12552 7715 12586 7749
rect 12620 7715 12654 7749
rect 12688 7715 12722 7749
rect 12756 7715 12790 7749
rect 12824 7715 12858 7749
rect 12892 7715 12926 7749
rect 12960 7715 12994 7749
rect 13028 7715 13062 7749
rect 13096 7715 13130 7749
rect 13164 7715 13198 7749
rect 13232 7715 13266 7749
rect 13300 7715 13334 7749
rect 13368 7715 13402 7749
rect 13436 7715 13470 7749
rect 13504 7715 13538 7749
rect 13572 7715 13606 7749
rect 13640 7715 13674 7749
rect 13708 7715 13742 7749
rect 13776 7715 13810 7749
rect 13844 7715 13878 7749
rect 13912 7715 13946 7749
rect 13980 7715 14014 7749
rect 14048 7715 14082 7749
rect 14116 7715 14150 7749
rect 14184 7715 14218 7749
rect 14252 7715 14286 7749
rect 14320 7715 14354 7749
rect 14388 7715 14422 7749
rect 14456 7715 14490 7749
rect 14524 7715 14558 7749
rect 14592 7715 14626 7749
rect 14660 7715 14694 7749
rect 14728 7715 14762 7749
rect 14796 7715 14830 7749
rect 14864 7715 14898 7749
rect 14932 7679 14966 7713
rect 15000 7679 15034 7713
rect 15068 7679 15102 7713
rect 68 7608 102 7642
rect 137 7608 171 7642
rect 206 7608 240 7642
rect 275 7608 309 7642
rect 344 7608 378 7642
rect 413 7608 447 7642
rect 482 7608 516 7642
rect 551 7608 585 7642
rect 620 7608 654 7642
rect 689 7608 723 7642
rect 758 7608 792 7642
rect 827 7608 861 7642
rect 896 7608 930 7642
rect 965 7608 999 7642
rect 1033 7608 1067 7642
rect 1101 7608 1135 7642
rect 1169 7608 1203 7642
rect 1237 7608 1271 7642
rect 1305 7608 1339 7642
rect 1373 7608 1407 7642
rect 1441 7608 1475 7642
rect 1509 7608 1543 7642
rect 1577 7608 1611 7642
rect 1645 7608 1679 7642
rect 1713 7608 1747 7642
rect 1781 7608 1815 7642
rect 1849 7608 1883 7642
rect 1917 7608 1951 7642
rect 1985 7608 2019 7642
rect 2053 7608 2087 7642
rect 2121 7608 2155 7642
rect 2189 7608 2223 7642
rect 2257 7608 2291 7642
rect 2325 7608 2359 7642
rect 2393 7608 2427 7642
rect 2461 7608 2495 7642
rect 2529 7608 2563 7642
rect 2597 7608 2631 7642
rect 2665 7608 2699 7642
rect 68 7536 102 7570
rect 137 7536 171 7570
rect 206 7536 240 7570
rect 275 7536 309 7570
rect 344 7536 378 7570
rect 413 7536 447 7570
rect 482 7536 516 7570
rect 551 7536 585 7570
rect 620 7536 654 7570
rect 689 7536 723 7570
rect 758 7536 792 7570
rect 827 7536 861 7570
rect 896 7536 930 7570
rect 965 7536 999 7570
rect 1033 7536 1067 7570
rect 1101 7536 1135 7570
rect 1169 7536 1203 7570
rect 1237 7536 1271 7570
rect 1305 7536 1339 7570
rect 1373 7536 1407 7570
rect 1441 7536 1475 7570
rect 1509 7536 1543 7570
rect 1577 7536 1611 7570
rect 1645 7536 1679 7570
rect 1713 7536 1747 7570
rect 1781 7536 1815 7570
rect 1849 7536 1883 7570
rect 1917 7536 1951 7570
rect 1985 7536 2019 7570
rect 2053 7536 2087 7570
rect 2121 7536 2155 7570
rect 2189 7536 2223 7570
rect 2257 7536 2291 7570
rect 2325 7536 2359 7570
rect 2393 7536 2427 7570
rect 2461 7536 2495 7570
rect 2529 7536 2563 7570
rect 2597 7536 2631 7570
rect 2665 7536 2699 7570
rect 68 7464 102 7498
rect 137 7464 171 7498
rect 206 7464 240 7498
rect 275 7464 309 7498
rect 344 7464 378 7498
rect 413 7464 447 7498
rect 482 7464 516 7498
rect 551 7464 585 7498
rect 620 7464 654 7498
rect 689 7464 723 7498
rect 758 7464 792 7498
rect 827 7464 861 7498
rect 896 7464 930 7498
rect 965 7464 999 7498
rect 1033 7464 1067 7498
rect 1101 7464 1135 7498
rect 1169 7464 1203 7498
rect 1237 7464 1271 7498
rect 1305 7464 1339 7498
rect 1373 7464 1407 7498
rect 1441 7464 1475 7498
rect 1509 7464 1543 7498
rect 1577 7464 1611 7498
rect 1645 7464 1679 7498
rect 1713 7464 1747 7498
rect 1781 7464 1815 7498
rect 1849 7464 1883 7498
rect 1917 7464 1951 7498
rect 1985 7464 2019 7498
rect 2053 7464 2087 7498
rect 2121 7464 2155 7498
rect 2189 7464 2223 7498
rect 2257 7464 2291 7498
rect 2325 7464 2359 7498
rect 2393 7464 2427 7498
rect 2461 7464 2495 7498
rect 2529 7464 2563 7498
rect 2597 7464 2631 7498
rect 2665 7464 2699 7498
rect 68 7392 102 7426
rect 137 7392 171 7426
rect 206 7392 240 7426
rect 275 7392 309 7426
rect 344 7392 378 7426
rect 413 7392 447 7426
rect 482 7392 516 7426
rect 551 7392 585 7426
rect 620 7392 654 7426
rect 689 7392 723 7426
rect 758 7392 792 7426
rect 827 7392 861 7426
rect 896 7392 930 7426
rect 965 7392 999 7426
rect 1033 7392 1067 7426
rect 1101 7392 1135 7426
rect 1169 7392 1203 7426
rect 1237 7392 1271 7426
rect 1305 7392 1339 7426
rect 1373 7392 1407 7426
rect 1441 7392 1475 7426
rect 1509 7392 1543 7426
rect 1577 7392 1611 7426
rect 1645 7392 1679 7426
rect 1713 7392 1747 7426
rect 1781 7392 1815 7426
rect 1849 7392 1883 7426
rect 1917 7392 1951 7426
rect 1985 7392 2019 7426
rect 2053 7392 2087 7426
rect 2121 7392 2155 7426
rect 2189 7392 2223 7426
rect 2257 7392 2291 7426
rect 2325 7392 2359 7426
rect 2393 7392 2427 7426
rect 2461 7392 2495 7426
rect 2529 7392 2563 7426
rect 2597 7392 2631 7426
rect 2665 7392 2699 7426
rect 68 7320 102 7354
rect 137 7320 171 7354
rect 206 7320 240 7354
rect 275 7320 309 7354
rect 344 7320 378 7354
rect 413 7320 447 7354
rect 482 7320 516 7354
rect 551 7320 585 7354
rect 620 7320 654 7354
rect 689 7320 723 7354
rect 758 7320 792 7354
rect 827 7320 861 7354
rect 896 7320 930 7354
rect 965 7320 999 7354
rect 1033 7320 1067 7354
rect 1101 7320 1135 7354
rect 1169 7320 1203 7354
rect 1237 7320 1271 7354
rect 1305 7320 1339 7354
rect 1373 7320 1407 7354
rect 1441 7320 1475 7354
rect 1509 7320 1543 7354
rect 1577 7320 1611 7354
rect 1645 7320 1679 7354
rect 1713 7320 1747 7354
rect 1781 7320 1815 7354
rect 1849 7320 1883 7354
rect 1917 7320 1951 7354
rect 1985 7320 2019 7354
rect 2053 7320 2087 7354
rect 2121 7320 2155 7354
rect 2189 7320 2223 7354
rect 2257 7320 2291 7354
rect 2325 7320 2359 7354
rect 2393 7320 2427 7354
rect 2461 7320 2495 7354
rect 2529 7320 2563 7354
rect 2597 7320 2631 7354
rect 2665 7320 2699 7354
rect 12524 7606 12558 7640
rect 12593 7606 12627 7640
rect 12662 7606 12696 7640
rect 12731 7606 12765 7640
rect 12800 7606 12834 7640
rect 12869 7606 12903 7640
rect 12938 7606 12972 7640
rect 13007 7606 13041 7640
rect 13076 7606 13110 7640
rect 13145 7606 13179 7640
rect 13214 7606 13248 7640
rect 13283 7606 13317 7640
rect 13352 7606 13386 7640
rect 13421 7606 13455 7640
rect 13490 7606 13524 7640
rect 13559 7606 13593 7640
rect 13628 7606 13662 7640
rect 13697 7606 13731 7640
rect 13766 7606 13800 7640
rect 13835 7606 13869 7640
rect 13904 7606 13938 7640
rect 13973 7606 14007 7640
rect 14042 7606 14076 7640
rect 14111 7606 14145 7640
rect 14180 7606 14214 7640
rect 14249 7606 14283 7640
rect 14318 7606 14352 7640
rect 14387 7606 14421 7640
rect 14456 7606 14490 7640
rect 14524 7606 14558 7640
rect 14592 7606 14626 7640
rect 14660 7606 14694 7640
rect 14728 7606 14762 7640
rect 14796 7606 14830 7640
rect 14864 7606 14898 7640
rect 14932 7607 14966 7641
rect 15000 7607 15034 7641
rect 15068 7607 15102 7641
rect 12524 7522 12558 7556
rect 12593 7522 12627 7556
rect 12662 7522 12696 7556
rect 12731 7522 12765 7556
rect 12800 7522 12834 7556
rect 12869 7522 12903 7556
rect 12938 7522 12972 7556
rect 13007 7522 13041 7556
rect 13076 7522 13110 7556
rect 13145 7522 13179 7556
rect 13214 7522 13248 7556
rect 13283 7522 13317 7556
rect 13352 7522 13386 7556
rect 13421 7522 13455 7556
rect 13490 7522 13524 7556
rect 13559 7522 13593 7556
rect 13628 7522 13662 7556
rect 13697 7522 13731 7556
rect 13766 7522 13800 7556
rect 13835 7522 13869 7556
rect 13904 7522 13938 7556
rect 13973 7522 14007 7556
rect 14042 7522 14076 7556
rect 14111 7522 14145 7556
rect 14180 7522 14214 7556
rect 14249 7522 14283 7556
rect 14318 7522 14352 7556
rect 14387 7522 14421 7556
rect 14456 7522 14490 7556
rect 14524 7522 14558 7556
rect 14592 7522 14626 7556
rect 14660 7522 14694 7556
rect 14728 7522 14762 7556
rect 14796 7522 14830 7556
rect 14864 7522 14898 7556
rect 14932 7535 14966 7569
rect 15000 7535 15034 7569
rect 15068 7535 15102 7569
rect 12524 7438 12558 7472
rect 12593 7438 12627 7472
rect 12662 7438 12696 7472
rect 12731 7438 12765 7472
rect 12800 7438 12834 7472
rect 12869 7438 12903 7472
rect 12938 7438 12972 7472
rect 13007 7438 13041 7472
rect 13076 7438 13110 7472
rect 13145 7438 13179 7472
rect 13214 7438 13248 7472
rect 13283 7438 13317 7472
rect 13352 7438 13386 7472
rect 13421 7438 13455 7472
rect 13490 7438 13524 7472
rect 13559 7438 13593 7472
rect 13628 7438 13662 7472
rect 13697 7438 13731 7472
rect 13766 7438 13800 7472
rect 13835 7438 13869 7472
rect 13904 7438 13938 7472
rect 13973 7438 14007 7472
rect 14042 7438 14076 7472
rect 14111 7438 14145 7472
rect 14180 7438 14214 7472
rect 14249 7438 14283 7472
rect 14318 7438 14352 7472
rect 14387 7438 14421 7472
rect 14456 7438 14490 7472
rect 14524 7438 14558 7472
rect 14592 7438 14626 7472
rect 14660 7438 14694 7472
rect 14728 7438 14762 7472
rect 14796 7438 14830 7472
rect 14864 7438 14898 7472
rect 14932 7463 14966 7497
rect 15000 7463 15034 7497
rect 15068 7463 15102 7497
rect 14932 7391 14966 7425
rect 15000 7391 15034 7425
rect 15068 7391 15102 7425
rect 12524 7354 12558 7388
rect 12593 7354 12627 7388
rect 12662 7354 12696 7388
rect 12731 7354 12765 7388
rect 12800 7354 12834 7388
rect 12869 7354 12903 7388
rect 12938 7354 12972 7388
rect 13007 7354 13041 7388
rect 13076 7354 13110 7388
rect 13145 7354 13179 7388
rect 13214 7354 13248 7388
rect 13283 7354 13317 7388
rect 13352 7354 13386 7388
rect 13421 7354 13455 7388
rect 13490 7354 13524 7388
rect 13559 7354 13593 7388
rect 13628 7354 13662 7388
rect 13697 7354 13731 7388
rect 13766 7354 13800 7388
rect 13835 7354 13869 7388
rect 13904 7354 13938 7388
rect 13973 7354 14007 7388
rect 14042 7354 14076 7388
rect 14111 7354 14145 7388
rect 14180 7354 14214 7388
rect 14249 7354 14283 7388
rect 14318 7354 14352 7388
rect 14387 7354 14421 7388
rect 14456 7354 14490 7388
rect 14524 7354 14558 7388
rect 14592 7354 14626 7388
rect 14660 7354 14694 7388
rect 14728 7354 14762 7388
rect 14796 7354 14830 7388
rect 14864 7354 14898 7388
rect 14932 7319 14966 7353
rect 15000 7319 15034 7353
rect 15068 7319 15102 7353
rect 68 7248 102 7282
rect 137 7248 171 7282
rect 206 7248 240 7282
rect 275 7248 309 7282
rect 344 7248 378 7282
rect 413 7248 447 7282
rect 482 7248 516 7282
rect 551 7248 585 7282
rect 620 7248 654 7282
rect 689 7248 723 7282
rect 758 7248 792 7282
rect 827 7248 861 7282
rect 896 7248 930 7282
rect 965 7248 999 7282
rect 1033 7248 1067 7282
rect 1101 7248 1135 7282
rect 1169 7248 1203 7282
rect 1237 7248 1271 7282
rect 1305 7248 1339 7282
rect 1373 7248 1407 7282
rect 1441 7248 1475 7282
rect 1509 7248 1543 7282
rect 1577 7248 1611 7282
rect 1645 7248 1679 7282
rect 1713 7248 1747 7282
rect 1781 7248 1815 7282
rect 1849 7248 1883 7282
rect 1917 7248 1951 7282
rect 1985 7248 2019 7282
rect 2053 7248 2087 7282
rect 2121 7248 2155 7282
rect 2189 7248 2223 7282
rect 2257 7248 2291 7282
rect 2325 7248 2359 7282
rect 2393 7248 2427 7282
rect 2461 7248 2495 7282
rect 2529 7248 2563 7282
rect 2597 7248 2631 7282
rect 2665 7248 2699 7282
rect 68 7176 102 7210
rect 137 7176 171 7210
rect 206 7176 240 7210
rect 275 7176 309 7210
rect 344 7176 378 7210
rect 413 7176 447 7210
rect 482 7176 516 7210
rect 551 7176 585 7210
rect 620 7176 654 7210
rect 689 7176 723 7210
rect 758 7176 792 7210
rect 827 7176 861 7210
rect 896 7176 930 7210
rect 965 7176 999 7210
rect 1033 7176 1067 7210
rect 1101 7176 1135 7210
rect 1169 7176 1203 7210
rect 1237 7176 1271 7210
rect 1305 7176 1339 7210
rect 1373 7176 1407 7210
rect 1441 7176 1475 7210
rect 1509 7176 1543 7210
rect 1577 7176 1611 7210
rect 1645 7176 1679 7210
rect 1713 7176 1747 7210
rect 1781 7176 1815 7210
rect 1849 7176 1883 7210
rect 1917 7176 1951 7210
rect 1985 7176 2019 7210
rect 2053 7176 2087 7210
rect 2121 7176 2155 7210
rect 2189 7176 2223 7210
rect 2257 7176 2291 7210
rect 2325 7176 2359 7210
rect 2393 7176 2427 7210
rect 2461 7176 2495 7210
rect 2529 7176 2563 7210
rect 2597 7176 2631 7210
rect 2665 7176 2699 7210
rect 68 7104 102 7138
rect 137 7104 171 7138
rect 206 7104 240 7138
rect 275 7104 309 7138
rect 344 7104 378 7138
rect 413 7104 447 7138
rect 482 7104 516 7138
rect 551 7104 585 7138
rect 620 7104 654 7138
rect 689 7104 723 7138
rect 758 7104 792 7138
rect 827 7104 861 7138
rect 896 7104 930 7138
rect 965 7104 999 7138
rect 1033 7104 1067 7138
rect 1101 7104 1135 7138
rect 1169 7104 1203 7138
rect 1237 7104 1271 7138
rect 1305 7104 1339 7138
rect 1373 7104 1407 7138
rect 1441 7104 1475 7138
rect 1509 7104 1543 7138
rect 1577 7104 1611 7138
rect 1645 7104 1679 7138
rect 1713 7104 1747 7138
rect 1781 7104 1815 7138
rect 1849 7104 1883 7138
rect 1917 7104 1951 7138
rect 1985 7104 2019 7138
rect 2053 7104 2087 7138
rect 2121 7104 2155 7138
rect 2189 7104 2223 7138
rect 2257 7104 2291 7138
rect 2325 7104 2359 7138
rect 2393 7104 2427 7138
rect 2461 7104 2495 7138
rect 2529 7104 2563 7138
rect 2597 7104 2631 7138
rect 2665 7104 2699 7138
rect 68 7032 102 7066
rect 137 7032 171 7066
rect 206 7032 240 7066
rect 275 7032 309 7066
rect 344 7032 378 7066
rect 413 7032 447 7066
rect 482 7032 516 7066
rect 551 7032 585 7066
rect 620 7032 654 7066
rect 689 7032 723 7066
rect 758 7032 792 7066
rect 827 7032 861 7066
rect 896 7032 930 7066
rect 965 7032 999 7066
rect 1033 7032 1067 7066
rect 1101 7032 1135 7066
rect 1169 7032 1203 7066
rect 1237 7032 1271 7066
rect 1305 7032 1339 7066
rect 1373 7032 1407 7066
rect 1441 7032 1475 7066
rect 1509 7032 1543 7066
rect 1577 7032 1611 7066
rect 1645 7032 1679 7066
rect 1713 7032 1747 7066
rect 1781 7032 1815 7066
rect 1849 7032 1883 7066
rect 1917 7032 1951 7066
rect 1985 7032 2019 7066
rect 2053 7032 2087 7066
rect 2121 7032 2155 7066
rect 2189 7032 2223 7066
rect 2257 7032 2291 7066
rect 2325 7032 2359 7066
rect 2393 7032 2427 7066
rect 2461 7032 2495 7066
rect 2529 7032 2563 7066
rect 2597 7032 2631 7066
rect 2665 7032 2699 7066
rect 8210 7248 8244 7282
rect 8279 7248 8313 7282
rect 8348 7248 8382 7282
rect 8417 7248 8451 7282
rect 8486 7248 8520 7282
rect 8555 7248 8589 7282
rect 8624 7248 8658 7282
rect 8693 7248 8727 7282
rect 8762 7248 8796 7282
rect 8831 7248 8865 7282
rect 8900 7248 8934 7282
rect 8969 7248 9003 7282
rect 9038 7248 9072 7282
rect 9107 7248 9141 7282
rect 9176 7248 9210 7282
rect 9245 7248 9279 7282
rect 9314 7248 9348 7282
rect 9383 7248 9417 7282
rect 9452 7248 9486 7282
rect 9521 7248 9555 7282
rect 9590 7248 9624 7282
rect 9659 7248 9693 7282
rect 9728 7248 9762 7282
rect 9797 7248 9831 7282
rect 9866 7248 9900 7282
rect 9935 7248 9969 7282
rect 10004 7248 10038 7282
rect 10073 7248 10107 7282
rect 10142 7248 10176 7282
rect 10211 7248 10245 7282
rect 10280 7248 10314 7282
rect 10349 7248 10383 7282
rect 10418 7248 10452 7282
rect 10487 7248 10521 7282
rect 10556 7248 10590 7282
rect 10625 7248 10659 7282
rect 10694 7248 10728 7282
rect 10763 7248 10797 7282
rect 10832 7248 10866 7282
rect 10901 7248 10935 7282
rect 10970 7248 11004 7282
rect 11039 7248 11073 7282
rect 11108 7248 11142 7282
rect 11177 7248 11211 7282
rect 11246 7248 11280 7282
rect 11315 7248 11349 7282
rect 11384 7248 11418 7282
rect 11453 7248 11487 7282
rect 11522 7248 11556 7282
rect 11591 7248 11625 7282
rect 11660 7248 11694 7282
rect 11729 7248 11763 7282
rect 11798 7248 11832 7282
rect 11867 7248 11901 7282
rect 11936 7248 11970 7282
rect 12005 7248 12039 7282
rect 12074 7248 12108 7282
rect 12143 7248 12177 7282
rect 12212 7248 12246 7282
rect 12280 7248 12314 7282
rect 12348 7248 12382 7282
rect 12416 7248 12450 7282
rect 12484 7248 12518 7282
rect 12552 7248 12586 7282
rect 12620 7248 12654 7282
rect 12688 7248 12722 7282
rect 12756 7248 12790 7282
rect 12824 7248 12858 7282
rect 12892 7248 12926 7282
rect 12960 7248 12994 7282
rect 13028 7248 13062 7282
rect 13096 7248 13130 7282
rect 13164 7248 13198 7282
rect 13232 7248 13266 7282
rect 13300 7248 13334 7282
rect 13368 7248 13402 7282
rect 13436 7248 13470 7282
rect 13504 7248 13538 7282
rect 13572 7248 13606 7282
rect 13640 7248 13674 7282
rect 13708 7248 13742 7282
rect 13776 7248 13810 7282
rect 13844 7248 13878 7282
rect 13912 7248 13946 7282
rect 13980 7248 14014 7282
rect 14048 7248 14082 7282
rect 14116 7248 14150 7282
rect 14184 7248 14218 7282
rect 14252 7248 14286 7282
rect 14320 7248 14354 7282
rect 14388 7248 14422 7282
rect 14456 7248 14490 7282
rect 14524 7248 14558 7282
rect 14592 7248 14626 7282
rect 14660 7248 14694 7282
rect 14728 7248 14762 7282
rect 14796 7248 14830 7282
rect 14864 7248 14898 7282
rect 14932 7247 14966 7281
rect 15000 7247 15034 7281
rect 15068 7247 15102 7281
rect 8210 7176 8244 7210
rect 8279 7176 8313 7210
rect 8348 7176 8382 7210
rect 8417 7176 8451 7210
rect 8486 7176 8520 7210
rect 8555 7176 8589 7210
rect 8624 7176 8658 7210
rect 8693 7176 8727 7210
rect 8762 7176 8796 7210
rect 8831 7176 8865 7210
rect 8900 7176 8934 7210
rect 8969 7176 9003 7210
rect 9038 7176 9072 7210
rect 9107 7176 9141 7210
rect 9176 7176 9210 7210
rect 9245 7176 9279 7210
rect 9314 7176 9348 7210
rect 9383 7176 9417 7210
rect 9452 7176 9486 7210
rect 9521 7176 9555 7210
rect 9590 7176 9624 7210
rect 9659 7176 9693 7210
rect 9728 7176 9762 7210
rect 9797 7176 9831 7210
rect 9866 7176 9900 7210
rect 9935 7176 9969 7210
rect 10004 7176 10038 7210
rect 10073 7176 10107 7210
rect 10142 7176 10176 7210
rect 10211 7176 10245 7210
rect 10280 7176 10314 7210
rect 10349 7176 10383 7210
rect 10418 7176 10452 7210
rect 10487 7176 10521 7210
rect 10556 7176 10590 7210
rect 10625 7176 10659 7210
rect 10694 7176 10728 7210
rect 10763 7176 10797 7210
rect 10832 7176 10866 7210
rect 10901 7176 10935 7210
rect 10970 7176 11004 7210
rect 11039 7176 11073 7210
rect 11108 7176 11142 7210
rect 11177 7176 11211 7210
rect 11246 7176 11280 7210
rect 11315 7176 11349 7210
rect 11384 7176 11418 7210
rect 11453 7176 11487 7210
rect 11522 7176 11556 7210
rect 11591 7176 11625 7210
rect 11660 7176 11694 7210
rect 11729 7176 11763 7210
rect 11798 7176 11832 7210
rect 11867 7176 11901 7210
rect 11936 7176 11970 7210
rect 12005 7176 12039 7210
rect 12074 7176 12108 7210
rect 12143 7176 12177 7210
rect 12212 7176 12246 7210
rect 12280 7176 12314 7210
rect 12348 7176 12382 7210
rect 12416 7176 12450 7210
rect 12484 7176 12518 7210
rect 12552 7176 12586 7210
rect 12620 7176 12654 7210
rect 12688 7176 12722 7210
rect 12756 7176 12790 7210
rect 12824 7176 12858 7210
rect 12892 7176 12926 7210
rect 12960 7176 12994 7210
rect 13028 7176 13062 7210
rect 13096 7176 13130 7210
rect 13164 7176 13198 7210
rect 13232 7176 13266 7210
rect 13300 7176 13334 7210
rect 13368 7176 13402 7210
rect 13436 7176 13470 7210
rect 13504 7176 13538 7210
rect 13572 7176 13606 7210
rect 13640 7176 13674 7210
rect 13708 7176 13742 7210
rect 13776 7176 13810 7210
rect 13844 7176 13878 7210
rect 13912 7176 13946 7210
rect 13980 7176 14014 7210
rect 14048 7176 14082 7210
rect 14116 7176 14150 7210
rect 14184 7176 14218 7210
rect 14252 7176 14286 7210
rect 14320 7176 14354 7210
rect 14388 7176 14422 7210
rect 14456 7176 14490 7210
rect 14524 7176 14558 7210
rect 14592 7176 14626 7210
rect 14660 7176 14694 7210
rect 14728 7176 14762 7210
rect 14796 7176 14830 7210
rect 14864 7176 14898 7210
rect 14932 7175 14966 7209
rect 15000 7175 15034 7209
rect 15068 7175 15102 7209
rect 8210 7104 8244 7138
rect 8279 7104 8313 7138
rect 8348 7104 8382 7138
rect 8417 7104 8451 7138
rect 8486 7104 8520 7138
rect 8555 7104 8589 7138
rect 8624 7104 8658 7138
rect 8693 7104 8727 7138
rect 8762 7104 8796 7138
rect 8831 7104 8865 7138
rect 8900 7104 8934 7138
rect 8969 7104 9003 7138
rect 9038 7104 9072 7138
rect 9107 7104 9141 7138
rect 9176 7104 9210 7138
rect 9245 7104 9279 7138
rect 9314 7104 9348 7138
rect 9383 7104 9417 7138
rect 9452 7104 9486 7138
rect 9521 7104 9555 7138
rect 9590 7104 9624 7138
rect 9659 7104 9693 7138
rect 9728 7104 9762 7138
rect 9797 7104 9831 7138
rect 9866 7104 9900 7138
rect 9935 7104 9969 7138
rect 10004 7104 10038 7138
rect 10073 7104 10107 7138
rect 10142 7104 10176 7138
rect 10211 7104 10245 7138
rect 10280 7104 10314 7138
rect 10349 7104 10383 7138
rect 10418 7104 10452 7138
rect 10487 7104 10521 7138
rect 10556 7104 10590 7138
rect 10625 7104 10659 7138
rect 10694 7104 10728 7138
rect 10763 7104 10797 7138
rect 10832 7104 10866 7138
rect 10901 7104 10935 7138
rect 10970 7104 11004 7138
rect 11039 7104 11073 7138
rect 11108 7104 11142 7138
rect 11177 7104 11211 7138
rect 11246 7104 11280 7138
rect 11315 7104 11349 7138
rect 11384 7104 11418 7138
rect 11453 7104 11487 7138
rect 11522 7104 11556 7138
rect 11591 7104 11625 7138
rect 11660 7104 11694 7138
rect 11729 7104 11763 7138
rect 11798 7104 11832 7138
rect 11867 7104 11901 7138
rect 11936 7104 11970 7138
rect 12005 7104 12039 7138
rect 12074 7104 12108 7138
rect 12143 7104 12177 7138
rect 12212 7104 12246 7138
rect 12280 7104 12314 7138
rect 12348 7104 12382 7138
rect 12416 7104 12450 7138
rect 12484 7104 12518 7138
rect 12552 7104 12586 7138
rect 12620 7104 12654 7138
rect 12688 7104 12722 7138
rect 12756 7104 12790 7138
rect 12824 7104 12858 7138
rect 12892 7104 12926 7138
rect 12960 7104 12994 7138
rect 13028 7104 13062 7138
rect 13096 7104 13130 7138
rect 13164 7104 13198 7138
rect 13232 7104 13266 7138
rect 13300 7104 13334 7138
rect 13368 7104 13402 7138
rect 13436 7104 13470 7138
rect 13504 7104 13538 7138
rect 13572 7104 13606 7138
rect 13640 7104 13674 7138
rect 13708 7104 13742 7138
rect 13776 7104 13810 7138
rect 13844 7104 13878 7138
rect 13912 7104 13946 7138
rect 13980 7104 14014 7138
rect 14048 7104 14082 7138
rect 14116 7104 14150 7138
rect 14184 7104 14218 7138
rect 14252 7104 14286 7138
rect 14320 7104 14354 7138
rect 14388 7104 14422 7138
rect 14456 7104 14490 7138
rect 14524 7104 14558 7138
rect 14592 7104 14626 7138
rect 14660 7104 14694 7138
rect 14728 7104 14762 7138
rect 14796 7104 14830 7138
rect 14864 7104 14898 7138
rect 14932 7103 14966 7137
rect 15000 7103 15034 7137
rect 15068 7103 15102 7137
rect 2757 7013 2791 7047
rect 2825 7013 2859 7047
rect 2893 7013 2927 7047
rect 2961 7013 2995 7047
rect 3029 7013 3063 7047
rect 3097 7013 3131 7047
rect 3165 7013 3199 7047
rect 3233 7013 3267 7047
rect 3301 7013 3335 7047
rect 3369 7013 3403 7047
rect 3437 7013 3471 7047
rect 3505 7013 3539 7047
rect 3573 7013 3607 7047
rect 3641 7013 3675 7047
rect 3709 7013 3743 7047
rect 3777 7013 3811 7047
rect 3845 7013 3879 7047
rect 3913 7013 3947 7047
rect 3981 7013 4015 7047
rect 4049 7013 4083 7047
rect 4117 7013 4151 7047
rect 4185 7013 4219 7047
rect 4253 7013 4287 7047
rect 4321 7013 4355 7047
rect 4389 7013 4423 7047
rect 4457 7013 4491 7047
rect 4525 7013 4559 7047
rect 4593 7013 4627 7047
rect 4661 7013 4695 7047
rect 4729 7013 4763 7047
rect 4797 7013 4831 7047
rect 4865 7013 4899 7047
rect 4933 7013 4967 7047
rect 5001 7013 5035 7047
rect 5069 7013 5103 7047
rect 5137 7013 5171 7047
rect 5205 7013 5239 7047
rect 5273 7013 5307 7047
rect 5341 7013 5375 7047
rect 5409 7013 5443 7047
rect 5477 7013 5511 7047
rect 5545 7013 5579 7047
rect 5613 7013 5647 7047
rect 5681 7013 5715 7047
rect 5749 7013 5783 7047
rect 5817 7013 5851 7047
rect 5885 7013 5919 7047
rect 5953 7013 5987 7047
rect 6021 7013 6055 7047
rect 6089 7013 6123 7047
rect 6157 7013 6191 7047
rect 6225 7013 6259 7047
rect 6293 7013 6327 7047
rect 6361 7013 6395 7047
rect 6429 7013 6463 7047
rect 6497 7013 6531 7047
rect 6565 7013 6599 7047
rect 6633 7013 6667 7047
rect 6701 7013 6735 7047
rect 6769 7013 6803 7047
rect 6837 7013 6871 7047
rect 6905 7013 6939 7047
rect 6973 7013 7007 7047
rect 7041 7013 7075 7047
rect 7109 7013 7143 7047
rect 7177 7013 7211 7047
rect 7245 7013 7279 7047
rect 7313 7013 7347 7047
rect 7381 7013 7415 7047
rect 7449 7013 7483 7047
rect 7517 7013 7551 7047
rect 7585 7013 7619 7047
rect 7653 7013 7687 7047
rect 8210 7032 8244 7066
rect 8279 7032 8313 7066
rect 8348 7032 8382 7066
rect 8417 7032 8451 7066
rect 8486 7032 8520 7066
rect 8555 7032 8589 7066
rect 8624 7032 8658 7066
rect 8693 7032 8727 7066
rect 8762 7032 8796 7066
rect 8831 7032 8865 7066
rect 8900 7032 8934 7066
rect 8969 7032 9003 7066
rect 9038 7032 9072 7066
rect 9107 7032 9141 7066
rect 9176 7032 9210 7066
rect 9245 7032 9279 7066
rect 9314 7032 9348 7066
rect 9383 7032 9417 7066
rect 9452 7032 9486 7066
rect 9521 7032 9555 7066
rect 9590 7032 9624 7066
rect 9659 7032 9693 7066
rect 9728 7032 9762 7066
rect 9797 7032 9831 7066
rect 9866 7032 9900 7066
rect 9935 7032 9969 7066
rect 10004 7032 10038 7066
rect 10073 7032 10107 7066
rect 10142 7032 10176 7066
rect 10211 7032 10245 7066
rect 10280 7032 10314 7066
rect 10349 7032 10383 7066
rect 10418 7032 10452 7066
rect 10487 7032 10521 7066
rect 10556 7032 10590 7066
rect 10625 7032 10659 7066
rect 10694 7032 10728 7066
rect 10763 7032 10797 7066
rect 10832 7032 10866 7066
rect 10901 7032 10935 7066
rect 10970 7032 11004 7066
rect 11039 7032 11073 7066
rect 11108 7032 11142 7066
rect 11177 7032 11211 7066
rect 11246 7032 11280 7066
rect 11315 7032 11349 7066
rect 11384 7032 11418 7066
rect 11453 7032 11487 7066
rect 11522 7032 11556 7066
rect 11591 7032 11625 7066
rect 11660 7032 11694 7066
rect 11729 7032 11763 7066
rect 11798 7032 11832 7066
rect 11867 7032 11901 7066
rect 11936 7032 11970 7066
rect 12005 7032 12039 7066
rect 12074 7032 12108 7066
rect 12143 7032 12177 7066
rect 12212 7032 12246 7066
rect 12280 7032 12314 7066
rect 12348 7032 12382 7066
rect 12416 7032 12450 7066
rect 12484 7032 12518 7066
rect 12552 7032 12586 7066
rect 12620 7032 12654 7066
rect 12688 7032 12722 7066
rect 12756 7032 12790 7066
rect 12824 7032 12858 7066
rect 12892 7032 12926 7066
rect 12960 7032 12994 7066
rect 13028 7032 13062 7066
rect 13096 7032 13130 7066
rect 13164 7032 13198 7066
rect 13232 7032 13266 7066
rect 13300 7032 13334 7066
rect 13368 7032 13402 7066
rect 13436 7032 13470 7066
rect 13504 7032 13538 7066
rect 13572 7032 13606 7066
rect 13640 7032 13674 7066
rect 13708 7032 13742 7066
rect 13776 7032 13810 7066
rect 13844 7032 13878 7066
rect 13912 7032 13946 7066
rect 13980 7032 14014 7066
rect 14048 7032 14082 7066
rect 14116 7032 14150 7066
rect 14184 7032 14218 7066
rect 14252 7032 14286 7066
rect 14320 7032 14354 7066
rect 14388 7032 14422 7066
rect 14456 7032 14490 7066
rect 14524 7032 14558 7066
rect 14592 7032 14626 7066
rect 14660 7032 14694 7066
rect 14728 7032 14762 7066
rect 14796 7032 14830 7066
rect 14864 7032 14898 7066
rect 14932 7031 14966 7065
rect 15000 7031 15034 7065
rect 15068 7031 15102 7065
<< poly >>
rect 8490 8239 8612 8286
rect 8490 7933 8510 8239
rect 8490 7886 8612 7933
rect 9612 8239 9714 8286
rect 9612 7886 9714 7933
rect 10314 8239 10416 8286
rect 10314 7886 10416 7933
rect 10816 8239 10934 8286
rect 10918 7933 10934 8239
rect 10816 7886 10934 7933
<< polycont >>
rect 8510 7933 8612 8239
rect 9612 7933 9714 8239
rect 10314 7933 10416 8239
rect 10816 7933 10918 8239
<< npolyres >>
rect 8612 7886 9612 8286
rect 9714 7886 10314 8286
rect 10416 7886 10816 8286
<< locali >>
rect 12580 15655 12636 15661
rect 14376 15655 14416 15661
rect 12580 15651 14416 15655
rect 12580 15617 12660 15651
rect 12694 15617 12730 15651
rect 12764 15617 12800 15651
rect 12834 15617 12869 15651
rect 12903 15617 12938 15651
rect 12972 15617 13007 15651
rect 13041 15617 13076 15651
rect 13110 15617 13145 15651
rect 13179 15617 13214 15651
rect 13248 15617 13283 15651
rect 13317 15617 13352 15651
rect 13386 15617 13421 15651
rect 13455 15617 13490 15651
rect 13524 15617 13559 15651
rect 13593 15617 13628 15651
rect 13662 15617 13697 15651
rect 13731 15617 13766 15651
rect 13800 15617 13835 15651
rect 13869 15617 13904 15651
rect 13938 15617 13973 15651
rect 14007 15617 14042 15651
rect 14076 15617 14111 15651
rect 14145 15617 14180 15651
rect 14214 15617 14249 15651
rect 14283 15617 14318 15651
rect 14352 15617 14416 15651
rect 12580 15581 14416 15617
rect 12580 15547 12660 15581
rect 12694 15547 12730 15581
rect 12764 15547 12800 15581
rect 12834 15547 12869 15581
rect 12903 15547 12938 15581
rect 12972 15547 13007 15581
rect 13041 15547 13076 15581
rect 13110 15547 13145 15581
rect 13179 15547 13214 15581
rect 13248 15547 13283 15581
rect 13317 15547 13352 15581
rect 13386 15547 13421 15581
rect 13455 15547 13490 15581
rect 13524 15547 13559 15581
rect 13593 15547 13628 15581
rect 13662 15547 13697 15581
rect 13731 15547 13766 15581
rect 13800 15547 13835 15581
rect 13869 15547 13904 15581
rect 13938 15547 13973 15581
rect 14007 15547 14042 15581
rect 14076 15547 14111 15581
rect 14145 15547 14180 15581
rect 14214 15547 14249 15581
rect 14283 15547 14318 15581
rect 14352 15547 14416 15581
rect 12580 15511 14416 15547
rect 12580 15477 12660 15511
rect 12694 15477 12730 15511
rect 12764 15477 12800 15511
rect 12834 15477 12869 15511
rect 12903 15477 12938 15511
rect 12972 15477 13007 15511
rect 13041 15477 13076 15511
rect 13110 15477 13145 15511
rect 13179 15477 13214 15511
rect 13248 15477 13283 15511
rect 13317 15477 13352 15511
rect 13386 15477 13421 15511
rect 13455 15477 13490 15511
rect 13524 15477 13559 15511
rect 13593 15477 13628 15511
rect 13662 15477 13697 15511
rect 13731 15477 13766 15511
rect 13800 15477 13835 15511
rect 13869 15477 13904 15511
rect 13938 15477 13973 15511
rect 14007 15477 14042 15511
rect 14076 15477 14111 15511
rect 14145 15477 14180 15511
rect 14214 15477 14249 15511
rect 14283 15477 14318 15511
rect 14352 15477 14416 15511
rect 12580 15441 14416 15477
rect 12580 15407 12660 15441
rect 12694 15407 12730 15441
rect 12764 15407 12800 15441
rect 12834 15407 12869 15441
rect 12903 15407 12938 15441
rect 12972 15407 13007 15441
rect 13041 15407 13076 15441
rect 13110 15407 13145 15441
rect 13179 15407 13214 15441
rect 13248 15407 13283 15441
rect 13317 15407 13352 15441
rect 13386 15407 13421 15441
rect 13455 15407 13490 15441
rect 13524 15407 13559 15441
rect 13593 15407 13628 15441
rect 13662 15407 13697 15441
rect 13731 15407 13766 15441
rect 13800 15407 13835 15441
rect 13869 15407 13904 15441
rect 13938 15407 13973 15441
rect 14007 15407 14042 15441
rect 14076 15407 14111 15441
rect 14145 15407 14180 15441
rect 14214 15407 14249 15441
rect 14283 15407 14318 15441
rect 14352 15407 14416 15441
rect 12580 15371 14416 15407
rect 12580 15337 12660 15371
rect 12694 15337 12730 15371
rect 12764 15337 12800 15371
rect 12834 15337 12869 15371
rect 12903 15337 12938 15371
rect 12972 15337 13007 15371
rect 13041 15337 13076 15371
rect 13110 15337 13145 15371
rect 13179 15337 13214 15371
rect 13248 15337 13283 15371
rect 13317 15337 13352 15371
rect 13386 15337 13421 15371
rect 13455 15337 13490 15371
rect 13524 15337 13559 15371
rect 13593 15337 13628 15371
rect 13662 15337 13697 15371
rect 13731 15337 13766 15371
rect 13800 15337 13835 15371
rect 13869 15337 13904 15371
rect 13938 15337 13973 15371
rect 14007 15337 14042 15371
rect 14076 15337 14111 15371
rect 14145 15337 14180 15371
rect 14214 15337 14249 15371
rect 14283 15337 14318 15371
rect 14352 15337 14416 15371
rect 12580 15301 14416 15337
rect 12580 15267 12660 15301
rect 12694 15267 12730 15301
rect 12764 15267 12800 15301
rect 12834 15267 12869 15301
rect 12903 15267 12938 15301
rect 12972 15267 13007 15301
rect 13041 15267 13076 15301
rect 13110 15267 13145 15301
rect 13179 15267 13214 15301
rect 13248 15267 13283 15301
rect 13317 15267 13352 15301
rect 13386 15267 13421 15301
rect 13455 15267 13490 15301
rect 13524 15267 13559 15301
rect 13593 15267 13628 15301
rect 13662 15267 13697 15301
rect 13731 15267 13766 15301
rect 13800 15267 13835 15301
rect 13869 15267 13904 15301
rect 13938 15267 13973 15301
rect 14007 15267 14042 15301
rect 14076 15267 14111 15301
rect 14145 15267 14180 15301
rect 14214 15267 14249 15301
rect 14283 15267 14318 15301
rect 14352 15267 14416 15301
rect 12580 15231 14416 15267
rect 12580 15197 12660 15231
rect 12694 15197 12730 15231
rect 12764 15197 12800 15231
rect 12834 15197 12869 15231
rect 12903 15197 12938 15231
rect 12972 15197 13007 15231
rect 13041 15197 13076 15231
rect 13110 15197 13145 15231
rect 13179 15197 13214 15231
rect 13248 15197 13283 15231
rect 13317 15197 13352 15231
rect 13386 15197 13421 15231
rect 13455 15197 13490 15231
rect 13524 15197 13559 15231
rect 13593 15197 13628 15231
rect 13662 15197 13697 15231
rect 13731 15197 13766 15231
rect 13800 15197 13835 15231
rect 13869 15197 13904 15231
rect 13938 15197 13973 15231
rect 14007 15197 14042 15231
rect 14076 15197 14111 15231
rect 14145 15197 14180 15231
rect 14214 15197 14249 15231
rect 14283 15197 14318 15231
rect 14352 15197 14416 15231
rect 12580 15161 14416 15197
rect 12580 15127 12660 15161
rect 12694 15127 12730 15161
rect 12764 15127 12800 15161
rect 12834 15127 12869 15161
rect 12903 15127 12938 15161
rect 12972 15127 13007 15161
rect 13041 15127 13076 15161
rect 13110 15127 13145 15161
rect 13179 15127 13214 15161
rect 13248 15127 13283 15161
rect 13317 15127 13352 15161
rect 13386 15127 13421 15161
rect 13455 15127 13490 15161
rect 13524 15127 13559 15161
rect 13593 15127 13628 15161
rect 13662 15127 13697 15161
rect 13731 15127 13766 15161
rect 13800 15127 13835 15161
rect 13869 15127 13904 15161
rect 13938 15127 13973 15161
rect 14007 15127 14042 15161
rect 14076 15127 14111 15161
rect 14145 15127 14180 15161
rect 14214 15127 14249 15161
rect 14283 15127 14318 15161
rect 14352 15127 14416 15161
rect 12580 15091 14416 15127
rect 12580 15057 12660 15091
rect 12694 15057 12730 15091
rect 12764 15057 12800 15091
rect 12834 15057 12869 15091
rect 12903 15057 12938 15091
rect 12972 15057 13007 15091
rect 13041 15057 13076 15091
rect 13110 15057 13145 15091
rect 13179 15057 13214 15091
rect 13248 15057 13283 15091
rect 13317 15057 13352 15091
rect 13386 15057 13421 15091
rect 13455 15057 13490 15091
rect 13524 15057 13559 15091
rect 13593 15057 13628 15091
rect 13662 15057 13697 15091
rect 13731 15057 13766 15091
rect 13800 15057 13835 15091
rect 13869 15057 13904 15091
rect 13938 15057 13973 15091
rect 14007 15057 14042 15091
rect 14076 15057 14111 15091
rect 14145 15057 14180 15091
rect 14214 15057 14249 15091
rect 14283 15057 14318 15091
rect 14352 15057 14416 15091
rect 12580 15021 14416 15057
rect 12580 14987 12660 15021
rect 12694 14987 12730 15021
rect 12764 14987 12800 15021
rect 12834 14987 12869 15021
rect 12903 14987 12938 15021
rect 12972 14987 13007 15021
rect 13041 14987 13076 15021
rect 13110 14987 13145 15021
rect 13179 14987 13214 15021
rect 13248 14987 13283 15021
rect 13317 14987 13352 15021
rect 13386 14987 13421 15021
rect 13455 14987 13490 15021
rect 13524 14987 13559 15021
rect 13593 14987 13628 15021
rect 13662 14987 13697 15021
rect 13731 14987 13766 15021
rect 13800 14987 13835 15021
rect 13869 14987 13904 15021
rect 13938 14987 13973 15021
rect 14007 14987 14042 15021
rect 14076 14987 14111 15021
rect 14145 14987 14180 15021
rect 14214 14987 14249 15021
rect 14283 14987 14318 15021
rect 14352 14987 14416 15021
rect 12580 14951 14416 14987
rect 12580 14917 12660 14951
rect 12694 14917 12730 14951
rect 12764 14917 12800 14951
rect 12834 14917 12869 14951
rect 12903 14917 12938 14951
rect 12972 14917 13007 14951
rect 13041 14917 13076 14951
rect 13110 14917 13145 14951
rect 13179 14917 13214 14951
rect 13248 14917 13283 14951
rect 13317 14917 13352 14951
rect 13386 14917 13421 14951
rect 13455 14917 13490 14951
rect 13524 14917 13559 14951
rect 13593 14917 13628 14951
rect 13662 14917 13697 14951
rect 13731 14917 13766 14951
rect 13800 14917 13835 14951
rect 13869 14917 13904 14951
rect 13938 14917 13973 14951
rect 14007 14917 14042 14951
rect 14076 14917 14111 14951
rect 14145 14917 14180 14951
rect 14214 14917 14249 14951
rect 14283 14917 14318 14951
rect 14352 14917 14416 14951
rect 12580 14881 14416 14917
rect 12580 14847 12660 14881
rect 12694 14847 12730 14881
rect 12764 14847 12800 14881
rect 12834 14847 12869 14881
rect 12903 14847 12938 14881
rect 12972 14847 13007 14881
rect 13041 14847 13076 14881
rect 13110 14847 13145 14881
rect 13179 14847 13214 14881
rect 13248 14847 13283 14881
rect 13317 14847 13352 14881
rect 13386 14847 13421 14881
rect 13455 14847 13490 14881
rect 13524 14847 13559 14881
rect 13593 14847 13628 14881
rect 13662 14847 13697 14881
rect 13731 14847 13766 14881
rect 13800 14847 13835 14881
rect 13869 14847 13904 14881
rect 13938 14847 13973 14881
rect 14007 14847 14042 14881
rect 14076 14847 14111 14881
rect 14145 14847 14180 14881
rect 14214 14847 14249 14881
rect 14283 14847 14318 14881
rect 14352 14847 14416 14881
rect 12580 14777 14416 14847
rect -947 9680 15117 9685
rect -947 9647 -723 9680
rect -947 9613 -932 9647
rect -898 9613 -864 9647
rect -830 9613 -796 9647
rect -762 9646 -723 9647
rect -689 9646 -654 9680
rect -620 9646 -585 9680
rect -551 9646 -516 9680
rect -482 9646 -447 9680
rect -413 9646 -378 9680
rect -344 9646 -309 9680
rect -275 9646 -240 9680
rect -206 9646 -171 9680
rect -137 9646 -102 9680
rect -68 9646 -33 9680
rect -762 9613 -33 9646
rect -947 9612 -33 9613
rect -947 9578 -723 9612
rect -689 9578 -654 9612
rect -620 9578 -585 9612
rect -551 9578 -516 9612
rect -482 9578 -447 9612
rect -413 9578 -378 9612
rect -344 9578 -309 9612
rect -275 9578 -240 9612
rect -206 9578 -171 9612
rect -137 9578 -102 9612
rect -68 9578 -33 9612
rect -947 9571 -33 9578
rect -947 9537 -932 9571
rect -898 9537 -864 9571
rect -830 9537 -796 9571
rect -762 9544 -33 9571
rect -762 9537 -723 9544
rect -947 9510 -723 9537
rect -689 9510 -654 9544
rect -620 9510 -585 9544
rect -551 9510 -516 9544
rect -482 9514 -447 9544
rect -450 9510 -447 9514
rect -413 9514 -378 9544
rect -344 9514 -309 9544
rect -275 9514 -240 9544
rect -206 9514 -171 9544
rect -137 9514 -102 9544
rect -68 9514 -33 9544
rect 14893 9647 15117 9680
rect 14893 9613 14932 9647
rect 14966 9613 15000 9647
rect 15034 9613 15068 9647
rect 15102 9613 15117 9647
rect 14893 9571 15117 9613
rect 14893 9537 14932 9571
rect 14966 9537 15000 9571
rect 15034 9537 15068 9571
rect 15102 9537 15117 9571
rect -413 9510 -411 9514
rect -344 9510 -338 9514
rect -275 9510 -265 9514
rect -206 9510 -192 9514
rect -137 9510 -119 9514
rect -68 9510 -46 9514
rect -947 9495 -484 9510
rect -947 9461 -932 9495
rect -898 9461 -864 9495
rect -830 9461 -796 9495
rect -762 9480 -484 9495
rect -450 9480 -411 9510
rect -377 9480 -338 9510
rect -304 9480 -265 9510
rect -231 9480 -192 9510
rect -158 9480 -119 9510
rect -85 9480 -46 9510
rect 14893 9495 15117 9537
rect -762 9476 -33 9480
rect -762 9461 -723 9476
rect -947 9442 -723 9461
rect -689 9442 -654 9476
rect -620 9442 -585 9476
rect -551 9442 -516 9476
rect -482 9442 -447 9476
rect -413 9442 -378 9476
rect -344 9442 -309 9476
rect -275 9442 -240 9476
rect -206 9442 -171 9476
rect -137 9442 -102 9476
rect -68 9442 -33 9476
rect -947 9428 -33 9442
rect 14893 9461 14932 9495
rect 14966 9461 15000 9495
rect 15034 9461 15068 9495
rect 15102 9461 15117 9495
rect -947 9418 -484 9428
rect -947 9384 -932 9418
rect -898 9384 -864 9418
rect -830 9384 -796 9418
rect -762 9408 -484 9418
rect -450 9408 -411 9428
rect -377 9408 -338 9428
rect -304 9408 -265 9428
rect -231 9408 -192 9428
rect -158 9408 -119 9428
rect -85 9408 -46 9428
rect -762 9384 -723 9408
rect -947 9374 -723 9384
rect -689 9374 -654 9408
rect -620 9374 -585 9408
rect -551 9374 -516 9408
rect -450 9394 -447 9408
rect -482 9374 -447 9394
rect -413 9394 -411 9408
rect -344 9394 -338 9408
rect -275 9394 -265 9408
rect -206 9394 -192 9408
rect -137 9394 -119 9408
rect -68 9394 -46 9408
rect 14893 9418 15117 9461
rect -413 9374 -378 9394
rect -344 9374 -309 9394
rect -275 9374 -240 9394
rect -206 9374 -171 9394
rect -137 9374 -102 9394
rect -68 9374 -33 9394
rect -947 9342 -33 9374
rect 14893 9384 14932 9418
rect 14966 9384 15000 9418
rect 15034 9384 15068 9418
rect 15102 9384 15117 9418
rect -947 9341 -484 9342
rect -947 9307 -932 9341
rect -898 9307 -864 9341
rect -830 9307 -796 9341
rect -762 9340 -484 9341
rect -450 9340 -411 9342
rect -377 9340 -338 9342
rect -304 9340 -265 9342
rect -231 9340 -192 9342
rect -158 9340 -119 9342
rect -85 9340 -46 9342
rect -762 9307 -723 9340
rect -947 9306 -723 9307
rect -689 9306 -654 9340
rect -620 9306 -585 9340
rect -551 9306 -516 9340
rect -450 9308 -447 9340
rect -482 9306 -447 9308
rect -413 9308 -411 9340
rect -344 9308 -338 9340
rect -275 9308 -265 9340
rect -206 9308 -192 9340
rect -137 9308 -119 9340
rect -68 9308 -46 9340
rect 14893 9341 15117 9384
rect -413 9306 -378 9308
rect -344 9306 -309 9308
rect -275 9306 -240 9308
rect -206 9306 -171 9308
rect -137 9306 -102 9308
rect -68 9306 -33 9308
rect -947 9272 -33 9306
rect -947 9264 -723 9272
rect -947 9230 -932 9264
rect -898 9230 -864 9264
rect -830 9230 -796 9264
rect -762 9238 -723 9264
rect -689 9238 -654 9272
rect -620 9238 -585 9272
rect -551 9238 -516 9272
rect -482 9256 -447 9272
rect -450 9238 -447 9256
rect -413 9256 -378 9272
rect -344 9256 -309 9272
rect -275 9256 -240 9272
rect -206 9256 -171 9272
rect -137 9256 -102 9272
rect -68 9256 -33 9272
rect 14893 9307 14932 9341
rect 14966 9307 15000 9341
rect 15034 9307 15068 9341
rect 15102 9307 15117 9341
rect 14893 9264 15117 9307
rect -413 9238 -411 9256
rect -344 9238 -338 9256
rect -275 9238 -265 9256
rect -206 9238 -192 9256
rect -137 9238 -119 9256
rect -68 9238 -46 9256
rect -762 9230 -484 9238
rect -947 9222 -484 9230
rect -450 9222 -411 9238
rect -377 9222 -338 9238
rect -304 9222 -265 9238
rect -231 9222 -192 9238
rect -158 9222 -119 9238
rect -85 9222 -46 9238
rect 14893 9230 14932 9264
rect 14966 9230 15000 9264
rect 15034 9230 15068 9264
rect 15102 9230 15117 9264
rect -947 9204 -33 9222
rect -947 9187 -723 9204
rect -947 9153 -932 9187
rect -898 9153 -864 9187
rect -830 9153 -796 9187
rect -762 9170 -723 9187
rect -689 9170 -654 9204
rect -620 9170 -585 9204
rect -551 9170 -516 9204
rect -482 9170 -447 9204
rect -413 9170 -378 9204
rect -344 9170 -309 9204
rect -275 9170 -240 9204
rect -206 9170 -171 9204
rect -137 9170 -102 9204
rect -68 9170 -33 9204
rect 14893 9187 15117 9230
rect -762 9153 -484 9170
rect -947 9136 -484 9153
rect -450 9136 -411 9170
rect -377 9136 -338 9170
rect -304 9136 -265 9170
rect -231 9136 -192 9170
rect -158 9136 -119 9170
rect -85 9136 -46 9170
rect 14893 9153 14932 9187
rect 14966 9153 15000 9187
rect 15034 9153 15068 9187
rect 15102 9153 15117 9187
rect -947 9110 -723 9136
rect -947 9076 -932 9110
rect -898 9076 -864 9110
rect -830 9076 -796 9110
rect -762 9102 -723 9110
rect -689 9102 -654 9136
rect -620 9102 -585 9136
rect -551 9102 -516 9136
rect -482 9102 -447 9136
rect -413 9102 -378 9136
rect -344 9102 -309 9136
rect -275 9102 -240 9136
rect -206 9102 -171 9136
rect -137 9102 -102 9136
rect -68 9102 -33 9136
rect -762 9076 -33 9102
rect -947 9068 -33 9076
rect -947 9034 -723 9068
rect -689 9034 -654 9068
rect -620 9034 -585 9068
rect -551 9034 -516 9068
rect -482 9034 -447 9068
rect -413 9034 -378 9068
rect -344 9034 -309 9068
rect -275 9034 -240 9068
rect -206 9034 -171 9068
rect -137 9034 -102 9068
rect -68 9034 -33 9068
rect -947 9033 -33 9034
rect -947 8999 -932 9033
rect -898 8999 -864 9033
rect -830 8999 -796 9033
rect -762 9000 -33 9033
rect -762 8999 -723 9000
rect -947 8966 -723 8999
rect -689 8966 -654 9000
rect -620 8966 -585 9000
rect -551 8966 -516 9000
rect -482 8966 -447 9000
rect -413 8966 -378 9000
rect -344 8966 -309 9000
rect -275 8966 -240 9000
rect -206 8966 -171 9000
rect -137 8966 -102 9000
rect -68 8966 -33 9000
rect 14893 9110 15117 9153
rect 14893 9076 14932 9110
rect 14966 9076 15000 9110
rect 15034 9076 15068 9110
rect 15102 9076 15117 9110
rect 14893 9033 15117 9076
rect 14893 8999 14932 9033
rect 14966 8999 15000 9033
rect 15034 8999 15068 9033
rect 15102 8999 15117 9033
rect 14893 8966 15117 8999
rect -947 8961 15117 8966
rect 8367 8808 15102 8809
rect 42 8774 15102 8808
rect 42 8740 68 8774
rect 102 8740 138 8774
rect 172 8740 208 8774
rect 242 8753 278 8774
rect 312 8753 348 8774
rect 382 8753 418 8774
rect 452 8753 488 8774
rect 522 8753 558 8774
rect 592 8753 628 8774
rect 662 8753 698 8774
rect 732 8753 768 8774
rect 802 8753 838 8774
rect 242 8740 248 8753
rect 312 8740 322 8753
rect 382 8740 396 8753
rect 452 8740 470 8753
rect 522 8740 544 8753
rect 592 8740 618 8753
rect 662 8740 691 8753
rect 732 8740 764 8753
rect 802 8740 837 8753
rect 872 8740 908 8774
rect 942 8760 978 8774
rect 1012 8760 1048 8774
rect 1082 8760 1118 8774
rect 1152 8760 1188 8774
rect 1222 8760 1258 8774
rect 1292 8760 1328 8774
rect 1362 8760 1398 8774
rect 1432 8760 1467 8774
rect 1501 8760 1536 8774
rect 1570 8760 1605 8774
rect 1639 8760 1674 8774
rect 1708 8760 1743 8774
rect 1777 8760 1812 8774
rect 946 8740 978 8760
rect 1018 8740 1048 8760
rect 1090 8740 1118 8760
rect 1162 8740 1188 8760
rect 1234 8740 1258 8760
rect 1306 8740 1328 8760
rect 1378 8740 1398 8760
rect 1450 8740 1467 8760
rect 1522 8740 1536 8760
rect 1594 8740 1605 8760
rect 1666 8740 1674 8760
rect 1738 8740 1743 8760
rect 1810 8740 1812 8760
rect 1846 8760 1881 8774
rect 1915 8760 1950 8774
rect 1984 8760 2019 8774
rect 2053 8760 2088 8774
rect 2122 8760 2157 8774
rect 1846 8740 1849 8760
rect 1915 8740 1922 8760
rect 1984 8740 1995 8760
rect 2053 8740 2068 8760
rect 2122 8740 2141 8760
rect 2191 8740 2226 8774
rect 2260 8753 2295 8774
rect 2329 8753 2364 8774
rect 2398 8753 2433 8774
rect 2467 8753 2502 8774
rect 2261 8740 2295 8753
rect 2340 8740 2364 8753
rect 2419 8740 2433 8753
rect 2498 8740 2502 8753
rect 2536 8753 2571 8774
rect 2605 8753 2640 8774
rect 2674 8753 2709 8774
rect 2743 8753 2778 8774
rect 2536 8740 2543 8753
rect 2605 8740 2621 8753
rect 2674 8740 2699 8753
rect 2743 8740 2777 8753
rect 2812 8740 2847 8774
rect 2881 8773 15102 8774
rect 2881 8770 8393 8773
rect 2881 8753 2933 8770
rect 42 8719 248 8740
rect 282 8719 322 8740
rect 356 8719 396 8740
rect 430 8719 470 8740
rect 504 8719 544 8740
rect 578 8719 618 8740
rect 652 8719 691 8740
rect 725 8719 764 8740
rect 798 8719 837 8740
rect 871 8726 912 8740
rect 946 8726 984 8740
rect 1018 8726 1056 8740
rect 1090 8726 1128 8740
rect 1162 8726 1200 8740
rect 1234 8726 1272 8740
rect 1306 8726 1344 8740
rect 1378 8726 1416 8740
rect 1450 8726 1488 8740
rect 1522 8726 1560 8740
rect 1594 8726 1632 8740
rect 1666 8726 1704 8740
rect 1738 8726 1776 8740
rect 1810 8726 1849 8740
rect 1883 8726 1922 8740
rect 1956 8726 1995 8740
rect 2029 8726 2068 8740
rect 2102 8726 2141 8740
rect 2175 8726 2227 8740
rect 871 8719 2227 8726
rect 2261 8719 2306 8740
rect 2340 8719 2385 8740
rect 2419 8719 2464 8740
rect 2498 8719 2543 8740
rect 2577 8719 2621 8740
rect 2655 8719 2699 8740
rect 2733 8719 2777 8740
rect 2811 8719 2855 8740
rect 2889 8719 2933 8753
rect 2967 8736 3002 8770
rect 3036 8753 3071 8770
rect 3045 8736 3071 8753
rect 3105 8736 3139 8770
rect 3173 8736 3207 8770
rect 3241 8736 3275 8770
rect 3309 8736 3343 8770
rect 3377 8736 3411 8770
rect 3445 8760 3479 8770
rect 3445 8736 3477 8760
rect 3513 8736 3547 8770
rect 3581 8760 3615 8770
rect 3649 8760 3683 8770
rect 3717 8760 3751 8770
rect 3785 8760 3819 8770
rect 3853 8760 3887 8770
rect 3921 8760 3955 8770
rect 3989 8760 4023 8770
rect 3584 8736 3615 8760
rect 3657 8736 3683 8760
rect 3730 8736 3751 8760
rect 3803 8736 3819 8760
rect 3876 8736 3887 8760
rect 3949 8736 3955 8760
rect 4022 8736 4023 8760
rect 4057 8760 4091 8770
rect 4125 8760 4159 8770
rect 4193 8760 4227 8770
rect 4261 8760 4295 8770
rect 4329 8760 4363 8770
rect 4397 8760 4431 8770
rect 4057 8736 4061 8760
rect 4125 8736 4134 8760
rect 4193 8736 4207 8760
rect 4261 8736 4280 8760
rect 4329 8736 4353 8760
rect 4397 8736 4426 8760
rect 4465 8736 4499 8770
rect 4533 8736 4567 8770
rect 4601 8760 4635 8770
rect 4669 8760 4703 8770
rect 4737 8760 4771 8770
rect 4805 8760 4839 8770
rect 4873 8760 4907 8770
rect 4941 8760 4975 8770
rect 4606 8736 4635 8760
rect 4679 8736 4703 8760
rect 4752 8736 4771 8760
rect 4825 8736 4839 8760
rect 4898 8736 4907 8760
rect 4971 8736 4975 8760
rect 5009 8760 5043 8770
rect 5077 8760 5111 8770
rect 5145 8760 5179 8770
rect 5213 8760 5247 8770
rect 5281 8760 5315 8770
rect 5349 8760 5383 8770
rect 5417 8760 5451 8770
rect 5009 8736 5010 8760
rect 5077 8736 5083 8760
rect 5145 8736 5156 8760
rect 5213 8736 5229 8760
rect 5281 8736 5302 8760
rect 5349 8736 5375 8760
rect 5417 8736 5448 8760
rect 5485 8736 5519 8770
rect 5553 8760 5587 8770
rect 5621 8760 5655 8770
rect 5689 8760 5723 8770
rect 5757 8760 5791 8770
rect 5825 8760 5859 8770
rect 5893 8760 5927 8770
rect 5961 8760 5995 8770
rect 5555 8736 5587 8760
rect 5628 8736 5655 8760
rect 5701 8736 5723 8760
rect 5774 8736 5791 8760
rect 5847 8736 5859 8760
rect 5920 8736 5927 8760
rect 5993 8736 5995 8760
rect 6029 8760 6063 8770
rect 6097 8760 6131 8770
rect 6165 8760 6199 8770
rect 6233 8760 6267 8770
rect 6301 8760 6335 8770
rect 6369 8760 6403 8770
rect 6437 8760 6471 8770
rect 6029 8736 6032 8760
rect 6097 8736 6105 8760
rect 6165 8736 6178 8760
rect 6233 8736 6251 8760
rect 6301 8736 6324 8760
rect 6369 8736 6397 8760
rect 6437 8736 6470 8760
rect 6505 8736 6539 8770
rect 6573 8760 6607 8770
rect 6641 8760 6675 8770
rect 6709 8760 6743 8770
rect 6777 8760 6811 8770
rect 6845 8760 6879 8770
rect 6913 8760 6947 8770
rect 6577 8736 6607 8760
rect 6650 8736 6675 8760
rect 6723 8736 6743 8760
rect 6796 8736 6811 8760
rect 6869 8736 6879 8760
rect 6942 8736 6947 8760
rect 6981 8760 7015 8770
rect 2967 8719 3011 8736
rect 3045 8726 3477 8736
rect 3511 8726 3550 8736
rect 3584 8726 3623 8736
rect 3657 8726 3696 8736
rect 3730 8726 3769 8736
rect 3803 8726 3842 8736
rect 3876 8726 3915 8736
rect 3949 8726 3988 8736
rect 4022 8726 4061 8736
rect 4095 8726 4134 8736
rect 4168 8726 4207 8736
rect 4241 8726 4280 8736
rect 4314 8726 4353 8736
rect 4387 8726 4426 8736
rect 4460 8726 4499 8736
rect 4533 8726 4572 8736
rect 4606 8726 4645 8736
rect 4679 8726 4718 8736
rect 4752 8726 4791 8736
rect 4825 8726 4864 8736
rect 4898 8726 4937 8736
rect 4971 8726 5010 8736
rect 5044 8726 5083 8736
rect 5117 8726 5156 8736
rect 5190 8726 5229 8736
rect 5263 8726 5302 8736
rect 5336 8726 5375 8736
rect 5409 8726 5448 8736
rect 5482 8726 5521 8736
rect 5555 8726 5594 8736
rect 5628 8726 5667 8736
rect 5701 8726 5740 8736
rect 5774 8726 5813 8736
rect 5847 8726 5886 8736
rect 5920 8726 5959 8736
rect 5993 8726 6032 8736
rect 6066 8726 6105 8736
rect 6139 8726 6178 8736
rect 6212 8726 6251 8736
rect 6285 8726 6324 8736
rect 6358 8726 6397 8736
rect 6431 8726 6470 8736
rect 6504 8726 6543 8736
rect 6577 8726 6616 8736
rect 6650 8726 6689 8736
rect 6723 8726 6762 8736
rect 6796 8726 6835 8736
rect 6869 8726 6908 8736
rect 6942 8726 6981 8736
rect 7049 8760 7083 8770
rect 7117 8760 7151 8770
rect 7185 8760 7219 8770
rect 7253 8760 7287 8770
rect 7321 8760 7355 8770
rect 7389 8760 7423 8770
rect 7049 8736 7054 8760
rect 7117 8736 7127 8760
rect 7185 8736 7200 8760
rect 7253 8736 7273 8760
rect 7321 8736 7346 8760
rect 7389 8736 7419 8760
rect 7457 8736 7491 8770
rect 7525 8760 7559 8770
rect 7593 8760 7627 8770
rect 7661 8760 7695 8770
rect 7729 8760 7763 8770
rect 7797 8760 7831 8770
rect 7865 8760 7899 8770
rect 7933 8760 7967 8770
rect 7526 8736 7559 8760
rect 7599 8736 7627 8760
rect 7672 8736 7695 8760
rect 7745 8736 7763 8760
rect 7818 8736 7831 8760
rect 7891 8736 7899 8760
rect 7964 8736 7967 8760
rect 8001 8760 8035 8770
rect 8069 8760 8103 8770
rect 8137 8760 8171 8770
rect 8205 8760 8239 8770
rect 8273 8760 8307 8770
rect 8341 8760 8393 8770
rect 8427 8760 8462 8773
rect 8496 8760 8531 8773
rect 8565 8760 8600 8773
rect 8634 8760 8669 8773
rect 8703 8760 8738 8773
rect 8772 8760 8807 8773
rect 8841 8760 8876 8773
rect 8910 8760 8945 8773
rect 8979 8760 9014 8773
rect 8001 8736 8003 8760
rect 8069 8736 8075 8760
rect 8137 8736 8147 8760
rect 8205 8736 8219 8760
rect 8273 8736 8291 8760
rect 8341 8736 8363 8760
rect 8427 8739 8435 8760
rect 8496 8739 8507 8760
rect 8565 8739 8579 8760
rect 8634 8739 8651 8760
rect 8703 8739 8723 8760
rect 8772 8739 8795 8760
rect 8841 8739 8867 8760
rect 8910 8739 8939 8760
rect 8979 8739 9011 8760
rect 9048 8739 9083 8773
rect 9117 8739 9152 8773
rect 9186 8760 9220 8773
rect 9254 8760 9288 8773
rect 9322 8760 9356 8773
rect 9390 8760 9424 8773
rect 9458 8760 9492 8773
rect 9526 8760 9560 8773
rect 9594 8760 9628 8773
rect 9662 8760 9696 8773
rect 9189 8739 9220 8760
rect 9261 8739 9288 8760
rect 9333 8739 9356 8760
rect 9405 8739 9424 8760
rect 9477 8739 9492 8760
rect 9549 8739 9560 8760
rect 9621 8739 9628 8760
rect 9693 8739 9696 8760
rect 9730 8760 9764 8773
rect 9798 8760 9832 8773
rect 9866 8760 9900 8773
rect 9934 8760 9968 8773
rect 10002 8760 10036 8773
rect 10070 8760 10104 8773
rect 10138 8760 10172 8773
rect 10206 8760 10240 8773
rect 10274 8760 10308 8773
rect 9730 8739 9731 8760
rect 9798 8739 9803 8760
rect 9866 8739 9875 8760
rect 9934 8739 9947 8760
rect 10002 8739 10019 8760
rect 10070 8739 10091 8760
rect 10138 8739 10163 8760
rect 10206 8739 10235 8760
rect 10274 8739 10307 8760
rect 10342 8739 10376 8773
rect 10410 8760 10444 8773
rect 10478 8760 10512 8773
rect 10546 8760 10580 8773
rect 10614 8760 10648 8773
rect 10682 8760 10716 8773
rect 10750 8760 10784 8773
rect 10818 8760 10852 8773
rect 10886 8760 10920 8773
rect 10413 8739 10444 8760
rect 10485 8739 10512 8760
rect 10557 8739 10580 8760
rect 10629 8739 10648 8760
rect 10701 8739 10716 8760
rect 10773 8739 10784 8760
rect 10845 8739 10852 8760
rect 10917 8739 10920 8760
rect 10954 8760 10988 8773
rect 11022 8760 11056 8773
rect 11090 8760 11124 8773
rect 11158 8760 11192 8773
rect 11226 8760 11260 8773
rect 11294 8760 11328 8773
rect 11362 8760 11396 8773
rect 11430 8760 11464 8773
rect 11498 8760 11532 8773
rect 10954 8739 10955 8760
rect 11022 8739 11027 8760
rect 11090 8739 11099 8760
rect 11158 8739 11171 8760
rect 11226 8739 11243 8760
rect 11294 8739 11315 8760
rect 11362 8739 11387 8760
rect 11430 8739 11459 8760
rect 11498 8739 11531 8760
rect 11566 8739 11600 8773
rect 11634 8760 11668 8773
rect 11702 8760 11736 8773
rect 11770 8760 11804 8773
rect 11838 8760 11872 8773
rect 11906 8760 11940 8773
rect 11974 8760 12008 8773
rect 12042 8760 12076 8773
rect 12110 8760 12144 8773
rect 11637 8739 11668 8760
rect 11709 8739 11736 8760
rect 11781 8739 11804 8760
rect 11853 8739 11872 8760
rect 11925 8739 11940 8760
rect 11997 8739 12008 8760
rect 12069 8739 12076 8760
rect 12141 8739 12144 8760
rect 12178 8760 12212 8773
rect 12246 8760 12280 8773
rect 12314 8760 12348 8773
rect 12382 8760 12416 8773
rect 12450 8760 12484 8773
rect 12518 8760 12552 8773
rect 12586 8760 12620 8773
rect 12654 8760 12688 8773
rect 12722 8760 12756 8773
rect 12178 8739 12179 8760
rect 12246 8739 12251 8760
rect 12314 8739 12323 8760
rect 12382 8739 12395 8760
rect 12450 8739 12467 8760
rect 12518 8739 12539 8760
rect 12586 8739 12611 8760
rect 12654 8739 12683 8760
rect 12722 8739 12755 8760
rect 12790 8739 12824 8773
rect 12858 8760 12892 8773
rect 12926 8760 12960 8773
rect 12994 8760 13028 8773
rect 13062 8760 13096 8773
rect 13130 8760 13164 8773
rect 13198 8760 13232 8773
rect 13266 8760 13300 8773
rect 13334 8760 13368 8773
rect 12861 8739 12892 8760
rect 12933 8739 12960 8760
rect 13005 8739 13028 8760
rect 13077 8739 13096 8760
rect 13149 8739 13164 8760
rect 13221 8739 13232 8760
rect 13293 8739 13300 8760
rect 13365 8739 13368 8760
rect 13402 8760 13436 8773
rect 13470 8760 13504 8773
rect 13538 8760 13572 8773
rect 13606 8760 13640 8773
rect 13674 8760 13708 8773
rect 13742 8760 13776 8773
rect 13810 8760 13844 8773
rect 13878 8760 13912 8773
rect 13946 8760 13980 8773
rect 13402 8739 13403 8760
rect 13470 8739 13475 8760
rect 13538 8739 13547 8760
rect 13606 8739 13619 8760
rect 13674 8739 13691 8760
rect 13742 8739 13763 8760
rect 13810 8739 13835 8760
rect 13878 8739 13907 8760
rect 13946 8739 13979 8760
rect 14014 8739 14048 8773
rect 14082 8760 14116 8773
rect 14150 8760 14184 8773
rect 14218 8760 14252 8773
rect 14286 8760 14320 8773
rect 14354 8760 14388 8773
rect 14422 8760 14456 8773
rect 14490 8760 14524 8773
rect 14558 8760 14592 8773
rect 14085 8739 14116 8760
rect 14157 8739 14184 8760
rect 14229 8739 14252 8760
rect 14301 8739 14320 8760
rect 14373 8739 14388 8760
rect 14445 8739 14456 8760
rect 14517 8739 14524 8760
rect 14589 8739 14592 8760
rect 14626 8760 14660 8773
rect 14694 8760 14728 8773
rect 14762 8760 14796 8773
rect 14830 8760 14864 8773
rect 14626 8739 14627 8760
rect 14694 8739 14699 8760
rect 14762 8739 14771 8760
rect 14830 8739 14843 8760
rect 14898 8739 15102 8773
rect 7015 8726 7054 8736
rect 7088 8726 7127 8736
rect 7161 8726 7200 8736
rect 7234 8726 7273 8736
rect 7307 8726 7346 8736
rect 7380 8726 7419 8736
rect 7453 8726 7492 8736
rect 7526 8726 7565 8736
rect 7599 8726 7638 8736
rect 7672 8726 7711 8736
rect 7745 8726 7784 8736
rect 7818 8726 7857 8736
rect 7891 8726 7930 8736
rect 7964 8726 8003 8736
rect 8037 8726 8075 8736
rect 8109 8726 8147 8736
rect 8181 8726 8219 8736
rect 8253 8726 8291 8736
rect 8325 8726 8363 8736
rect 8397 8726 8435 8739
rect 8469 8726 8507 8739
rect 8541 8726 8579 8739
rect 8613 8726 8651 8739
rect 8685 8726 8723 8739
rect 8757 8726 8795 8739
rect 8829 8726 8867 8739
rect 8901 8726 8939 8739
rect 8973 8726 9011 8739
rect 9045 8726 9083 8739
rect 9117 8726 9155 8739
rect 9189 8726 9227 8739
rect 9261 8726 9299 8739
rect 9333 8726 9371 8739
rect 9405 8726 9443 8739
rect 9477 8726 9515 8739
rect 9549 8726 9587 8739
rect 9621 8726 9659 8739
rect 9693 8726 9731 8739
rect 9765 8726 9803 8739
rect 9837 8726 9875 8739
rect 9909 8726 9947 8739
rect 9981 8726 10019 8739
rect 10053 8726 10091 8739
rect 10125 8726 10163 8739
rect 10197 8726 10235 8739
rect 10269 8726 10307 8739
rect 10341 8726 10379 8739
rect 10413 8726 10451 8739
rect 10485 8726 10523 8739
rect 10557 8726 10595 8739
rect 10629 8726 10667 8739
rect 10701 8726 10739 8739
rect 10773 8726 10811 8739
rect 10845 8726 10883 8739
rect 10917 8726 10955 8739
rect 10989 8726 11027 8739
rect 11061 8726 11099 8739
rect 11133 8726 11171 8739
rect 11205 8726 11243 8739
rect 11277 8726 11315 8739
rect 11349 8726 11387 8739
rect 11421 8726 11459 8739
rect 11493 8726 11531 8739
rect 11565 8726 11603 8739
rect 11637 8726 11675 8739
rect 11709 8726 11747 8739
rect 11781 8726 11819 8739
rect 11853 8726 11891 8739
rect 11925 8726 11963 8739
rect 11997 8726 12035 8739
rect 12069 8726 12107 8739
rect 12141 8726 12179 8739
rect 12213 8726 12251 8739
rect 12285 8726 12323 8739
rect 12357 8726 12395 8739
rect 12429 8726 12467 8739
rect 12501 8726 12539 8739
rect 12573 8726 12611 8739
rect 12645 8726 12683 8739
rect 12717 8726 12755 8739
rect 12789 8726 12827 8739
rect 12861 8726 12899 8739
rect 12933 8726 12971 8739
rect 13005 8726 13043 8739
rect 13077 8726 13115 8739
rect 13149 8726 13187 8739
rect 13221 8726 13259 8739
rect 13293 8726 13331 8739
rect 13365 8726 13403 8739
rect 13437 8726 13475 8739
rect 13509 8726 13547 8739
rect 13581 8726 13619 8739
rect 13653 8726 13691 8739
rect 13725 8726 13763 8739
rect 13797 8726 13835 8739
rect 13869 8726 13907 8739
rect 13941 8726 13979 8739
rect 14013 8726 14051 8739
rect 14085 8726 14123 8739
rect 14157 8726 14195 8739
rect 14229 8726 14267 8739
rect 14301 8726 14339 8739
rect 14373 8726 14411 8739
rect 14445 8726 14483 8739
rect 14517 8726 14555 8739
rect 14589 8726 14627 8739
rect 14661 8726 14699 8739
rect 14733 8726 14771 8739
rect 14805 8726 14843 8739
rect 14877 8726 15102 8739
rect 3045 8721 15102 8726
rect 3045 8719 14932 8721
rect 42 8700 14932 8719
rect 42 8666 68 8700
rect 102 8666 138 8700
rect 172 8666 208 8700
rect 242 8666 278 8700
rect 312 8666 348 8700
rect 382 8666 418 8700
rect 452 8666 488 8700
rect 522 8666 558 8700
rect 592 8666 628 8700
rect 662 8666 698 8700
rect 732 8666 768 8700
rect 802 8666 838 8700
rect 872 8666 908 8700
rect 942 8666 978 8700
rect 1012 8666 1048 8700
rect 1082 8666 1118 8700
rect 1152 8666 1188 8700
rect 1222 8666 1258 8700
rect 1292 8666 1328 8700
rect 1362 8666 1398 8700
rect 1432 8666 1467 8700
rect 1501 8666 1536 8700
rect 1570 8666 1605 8700
rect 1639 8666 1674 8700
rect 1708 8666 1743 8700
rect 1777 8666 1812 8700
rect 1846 8666 1881 8700
rect 1915 8666 1950 8700
rect 1984 8666 2019 8700
rect 2053 8666 2088 8700
rect 2122 8666 2157 8700
rect 2191 8666 2226 8700
rect 2260 8666 2295 8700
rect 2329 8666 2364 8700
rect 2398 8666 2433 8700
rect 2467 8666 2502 8700
rect 2536 8666 2571 8700
rect 2605 8666 2640 8700
rect 2674 8666 2709 8700
rect 2743 8666 2778 8700
rect 2812 8666 2847 8700
rect 2881 8666 2933 8700
rect 2967 8666 3002 8700
rect 3036 8666 3071 8700
rect 3105 8666 3139 8700
rect 3173 8666 3207 8700
rect 3241 8666 3275 8700
rect 3309 8666 3343 8700
rect 3377 8666 3411 8700
rect 3445 8666 3479 8700
rect 3513 8666 3547 8700
rect 3581 8666 3615 8700
rect 3649 8666 3683 8700
rect 3717 8666 3751 8700
rect 3785 8666 3819 8700
rect 3853 8666 3887 8700
rect 3921 8666 3955 8700
rect 3989 8666 4023 8700
rect 4057 8666 4091 8700
rect 4125 8666 4159 8700
rect 4193 8666 4227 8700
rect 4261 8666 4295 8700
rect 4329 8666 4363 8700
rect 4397 8666 4431 8700
rect 4465 8666 4499 8700
rect 4533 8666 4567 8700
rect 4601 8666 4635 8700
rect 4669 8666 4703 8700
rect 4737 8666 4771 8700
rect 4805 8666 4839 8700
rect 4873 8666 4907 8700
rect 4941 8666 4975 8700
rect 5009 8666 5043 8700
rect 5077 8666 5111 8700
rect 5145 8666 5179 8700
rect 5213 8666 5247 8700
rect 5281 8666 5315 8700
rect 5349 8666 5383 8700
rect 5417 8666 5451 8700
rect 5485 8666 5519 8700
rect 5553 8666 5587 8700
rect 5621 8666 5655 8700
rect 5689 8666 5723 8700
rect 5757 8666 5791 8700
rect 5825 8666 5859 8700
rect 5893 8666 5927 8700
rect 5961 8666 5995 8700
rect 6029 8666 6063 8700
rect 6097 8666 6131 8700
rect 6165 8666 6199 8700
rect 6233 8666 6267 8700
rect 6301 8666 6335 8700
rect 6369 8666 6403 8700
rect 6437 8666 6471 8700
rect 6505 8666 6539 8700
rect 6573 8666 6607 8700
rect 6641 8666 6675 8700
rect 6709 8666 6743 8700
rect 6777 8666 6811 8700
rect 6845 8666 6879 8700
rect 6913 8666 6947 8700
rect 6981 8666 7015 8700
rect 7049 8666 7083 8700
rect 7117 8666 7151 8700
rect 7185 8666 7219 8700
rect 7253 8666 7287 8700
rect 7321 8666 7355 8700
rect 7389 8666 7423 8700
rect 7457 8666 7491 8700
rect 7525 8666 7559 8700
rect 7593 8666 7627 8700
rect 7661 8666 7695 8700
rect 7729 8666 7763 8700
rect 7797 8666 7831 8700
rect 7865 8666 7899 8700
rect 7933 8666 7967 8700
rect 8001 8666 8035 8700
rect 8069 8666 8103 8700
rect 8137 8666 8171 8700
rect 8205 8666 8239 8700
rect 8273 8666 8307 8700
rect 8341 8693 14932 8700
rect 8341 8666 8393 8693
rect 42 8659 8393 8666
rect 8427 8659 8462 8693
rect 8496 8659 8531 8693
rect 8565 8659 8600 8693
rect 8634 8659 8669 8693
rect 8703 8659 8738 8693
rect 8772 8659 8807 8693
rect 8841 8659 8876 8693
rect 8910 8659 8945 8693
rect 8979 8659 9014 8693
rect 9048 8659 9083 8693
rect 9117 8659 9152 8693
rect 9186 8659 9220 8693
rect 9254 8659 9288 8693
rect 9322 8659 9356 8693
rect 9390 8659 9424 8693
rect 9458 8659 9492 8693
rect 9526 8659 9560 8693
rect 9594 8659 9628 8693
rect 9662 8659 9696 8693
rect 9730 8659 9764 8693
rect 9798 8659 9832 8693
rect 9866 8659 9900 8693
rect 9934 8659 9968 8693
rect 10002 8659 10036 8693
rect 10070 8659 10104 8693
rect 10138 8659 10172 8693
rect 10206 8659 10240 8693
rect 10274 8659 10308 8693
rect 10342 8659 10376 8693
rect 10410 8659 10444 8693
rect 10478 8659 10512 8693
rect 10546 8659 10580 8693
rect 10614 8659 10648 8693
rect 10682 8659 10716 8693
rect 10750 8659 10784 8693
rect 10818 8659 10852 8693
rect 10886 8659 10920 8693
rect 10954 8659 10988 8693
rect 11022 8659 11056 8693
rect 11090 8659 11124 8693
rect 11158 8659 11192 8693
rect 11226 8659 11260 8693
rect 11294 8659 11328 8693
rect 11362 8659 11396 8693
rect 11430 8659 11464 8693
rect 11498 8659 11532 8693
rect 11566 8659 11600 8693
rect 11634 8659 11668 8693
rect 11702 8659 11736 8693
rect 11770 8659 11804 8693
rect 11838 8659 11872 8693
rect 11906 8659 11940 8693
rect 11974 8659 12008 8693
rect 12042 8659 12076 8693
rect 12110 8659 12144 8693
rect 12178 8659 12212 8693
rect 12246 8659 12280 8693
rect 12314 8659 12348 8693
rect 12382 8659 12416 8693
rect 12450 8659 12484 8693
rect 12518 8659 12552 8693
rect 12586 8659 12620 8693
rect 12654 8659 12688 8693
rect 12722 8659 12756 8693
rect 12790 8659 12824 8693
rect 12858 8659 12892 8693
rect 12926 8659 12960 8693
rect 12994 8659 13028 8693
rect 13062 8659 13096 8693
rect 13130 8659 13164 8693
rect 13198 8659 13232 8693
rect 13266 8659 13300 8693
rect 13334 8659 13368 8693
rect 13402 8659 13436 8693
rect 13470 8659 13504 8693
rect 13538 8659 13572 8693
rect 13606 8659 13640 8693
rect 13674 8659 13708 8693
rect 13742 8659 13776 8693
rect 13810 8659 13844 8693
rect 13878 8659 13912 8693
rect 13946 8659 13980 8693
rect 14014 8659 14048 8693
rect 14082 8659 14116 8693
rect 14150 8659 14184 8693
rect 14218 8659 14252 8693
rect 14286 8659 14320 8693
rect 14354 8659 14388 8693
rect 14422 8659 14456 8693
rect 14490 8659 14524 8693
rect 14558 8659 14592 8693
rect 14626 8659 14660 8693
rect 14694 8659 14728 8693
rect 14762 8659 14796 8693
rect 14830 8659 14864 8693
rect 14898 8687 14932 8693
rect 14966 8687 15000 8721
rect 15034 8687 15068 8721
rect 14898 8659 15102 8687
rect 42 8649 15102 8659
rect 42 8636 14932 8649
rect 42 8626 912 8636
rect 946 8626 984 8636
rect 1018 8626 1056 8636
rect 1090 8626 1128 8636
rect 1162 8626 1200 8636
rect 1234 8626 1272 8636
rect 1306 8626 1344 8636
rect 1378 8626 1416 8636
rect 1450 8626 1488 8636
rect 1522 8626 1560 8636
rect 1594 8626 1632 8636
rect 1666 8626 1704 8636
rect 1738 8626 1776 8636
rect 1810 8626 1849 8636
rect 1883 8626 1922 8636
rect 1956 8626 1995 8636
rect 2029 8626 2068 8636
rect 2102 8626 2141 8636
rect 2175 8630 3477 8636
rect 3511 8630 3550 8636
rect 3584 8630 3623 8636
rect 3657 8630 3696 8636
rect 3730 8630 3769 8636
rect 3803 8630 3842 8636
rect 3876 8630 3915 8636
rect 3949 8630 3988 8636
rect 4022 8630 4061 8636
rect 4095 8630 4134 8636
rect 4168 8630 4207 8636
rect 4241 8630 4280 8636
rect 4314 8630 4353 8636
rect 4387 8630 4426 8636
rect 4460 8630 4499 8636
rect 4533 8630 4572 8636
rect 4606 8630 4645 8636
rect 4679 8630 4718 8636
rect 4752 8630 4791 8636
rect 4825 8630 4864 8636
rect 4898 8630 4937 8636
rect 4971 8630 5010 8636
rect 5044 8630 5083 8636
rect 5117 8630 5156 8636
rect 5190 8630 5229 8636
rect 5263 8630 5302 8636
rect 5336 8630 5375 8636
rect 5409 8630 5448 8636
rect 5482 8630 5521 8636
rect 5555 8630 5594 8636
rect 5628 8630 5667 8636
rect 5701 8630 5740 8636
rect 5774 8630 5813 8636
rect 5847 8630 5886 8636
rect 5920 8630 5959 8636
rect 5993 8630 6032 8636
rect 6066 8630 6105 8636
rect 6139 8630 6178 8636
rect 6212 8630 6251 8636
rect 6285 8630 6324 8636
rect 6358 8630 6397 8636
rect 6431 8630 6470 8636
rect 6504 8630 6543 8636
rect 6577 8630 6616 8636
rect 6650 8630 6689 8636
rect 6723 8630 6762 8636
rect 6796 8630 6835 8636
rect 6869 8630 6908 8636
rect 6942 8630 6981 8636
rect 2175 8626 2933 8630
rect 42 8592 68 8626
rect 102 8592 138 8626
rect 172 8592 208 8626
rect 242 8592 278 8626
rect 312 8592 348 8626
rect 382 8592 418 8626
rect 452 8592 488 8626
rect 522 8592 558 8626
rect 592 8592 628 8626
rect 662 8592 698 8626
rect 732 8592 768 8626
rect 802 8592 838 8626
rect 872 8592 908 8626
rect 946 8602 978 8626
rect 1018 8602 1048 8626
rect 1090 8602 1118 8626
rect 1162 8602 1188 8626
rect 1234 8602 1258 8626
rect 1306 8602 1328 8626
rect 1378 8602 1398 8626
rect 1450 8602 1467 8626
rect 1522 8602 1536 8626
rect 1594 8602 1605 8626
rect 1666 8602 1674 8626
rect 1738 8602 1743 8626
rect 1810 8602 1812 8626
rect 942 8592 978 8602
rect 1012 8592 1048 8602
rect 1082 8592 1118 8602
rect 1152 8592 1188 8602
rect 1222 8592 1258 8602
rect 1292 8592 1328 8602
rect 1362 8592 1398 8602
rect 1432 8592 1467 8602
rect 1501 8592 1536 8602
rect 1570 8592 1605 8602
rect 1639 8592 1674 8602
rect 1708 8592 1743 8602
rect 1777 8592 1812 8602
rect 1846 8602 1849 8626
rect 1915 8602 1922 8626
rect 1984 8602 1995 8626
rect 2053 8602 2068 8626
rect 2122 8602 2141 8626
rect 1846 8592 1881 8602
rect 1915 8592 1950 8602
rect 1984 8592 2019 8602
rect 2053 8592 2088 8602
rect 2122 8592 2157 8602
rect 2191 8592 2226 8626
rect 2260 8592 2295 8626
rect 2329 8592 2364 8626
rect 2398 8592 2433 8626
rect 2467 8592 2502 8626
rect 2536 8592 2571 8626
rect 2605 8592 2640 8626
rect 2674 8592 2709 8626
rect 2743 8592 2778 8626
rect 2812 8592 2847 8626
rect 2881 8596 2933 8626
rect 2967 8596 3002 8630
rect 3036 8596 3071 8630
rect 3105 8596 3139 8630
rect 3173 8596 3207 8630
rect 3241 8596 3275 8630
rect 3309 8596 3343 8630
rect 3377 8596 3411 8630
rect 3445 8602 3477 8630
rect 3445 8596 3479 8602
rect 3513 8596 3547 8630
rect 3584 8602 3615 8630
rect 3657 8602 3683 8630
rect 3730 8602 3751 8630
rect 3803 8602 3819 8630
rect 3876 8602 3887 8630
rect 3949 8602 3955 8630
rect 4022 8602 4023 8630
rect 3581 8596 3615 8602
rect 3649 8596 3683 8602
rect 3717 8596 3751 8602
rect 3785 8596 3819 8602
rect 3853 8596 3887 8602
rect 3921 8596 3955 8602
rect 3989 8596 4023 8602
rect 4057 8602 4061 8630
rect 4125 8602 4134 8630
rect 4193 8602 4207 8630
rect 4261 8602 4280 8630
rect 4329 8602 4353 8630
rect 4397 8602 4426 8630
rect 4057 8596 4091 8602
rect 4125 8596 4159 8602
rect 4193 8596 4227 8602
rect 4261 8596 4295 8602
rect 4329 8596 4363 8602
rect 4397 8596 4431 8602
rect 4465 8596 4499 8630
rect 4533 8596 4567 8630
rect 4606 8602 4635 8630
rect 4679 8602 4703 8630
rect 4752 8602 4771 8630
rect 4825 8602 4839 8630
rect 4898 8602 4907 8630
rect 4971 8602 4975 8630
rect 4601 8596 4635 8602
rect 4669 8596 4703 8602
rect 4737 8596 4771 8602
rect 4805 8596 4839 8602
rect 4873 8596 4907 8602
rect 4941 8596 4975 8602
rect 5009 8602 5010 8630
rect 5077 8602 5083 8630
rect 5145 8602 5156 8630
rect 5213 8602 5229 8630
rect 5281 8602 5302 8630
rect 5349 8602 5375 8630
rect 5417 8602 5448 8630
rect 5009 8596 5043 8602
rect 5077 8596 5111 8602
rect 5145 8596 5179 8602
rect 5213 8596 5247 8602
rect 5281 8596 5315 8602
rect 5349 8596 5383 8602
rect 5417 8596 5451 8602
rect 5485 8596 5519 8630
rect 5555 8602 5587 8630
rect 5628 8602 5655 8630
rect 5701 8602 5723 8630
rect 5774 8602 5791 8630
rect 5847 8602 5859 8630
rect 5920 8602 5927 8630
rect 5993 8602 5995 8630
rect 5553 8596 5587 8602
rect 5621 8596 5655 8602
rect 5689 8596 5723 8602
rect 5757 8596 5791 8602
rect 5825 8596 5859 8602
rect 5893 8596 5927 8602
rect 5961 8596 5995 8602
rect 6029 8602 6032 8630
rect 6097 8602 6105 8630
rect 6165 8602 6178 8630
rect 6233 8602 6251 8630
rect 6301 8602 6324 8630
rect 6369 8602 6397 8630
rect 6437 8602 6470 8630
rect 6029 8596 6063 8602
rect 6097 8596 6131 8602
rect 6165 8596 6199 8602
rect 6233 8596 6267 8602
rect 6301 8596 6335 8602
rect 6369 8596 6403 8602
rect 6437 8596 6471 8602
rect 6505 8596 6539 8630
rect 6577 8602 6607 8630
rect 6650 8602 6675 8630
rect 6723 8602 6743 8630
rect 6796 8602 6811 8630
rect 6869 8602 6879 8630
rect 6942 8602 6947 8630
rect 6573 8596 6607 8602
rect 6641 8596 6675 8602
rect 6709 8596 6743 8602
rect 6777 8596 6811 8602
rect 6845 8596 6879 8602
rect 6913 8596 6947 8602
rect 7015 8630 7054 8636
rect 7088 8630 7127 8636
rect 7161 8630 7200 8636
rect 7234 8630 7273 8636
rect 7307 8630 7346 8636
rect 7380 8630 7419 8636
rect 7453 8630 7492 8636
rect 7526 8630 7565 8636
rect 7599 8630 7638 8636
rect 7672 8630 7711 8636
rect 7745 8630 7784 8636
rect 7818 8630 7857 8636
rect 7891 8630 7930 8636
rect 7964 8630 8003 8636
rect 8037 8630 8075 8636
rect 8109 8630 8147 8636
rect 8181 8630 8219 8636
rect 8253 8630 8291 8636
rect 8325 8630 8363 8636
rect 6981 8596 7015 8602
rect 7049 8602 7054 8630
rect 7117 8602 7127 8630
rect 7185 8602 7200 8630
rect 7253 8602 7273 8630
rect 7321 8602 7346 8630
rect 7389 8602 7419 8630
rect 7049 8596 7083 8602
rect 7117 8596 7151 8602
rect 7185 8596 7219 8602
rect 7253 8596 7287 8602
rect 7321 8596 7355 8602
rect 7389 8596 7423 8602
rect 7457 8596 7491 8630
rect 7526 8602 7559 8630
rect 7599 8602 7627 8630
rect 7672 8602 7695 8630
rect 7745 8602 7763 8630
rect 7818 8602 7831 8630
rect 7891 8602 7899 8630
rect 7964 8602 7967 8630
rect 7525 8596 7559 8602
rect 7593 8596 7627 8602
rect 7661 8596 7695 8602
rect 7729 8596 7763 8602
rect 7797 8596 7831 8602
rect 7865 8596 7899 8602
rect 7933 8596 7967 8602
rect 8001 8602 8003 8630
rect 8069 8602 8075 8630
rect 8137 8602 8147 8630
rect 8205 8602 8219 8630
rect 8273 8602 8291 8630
rect 8341 8602 8363 8630
rect 8397 8613 8435 8636
rect 8469 8613 8507 8636
rect 8541 8613 8579 8636
rect 8613 8613 8651 8636
rect 8685 8613 8723 8636
rect 8757 8613 8795 8636
rect 8829 8613 8867 8636
rect 8901 8613 8939 8636
rect 8973 8613 9011 8636
rect 9045 8613 9083 8636
rect 9117 8613 9155 8636
rect 9189 8613 9227 8636
rect 9261 8613 9299 8636
rect 9333 8613 9371 8636
rect 9405 8613 9443 8636
rect 9477 8613 9515 8636
rect 9549 8613 9587 8636
rect 9621 8613 9659 8636
rect 9693 8613 9731 8636
rect 9765 8613 9803 8636
rect 9837 8613 9875 8636
rect 9909 8613 9947 8636
rect 9981 8613 10019 8636
rect 10053 8613 10091 8636
rect 10125 8613 10163 8636
rect 10197 8613 10235 8636
rect 10269 8613 10307 8636
rect 10341 8613 10379 8636
rect 10413 8613 10451 8636
rect 10485 8613 10523 8636
rect 10557 8613 10595 8636
rect 10629 8613 10667 8636
rect 10701 8613 10739 8636
rect 10773 8613 10811 8636
rect 10845 8613 10883 8636
rect 10917 8613 10955 8636
rect 10989 8613 11027 8636
rect 11061 8613 11099 8636
rect 11133 8613 11171 8636
rect 11205 8613 11243 8636
rect 11277 8613 11315 8636
rect 11349 8613 11387 8636
rect 11421 8613 11459 8636
rect 11493 8613 11531 8636
rect 11565 8613 11603 8636
rect 11637 8613 11675 8636
rect 11709 8613 11747 8636
rect 11781 8613 11819 8636
rect 11853 8613 11891 8636
rect 11925 8613 11963 8636
rect 11997 8613 12035 8636
rect 12069 8613 12107 8636
rect 12141 8613 12179 8636
rect 12213 8613 12251 8636
rect 12285 8613 12323 8636
rect 12357 8613 12395 8636
rect 12429 8613 12467 8636
rect 12501 8613 12539 8636
rect 12573 8613 12611 8636
rect 12645 8613 12683 8636
rect 12717 8613 12755 8636
rect 12789 8613 12827 8636
rect 12861 8613 12899 8636
rect 12933 8613 12971 8636
rect 13005 8613 13043 8636
rect 13077 8613 13115 8636
rect 13149 8613 13187 8636
rect 13221 8613 13259 8636
rect 13293 8613 13331 8636
rect 13365 8613 13403 8636
rect 13437 8613 13475 8636
rect 13509 8613 13547 8636
rect 13581 8613 13619 8636
rect 13653 8613 13691 8636
rect 13725 8613 13763 8636
rect 13797 8613 13835 8636
rect 13869 8613 13907 8636
rect 13941 8613 13979 8636
rect 14013 8613 14051 8636
rect 14085 8613 14123 8636
rect 14157 8613 14195 8636
rect 14229 8613 14267 8636
rect 14301 8613 14339 8636
rect 14373 8613 14411 8636
rect 14445 8613 14483 8636
rect 14517 8613 14555 8636
rect 14589 8613 14627 8636
rect 14661 8613 14699 8636
rect 14733 8613 14771 8636
rect 14805 8613 14843 8636
rect 14877 8615 14932 8636
rect 14966 8615 15000 8649
rect 15034 8615 15068 8649
rect 14877 8613 15102 8615
rect 8427 8602 8435 8613
rect 8496 8602 8507 8613
rect 8565 8602 8579 8613
rect 8634 8602 8651 8613
rect 8703 8602 8723 8613
rect 8772 8602 8795 8613
rect 8841 8602 8867 8613
rect 8910 8602 8939 8613
rect 8979 8602 9011 8613
rect 8001 8596 8035 8602
rect 8069 8596 8103 8602
rect 8137 8596 8171 8602
rect 8205 8596 8239 8602
rect 8273 8596 8307 8602
rect 8341 8596 8393 8602
rect 2881 8592 8393 8596
rect 42 8579 8393 8592
rect 8427 8579 8462 8602
rect 8496 8579 8531 8602
rect 8565 8579 8600 8602
rect 8634 8579 8669 8602
rect 8703 8579 8738 8602
rect 8772 8579 8807 8602
rect 8841 8579 8876 8602
rect 8910 8579 8945 8602
rect 8979 8579 9014 8602
rect 9048 8579 9083 8613
rect 9117 8579 9152 8613
rect 9189 8602 9220 8613
rect 9261 8602 9288 8613
rect 9333 8602 9356 8613
rect 9405 8602 9424 8613
rect 9477 8602 9492 8613
rect 9549 8602 9560 8613
rect 9621 8602 9628 8613
rect 9693 8602 9696 8613
rect 9186 8579 9220 8602
rect 9254 8579 9288 8602
rect 9322 8579 9356 8602
rect 9390 8579 9424 8602
rect 9458 8579 9492 8602
rect 9526 8579 9560 8602
rect 9594 8579 9628 8602
rect 9662 8579 9696 8602
rect 9730 8602 9731 8613
rect 9798 8602 9803 8613
rect 9866 8602 9875 8613
rect 9934 8602 9947 8613
rect 10002 8602 10019 8613
rect 10070 8602 10091 8613
rect 10138 8602 10163 8613
rect 10206 8602 10235 8613
rect 10274 8602 10307 8613
rect 9730 8579 9764 8602
rect 9798 8579 9832 8602
rect 9866 8579 9900 8602
rect 9934 8579 9968 8602
rect 10002 8579 10036 8602
rect 10070 8579 10104 8602
rect 10138 8579 10172 8602
rect 10206 8579 10240 8602
rect 10274 8579 10308 8602
rect 10342 8579 10376 8613
rect 10413 8602 10444 8613
rect 10485 8602 10512 8613
rect 10557 8602 10580 8613
rect 10629 8602 10648 8613
rect 10701 8602 10716 8613
rect 10773 8602 10784 8613
rect 10845 8602 10852 8613
rect 10917 8602 10920 8613
rect 10410 8579 10444 8602
rect 10478 8579 10512 8602
rect 10546 8579 10580 8602
rect 10614 8579 10648 8602
rect 10682 8579 10716 8602
rect 10750 8579 10784 8602
rect 10818 8579 10852 8602
rect 10886 8579 10920 8602
rect 10954 8602 10955 8613
rect 11022 8602 11027 8613
rect 11090 8602 11099 8613
rect 11158 8602 11171 8613
rect 11226 8602 11243 8613
rect 11294 8602 11315 8613
rect 11362 8602 11387 8613
rect 11430 8602 11459 8613
rect 11498 8602 11531 8613
rect 10954 8579 10988 8602
rect 11022 8579 11056 8602
rect 11090 8579 11124 8602
rect 11158 8579 11192 8602
rect 11226 8579 11260 8602
rect 11294 8579 11328 8602
rect 11362 8579 11396 8602
rect 11430 8579 11464 8602
rect 11498 8579 11532 8602
rect 11566 8579 11600 8613
rect 11637 8602 11668 8613
rect 11709 8602 11736 8613
rect 11781 8602 11804 8613
rect 11853 8602 11872 8613
rect 11925 8602 11940 8613
rect 11997 8602 12008 8613
rect 12069 8602 12076 8613
rect 12141 8602 12144 8613
rect 11634 8579 11668 8602
rect 11702 8579 11736 8602
rect 11770 8579 11804 8602
rect 11838 8579 11872 8602
rect 11906 8579 11940 8602
rect 11974 8579 12008 8602
rect 12042 8579 12076 8602
rect 12110 8579 12144 8602
rect 12178 8602 12179 8613
rect 12246 8602 12251 8613
rect 12314 8602 12323 8613
rect 12382 8602 12395 8613
rect 12450 8602 12467 8613
rect 12518 8602 12539 8613
rect 12586 8602 12611 8613
rect 12654 8602 12683 8613
rect 12722 8602 12755 8613
rect 12178 8579 12212 8602
rect 12246 8579 12280 8602
rect 12314 8579 12348 8602
rect 12382 8579 12416 8602
rect 12450 8579 12484 8602
rect 12518 8579 12552 8602
rect 12586 8579 12620 8602
rect 12654 8579 12688 8602
rect 12722 8579 12756 8602
rect 12790 8579 12824 8613
rect 12861 8602 12892 8613
rect 12933 8602 12960 8613
rect 13005 8602 13028 8613
rect 13077 8602 13096 8613
rect 13149 8602 13164 8613
rect 13221 8602 13232 8613
rect 13293 8602 13300 8613
rect 13365 8602 13368 8613
rect 12858 8579 12892 8602
rect 12926 8579 12960 8602
rect 12994 8579 13028 8602
rect 13062 8579 13096 8602
rect 13130 8579 13164 8602
rect 13198 8579 13232 8602
rect 13266 8579 13300 8602
rect 13334 8579 13368 8602
rect 13402 8602 13403 8613
rect 13470 8602 13475 8613
rect 13538 8602 13547 8613
rect 13606 8602 13619 8613
rect 13674 8602 13691 8613
rect 13742 8602 13763 8613
rect 13810 8602 13835 8613
rect 13878 8602 13907 8613
rect 13946 8602 13979 8613
rect 13402 8579 13436 8602
rect 13470 8579 13504 8602
rect 13538 8579 13572 8602
rect 13606 8579 13640 8602
rect 13674 8579 13708 8602
rect 13742 8579 13776 8602
rect 13810 8579 13844 8602
rect 13878 8579 13912 8602
rect 13946 8579 13980 8602
rect 14014 8579 14048 8613
rect 14085 8602 14116 8613
rect 14157 8602 14184 8613
rect 14229 8602 14252 8613
rect 14301 8602 14320 8613
rect 14373 8602 14388 8613
rect 14445 8602 14456 8613
rect 14517 8602 14524 8613
rect 14589 8602 14592 8613
rect 14082 8579 14116 8602
rect 14150 8579 14184 8602
rect 14218 8579 14252 8602
rect 14286 8579 14320 8602
rect 14354 8579 14388 8602
rect 14422 8579 14456 8602
rect 14490 8579 14524 8602
rect 14558 8579 14592 8602
rect 14626 8602 14627 8613
rect 14694 8602 14699 8613
rect 14762 8602 14771 8613
rect 14830 8602 14843 8613
rect 14626 8579 14660 8602
rect 14694 8579 14728 8602
rect 14762 8579 14796 8602
rect 14830 8579 14864 8602
rect 14898 8579 15102 8613
rect 42 8577 15102 8579
rect 42 8560 14932 8577
rect 42 8552 2933 8560
rect 42 8518 68 8552
rect 102 8518 138 8552
rect 172 8518 208 8552
rect 242 8518 278 8552
rect 312 8518 348 8552
rect 382 8518 418 8552
rect 452 8518 488 8552
rect 522 8518 558 8552
rect 592 8518 628 8552
rect 662 8518 698 8552
rect 732 8518 768 8552
rect 802 8518 838 8552
rect 872 8518 908 8552
rect 942 8518 978 8552
rect 1012 8518 1048 8552
rect 1082 8518 1118 8552
rect 1152 8518 1188 8552
rect 1222 8518 1258 8552
rect 1292 8518 1328 8552
rect 1362 8518 1398 8552
rect 1432 8518 1467 8552
rect 1501 8518 1536 8552
rect 1570 8518 1605 8552
rect 1639 8518 1674 8552
rect 1708 8518 1743 8552
rect 1777 8518 1812 8552
rect 1846 8518 1881 8552
rect 1915 8518 1950 8552
rect 1984 8518 2019 8552
rect 2053 8518 2088 8552
rect 2122 8518 2157 8552
rect 2191 8518 2226 8552
rect 2260 8518 2295 8552
rect 2329 8518 2364 8552
rect 2398 8518 2433 8552
rect 2467 8518 2502 8552
rect 2536 8518 2571 8552
rect 2605 8518 2640 8552
rect 2674 8518 2709 8552
rect 2743 8518 2778 8552
rect 2812 8518 2847 8552
rect 2881 8526 2933 8552
rect 2967 8526 3002 8560
rect 3036 8526 3071 8560
rect 3105 8526 3139 8560
rect 3173 8526 3207 8560
rect 3241 8526 3275 8560
rect 3309 8526 3343 8560
rect 3377 8526 3411 8560
rect 3445 8526 3479 8560
rect 3513 8526 3547 8560
rect 3581 8526 3615 8560
rect 3649 8526 3683 8560
rect 3717 8526 3751 8560
rect 3785 8526 3819 8560
rect 3853 8526 3887 8560
rect 3921 8526 3955 8560
rect 3989 8526 4023 8560
rect 4057 8526 4091 8560
rect 4125 8526 4159 8560
rect 4193 8526 4227 8560
rect 4261 8526 4295 8560
rect 4329 8526 4363 8560
rect 4397 8526 4431 8560
rect 4465 8526 4499 8560
rect 4533 8526 4567 8560
rect 4601 8526 4635 8560
rect 4669 8526 4703 8560
rect 4737 8526 4771 8560
rect 4805 8526 4839 8560
rect 4873 8526 4907 8560
rect 4941 8526 4975 8560
rect 5009 8526 5043 8560
rect 5077 8526 5111 8560
rect 5145 8526 5179 8560
rect 5213 8526 5247 8560
rect 5281 8526 5315 8560
rect 5349 8526 5383 8560
rect 5417 8526 5451 8560
rect 5485 8526 5519 8560
rect 5553 8526 5587 8560
rect 5621 8526 5655 8560
rect 5689 8526 5723 8560
rect 5757 8526 5791 8560
rect 5825 8526 5859 8560
rect 5893 8526 5927 8560
rect 5961 8526 5995 8560
rect 6029 8526 6063 8560
rect 6097 8526 6131 8560
rect 6165 8526 6199 8560
rect 6233 8526 6267 8560
rect 6301 8526 6335 8560
rect 6369 8526 6403 8560
rect 6437 8526 6471 8560
rect 6505 8526 6539 8560
rect 6573 8526 6607 8560
rect 6641 8526 6675 8560
rect 6709 8526 6743 8560
rect 6777 8526 6811 8560
rect 6845 8526 6879 8560
rect 6913 8526 6947 8560
rect 6981 8526 7015 8560
rect 7049 8526 7083 8560
rect 7117 8526 7151 8560
rect 7185 8526 7219 8560
rect 7253 8526 7287 8560
rect 7321 8526 7355 8560
rect 7389 8526 7423 8560
rect 7457 8526 7491 8560
rect 7525 8526 7559 8560
rect 7593 8526 7627 8560
rect 7661 8526 7695 8560
rect 7729 8526 7763 8560
rect 7797 8526 7831 8560
rect 7865 8526 7899 8560
rect 7933 8526 7967 8560
rect 8001 8526 8035 8560
rect 8069 8526 8103 8560
rect 8137 8526 8171 8560
rect 8205 8526 8239 8560
rect 8273 8526 8307 8560
rect 8341 8546 14932 8560
rect 8341 8533 13992 8546
rect 14026 8533 14076 8546
rect 14110 8543 14932 8546
rect 14966 8543 15000 8577
rect 15034 8543 15068 8577
rect 14110 8533 15102 8543
rect 8341 8526 8393 8533
rect 2881 8518 8393 8526
rect 42 8499 8393 8518
rect 8427 8499 8462 8533
rect 8496 8499 8531 8533
rect 8565 8499 8600 8533
rect 8634 8499 8669 8533
rect 8703 8499 8738 8533
rect 8772 8499 8807 8533
rect 8841 8499 8876 8533
rect 8910 8499 8945 8533
rect 8979 8499 9014 8533
rect 9048 8499 9083 8533
rect 9117 8499 9152 8533
rect 9186 8499 9220 8533
rect 9254 8499 9288 8533
rect 9322 8499 9356 8533
rect 9390 8499 9424 8533
rect 9458 8499 9492 8533
rect 9526 8499 9560 8533
rect 9594 8499 9628 8533
rect 9662 8499 9696 8533
rect 9730 8499 9764 8533
rect 9798 8499 9832 8533
rect 9866 8499 9900 8533
rect 9934 8499 9968 8533
rect 10002 8499 10036 8533
rect 10070 8499 10104 8533
rect 10138 8499 10172 8533
rect 10206 8499 10240 8533
rect 10274 8499 10308 8533
rect 10342 8499 10376 8533
rect 10410 8499 10444 8533
rect 10478 8499 10512 8533
rect 10546 8499 10580 8533
rect 10614 8499 10648 8533
rect 10682 8499 10716 8533
rect 10750 8499 10784 8533
rect 10818 8499 10852 8533
rect 10886 8499 10920 8533
rect 10954 8499 10988 8533
rect 11022 8499 11056 8533
rect 11090 8499 11124 8533
rect 11158 8499 11192 8533
rect 11226 8499 11260 8533
rect 11294 8499 11328 8533
rect 11362 8499 11396 8533
rect 11430 8499 11464 8533
rect 11498 8499 11532 8533
rect 11566 8499 11600 8533
rect 11634 8499 11668 8533
rect 11702 8499 11736 8533
rect 11770 8499 11804 8533
rect 11838 8499 11872 8533
rect 11906 8499 11940 8533
rect 11974 8499 12008 8533
rect 12042 8499 12076 8533
rect 12110 8499 12144 8533
rect 12178 8499 12212 8533
rect 12246 8499 12280 8533
rect 12314 8499 12348 8533
rect 12382 8499 12416 8533
rect 12450 8499 12484 8533
rect 12518 8499 12552 8533
rect 12586 8499 12620 8533
rect 12654 8499 12688 8533
rect 12722 8499 12756 8533
rect 12790 8499 12824 8533
rect 12858 8499 12892 8533
rect 12926 8499 12960 8533
rect 12994 8499 13028 8533
rect 13062 8499 13096 8533
rect 13130 8499 13164 8533
rect 13198 8499 13232 8533
rect 13266 8499 13300 8533
rect 13334 8499 13368 8533
rect 13402 8499 13436 8533
rect 13470 8499 13504 8533
rect 13538 8499 13572 8533
rect 13606 8499 13640 8533
rect 13674 8499 13708 8533
rect 13742 8499 13776 8533
rect 13810 8499 13844 8533
rect 13878 8499 13912 8533
rect 13946 8499 13980 8533
rect 14026 8512 14048 8533
rect 14110 8512 14116 8533
rect 14014 8499 14048 8512
rect 14082 8499 14116 8512
rect 14150 8499 14184 8533
rect 14218 8512 14252 8533
rect 14286 8512 14320 8533
rect 14354 8512 14388 8533
rect 14422 8512 14456 8533
rect 14490 8512 14524 8533
rect 14219 8499 14252 8512
rect 14291 8499 14320 8512
rect 14363 8499 14388 8512
rect 14435 8499 14456 8512
rect 14507 8499 14524 8512
rect 14558 8499 14592 8533
rect 14626 8499 14660 8533
rect 14694 8499 14728 8533
rect 14762 8499 14796 8533
rect 14830 8499 14864 8533
rect 14898 8505 15102 8533
rect 14898 8499 14932 8505
rect 42 8490 14185 8499
rect 42 8484 2933 8490
rect 34 8460 136 8484
rect 34 8426 68 8460
rect 102 8426 136 8460
rect 34 8392 136 8426
rect 34 8358 68 8392
rect 102 8358 136 8392
rect 34 8324 136 8358
rect 34 8290 68 8324
rect 102 8290 136 8324
rect 34 8256 136 8290
rect 34 8222 68 8256
rect 102 8222 136 8256
rect 34 8192 136 8222
rect 2907 8456 2933 8484
rect 2967 8456 3002 8490
rect 3036 8456 3071 8490
rect 3105 8456 3139 8490
rect 3173 8456 3207 8490
rect 3241 8456 3275 8490
rect 3309 8456 3343 8490
rect 3377 8456 3411 8490
rect 3445 8456 3479 8490
rect 3513 8456 3547 8490
rect 3581 8456 3615 8490
rect 3649 8456 3683 8490
rect 3717 8456 3751 8490
rect 3785 8456 3819 8490
rect 3853 8456 3887 8490
rect 3921 8456 3955 8490
rect 3989 8456 4023 8490
rect 4057 8456 4091 8490
rect 4125 8456 4159 8490
rect 4193 8456 4227 8490
rect 4261 8456 4295 8490
rect 4329 8456 4363 8490
rect 4397 8456 4431 8490
rect 4465 8456 4499 8490
rect 4533 8456 4567 8490
rect 4601 8456 4635 8490
rect 4669 8456 4703 8490
rect 4737 8456 4771 8490
rect 4805 8456 4839 8490
rect 4873 8456 4907 8490
rect 4941 8456 4975 8490
rect 5009 8456 5043 8490
rect 5077 8456 5111 8490
rect 5145 8456 5179 8490
rect 5213 8456 5247 8490
rect 5281 8456 5315 8490
rect 5349 8456 5383 8490
rect 5417 8456 5451 8490
rect 5485 8456 5519 8490
rect 5553 8456 5587 8490
rect 5621 8456 5655 8490
rect 5689 8456 5723 8490
rect 5757 8456 5791 8490
rect 5825 8456 5859 8490
rect 5893 8456 5927 8490
rect 5961 8456 5995 8490
rect 6029 8456 6063 8490
rect 6097 8456 6131 8490
rect 6165 8456 6199 8490
rect 6233 8456 6267 8490
rect 6301 8456 6335 8490
rect 6369 8456 6403 8490
rect 6437 8456 6471 8490
rect 6505 8456 6539 8490
rect 6573 8456 6607 8490
rect 6641 8456 6675 8490
rect 6709 8456 6743 8490
rect 6777 8456 6811 8490
rect 6845 8456 6879 8490
rect 6913 8456 6947 8490
rect 6981 8456 7015 8490
rect 7049 8456 7083 8490
rect 7117 8456 7151 8490
rect 7185 8456 7219 8490
rect 7253 8456 7287 8490
rect 7321 8456 7355 8490
rect 7389 8456 7423 8490
rect 7457 8456 7491 8490
rect 7525 8456 7559 8490
rect 7593 8456 7627 8490
rect 7661 8456 7695 8490
rect 7729 8456 7763 8490
rect 7797 8456 7831 8490
rect 7865 8456 7899 8490
rect 7933 8456 7967 8490
rect 8001 8456 8035 8490
rect 8069 8456 8103 8490
rect 8137 8456 8171 8490
rect 8205 8456 8239 8490
rect 8273 8456 8307 8490
rect 8341 8478 14185 8490
rect 14219 8478 14257 8499
rect 14291 8478 14329 8499
rect 14363 8478 14401 8499
rect 14435 8478 14473 8499
rect 14507 8478 14932 8499
rect 8341 8474 14932 8478
rect 8341 8456 13992 8474
rect 2907 8453 13992 8456
rect 14026 8453 14076 8474
rect 14110 8471 14932 8474
rect 14966 8471 15000 8505
rect 15034 8471 15068 8505
rect 14110 8462 15102 8471
rect 14110 8453 14614 8462
rect 14648 8453 14692 8462
rect 14726 8453 14770 8462
rect 14804 8453 14848 8462
rect 14882 8453 14926 8462
rect 2907 8420 8393 8453
rect 2907 8386 2933 8420
rect 2967 8386 3002 8420
rect 3036 8386 3071 8420
rect 3105 8386 3139 8420
rect 3173 8386 3207 8420
rect 3241 8386 3275 8420
rect 3309 8386 3343 8420
rect 3377 8386 3411 8420
rect 3445 8386 3479 8420
rect 3513 8386 3547 8420
rect 3581 8386 3615 8420
rect 3649 8386 3683 8420
rect 3717 8386 3751 8420
rect 3785 8386 3819 8420
rect 3853 8386 3887 8420
rect 3921 8386 3955 8420
rect 3989 8386 4023 8420
rect 4057 8386 4091 8420
rect 4125 8386 4159 8420
rect 4193 8386 4227 8420
rect 4261 8386 4295 8420
rect 4329 8386 4363 8420
rect 4397 8386 4431 8420
rect 4465 8386 4499 8420
rect 4533 8386 4567 8420
rect 4601 8386 4635 8420
rect 4669 8386 4703 8420
rect 4737 8386 4771 8420
rect 4805 8386 4839 8420
rect 4873 8386 4907 8420
rect 4941 8386 4975 8420
rect 5009 8386 5043 8420
rect 5077 8386 5111 8420
rect 5145 8386 5179 8420
rect 5213 8386 5247 8420
rect 5281 8386 5315 8420
rect 5349 8386 5383 8420
rect 5417 8386 5451 8420
rect 5485 8386 5519 8420
rect 5553 8386 5587 8420
rect 5621 8386 5655 8420
rect 5689 8386 5723 8420
rect 5757 8386 5791 8420
rect 5825 8386 5859 8420
rect 5893 8386 5927 8420
rect 5961 8386 5995 8420
rect 6029 8386 6063 8420
rect 6097 8386 6131 8420
rect 6165 8386 6199 8420
rect 6233 8386 6267 8420
rect 6301 8386 6335 8420
rect 6369 8386 6403 8420
rect 6437 8386 6471 8420
rect 6505 8386 6539 8420
rect 6573 8386 6607 8420
rect 6641 8386 6675 8420
rect 6709 8386 6743 8420
rect 6777 8386 6811 8420
rect 6845 8386 6879 8420
rect 6913 8386 6947 8420
rect 6981 8386 7015 8420
rect 7049 8386 7083 8420
rect 7117 8386 7151 8420
rect 7185 8386 7219 8420
rect 7253 8386 7287 8420
rect 7321 8386 7355 8420
rect 7389 8386 7423 8420
rect 7457 8386 7491 8420
rect 7525 8386 7559 8420
rect 7593 8386 7627 8420
rect 7661 8386 7695 8420
rect 7729 8386 7763 8420
rect 7797 8386 7831 8420
rect 7865 8386 7899 8420
rect 7933 8386 7967 8420
rect 8001 8386 8035 8420
rect 8069 8386 8103 8420
rect 8137 8386 8171 8420
rect 8205 8386 8239 8420
rect 8273 8386 8307 8420
rect 8341 8419 8393 8420
rect 8427 8419 8462 8453
rect 8496 8419 8531 8453
rect 8565 8419 8600 8453
rect 8634 8419 8669 8453
rect 8703 8419 8738 8453
rect 8772 8419 8807 8453
rect 8841 8419 8876 8453
rect 8910 8419 8945 8453
rect 8979 8419 9014 8453
rect 9048 8419 9083 8453
rect 9117 8419 9152 8453
rect 9186 8419 9220 8453
rect 9254 8419 9288 8453
rect 9322 8419 9356 8453
rect 9390 8419 9424 8453
rect 9458 8419 9492 8453
rect 9526 8419 9560 8453
rect 9594 8419 9628 8453
rect 9662 8419 9696 8453
rect 9730 8419 9764 8453
rect 9798 8419 9832 8453
rect 9866 8419 9900 8453
rect 9934 8419 9968 8453
rect 10002 8419 10036 8453
rect 10070 8419 10104 8453
rect 10138 8419 10172 8453
rect 10206 8419 10240 8453
rect 10274 8419 10308 8453
rect 10342 8419 10376 8453
rect 10410 8419 10444 8453
rect 10478 8419 10512 8453
rect 10546 8419 10580 8453
rect 10614 8419 10648 8453
rect 10682 8419 10716 8453
rect 10750 8419 10784 8453
rect 10818 8419 10852 8453
rect 10886 8419 10920 8453
rect 10954 8419 10988 8453
rect 11022 8419 11056 8453
rect 11090 8419 11124 8453
rect 11158 8419 11192 8453
rect 11226 8419 11260 8453
rect 11294 8419 11328 8453
rect 11362 8419 11396 8453
rect 11430 8419 11464 8453
rect 11498 8419 11532 8453
rect 11566 8419 11600 8453
rect 11634 8419 11668 8453
rect 11702 8419 11736 8453
rect 11770 8419 11804 8453
rect 11838 8419 11872 8453
rect 11906 8419 11940 8453
rect 11974 8419 12008 8453
rect 12042 8419 12076 8453
rect 12110 8419 12144 8453
rect 12178 8419 12212 8453
rect 12246 8419 12280 8453
rect 12314 8419 12348 8453
rect 12382 8419 12416 8453
rect 12450 8419 12484 8453
rect 12518 8419 12552 8453
rect 12586 8419 12620 8453
rect 12654 8419 12688 8453
rect 12722 8419 12756 8453
rect 12790 8419 12824 8453
rect 12858 8419 12892 8453
rect 12926 8419 12960 8453
rect 12994 8419 13028 8453
rect 13062 8419 13096 8453
rect 13130 8419 13164 8453
rect 13198 8419 13232 8453
rect 13266 8419 13300 8453
rect 13334 8419 13368 8453
rect 13402 8419 13436 8453
rect 13470 8419 13504 8453
rect 13538 8419 13572 8453
rect 13606 8419 13640 8453
rect 13674 8419 13708 8453
rect 13742 8419 13776 8453
rect 13810 8419 13844 8453
rect 13878 8419 13912 8453
rect 13946 8419 13980 8453
rect 14026 8440 14048 8453
rect 14110 8440 14116 8453
rect 14014 8419 14048 8440
rect 14082 8419 14116 8440
rect 14150 8419 14184 8453
rect 14218 8435 14252 8453
rect 14286 8435 14320 8453
rect 14354 8435 14388 8453
rect 14422 8435 14456 8453
rect 14490 8435 14524 8453
rect 14219 8419 14252 8435
rect 14291 8419 14320 8435
rect 14363 8419 14388 8435
rect 14435 8419 14456 8435
rect 14507 8419 14524 8435
rect 14558 8419 14592 8453
rect 14648 8428 14660 8453
rect 14726 8428 14728 8453
rect 14626 8419 14660 8428
rect 14694 8419 14728 8428
rect 14762 8428 14770 8453
rect 14830 8428 14848 8453
rect 14898 8428 14926 8453
rect 14960 8433 15004 8462
rect 15038 8433 15102 8462
rect 14762 8419 14796 8428
rect 14830 8419 14864 8428
rect 14898 8419 14932 8428
rect 8341 8401 14185 8419
rect 14219 8401 14257 8419
rect 14291 8401 14329 8419
rect 14363 8401 14401 8419
rect 14435 8401 14473 8419
rect 14507 8401 14932 8419
rect 8341 8386 13992 8401
rect 2907 8383 13992 8386
rect 2907 8350 8367 8383
rect 2907 8316 2933 8350
rect 2967 8316 3002 8350
rect 3036 8316 3071 8350
rect 3105 8316 3139 8350
rect 3173 8316 3207 8350
rect 3241 8316 3275 8350
rect 3309 8316 3343 8350
rect 3377 8316 3411 8350
rect 3445 8316 3479 8350
rect 3513 8316 3547 8350
rect 3581 8316 3615 8350
rect 3649 8316 3683 8350
rect 3717 8316 3751 8350
rect 3785 8316 3819 8350
rect 3853 8316 3887 8350
rect 3921 8316 3955 8350
rect 3989 8316 4023 8350
rect 4057 8316 4091 8350
rect 4125 8316 4159 8350
rect 4193 8316 4227 8350
rect 4261 8316 4295 8350
rect 4329 8316 4363 8350
rect 4397 8316 4431 8350
rect 4465 8316 4499 8350
rect 4533 8316 4567 8350
rect 4601 8316 4635 8350
rect 4669 8316 4703 8350
rect 4737 8316 4771 8350
rect 4805 8316 4839 8350
rect 4873 8316 4907 8350
rect 4941 8316 4975 8350
rect 5009 8316 5043 8350
rect 5077 8316 5111 8350
rect 5145 8316 5179 8350
rect 5213 8316 5247 8350
rect 5281 8316 5315 8350
rect 5349 8316 5383 8350
rect 5417 8316 5451 8350
rect 5485 8316 5519 8350
rect 5553 8316 5587 8350
rect 5621 8316 5655 8350
rect 5689 8316 5723 8350
rect 5757 8316 5791 8350
rect 5825 8316 5859 8350
rect 5893 8316 5927 8350
rect 5961 8316 5995 8350
rect 6029 8316 6063 8350
rect 6097 8316 6131 8350
rect 6165 8316 6199 8350
rect 6233 8316 6267 8350
rect 6301 8316 6335 8350
rect 6369 8316 6403 8350
rect 6437 8316 6471 8350
rect 6505 8316 6539 8350
rect 6573 8316 6607 8350
rect 6641 8316 6675 8350
rect 6709 8316 6743 8350
rect 6777 8316 6811 8350
rect 6845 8316 6879 8350
rect 6913 8316 6947 8350
rect 6981 8316 7015 8350
rect 7049 8316 7083 8350
rect 7117 8316 7151 8350
rect 7185 8316 7219 8350
rect 7253 8316 7287 8350
rect 7321 8316 7355 8350
rect 7389 8316 7423 8350
rect 7457 8316 7491 8350
rect 7525 8316 7559 8350
rect 7593 8316 7627 8350
rect 7661 8316 7695 8350
rect 7729 8316 7763 8350
rect 7797 8316 7831 8350
rect 7865 8316 7899 8350
rect 7933 8316 7967 8350
rect 8001 8316 8035 8350
rect 8069 8316 8103 8350
rect 8137 8316 8171 8350
rect 8205 8316 8239 8350
rect 8273 8316 8307 8350
rect 8341 8316 8367 8350
rect 2907 8280 8367 8316
rect 2907 8246 2933 8280
rect 2967 8246 3002 8280
rect 3036 8246 3071 8280
rect 3105 8246 3139 8280
rect 3173 8246 3207 8280
rect 3241 8246 3275 8280
rect 3309 8246 3343 8280
rect 3377 8246 3411 8280
rect 3445 8246 3479 8280
rect 3513 8246 3547 8280
rect 3581 8246 3615 8280
rect 3649 8246 3683 8280
rect 3717 8246 3751 8280
rect 3785 8246 3819 8280
rect 3853 8246 3887 8280
rect 3921 8246 3955 8280
rect 3989 8246 4023 8280
rect 4057 8246 4091 8280
rect 4125 8246 4159 8280
rect 4193 8246 4227 8280
rect 4261 8246 4295 8280
rect 4329 8246 4363 8280
rect 4397 8246 4431 8280
rect 4465 8246 4499 8280
rect 4533 8246 4567 8280
rect 4601 8246 4635 8280
rect 4669 8246 4703 8280
rect 4737 8246 4771 8280
rect 4805 8246 4839 8280
rect 4873 8246 4907 8280
rect 4941 8246 4975 8280
rect 5009 8246 5043 8280
rect 5077 8246 5111 8280
rect 5145 8246 5179 8280
rect 5213 8246 5247 8280
rect 5281 8246 5315 8280
rect 5349 8246 5383 8280
rect 5417 8246 5451 8280
rect 5485 8246 5519 8280
rect 5553 8246 5587 8280
rect 5621 8246 5655 8280
rect 5689 8246 5723 8280
rect 5757 8246 5791 8280
rect 5825 8246 5859 8280
rect 5893 8246 5927 8280
rect 5961 8246 5995 8280
rect 6029 8246 6063 8280
rect 6097 8246 6131 8280
rect 6165 8246 6199 8280
rect 6233 8246 6267 8280
rect 6301 8246 6335 8280
rect 6369 8246 6403 8280
rect 6437 8246 6471 8280
rect 6505 8246 6539 8280
rect 6573 8246 6607 8280
rect 6641 8246 6675 8280
rect 6709 8246 6743 8280
rect 6777 8246 6811 8280
rect 6845 8246 6879 8280
rect 6913 8246 6947 8280
rect 6981 8246 7015 8280
rect 7049 8246 7083 8280
rect 7117 8246 7151 8280
rect 7185 8246 7219 8280
rect 7253 8246 7287 8280
rect 7321 8246 7355 8280
rect 7389 8246 7423 8280
rect 7457 8246 7491 8280
rect 7525 8246 7559 8280
rect 7593 8246 7627 8280
rect 7661 8246 7695 8280
rect 7729 8246 7763 8280
rect 7797 8246 7831 8280
rect 7865 8246 7899 8280
rect 7933 8246 7967 8280
rect 8001 8246 8035 8280
rect 8069 8246 8103 8280
rect 8137 8246 8171 8280
rect 8205 8246 8239 8280
rect 8273 8246 8307 8280
rect 8341 8246 8367 8280
rect 13506 8367 13992 8383
rect 14026 8367 14076 8401
rect 14110 8399 14932 8401
rect 14966 8399 15000 8433
rect 15038 8428 15068 8433
rect 15034 8399 15068 8428
rect 14110 8388 15102 8399
rect 14110 8367 14614 8388
rect 13506 8358 14614 8367
rect 13506 8357 14185 8358
rect 14219 8357 14257 8358
rect 14291 8357 14329 8358
rect 14363 8357 14401 8358
rect 14435 8357 14473 8358
rect 14507 8357 14614 8358
rect 14648 8357 14692 8388
rect 14726 8357 14770 8388
rect 14804 8357 14848 8388
rect 14882 8357 14926 8388
rect 14960 8361 15004 8388
rect 15038 8361 15102 8388
rect 13506 8323 13532 8357
rect 13566 8323 13603 8357
rect 13637 8323 13674 8357
rect 13708 8323 13744 8357
rect 13778 8323 13814 8357
rect 13848 8323 13884 8357
rect 13918 8323 13954 8357
rect 13988 8323 14024 8357
rect 14058 8323 14094 8357
rect 14128 8323 14164 8357
rect 14219 8324 14234 8357
rect 14291 8324 14304 8357
rect 14363 8324 14374 8357
rect 14435 8324 14444 8357
rect 14507 8324 14514 8357
rect 14198 8323 14234 8324
rect 14268 8323 14304 8324
rect 14338 8323 14374 8324
rect 14408 8323 14444 8324
rect 14478 8323 14514 8324
rect 14548 8323 14584 8357
rect 14648 8354 14654 8357
rect 14618 8323 14654 8354
rect 14688 8354 14692 8357
rect 14758 8354 14770 8357
rect 14828 8354 14848 8357
rect 14898 8354 14926 8357
rect 14688 8323 14724 8354
rect 14758 8323 14794 8354
rect 14828 8323 14864 8354
rect 14898 8327 14932 8354
rect 14966 8327 15000 8361
rect 15038 8354 15068 8361
rect 15034 8327 15068 8354
rect 14898 8323 15102 8327
rect 13506 8314 15102 8323
rect 13506 8283 14614 8314
rect 14648 8283 14692 8314
rect 14726 8283 14770 8314
rect 14804 8283 14848 8314
rect 14882 8283 14926 8314
rect 14960 8289 15004 8314
rect 15038 8289 15102 8314
rect 2907 8210 8367 8246
rect 2907 8192 2933 8210
rect 42 8176 2933 8192
rect 2967 8176 3002 8210
rect 3036 8176 3071 8210
rect 3105 8176 3139 8210
rect 3173 8176 3207 8210
rect 3241 8176 3275 8210
rect 3309 8176 3343 8210
rect 3377 8176 3411 8210
rect 3445 8176 3479 8210
rect 3513 8176 3547 8210
rect 3581 8176 3615 8210
rect 3649 8176 3683 8210
rect 3717 8176 3751 8210
rect 3785 8176 3819 8210
rect 3853 8176 3887 8210
rect 3921 8176 3955 8210
rect 3989 8176 4023 8210
rect 4057 8176 4091 8210
rect 4125 8176 4159 8210
rect 4193 8176 4227 8210
rect 4261 8176 4295 8210
rect 4329 8176 4363 8210
rect 4397 8176 4431 8210
rect 4465 8176 4499 8210
rect 4533 8176 4567 8210
rect 4601 8176 4635 8210
rect 4669 8176 4703 8210
rect 4737 8176 4771 8210
rect 4805 8176 4839 8210
rect 4873 8176 4907 8210
rect 4941 8176 4975 8210
rect 5009 8176 5043 8210
rect 5077 8176 5111 8210
rect 5145 8176 5179 8210
rect 5213 8176 5247 8210
rect 5281 8176 5315 8210
rect 5349 8176 5383 8210
rect 5417 8176 5451 8210
rect 5485 8176 5519 8210
rect 5553 8176 5587 8210
rect 5621 8176 5655 8210
rect 5689 8176 5723 8210
rect 5757 8176 5791 8210
rect 5825 8176 5859 8210
rect 5893 8176 5927 8210
rect 5961 8176 5995 8210
rect 6029 8176 6063 8210
rect 6097 8176 6131 8210
rect 6165 8176 6199 8210
rect 6233 8176 6267 8210
rect 6301 8176 6335 8210
rect 6369 8176 6403 8210
rect 6437 8176 6471 8210
rect 6505 8176 6539 8210
rect 6573 8176 6607 8210
rect 6641 8176 6675 8210
rect 6709 8176 6743 8210
rect 6777 8176 6811 8210
rect 6845 8176 6879 8210
rect 6913 8176 6947 8210
rect 6981 8176 7015 8210
rect 7049 8176 7083 8210
rect 7117 8176 7151 8210
rect 7185 8176 7219 8210
rect 7253 8176 7287 8210
rect 7321 8176 7355 8210
rect 7389 8176 7423 8210
rect 7457 8176 7491 8210
rect 7525 8176 7559 8210
rect 7593 8176 7627 8210
rect 7661 8176 7695 8210
rect 7729 8176 7763 8210
rect 7797 8176 7831 8210
rect 7865 8176 7899 8210
rect 7933 8176 7967 8210
rect 8001 8176 8035 8210
rect 8069 8176 8103 8210
rect 8137 8176 8171 8210
rect 8205 8176 8239 8210
rect 8273 8176 8307 8210
rect 8341 8176 8367 8210
rect 42 8157 8367 8176
rect 42 8123 68 8157
rect 102 8123 138 8157
rect 172 8123 208 8157
rect 242 8123 278 8157
rect 312 8123 348 8157
rect 382 8123 418 8157
rect 452 8123 488 8157
rect 522 8123 558 8157
rect 592 8123 628 8157
rect 662 8123 698 8157
rect 732 8123 768 8157
rect 802 8123 838 8157
rect 872 8123 908 8157
rect 942 8123 978 8157
rect 1012 8123 1048 8157
rect 1082 8123 1118 8157
rect 1152 8123 1188 8157
rect 1222 8123 1258 8157
rect 1292 8123 1328 8157
rect 1362 8123 1398 8157
rect 1432 8123 1467 8157
rect 1501 8123 1536 8157
rect 1570 8123 1605 8157
rect 1639 8123 1674 8157
rect 1708 8123 1743 8157
rect 1777 8123 1812 8157
rect 1846 8123 1881 8157
rect 1915 8123 1950 8157
rect 1984 8123 2019 8157
rect 2053 8123 2088 8157
rect 2122 8123 2157 8157
rect 2191 8123 2226 8157
rect 2260 8123 2295 8157
rect 2329 8123 2364 8157
rect 2398 8123 2433 8157
rect 2467 8123 2502 8157
rect 2536 8123 2571 8157
rect 2605 8123 2640 8157
rect 2674 8123 2709 8157
rect 2743 8123 2778 8157
rect 2812 8123 2847 8157
rect 2881 8140 8367 8157
rect 2881 8123 2933 8140
rect 42 8106 2933 8123
rect 2967 8106 3002 8140
rect 3036 8106 3071 8140
rect 3105 8106 3139 8140
rect 3173 8106 3207 8140
rect 3241 8106 3275 8140
rect 3309 8106 3343 8140
rect 3377 8106 3411 8140
rect 3445 8106 3479 8140
rect 3513 8106 3547 8140
rect 3581 8106 3615 8140
rect 3649 8106 3683 8140
rect 3717 8106 3751 8140
rect 3785 8106 3819 8140
rect 3853 8106 3887 8140
rect 3921 8106 3955 8140
rect 3989 8106 4023 8140
rect 4057 8106 4091 8140
rect 4125 8106 4159 8140
rect 4193 8106 4227 8140
rect 4261 8106 4295 8140
rect 4329 8106 4363 8140
rect 4397 8106 4431 8140
rect 4465 8106 4499 8140
rect 4533 8106 4567 8140
rect 4601 8106 4635 8140
rect 4669 8106 4703 8140
rect 4737 8106 4771 8140
rect 4805 8106 4839 8140
rect 4873 8106 4907 8140
rect 4941 8106 4975 8140
rect 5009 8106 5043 8140
rect 5077 8106 5111 8140
rect 5145 8106 5179 8140
rect 5213 8106 5247 8140
rect 5281 8106 5315 8140
rect 5349 8106 5383 8140
rect 5417 8106 5451 8140
rect 5485 8106 5519 8140
rect 5553 8106 5587 8140
rect 5621 8106 5655 8140
rect 5689 8106 5723 8140
rect 5757 8106 5791 8140
rect 5825 8106 5859 8140
rect 5893 8106 5927 8140
rect 5961 8106 5995 8140
rect 6029 8106 6063 8140
rect 6097 8106 6131 8140
rect 6165 8106 6199 8140
rect 6233 8106 6267 8140
rect 6301 8106 6335 8140
rect 6369 8106 6403 8140
rect 6437 8106 6471 8140
rect 6505 8106 6539 8140
rect 6573 8106 6607 8140
rect 6641 8106 6675 8140
rect 6709 8106 6743 8140
rect 6777 8106 6811 8140
rect 6845 8106 6879 8140
rect 6913 8106 6947 8140
rect 6981 8106 7015 8140
rect 7049 8106 7083 8140
rect 7117 8106 7151 8140
rect 7185 8106 7219 8140
rect 7253 8106 7287 8140
rect 7321 8106 7355 8140
rect 7389 8106 7423 8140
rect 7457 8106 7491 8140
rect 7525 8106 7559 8140
rect 7593 8106 7627 8140
rect 7661 8106 7695 8140
rect 7729 8106 7763 8140
rect 7797 8106 7831 8140
rect 7865 8106 7899 8140
rect 7933 8106 7967 8140
rect 8001 8106 8035 8140
rect 8069 8106 8103 8140
rect 8137 8106 8171 8140
rect 8205 8106 8239 8140
rect 8273 8106 8307 8140
rect 8341 8106 8367 8140
rect 42 8082 8367 8106
rect 42 8048 68 8082
rect 102 8048 138 8082
rect 172 8048 208 8082
rect 242 8048 278 8082
rect 312 8048 348 8082
rect 382 8048 418 8082
rect 452 8048 488 8082
rect 522 8048 558 8082
rect 592 8048 628 8082
rect 662 8048 698 8082
rect 732 8048 768 8082
rect 802 8048 838 8082
rect 872 8048 908 8082
rect 942 8048 978 8082
rect 1012 8048 1048 8082
rect 1082 8048 1118 8082
rect 1152 8048 1188 8082
rect 1222 8048 1258 8082
rect 1292 8048 1328 8082
rect 1362 8048 1398 8082
rect 1432 8048 1467 8082
rect 1501 8048 1536 8082
rect 1570 8048 1605 8082
rect 1639 8048 1674 8082
rect 1708 8048 1743 8082
rect 1777 8048 1812 8082
rect 1846 8048 1881 8082
rect 1915 8048 1950 8082
rect 1984 8048 2019 8082
rect 2053 8048 2088 8082
rect 2122 8048 2157 8082
rect 2191 8048 2226 8082
rect 2260 8048 2295 8082
rect 2329 8048 2364 8082
rect 2398 8048 2433 8082
rect 2467 8048 2502 8082
rect 2536 8048 2571 8082
rect 2605 8048 2640 8082
rect 2674 8048 2709 8082
rect 2743 8048 2778 8082
rect 2812 8048 2847 8082
rect 2881 8070 8367 8082
rect 2881 8048 2933 8070
rect 42 8036 2933 8048
rect 2967 8036 3002 8070
rect 3036 8036 3071 8070
rect 3105 8036 3139 8070
rect 3173 8036 3207 8070
rect 3241 8036 3275 8070
rect 3309 8036 3343 8070
rect 3377 8036 3411 8070
rect 3445 8036 3479 8070
rect 3513 8036 3547 8070
rect 3581 8036 3615 8070
rect 3649 8036 3683 8070
rect 3717 8036 3751 8070
rect 3785 8036 3819 8070
rect 3853 8036 3887 8070
rect 3921 8036 3955 8070
rect 3989 8036 4023 8070
rect 4057 8036 4091 8070
rect 4125 8036 4159 8070
rect 4193 8036 4227 8070
rect 4261 8036 4295 8070
rect 4329 8036 4363 8070
rect 4397 8036 4431 8070
rect 4465 8036 4499 8070
rect 4533 8036 4567 8070
rect 4601 8036 4635 8070
rect 4669 8036 4703 8070
rect 4737 8036 4771 8070
rect 4805 8036 4839 8070
rect 4873 8036 4907 8070
rect 4941 8036 4975 8070
rect 5009 8036 5043 8070
rect 5077 8036 5111 8070
rect 5145 8036 5179 8070
rect 5213 8036 5247 8070
rect 5281 8036 5315 8070
rect 5349 8036 5383 8070
rect 5417 8036 5451 8070
rect 5485 8036 5519 8070
rect 5553 8036 5587 8070
rect 5621 8036 5655 8070
rect 5689 8036 5723 8070
rect 5757 8036 5791 8070
rect 5825 8036 5859 8070
rect 5893 8036 5927 8070
rect 5961 8036 5995 8070
rect 6029 8036 6063 8070
rect 6097 8036 6131 8070
rect 6165 8036 6199 8070
rect 6233 8036 6267 8070
rect 6301 8036 6335 8070
rect 6369 8036 6403 8070
rect 6437 8036 6471 8070
rect 6505 8036 6539 8070
rect 6573 8036 6607 8070
rect 6641 8036 6675 8070
rect 6709 8036 6743 8070
rect 6777 8036 6811 8070
rect 6845 8036 6879 8070
rect 6913 8036 6947 8070
rect 6981 8036 7015 8070
rect 7049 8036 7083 8070
rect 7117 8036 7151 8070
rect 7185 8036 7219 8070
rect 7253 8036 7287 8070
rect 7321 8036 7355 8070
rect 7389 8036 7423 8070
rect 7457 8036 7491 8070
rect 7525 8036 7559 8070
rect 7593 8036 7627 8070
rect 7661 8036 7695 8070
rect 7729 8036 7763 8070
rect 7797 8036 7831 8070
rect 7865 8036 7899 8070
rect 7933 8036 7967 8070
rect 8001 8036 8035 8070
rect 8069 8036 8103 8070
rect 8137 8036 8171 8070
rect 8205 8036 8239 8070
rect 8273 8036 8307 8070
rect 8341 8036 8367 8070
rect 42 8007 8367 8036
rect 42 7973 68 8007
rect 102 7973 138 8007
rect 172 7973 208 8007
rect 242 7973 278 8007
rect 312 7973 348 8007
rect 382 7973 418 8007
rect 452 7973 488 8007
rect 522 7973 558 8007
rect 592 7973 628 8007
rect 662 7973 698 8007
rect 732 7973 768 8007
rect 802 7973 838 8007
rect 872 7973 908 8007
rect 942 7973 978 8007
rect 1012 7973 1048 8007
rect 1082 7973 1118 8007
rect 1152 7973 1188 8007
rect 1222 7973 1258 8007
rect 1292 7973 1328 8007
rect 1362 7973 1398 8007
rect 1432 7973 1467 8007
rect 1501 7973 1536 8007
rect 1570 7973 1605 8007
rect 1639 7973 1674 8007
rect 1708 7973 1743 8007
rect 1777 7973 1812 8007
rect 1846 7973 1881 8007
rect 1915 7973 1950 8007
rect 1984 7973 2019 8007
rect 2053 7973 2088 8007
rect 2122 7973 2157 8007
rect 2191 7973 2226 8007
rect 2260 7973 2295 8007
rect 2329 7973 2364 8007
rect 2398 7973 2433 8007
rect 2467 7973 2502 8007
rect 2536 7973 2571 8007
rect 2605 7973 2640 8007
rect 2674 7973 2709 8007
rect 2743 7973 2778 8007
rect 2812 7973 2847 8007
rect 2881 8000 8367 8007
rect 2881 7973 2933 8000
rect 42 7966 2933 7973
rect 2967 7966 3002 8000
rect 3036 7966 3071 8000
rect 3105 7966 3139 8000
rect 3173 7966 3207 8000
rect 3241 7966 3275 8000
rect 3309 7966 3343 8000
rect 3377 7966 3411 8000
rect 3445 7966 3479 8000
rect 3513 7966 3547 8000
rect 3581 7966 3615 8000
rect 3649 7966 3683 8000
rect 3717 7966 3751 8000
rect 3785 7966 3819 8000
rect 3853 7966 3887 8000
rect 3921 7966 3955 8000
rect 3989 7966 4023 8000
rect 4057 7966 4091 8000
rect 4125 7966 4159 8000
rect 4193 7966 4227 8000
rect 4261 7966 4295 8000
rect 4329 7966 4363 8000
rect 4397 7966 4431 8000
rect 4465 7966 4499 8000
rect 4533 7966 4567 8000
rect 4601 7966 4635 8000
rect 4669 7966 4703 8000
rect 4737 7966 4771 8000
rect 4805 7966 4839 8000
rect 4873 7966 4907 8000
rect 4941 7966 4975 8000
rect 5009 7966 5043 8000
rect 5077 7966 5111 8000
rect 5145 7966 5179 8000
rect 5213 7966 5247 8000
rect 5281 7966 5315 8000
rect 5349 7966 5383 8000
rect 5417 7966 5451 8000
rect 5485 7966 5519 8000
rect 5553 7966 5587 8000
rect 5621 7966 5655 8000
rect 5689 7966 5723 8000
rect 5757 7966 5791 8000
rect 5825 7966 5859 8000
rect 5893 7966 5927 8000
rect 5961 7966 5995 8000
rect 6029 7966 6063 8000
rect 6097 7966 6131 8000
rect 6165 7966 6199 8000
rect 6233 7966 6267 8000
rect 6301 7966 6335 8000
rect 6369 7966 6403 8000
rect 6437 7966 6471 8000
rect 6505 7966 6539 8000
rect 6573 7966 6607 8000
rect 6641 7966 6675 8000
rect 6709 7966 6743 8000
rect 6777 7966 6811 8000
rect 6845 7966 6879 8000
rect 6913 7966 6947 8000
rect 6981 7966 7015 8000
rect 7049 7966 7083 8000
rect 7117 7966 7151 8000
rect 7185 7966 7219 8000
rect 7253 7966 7287 8000
rect 7321 7966 7355 8000
rect 7389 7966 7423 8000
rect 7457 7966 7491 8000
rect 7525 7966 7559 8000
rect 7593 7966 7627 8000
rect 7661 7966 7695 8000
rect 7729 7966 7763 8000
rect 7797 7966 7831 8000
rect 7865 7966 7899 8000
rect 7933 7966 7967 8000
rect 8001 7966 8035 8000
rect 8069 7966 8103 8000
rect 8137 7966 8171 8000
rect 8205 7966 8239 8000
rect 8273 7966 8307 8000
rect 8341 7966 8367 8000
rect 42 7932 8367 7966
rect 42 7898 68 7932
rect 102 7898 138 7932
rect 172 7898 208 7932
rect 242 7898 278 7932
rect 312 7898 348 7932
rect 382 7898 418 7932
rect 452 7898 488 7932
rect 522 7898 558 7932
rect 592 7898 628 7932
rect 662 7898 698 7932
rect 732 7898 768 7932
rect 802 7898 838 7932
rect 872 7898 908 7932
rect 942 7898 978 7932
rect 1012 7898 1048 7932
rect 1082 7898 1118 7932
rect 1152 7898 1188 7932
rect 1222 7898 1258 7932
rect 1292 7898 1328 7932
rect 1362 7898 1398 7932
rect 1432 7898 1467 7932
rect 1501 7898 1536 7932
rect 1570 7898 1605 7932
rect 1639 7898 1674 7932
rect 1708 7898 1743 7932
rect 1777 7898 1812 7932
rect 1846 7898 1881 7932
rect 1915 7898 1950 7932
rect 1984 7898 2019 7932
rect 2053 7898 2088 7932
rect 2122 7898 2157 7932
rect 2191 7898 2226 7932
rect 2260 7898 2295 7932
rect 2329 7898 2364 7932
rect 2398 7898 2433 7932
rect 2467 7898 2502 7932
rect 2536 7898 2571 7932
rect 2605 7898 2640 7932
rect 2674 7898 2709 7932
rect 2743 7898 2778 7932
rect 2812 7898 2847 7932
rect 2881 7930 8367 7932
rect 2881 7898 2933 7930
rect 42 7896 2933 7898
rect 2967 7896 3002 7930
rect 3036 7896 3071 7930
rect 3105 7896 3139 7930
rect 3173 7896 3207 7930
rect 3241 7896 3275 7930
rect 3309 7896 3343 7930
rect 3377 7896 3411 7930
rect 3445 7896 3479 7930
rect 3513 7896 3547 7930
rect 3581 7896 3615 7930
rect 3649 7896 3683 7930
rect 3717 7896 3751 7930
rect 3785 7896 3819 7930
rect 3853 7896 3887 7930
rect 3921 7896 3955 7930
rect 3989 7896 4023 7930
rect 4057 7896 4091 7930
rect 4125 7896 4159 7930
rect 4193 7896 4227 7930
rect 4261 7896 4295 7930
rect 4329 7896 4363 7930
rect 4397 7896 4431 7930
rect 4465 7896 4499 7930
rect 4533 7896 4567 7930
rect 4601 7896 4635 7930
rect 4669 7896 4703 7930
rect 4737 7896 4771 7930
rect 4805 7896 4839 7930
rect 4873 7896 4907 7930
rect 4941 7896 4975 7930
rect 5009 7896 5043 7930
rect 5077 7896 5111 7930
rect 5145 7896 5179 7930
rect 5213 7896 5247 7930
rect 5281 7896 5315 7930
rect 5349 7896 5383 7930
rect 5417 7896 5451 7930
rect 5485 7896 5519 7930
rect 5553 7896 5587 7930
rect 5621 7896 5655 7930
rect 5689 7896 5723 7930
rect 5757 7896 5791 7930
rect 5825 7896 5859 7930
rect 5893 7896 5927 7930
rect 5961 7896 5995 7930
rect 6029 7896 6063 7930
rect 6097 7896 6131 7930
rect 6165 7896 6199 7930
rect 6233 7896 6267 7930
rect 6301 7896 6335 7930
rect 6369 7896 6403 7930
rect 6437 7896 6471 7930
rect 6505 7896 6539 7930
rect 6573 7896 6607 7930
rect 6641 7896 6675 7930
rect 6709 7896 6743 7930
rect 6777 7896 6811 7930
rect 6845 7896 6879 7930
rect 6913 7896 6947 7930
rect 6981 7896 7015 7930
rect 7049 7896 7083 7930
rect 7117 7896 7151 7930
rect 7185 7896 7219 7930
rect 7253 7896 7287 7930
rect 7321 7896 7355 7930
rect 7389 7896 7423 7930
rect 7457 7896 7491 7930
rect 7525 7896 7559 7930
rect 7593 7896 7627 7930
rect 7661 7896 7695 7930
rect 7729 7896 7763 7930
rect 7797 7896 7831 7930
rect 7865 7896 7899 7930
rect 7933 7896 7967 7930
rect 8001 7896 8035 7930
rect 8069 7896 8103 7930
rect 8137 7896 8171 7930
rect 8205 7896 8239 7930
rect 8273 7896 8307 7930
rect 8341 7896 8367 7930
rect 8494 8254 8628 8255
rect 8494 7932 8509 8254
rect 8615 7932 8628 8254
rect 8494 7917 8628 7932
rect 9596 8247 9714 8255
rect 9630 8239 9678 8247
rect 9712 8239 9714 8247
rect 9596 8144 9612 8213
rect 9596 8041 9612 8110
rect 9596 7933 9612 8007
rect 9596 7917 9714 7933
rect 10314 8247 10430 8255
rect 10348 8239 10396 8247
rect 10416 8144 10430 8213
rect 10416 8041 10430 8110
rect 10416 7933 10430 8007
rect 10314 7917 10430 7933
rect 10800 8254 10934 8255
rect 10800 8220 10804 8254
rect 10838 8239 10898 8254
rect 10932 8220 10934 8254
rect 10800 8179 10816 8220
rect 10918 8179 10934 8220
rect 10800 8145 10804 8179
rect 10932 8145 10934 8179
rect 10800 8104 10816 8145
rect 10918 8104 10934 8145
rect 10800 8070 10804 8104
rect 10932 8070 10934 8104
rect 10800 8028 10816 8070
rect 10918 8028 10934 8070
rect 10800 7994 10804 8028
rect 10932 7994 10934 8028
rect 10800 7952 10816 7994
rect 10918 7952 10934 7994
rect 10800 7918 10804 7952
rect 10838 7918 10898 7933
rect 10932 7918 10934 7952
rect 10800 7917 10934 7918
rect 13506 8249 13532 8283
rect 13566 8249 13603 8283
rect 13637 8249 13674 8283
rect 13708 8249 13744 8283
rect 13778 8249 13814 8283
rect 13848 8249 13884 8283
rect 13918 8249 13954 8283
rect 13988 8249 14024 8283
rect 14058 8249 14094 8283
rect 14128 8249 14164 8283
rect 14198 8280 14234 8283
rect 14268 8280 14304 8283
rect 14338 8280 14374 8283
rect 14408 8280 14444 8283
rect 14478 8280 14514 8283
rect 14219 8249 14234 8280
rect 14291 8249 14304 8280
rect 14363 8249 14374 8280
rect 14435 8249 14444 8280
rect 14507 8249 14514 8280
rect 14548 8249 14584 8283
rect 14648 8280 14654 8283
rect 14618 8249 14654 8280
rect 14688 8280 14692 8283
rect 14758 8280 14770 8283
rect 14828 8280 14848 8283
rect 14898 8280 14926 8283
rect 14688 8249 14724 8280
rect 14758 8249 14794 8280
rect 14828 8249 14864 8280
rect 14898 8255 14932 8280
rect 14966 8255 15000 8289
rect 15038 8280 15068 8289
rect 15034 8255 15068 8280
rect 14898 8249 15102 8255
rect 13506 8246 14185 8249
rect 14219 8246 14257 8249
rect 14291 8246 14329 8249
rect 14363 8246 14401 8249
rect 14435 8246 14473 8249
rect 14507 8246 15102 8249
rect 13506 8240 15102 8246
rect 13506 8209 14614 8240
rect 14648 8209 14692 8240
rect 14726 8209 14770 8240
rect 14804 8209 14848 8240
rect 14882 8209 14926 8240
rect 14960 8217 15004 8240
rect 15038 8217 15102 8240
rect 13506 8175 13532 8209
rect 13566 8175 13603 8209
rect 13637 8175 13674 8209
rect 13708 8175 13744 8209
rect 13778 8175 13814 8209
rect 13848 8175 13884 8209
rect 13918 8175 13954 8209
rect 13988 8175 14024 8209
rect 14058 8175 14094 8209
rect 14128 8175 14164 8209
rect 14198 8202 14234 8209
rect 14268 8202 14304 8209
rect 14338 8202 14374 8209
rect 14408 8202 14444 8209
rect 14478 8202 14514 8209
rect 14219 8175 14234 8202
rect 14291 8175 14304 8202
rect 14363 8175 14374 8202
rect 14435 8175 14444 8202
rect 14507 8175 14514 8202
rect 14548 8175 14584 8209
rect 14648 8206 14654 8209
rect 14618 8175 14654 8206
rect 14688 8206 14692 8209
rect 14758 8206 14770 8209
rect 14828 8206 14848 8209
rect 14898 8206 14926 8209
rect 14688 8175 14724 8206
rect 14758 8175 14794 8206
rect 14828 8175 14864 8206
rect 14898 8183 14932 8206
rect 14966 8183 15000 8217
rect 15038 8206 15068 8217
rect 15034 8183 15068 8206
rect 14898 8175 15102 8183
rect 13506 8168 14185 8175
rect 14219 8168 14257 8175
rect 14291 8168 14329 8175
rect 14363 8168 14401 8175
rect 14435 8168 14473 8175
rect 14507 8168 15102 8175
rect 13506 8166 15102 8168
rect 13506 8135 14614 8166
rect 14648 8135 14692 8166
rect 14726 8135 14770 8166
rect 14804 8135 14848 8166
rect 14882 8135 14926 8166
rect 14960 8145 15004 8166
rect 15038 8145 15102 8166
rect 13506 8101 13532 8135
rect 13566 8101 13603 8135
rect 13637 8101 13674 8135
rect 13708 8101 13744 8135
rect 13778 8101 13814 8135
rect 13848 8101 13884 8135
rect 13918 8101 13954 8135
rect 13988 8101 14024 8135
rect 14058 8101 14094 8135
rect 14128 8101 14164 8135
rect 14198 8101 14234 8135
rect 14268 8101 14304 8135
rect 14338 8101 14374 8135
rect 14408 8115 14444 8135
rect 14478 8115 14514 8135
rect 14408 8101 14431 8115
rect 14478 8101 14511 8115
rect 14548 8101 14584 8135
rect 14648 8132 14654 8135
rect 14618 8101 14654 8132
rect 14688 8132 14692 8135
rect 14758 8132 14770 8135
rect 14828 8132 14848 8135
rect 14898 8132 14926 8135
rect 14688 8101 14724 8132
rect 14758 8101 14794 8132
rect 14828 8101 14864 8132
rect 14898 8111 14932 8132
rect 14966 8111 15000 8145
rect 15038 8132 15068 8145
rect 15034 8111 15068 8132
rect 14898 8101 15102 8111
rect 13506 8081 14431 8101
rect 14465 8081 14511 8101
rect 14545 8092 15102 8101
rect 14545 8081 14614 8092
rect 13506 8061 14614 8081
rect 14648 8061 14692 8092
rect 14726 8061 14770 8092
rect 14804 8061 14848 8092
rect 14882 8061 14926 8092
rect 14960 8073 15004 8092
rect 15038 8073 15102 8092
rect 13506 8027 13532 8061
rect 13566 8027 13603 8061
rect 13637 8027 13674 8061
rect 13708 8027 13744 8061
rect 13778 8027 13814 8061
rect 13848 8027 13884 8061
rect 13918 8027 13954 8061
rect 13988 8027 14024 8061
rect 14058 8027 14094 8061
rect 14128 8027 14164 8061
rect 14198 8027 14234 8061
rect 14268 8027 14304 8061
rect 14338 8027 14374 8061
rect 14408 8033 14444 8061
rect 14478 8033 14514 8061
rect 14408 8027 14431 8033
rect 14478 8027 14511 8033
rect 14548 8027 14584 8061
rect 14648 8058 14654 8061
rect 14618 8027 14654 8058
rect 14688 8058 14692 8061
rect 14758 8058 14770 8061
rect 14828 8058 14848 8061
rect 14898 8058 14926 8061
rect 14688 8027 14724 8058
rect 14758 8027 14794 8058
rect 14828 8027 14864 8058
rect 14898 8039 14932 8058
rect 14966 8039 15000 8073
rect 15038 8058 15068 8073
rect 15034 8039 15068 8058
rect 14898 8027 15102 8039
rect 13506 7999 14431 8027
rect 14465 7999 14511 8027
rect 14545 8018 15102 8027
rect 14545 7999 14614 8018
rect 13506 7987 14614 7999
rect 14648 7987 14692 8018
rect 14726 7987 14770 8018
rect 14804 7987 14848 8018
rect 14882 7987 14926 8018
rect 14960 8001 15004 8018
rect 15038 8001 15102 8018
rect 13506 7953 13532 7987
rect 13566 7953 13603 7987
rect 13637 7953 13674 7987
rect 13708 7953 13744 7987
rect 13778 7953 13814 7987
rect 13848 7953 13884 7987
rect 13918 7953 13954 7987
rect 13988 7953 14024 7987
rect 14058 7953 14094 7987
rect 14128 7953 14164 7987
rect 14198 7953 14234 7987
rect 14268 7953 14304 7987
rect 14338 7953 14374 7987
rect 14408 7953 14444 7987
rect 14478 7953 14514 7987
rect 14548 7953 14584 7987
rect 14648 7984 14654 7987
rect 14618 7953 14654 7984
rect 14688 7984 14692 7987
rect 14758 7984 14770 7987
rect 14828 7984 14848 7987
rect 14898 7984 14926 7987
rect 14688 7953 14724 7984
rect 14758 7953 14794 7984
rect 14828 7953 14864 7984
rect 14898 7967 14932 7984
rect 14966 7967 15000 8001
rect 15038 7984 15068 8001
rect 15034 7967 15068 7984
rect 14898 7953 15102 7967
rect 13506 7950 15102 7953
rect 42 7860 8367 7896
rect 42 7857 2933 7860
rect 42 7823 68 7857
rect 102 7823 138 7857
rect 172 7823 208 7857
rect 242 7823 278 7857
rect 312 7823 348 7857
rect 382 7823 418 7857
rect 452 7823 488 7857
rect 522 7823 558 7857
rect 592 7823 628 7857
rect 662 7823 698 7857
rect 732 7823 768 7857
rect 802 7823 838 7857
rect 872 7823 908 7857
rect 942 7823 978 7857
rect 1012 7823 1048 7857
rect 1082 7823 1118 7857
rect 1152 7823 1188 7857
rect 1222 7823 1258 7857
rect 1292 7823 1328 7857
rect 1362 7823 1398 7857
rect 1432 7823 1467 7857
rect 1501 7823 1536 7857
rect 1570 7823 1605 7857
rect 1639 7823 1674 7857
rect 1708 7823 1743 7857
rect 1777 7823 1812 7857
rect 1846 7823 1881 7857
rect 1915 7823 1950 7857
rect 1984 7823 2019 7857
rect 2053 7823 2088 7857
rect 2122 7823 2157 7857
rect 2191 7823 2226 7857
rect 2260 7823 2295 7857
rect 2329 7823 2364 7857
rect 2398 7823 2433 7857
rect 2467 7823 2502 7857
rect 2536 7823 2571 7857
rect 2605 7823 2640 7857
rect 2674 7823 2709 7857
rect 2743 7823 2778 7857
rect 2812 7823 2847 7857
rect 2881 7826 2933 7857
rect 2967 7826 3002 7860
rect 3036 7826 3071 7860
rect 3105 7826 3139 7860
rect 3173 7826 3207 7860
rect 3241 7826 3275 7860
rect 3309 7826 3343 7860
rect 3377 7826 3411 7860
rect 3445 7826 3479 7860
rect 3513 7826 3547 7860
rect 3581 7826 3615 7860
rect 3649 7826 3683 7860
rect 3717 7826 3751 7860
rect 3785 7826 3819 7860
rect 3853 7826 3887 7860
rect 3921 7826 3955 7860
rect 3989 7826 4023 7860
rect 4057 7826 4091 7860
rect 4125 7826 4159 7860
rect 4193 7826 4227 7860
rect 4261 7826 4295 7860
rect 4329 7826 4363 7860
rect 4397 7826 4431 7860
rect 4465 7826 4499 7860
rect 4533 7826 4567 7860
rect 4601 7826 4635 7860
rect 4669 7826 4703 7860
rect 4737 7826 4771 7860
rect 4805 7826 4839 7860
rect 4873 7826 4907 7860
rect 4941 7826 4975 7860
rect 5009 7826 5043 7860
rect 5077 7826 5111 7860
rect 5145 7826 5179 7860
rect 5213 7826 5247 7860
rect 5281 7826 5315 7860
rect 5349 7826 5383 7860
rect 5417 7826 5451 7860
rect 5485 7826 5519 7860
rect 5553 7826 5587 7860
rect 5621 7826 5655 7860
rect 5689 7826 5723 7860
rect 5757 7826 5791 7860
rect 5825 7826 5859 7860
rect 5893 7826 5927 7860
rect 5961 7826 5995 7860
rect 6029 7826 6063 7860
rect 6097 7826 6131 7860
rect 6165 7826 6199 7860
rect 6233 7826 6267 7860
rect 6301 7826 6335 7860
rect 6369 7826 6403 7860
rect 6437 7826 6471 7860
rect 6505 7826 6539 7860
rect 6573 7826 6607 7860
rect 6641 7826 6675 7860
rect 6709 7826 6743 7860
rect 6777 7826 6811 7860
rect 6845 7826 6879 7860
rect 6913 7826 6947 7860
rect 6981 7826 7015 7860
rect 7049 7826 7083 7860
rect 7117 7826 7151 7860
rect 7185 7826 7219 7860
rect 7253 7826 7287 7860
rect 7321 7826 7355 7860
rect 7389 7826 7423 7860
rect 7457 7826 7491 7860
rect 7525 7826 7559 7860
rect 7593 7826 7627 7860
rect 7661 7826 7695 7860
rect 7729 7826 7763 7860
rect 7797 7826 7831 7860
rect 7865 7826 7899 7860
rect 7933 7826 7967 7860
rect 8001 7826 8035 7860
rect 8069 7826 8103 7860
rect 8137 7826 8171 7860
rect 8205 7826 8239 7860
rect 8273 7826 8307 7860
rect 8341 7826 8367 7860
rect 2881 7823 8367 7826
rect 42 7788 8367 7823
rect 13506 7916 14431 7950
rect 14465 7916 14511 7950
rect 14545 7944 15102 7950
rect 14545 7916 14614 7944
rect 13506 7913 14614 7916
rect 14648 7913 14692 7944
rect 14726 7913 14770 7944
rect 14804 7913 14848 7944
rect 14882 7913 14926 7944
rect 14960 7929 15004 7944
rect 15038 7929 15102 7944
rect 13506 7879 13532 7913
rect 13566 7879 13603 7913
rect 13637 7879 13674 7913
rect 13708 7879 13744 7913
rect 13778 7879 13814 7913
rect 13848 7879 13884 7913
rect 13918 7879 13954 7913
rect 13988 7879 14024 7913
rect 14058 7879 14094 7913
rect 14128 7879 14164 7913
rect 14198 7879 14234 7913
rect 14268 7879 14304 7913
rect 14338 7879 14374 7913
rect 14408 7879 14444 7913
rect 14478 7879 14514 7913
rect 14548 7879 14584 7913
rect 14648 7910 14654 7913
rect 14618 7879 14654 7910
rect 14688 7910 14692 7913
rect 14758 7910 14770 7913
rect 14828 7910 14848 7913
rect 14898 7910 14926 7913
rect 14688 7879 14724 7910
rect 14758 7879 14794 7910
rect 14828 7879 14864 7910
rect 14898 7895 14932 7910
rect 14966 7895 15000 7929
rect 15038 7910 15068 7929
rect 15034 7895 15068 7910
rect 14898 7879 15102 7895
rect 13506 7870 15102 7879
rect 13506 7839 14614 7870
rect 14648 7839 14692 7870
rect 14726 7839 14770 7870
rect 14804 7839 14848 7870
rect 14882 7839 14926 7870
rect 14960 7857 15004 7870
rect 15038 7857 15102 7870
rect 13506 7805 13532 7839
rect 13566 7805 13603 7839
rect 13637 7805 13674 7839
rect 13708 7805 13744 7839
rect 13778 7805 13814 7839
rect 13848 7805 13884 7839
rect 13918 7805 13954 7839
rect 13988 7805 14024 7839
rect 14058 7805 14094 7839
rect 14128 7805 14164 7839
rect 14198 7805 14234 7839
rect 14268 7805 14304 7839
rect 14338 7805 14374 7839
rect 14408 7805 14444 7839
rect 14478 7805 14514 7839
rect 14548 7805 14584 7839
rect 14648 7836 14654 7839
rect 14618 7805 14654 7836
rect 14688 7836 14692 7839
rect 14758 7836 14770 7839
rect 14828 7836 14848 7839
rect 14898 7836 14926 7839
rect 14688 7805 14724 7836
rect 14758 7805 14794 7836
rect 14828 7805 14864 7836
rect 14898 7823 14932 7836
rect 14966 7823 15000 7857
rect 15038 7836 15068 7857
rect 15034 7823 15068 7836
rect 14898 7805 15102 7823
rect 13506 7796 15102 7805
rect 13506 7788 14614 7796
rect 42 7762 14614 7788
rect 14648 7762 14692 7796
rect 14726 7762 14770 7796
rect 14804 7762 14848 7796
rect 14882 7762 14926 7796
rect 14960 7785 15004 7796
rect 15038 7785 15102 7796
rect 42 7751 14932 7762
rect 14966 7751 15000 7785
rect 15038 7762 15068 7785
rect 15034 7751 15068 7762
rect 42 7749 15102 7751
rect 42 7715 68 7749
rect 102 7715 137 7749
rect 171 7715 206 7749
rect 240 7715 275 7749
rect 309 7715 344 7749
rect 378 7715 413 7749
rect 447 7715 482 7749
rect 516 7715 551 7749
rect 585 7715 620 7749
rect 654 7715 689 7749
rect 723 7715 758 7749
rect 792 7715 827 7749
rect 861 7715 896 7749
rect 930 7715 965 7749
rect 999 7715 1034 7749
rect 1068 7715 1103 7749
rect 1137 7715 1172 7749
rect 1206 7715 1241 7749
rect 1275 7715 1310 7749
rect 1344 7715 1379 7749
rect 1413 7715 1448 7749
rect 1482 7715 1517 7749
rect 1551 7715 1586 7749
rect 1620 7715 1655 7749
rect 1689 7715 1724 7749
rect 1758 7715 1793 7749
rect 1827 7715 1862 7749
rect 1896 7715 1931 7749
rect 1965 7715 2000 7749
rect 2034 7715 2069 7749
rect 2103 7715 2138 7749
rect 2172 7715 2207 7749
rect 2241 7715 2276 7749
rect 2310 7715 2345 7749
rect 2379 7715 2414 7749
rect 2448 7715 2483 7749
rect 2517 7715 2552 7749
rect 2586 7715 2621 7749
rect 2655 7715 2690 7749
rect 2724 7715 2759 7749
rect 2793 7715 2828 7749
rect 2862 7715 2896 7749
rect 2930 7715 2964 7749
rect 2998 7715 3032 7749
rect 3066 7715 3100 7749
rect 3134 7715 3168 7749
rect 3202 7715 3236 7749
rect 3270 7715 3304 7749
rect 3338 7715 3372 7749
rect 3406 7715 3440 7749
rect 3474 7715 3508 7749
rect 3542 7715 3576 7749
rect 3610 7715 3644 7749
rect 3678 7715 3712 7749
rect 3746 7715 3780 7749
rect 3814 7715 3848 7749
rect 3882 7715 3916 7749
rect 3950 7715 3984 7749
rect 4018 7715 4052 7749
rect 4086 7715 4120 7749
rect 4154 7715 4188 7749
rect 4222 7715 4256 7749
rect 4290 7715 4324 7749
rect 4358 7715 4392 7749
rect 4426 7715 4460 7749
rect 4494 7715 4528 7749
rect 4562 7715 4596 7749
rect 4630 7715 4664 7749
rect 4698 7715 4732 7749
rect 4766 7715 4800 7749
rect 4834 7715 4868 7749
rect 4902 7715 4936 7749
rect 4970 7715 5004 7749
rect 5038 7715 5072 7749
rect 5106 7715 5140 7749
rect 5174 7715 5208 7749
rect 5242 7715 5276 7749
rect 5310 7715 5344 7749
rect 5378 7715 5412 7749
rect 5446 7715 5480 7749
rect 5514 7715 5548 7749
rect 5582 7715 5616 7749
rect 5650 7715 5684 7749
rect 5718 7715 5752 7749
rect 5786 7715 5820 7749
rect 5854 7715 5888 7749
rect 5922 7715 5956 7749
rect 5990 7715 6024 7749
rect 6058 7715 6092 7749
rect 6126 7715 6160 7749
rect 6194 7715 6228 7749
rect 6262 7715 6296 7749
rect 6330 7715 6364 7749
rect 6398 7715 6432 7749
rect 6466 7715 6500 7749
rect 6534 7715 6568 7749
rect 6602 7715 6636 7749
rect 6670 7715 6704 7749
rect 6738 7715 6772 7749
rect 6806 7715 6840 7749
rect 6874 7715 6908 7749
rect 6942 7715 6976 7749
rect 7010 7715 7044 7749
rect 7078 7715 7112 7749
rect 7146 7715 7180 7749
rect 7214 7715 7248 7749
rect 7282 7715 7316 7749
rect 7350 7715 7384 7749
rect 7418 7715 7452 7749
rect 7486 7715 7520 7749
rect 7554 7715 7588 7749
rect 7622 7715 7656 7749
rect 7690 7715 7724 7749
rect 7758 7715 7792 7749
rect 7826 7715 7860 7749
rect 7894 7715 7928 7749
rect 7962 7715 7996 7749
rect 8030 7715 8064 7749
rect 8098 7715 8132 7749
rect 8166 7715 8200 7749
rect 8234 7715 8268 7749
rect 8302 7715 8336 7749
rect 8370 7715 8404 7749
rect 8438 7715 8472 7749
rect 8506 7715 8540 7749
rect 8574 7715 8608 7749
rect 8642 7715 8676 7749
rect 8710 7715 8744 7749
rect 8778 7715 8812 7749
rect 8846 7715 8880 7749
rect 8914 7715 8948 7749
rect 8982 7715 9016 7749
rect 9050 7715 9084 7749
rect 9118 7715 9152 7749
rect 9186 7715 9220 7749
rect 9254 7715 9288 7749
rect 9322 7715 9356 7749
rect 9390 7715 9424 7749
rect 9458 7715 9492 7749
rect 9526 7715 9560 7749
rect 9594 7715 9628 7749
rect 9662 7715 9696 7749
rect 9730 7715 9764 7749
rect 9798 7715 9832 7749
rect 9866 7715 9900 7749
rect 9934 7715 9968 7749
rect 10002 7715 10036 7749
rect 10070 7715 10104 7749
rect 10138 7715 10172 7749
rect 10206 7715 10240 7749
rect 10274 7715 10308 7749
rect 10342 7715 10376 7749
rect 10410 7715 10444 7749
rect 10478 7715 10512 7749
rect 10546 7715 10580 7749
rect 10614 7715 10648 7749
rect 10682 7715 10716 7749
rect 10750 7715 10784 7749
rect 10818 7715 10852 7749
rect 10886 7715 10920 7749
rect 10954 7715 10988 7749
rect 11022 7715 11056 7749
rect 11090 7715 11124 7749
rect 11158 7715 11192 7749
rect 11226 7715 11260 7749
rect 11294 7715 11328 7749
rect 11362 7715 11396 7749
rect 11430 7715 11464 7749
rect 11498 7715 11532 7749
rect 11566 7715 11600 7749
rect 11634 7715 11668 7749
rect 11702 7715 11736 7749
rect 11770 7715 11804 7749
rect 11838 7715 11872 7749
rect 11906 7715 11940 7749
rect 11974 7715 12008 7749
rect 12042 7715 12076 7749
rect 12110 7715 12144 7749
rect 12178 7715 12212 7749
rect 12246 7715 12280 7749
rect 12314 7715 12348 7749
rect 12382 7715 12416 7749
rect 12450 7715 12484 7749
rect 12518 7715 12552 7749
rect 12586 7715 12620 7749
rect 12654 7715 12688 7749
rect 12722 7715 12756 7749
rect 12790 7715 12824 7749
rect 12858 7715 12892 7749
rect 12926 7715 12960 7749
rect 12994 7715 13028 7749
rect 13062 7715 13096 7749
rect 13130 7715 13164 7749
rect 13198 7715 13232 7749
rect 13266 7715 13300 7749
rect 13334 7715 13368 7749
rect 13402 7715 13436 7749
rect 13470 7715 13504 7749
rect 13538 7715 13572 7749
rect 13606 7715 13640 7749
rect 13674 7715 13708 7749
rect 13742 7715 13776 7749
rect 13810 7715 13844 7749
rect 13878 7715 13912 7749
rect 13946 7715 13980 7749
rect 14014 7715 14048 7749
rect 14082 7715 14116 7749
rect 14150 7715 14184 7749
rect 14218 7715 14252 7749
rect 14286 7715 14320 7749
rect 14354 7715 14388 7749
rect 14422 7715 14456 7749
rect 14490 7715 14524 7749
rect 14558 7715 14592 7749
rect 14626 7722 14660 7749
rect 14694 7722 14728 7749
rect 14648 7715 14660 7722
rect 14726 7715 14728 7722
rect 14762 7722 14796 7749
rect 14830 7722 14864 7749
rect 14898 7722 15102 7749
rect 14762 7715 14770 7722
rect 14830 7715 14848 7722
rect 14898 7715 14926 7722
rect 42 7688 14614 7715
rect 14648 7688 14692 7715
rect 14726 7688 14770 7715
rect 14804 7688 14848 7715
rect 14882 7688 14926 7715
rect 14960 7713 15004 7722
rect 15038 7713 15102 7722
rect 42 7679 14932 7688
rect 14966 7679 15000 7713
rect 15038 7688 15068 7713
rect 15034 7679 15068 7688
rect 42 7677 15102 7679
rect 34 7676 15102 7677
rect 34 7642 2733 7676
rect 34 7608 68 7642
rect 102 7608 137 7642
rect 171 7608 206 7642
rect 240 7608 275 7642
rect 309 7608 344 7642
rect 378 7608 413 7642
rect 447 7608 482 7642
rect 516 7608 551 7642
rect 585 7608 620 7642
rect 654 7608 689 7642
rect 723 7608 758 7642
rect 792 7608 827 7642
rect 861 7608 896 7642
rect 930 7608 965 7642
rect 999 7608 1033 7642
rect 1067 7608 1101 7642
rect 1135 7608 1169 7642
rect 1203 7608 1237 7642
rect 1271 7608 1305 7642
rect 1339 7608 1373 7642
rect 1407 7608 1441 7642
rect 1475 7608 1509 7642
rect 1543 7608 1577 7642
rect 1611 7608 1645 7642
rect 1679 7608 1713 7642
rect 1747 7608 1781 7642
rect 1815 7608 1849 7642
rect 1883 7608 1917 7642
rect 1951 7608 1985 7642
rect 2019 7608 2053 7642
rect 2087 7608 2121 7642
rect 2155 7608 2189 7642
rect 2223 7608 2257 7642
rect 2291 7608 2325 7642
rect 2359 7608 2393 7642
rect 2427 7608 2461 7642
rect 2495 7608 2529 7642
rect 2563 7608 2597 7642
rect 2631 7608 2665 7642
rect 2699 7608 2733 7642
rect 34 7570 2733 7608
rect 34 7536 68 7570
rect 102 7536 137 7570
rect 171 7536 206 7570
rect 240 7536 275 7570
rect 309 7536 344 7570
rect 378 7536 413 7570
rect 447 7536 482 7570
rect 516 7536 551 7570
rect 585 7536 620 7570
rect 654 7536 689 7570
rect 723 7536 758 7570
rect 792 7536 827 7570
rect 861 7536 896 7570
rect 930 7536 965 7570
rect 999 7536 1033 7570
rect 1067 7536 1101 7570
rect 1135 7536 1169 7570
rect 1203 7536 1237 7570
rect 1271 7536 1305 7570
rect 1339 7536 1373 7570
rect 1407 7536 1441 7570
rect 1475 7536 1509 7570
rect 1543 7536 1577 7570
rect 1611 7536 1645 7570
rect 1679 7536 1713 7570
rect 1747 7536 1781 7570
rect 1815 7536 1849 7570
rect 1883 7536 1917 7570
rect 1951 7536 1985 7570
rect 2019 7536 2053 7570
rect 2087 7536 2121 7570
rect 2155 7536 2189 7570
rect 2223 7536 2257 7570
rect 2291 7536 2325 7570
rect 2359 7536 2393 7570
rect 2427 7536 2461 7570
rect 2495 7536 2529 7570
rect 2563 7536 2597 7570
rect 2631 7536 2665 7570
rect 2699 7536 2733 7570
rect 34 7498 2733 7536
rect 34 7464 68 7498
rect 102 7464 137 7498
rect 171 7464 206 7498
rect 240 7464 275 7498
rect 309 7464 344 7498
rect 378 7464 413 7498
rect 447 7464 482 7498
rect 516 7464 551 7498
rect 585 7464 620 7498
rect 654 7464 689 7498
rect 723 7464 758 7498
rect 792 7464 827 7498
rect 861 7464 896 7498
rect 930 7464 965 7498
rect 999 7464 1033 7498
rect 1067 7464 1101 7498
rect 1135 7464 1169 7498
rect 1203 7464 1237 7498
rect 1271 7464 1305 7498
rect 1339 7464 1373 7498
rect 1407 7464 1441 7498
rect 1475 7464 1509 7498
rect 1543 7464 1577 7498
rect 1611 7464 1645 7498
rect 1679 7464 1713 7498
rect 1747 7464 1781 7498
rect 1815 7464 1849 7498
rect 1883 7464 1917 7498
rect 1951 7464 1985 7498
rect 2019 7464 2053 7498
rect 2087 7464 2121 7498
rect 2155 7464 2189 7498
rect 2223 7464 2257 7498
rect 2291 7464 2325 7498
rect 2359 7464 2393 7498
rect 2427 7464 2461 7498
rect 2495 7464 2529 7498
rect 2563 7464 2597 7498
rect 2631 7464 2665 7498
rect 2699 7464 2733 7498
rect 34 7426 2733 7464
rect 34 7392 68 7426
rect 102 7392 137 7426
rect 171 7392 206 7426
rect 240 7392 275 7426
rect 309 7392 344 7426
rect 378 7392 413 7426
rect 447 7392 482 7426
rect 516 7392 551 7426
rect 585 7392 620 7426
rect 654 7392 689 7426
rect 723 7392 758 7426
rect 792 7392 827 7426
rect 861 7392 896 7426
rect 930 7392 965 7426
rect 999 7392 1033 7426
rect 1067 7392 1101 7426
rect 1135 7392 1169 7426
rect 1203 7392 1237 7426
rect 1271 7392 1305 7426
rect 1339 7392 1373 7426
rect 1407 7392 1441 7426
rect 1475 7392 1509 7426
rect 1543 7392 1577 7426
rect 1611 7392 1645 7426
rect 1679 7392 1713 7426
rect 1747 7392 1781 7426
rect 1815 7392 1849 7426
rect 1883 7392 1917 7426
rect 1951 7392 1985 7426
rect 2019 7392 2053 7426
rect 2087 7392 2121 7426
rect 2155 7392 2189 7426
rect 2223 7392 2257 7426
rect 2291 7392 2325 7426
rect 2359 7392 2393 7426
rect 2427 7392 2461 7426
rect 2495 7392 2529 7426
rect 2563 7392 2597 7426
rect 2631 7392 2665 7426
rect 2699 7392 2733 7426
rect 34 7381 2733 7392
rect 12498 7648 15102 7676
rect 12498 7640 14614 7648
rect 14648 7640 14692 7648
rect 14726 7640 14770 7648
rect 14804 7640 14848 7648
rect 14882 7640 14926 7648
rect 14960 7641 15004 7648
rect 15038 7641 15102 7648
rect 12498 7606 12524 7640
rect 12558 7606 12593 7640
rect 12627 7606 12662 7640
rect 12696 7606 12731 7640
rect 12765 7606 12800 7640
rect 12834 7606 12869 7640
rect 12903 7606 12938 7640
rect 12972 7606 13007 7640
rect 13041 7606 13076 7640
rect 13110 7606 13145 7640
rect 13179 7606 13214 7640
rect 13248 7606 13283 7640
rect 13317 7606 13352 7640
rect 13386 7606 13421 7640
rect 13455 7606 13490 7640
rect 13524 7606 13559 7640
rect 13593 7606 13628 7640
rect 13662 7606 13697 7640
rect 13731 7606 13766 7640
rect 13800 7606 13835 7640
rect 13869 7606 13904 7640
rect 13938 7606 13973 7640
rect 14007 7606 14042 7640
rect 14076 7606 14111 7640
rect 14145 7606 14180 7640
rect 14214 7606 14249 7640
rect 14283 7606 14318 7640
rect 14352 7606 14387 7640
rect 14421 7606 14456 7640
rect 14490 7606 14524 7640
rect 14558 7606 14592 7640
rect 14648 7614 14660 7640
rect 14726 7614 14728 7640
rect 14626 7606 14660 7614
rect 14694 7606 14728 7614
rect 14762 7614 14770 7640
rect 14830 7614 14848 7640
rect 14898 7614 14926 7640
rect 14762 7606 14796 7614
rect 14830 7606 14864 7614
rect 14898 7607 14932 7614
rect 14966 7607 15000 7641
rect 15038 7614 15068 7641
rect 15034 7607 15068 7614
rect 14898 7606 15102 7607
rect 12498 7574 15102 7606
rect 12498 7556 14614 7574
rect 14648 7556 14692 7574
rect 14726 7556 14770 7574
rect 14804 7556 14848 7574
rect 14882 7556 14926 7574
rect 14960 7569 15004 7574
rect 15038 7569 15102 7574
rect 12498 7522 12524 7556
rect 12558 7522 12593 7556
rect 12627 7522 12662 7556
rect 12696 7522 12731 7556
rect 12765 7522 12800 7556
rect 12834 7522 12869 7556
rect 12903 7522 12938 7556
rect 12972 7522 13007 7556
rect 13041 7522 13076 7556
rect 13110 7522 13145 7556
rect 13179 7522 13214 7556
rect 13248 7522 13283 7556
rect 13317 7522 13352 7556
rect 13386 7522 13421 7556
rect 13455 7522 13490 7556
rect 13524 7522 13559 7556
rect 13593 7522 13628 7556
rect 13662 7522 13697 7556
rect 13731 7522 13766 7556
rect 13800 7522 13835 7556
rect 13869 7522 13904 7556
rect 13938 7522 13973 7556
rect 14007 7522 14042 7556
rect 14076 7522 14111 7556
rect 14145 7522 14180 7556
rect 14214 7522 14249 7556
rect 14283 7522 14318 7556
rect 14352 7522 14387 7556
rect 14421 7522 14456 7556
rect 14490 7522 14524 7556
rect 14558 7522 14592 7556
rect 14648 7540 14660 7556
rect 14726 7540 14728 7556
rect 14626 7522 14660 7540
rect 14694 7522 14728 7540
rect 14762 7540 14770 7556
rect 14830 7540 14848 7556
rect 14898 7540 14926 7556
rect 14762 7522 14796 7540
rect 14830 7522 14864 7540
rect 14898 7535 14932 7540
rect 14966 7535 15000 7569
rect 15038 7540 15068 7569
rect 15034 7535 15068 7540
rect 14898 7522 15102 7535
rect 12498 7499 15102 7522
rect 12498 7472 14614 7499
rect 14648 7472 14692 7499
rect 14726 7472 14770 7499
rect 14804 7472 14848 7499
rect 14882 7472 14926 7499
rect 14960 7497 15004 7499
rect 15038 7497 15102 7499
rect 12498 7438 12524 7472
rect 12558 7438 12593 7472
rect 12627 7438 12662 7472
rect 12696 7438 12731 7472
rect 12765 7438 12800 7472
rect 12834 7438 12869 7472
rect 12903 7438 12938 7472
rect 12972 7438 13007 7472
rect 13041 7438 13076 7472
rect 13110 7438 13145 7472
rect 13179 7438 13214 7472
rect 13248 7438 13283 7472
rect 13317 7438 13352 7472
rect 13386 7438 13421 7472
rect 13455 7438 13490 7472
rect 13524 7438 13559 7472
rect 13593 7438 13628 7472
rect 13662 7438 13697 7472
rect 13731 7438 13766 7472
rect 13800 7438 13835 7472
rect 13869 7438 13904 7472
rect 13938 7438 13973 7472
rect 14007 7438 14042 7472
rect 14076 7438 14111 7472
rect 14145 7438 14180 7472
rect 14214 7438 14249 7472
rect 14283 7438 14318 7472
rect 14352 7438 14387 7472
rect 14421 7438 14456 7472
rect 14490 7438 14524 7472
rect 14558 7438 14592 7472
rect 14648 7465 14660 7472
rect 14726 7465 14728 7472
rect 14626 7438 14660 7465
rect 14694 7438 14728 7465
rect 14762 7465 14770 7472
rect 14830 7465 14848 7472
rect 14898 7465 14926 7472
rect 14762 7438 14796 7465
rect 14830 7438 14864 7465
rect 14898 7463 14932 7465
rect 14966 7463 15000 7497
rect 15038 7465 15068 7497
rect 15034 7463 15068 7465
rect 14898 7438 15102 7463
rect 12498 7425 15102 7438
rect 12498 7424 14932 7425
rect 12498 7390 14614 7424
rect 14648 7390 14692 7424
rect 14726 7390 14770 7424
rect 14804 7390 14848 7424
rect 14882 7390 14926 7424
rect 14966 7391 15000 7425
rect 15034 7424 15068 7425
rect 15038 7391 15068 7424
rect 14960 7390 15004 7391
rect 15038 7390 15102 7391
rect 12498 7388 15102 7390
rect 25 7374 7756 7381
rect 25 7340 57 7374
rect 91 7354 132 7374
rect 166 7354 207 7374
rect 241 7354 282 7374
rect 316 7354 357 7374
rect 391 7354 432 7374
rect 466 7354 507 7374
rect 541 7354 582 7374
rect 616 7354 657 7374
rect 691 7354 732 7374
rect 766 7354 807 7374
rect 841 7354 882 7374
rect 916 7354 957 7374
rect 991 7354 1032 7374
rect 1066 7354 1107 7374
rect 1141 7354 1182 7374
rect 1216 7354 1256 7374
rect 1290 7354 1330 7374
rect 1364 7354 7756 7374
rect 102 7340 132 7354
rect 25 7320 68 7340
rect 102 7320 137 7340
rect 171 7320 206 7354
rect 241 7340 275 7354
rect 316 7340 344 7354
rect 391 7340 413 7354
rect 466 7340 482 7354
rect 541 7340 551 7354
rect 616 7340 620 7354
rect 240 7320 275 7340
rect 309 7320 344 7340
rect 378 7320 413 7340
rect 447 7320 482 7340
rect 516 7320 551 7340
rect 585 7320 620 7340
rect 654 7340 657 7354
rect 723 7340 732 7354
rect 792 7340 807 7354
rect 861 7340 882 7354
rect 930 7340 957 7354
rect 999 7340 1032 7354
rect 654 7320 689 7340
rect 723 7320 758 7340
rect 792 7320 827 7340
rect 861 7320 896 7340
rect 930 7320 965 7340
rect 999 7320 1033 7340
rect 1067 7320 1101 7354
rect 1141 7340 1169 7354
rect 1216 7340 1237 7354
rect 1290 7340 1305 7354
rect 1364 7340 1373 7354
rect 1135 7320 1169 7340
rect 1203 7320 1237 7340
rect 1271 7320 1305 7340
rect 1339 7320 1373 7340
rect 1407 7320 1441 7354
rect 1475 7320 1509 7354
rect 1543 7320 1577 7354
rect 1611 7320 1645 7354
rect 1679 7320 1713 7354
rect 1747 7320 1781 7354
rect 1815 7320 1849 7354
rect 1883 7320 1917 7354
rect 1951 7320 1985 7354
rect 2019 7320 2053 7354
rect 2087 7320 2121 7354
rect 2155 7320 2189 7354
rect 2223 7320 2257 7354
rect 2291 7320 2325 7354
rect 2359 7320 2393 7354
rect 2427 7320 2461 7354
rect 2495 7320 2529 7354
rect 2563 7320 2597 7354
rect 2631 7320 2665 7354
rect 2699 7320 7756 7354
rect 25 7290 7756 7320
rect 12498 7354 12524 7388
rect 12558 7354 12593 7388
rect 12627 7354 12662 7388
rect 12696 7354 12731 7388
rect 12765 7354 12800 7388
rect 12834 7354 12869 7388
rect 12903 7354 12938 7388
rect 12972 7354 13007 7388
rect 13041 7354 13076 7388
rect 13110 7354 13145 7388
rect 13179 7354 13214 7388
rect 13248 7354 13283 7388
rect 13317 7354 13352 7388
rect 13386 7354 13421 7388
rect 13455 7354 13490 7388
rect 13524 7354 13559 7388
rect 13593 7354 13628 7388
rect 13662 7354 13697 7388
rect 13731 7354 13766 7388
rect 13800 7354 13835 7388
rect 13869 7354 13904 7388
rect 13938 7354 13973 7388
rect 14007 7354 14042 7388
rect 14076 7354 14111 7388
rect 14145 7354 14180 7388
rect 14214 7354 14249 7388
rect 14283 7354 14318 7388
rect 14352 7354 14387 7388
rect 14421 7354 14456 7388
rect 14490 7354 14524 7388
rect 14558 7354 14592 7388
rect 14626 7354 14660 7388
rect 14694 7354 14728 7388
rect 14762 7354 14796 7388
rect 14830 7354 14864 7388
rect 14898 7354 15102 7388
rect 12498 7353 15102 7354
rect 12498 7349 14932 7353
rect 12498 7317 14614 7349
rect 25 7256 57 7290
rect 91 7282 132 7290
rect 166 7282 207 7290
rect 241 7282 282 7290
rect 316 7282 357 7290
rect 391 7282 432 7290
rect 466 7282 507 7290
rect 541 7282 582 7290
rect 616 7282 657 7290
rect 691 7282 732 7290
rect 766 7282 807 7290
rect 841 7282 882 7290
rect 916 7282 957 7290
rect 991 7282 1032 7290
rect 1066 7282 1107 7290
rect 1141 7282 1182 7290
rect 1216 7282 1256 7290
rect 1290 7282 1330 7290
rect 1364 7282 7756 7290
rect 102 7256 132 7282
rect 25 7248 68 7256
rect 102 7248 137 7256
rect 171 7248 206 7282
rect 241 7256 275 7282
rect 316 7256 344 7282
rect 391 7256 413 7282
rect 466 7256 482 7282
rect 541 7256 551 7282
rect 616 7256 620 7282
rect 240 7248 275 7256
rect 309 7248 344 7256
rect 378 7248 413 7256
rect 447 7248 482 7256
rect 516 7248 551 7256
rect 585 7248 620 7256
rect 654 7256 657 7282
rect 723 7256 732 7282
rect 792 7256 807 7282
rect 861 7256 882 7282
rect 930 7256 957 7282
rect 999 7256 1032 7282
rect 654 7248 689 7256
rect 723 7248 758 7256
rect 792 7248 827 7256
rect 861 7248 896 7256
rect 930 7248 965 7256
rect 999 7248 1033 7256
rect 1067 7248 1101 7282
rect 1141 7256 1169 7282
rect 1216 7256 1237 7282
rect 1290 7256 1305 7282
rect 1364 7256 1373 7282
rect 1135 7248 1169 7256
rect 1203 7248 1237 7256
rect 1271 7248 1305 7256
rect 1339 7248 1373 7256
rect 1407 7248 1441 7282
rect 1475 7248 1509 7282
rect 1543 7248 1577 7282
rect 1611 7248 1645 7282
rect 1679 7248 1713 7282
rect 1747 7248 1781 7282
rect 1815 7248 1849 7282
rect 1883 7248 1917 7282
rect 1951 7248 1985 7282
rect 2019 7248 2053 7282
rect 2087 7248 2121 7282
rect 2155 7248 2189 7282
rect 2223 7248 2257 7282
rect 2291 7248 2325 7282
rect 2359 7248 2393 7282
rect 2427 7248 2461 7282
rect 2495 7248 2529 7282
rect 2563 7248 2597 7282
rect 2631 7248 2665 7282
rect 2699 7248 7756 7282
rect 25 7220 7756 7248
rect 25 7210 1431 7220
rect 1465 7210 1504 7220
rect 1538 7210 1577 7220
rect 1611 7210 1650 7220
rect 1684 7210 1723 7220
rect 1757 7210 1796 7220
rect 1830 7210 1869 7220
rect 1903 7210 1942 7220
rect 1976 7210 2015 7220
rect 2049 7210 2088 7220
rect 2122 7210 2161 7220
rect 2195 7210 2234 7220
rect 2268 7210 2307 7220
rect 2341 7210 2380 7220
rect 2414 7210 2453 7220
rect 2487 7210 2526 7220
rect 2560 7210 2599 7220
rect 2633 7210 2672 7220
rect 25 7206 68 7210
rect 102 7206 137 7210
rect 25 7172 57 7206
rect 102 7176 132 7206
rect 171 7176 206 7210
rect 240 7206 275 7210
rect 309 7206 344 7210
rect 378 7206 413 7210
rect 447 7206 482 7210
rect 516 7206 551 7210
rect 585 7206 620 7210
rect 241 7176 275 7206
rect 316 7176 344 7206
rect 391 7176 413 7206
rect 466 7176 482 7206
rect 541 7176 551 7206
rect 616 7176 620 7206
rect 654 7206 689 7210
rect 723 7206 758 7210
rect 792 7206 827 7210
rect 861 7206 896 7210
rect 930 7206 965 7210
rect 999 7206 1033 7210
rect 654 7176 657 7206
rect 723 7176 732 7206
rect 792 7176 807 7206
rect 861 7176 882 7206
rect 930 7176 957 7206
rect 999 7176 1032 7206
rect 1067 7176 1101 7210
rect 1135 7206 1169 7210
rect 1203 7206 1237 7210
rect 1271 7206 1305 7210
rect 1339 7206 1373 7210
rect 1141 7176 1169 7206
rect 1216 7176 1237 7206
rect 1290 7176 1305 7206
rect 1364 7176 1373 7206
rect 1407 7186 1431 7210
rect 1475 7186 1504 7210
rect 1407 7176 1441 7186
rect 1475 7176 1509 7186
rect 1543 7176 1577 7210
rect 1611 7176 1645 7210
rect 1684 7186 1713 7210
rect 1757 7186 1781 7210
rect 1830 7186 1849 7210
rect 1903 7186 1917 7210
rect 1976 7186 1985 7210
rect 2049 7186 2053 7210
rect 1679 7176 1713 7186
rect 1747 7176 1781 7186
rect 1815 7176 1849 7186
rect 1883 7176 1917 7186
rect 1951 7176 1985 7186
rect 2019 7176 2053 7186
rect 2087 7186 2088 7210
rect 2155 7186 2161 7210
rect 2223 7186 2234 7210
rect 2291 7186 2307 7210
rect 2359 7186 2380 7210
rect 2427 7186 2453 7210
rect 2495 7186 2526 7210
rect 2087 7176 2121 7186
rect 2155 7176 2189 7186
rect 2223 7176 2257 7186
rect 2291 7176 2325 7186
rect 2359 7176 2393 7186
rect 2427 7176 2461 7186
rect 2495 7176 2529 7186
rect 2563 7176 2597 7210
rect 2633 7186 2665 7210
rect 2706 7186 2745 7220
rect 2779 7186 2818 7220
rect 2852 7186 2891 7220
rect 2925 7186 2964 7220
rect 2998 7186 3037 7220
rect 3071 7186 3110 7220
rect 3144 7186 3183 7220
rect 3217 7186 3256 7220
rect 3290 7186 3329 7220
rect 3363 7186 3402 7220
rect 3436 7186 3475 7220
rect 3509 7186 3548 7220
rect 3582 7186 3621 7220
rect 3655 7186 3694 7220
rect 3728 7186 3767 7220
rect 3801 7186 3840 7220
rect 3874 7186 3913 7220
rect 3947 7186 3986 7220
rect 4020 7186 4059 7220
rect 4093 7186 4132 7220
rect 4166 7186 4205 7220
rect 4239 7186 4278 7220
rect 4312 7186 4351 7220
rect 4385 7186 4424 7220
rect 4458 7186 4497 7220
rect 4531 7186 4570 7220
rect 4604 7186 4643 7220
rect 4677 7186 4716 7220
rect 4750 7186 4789 7220
rect 4823 7186 4862 7220
rect 4896 7186 4935 7220
rect 4969 7186 5008 7220
rect 5042 7186 5081 7220
rect 5115 7186 5154 7220
rect 5188 7186 5227 7220
rect 5261 7186 5300 7220
rect 5334 7186 5373 7220
rect 5407 7186 5446 7220
rect 5480 7186 5519 7220
rect 5553 7186 5592 7220
rect 5626 7186 5665 7220
rect 5699 7186 5738 7220
rect 5772 7186 5811 7220
rect 5845 7186 5884 7220
rect 5918 7186 5957 7220
rect 5991 7186 6030 7220
rect 6064 7186 6103 7220
rect 6137 7186 6176 7220
rect 6210 7186 6249 7220
rect 6283 7186 6322 7220
rect 6356 7186 6395 7220
rect 6429 7186 6468 7220
rect 6502 7186 6540 7220
rect 6574 7186 6612 7220
rect 6646 7186 6684 7220
rect 6718 7186 6756 7220
rect 6790 7186 6828 7220
rect 6862 7186 6900 7220
rect 6934 7186 6972 7220
rect 7006 7186 7044 7220
rect 7078 7186 7116 7220
rect 7150 7186 7756 7220
rect 2631 7176 2665 7186
rect 2699 7176 7756 7186
rect 91 7172 132 7176
rect 166 7172 207 7176
rect 241 7172 282 7176
rect 316 7172 357 7176
rect 391 7172 432 7176
rect 466 7172 507 7176
rect 541 7172 582 7176
rect 616 7172 657 7176
rect 691 7172 732 7176
rect 766 7172 807 7176
rect 841 7172 882 7176
rect 916 7172 957 7176
rect 991 7172 1032 7176
rect 1066 7172 1107 7176
rect 1141 7172 1182 7176
rect 1216 7172 1256 7176
rect 1290 7172 1330 7176
rect 1364 7172 7756 7176
rect 25 7138 7756 7172
rect 25 7122 68 7138
rect 102 7122 137 7138
rect 25 7088 57 7122
rect 102 7104 132 7122
rect 171 7104 206 7138
rect 240 7122 275 7138
rect 309 7122 344 7138
rect 378 7122 413 7138
rect 447 7122 482 7138
rect 516 7122 551 7138
rect 585 7122 620 7138
rect 241 7104 275 7122
rect 316 7104 344 7122
rect 391 7104 413 7122
rect 466 7104 482 7122
rect 541 7104 551 7122
rect 616 7104 620 7122
rect 654 7122 689 7138
rect 723 7122 758 7138
rect 792 7122 827 7138
rect 861 7122 896 7138
rect 930 7122 965 7138
rect 999 7122 1033 7138
rect 654 7104 657 7122
rect 723 7104 732 7122
rect 792 7104 807 7122
rect 861 7104 882 7122
rect 930 7104 957 7122
rect 999 7104 1032 7122
rect 1067 7104 1101 7138
rect 1135 7122 1169 7138
rect 1203 7122 1237 7138
rect 1271 7122 1305 7138
rect 1339 7122 1373 7138
rect 1141 7104 1169 7122
rect 1216 7104 1237 7122
rect 1290 7104 1305 7122
rect 1364 7104 1373 7122
rect 1407 7104 1441 7138
rect 1475 7104 1509 7138
rect 1543 7104 1577 7138
rect 1611 7104 1645 7138
rect 1679 7104 1713 7138
rect 1747 7104 1781 7138
rect 1815 7104 1849 7138
rect 1883 7104 1917 7138
rect 1951 7104 1985 7138
rect 2019 7104 2053 7138
rect 2087 7104 2121 7138
rect 2155 7104 2189 7138
rect 2223 7104 2257 7138
rect 2291 7104 2325 7138
rect 2359 7104 2393 7138
rect 2427 7104 2461 7138
rect 2495 7104 2529 7138
rect 2563 7104 2597 7138
rect 2631 7104 2665 7138
rect 2699 7104 7756 7138
rect 91 7088 132 7104
rect 166 7088 207 7104
rect 241 7088 282 7104
rect 316 7088 357 7104
rect 391 7088 432 7104
rect 466 7088 507 7104
rect 541 7088 582 7104
rect 616 7088 657 7104
rect 691 7088 732 7104
rect 766 7088 807 7104
rect 841 7088 882 7104
rect 916 7088 957 7104
rect 991 7088 1032 7104
rect 1066 7088 1107 7104
rect 1141 7088 1182 7104
rect 1216 7088 1256 7104
rect 1290 7088 1330 7104
rect 1364 7088 7756 7104
rect 25 7066 7756 7088
rect 25 7038 68 7066
rect 102 7038 137 7066
rect 25 7004 57 7038
rect 102 7032 132 7038
rect 171 7032 206 7066
rect 240 7038 275 7066
rect 309 7038 344 7066
rect 378 7038 413 7066
rect 447 7038 482 7066
rect 516 7038 551 7066
rect 585 7038 620 7066
rect 241 7032 275 7038
rect 316 7032 344 7038
rect 391 7032 413 7038
rect 466 7032 482 7038
rect 541 7032 551 7038
rect 616 7032 620 7038
rect 654 7038 689 7066
rect 723 7038 758 7066
rect 792 7038 827 7066
rect 861 7038 896 7066
rect 930 7038 965 7066
rect 999 7038 1033 7066
rect 654 7032 657 7038
rect 723 7032 732 7038
rect 792 7032 807 7038
rect 861 7032 882 7038
rect 930 7032 957 7038
rect 999 7032 1032 7038
rect 1067 7032 1101 7066
rect 1135 7038 1169 7066
rect 1203 7038 1237 7066
rect 1271 7038 1305 7066
rect 1339 7038 1373 7066
rect 1141 7032 1169 7038
rect 1216 7032 1237 7038
rect 1290 7032 1305 7038
rect 1364 7032 1373 7038
rect 1407 7032 1441 7066
rect 1475 7032 1509 7066
rect 1543 7032 1577 7066
rect 1611 7032 1645 7066
rect 1679 7032 1713 7066
rect 1747 7032 1781 7066
rect 1815 7032 1849 7066
rect 1883 7032 1917 7066
rect 1951 7032 1985 7066
rect 2019 7032 2053 7066
rect 2087 7032 2121 7066
rect 2155 7032 2189 7066
rect 2223 7032 2257 7066
rect 2291 7032 2325 7066
rect 2359 7032 2393 7066
rect 2427 7032 2461 7066
rect 2495 7032 2529 7066
rect 2563 7032 2597 7066
rect 2631 7032 2665 7066
rect 2699 7047 7756 7066
rect 2699 7032 2757 7047
rect 91 7004 132 7032
rect 166 7004 207 7032
rect 241 7004 282 7032
rect 316 7004 357 7032
rect 391 7004 432 7032
rect 466 7004 507 7032
rect 541 7004 582 7032
rect 616 7004 657 7032
rect 691 7004 732 7032
rect 766 7004 807 7032
rect 841 7004 882 7032
rect 916 7004 957 7032
rect 991 7004 1032 7032
rect 1066 7004 1107 7032
rect 1141 7004 1182 7032
rect 1216 7004 1256 7032
rect 1290 7004 1330 7032
rect 1364 7013 2757 7032
rect 2791 7013 2825 7047
rect 2859 7013 2893 7047
rect 2927 7013 2961 7047
rect 2995 7013 3029 7047
rect 3063 7013 3097 7047
rect 3131 7013 3165 7047
rect 3199 7013 3233 7047
rect 3267 7013 3301 7047
rect 3335 7013 3369 7047
rect 3403 7013 3437 7047
rect 3471 7013 3505 7047
rect 3539 7013 3573 7047
rect 3607 7013 3641 7047
rect 3675 7013 3709 7047
rect 3743 7013 3777 7047
rect 3811 7013 3845 7047
rect 3879 7013 3913 7047
rect 3947 7013 3981 7047
rect 4015 7013 4049 7047
rect 4083 7013 4117 7047
rect 4151 7013 4185 7047
rect 4219 7013 4253 7047
rect 4287 7013 4321 7047
rect 4355 7013 4389 7047
rect 4423 7013 4457 7047
rect 4491 7013 4525 7047
rect 4559 7013 4593 7047
rect 4627 7013 4661 7047
rect 4695 7013 4729 7047
rect 4763 7013 4797 7047
rect 4831 7013 4865 7047
rect 4899 7013 4933 7047
rect 4967 7013 5001 7047
rect 5035 7013 5069 7047
rect 5103 7013 5137 7047
rect 5171 7013 5205 7047
rect 5239 7013 5273 7047
rect 5307 7013 5341 7047
rect 5375 7013 5409 7047
rect 5443 7013 5477 7047
rect 5511 7013 5545 7047
rect 5579 7013 5613 7047
rect 5647 7013 5681 7047
rect 5715 7013 5749 7047
rect 5783 7013 5817 7047
rect 5851 7013 5885 7047
rect 5919 7013 5953 7047
rect 5987 7013 6021 7047
rect 6055 7013 6089 7047
rect 6123 7013 6157 7047
rect 6191 7013 6225 7047
rect 6259 7013 6293 7047
rect 6327 7013 6361 7047
rect 6395 7013 6429 7047
rect 6463 7013 6497 7047
rect 6531 7013 6565 7047
rect 6599 7013 6633 7047
rect 6667 7013 6701 7047
rect 6735 7013 6769 7047
rect 6803 7013 6837 7047
rect 6871 7013 6905 7047
rect 6939 7013 6973 7047
rect 7007 7013 7041 7047
rect 7075 7013 7109 7047
rect 7143 7013 7177 7047
rect 7211 7013 7245 7047
rect 7279 7013 7313 7047
rect 7347 7013 7381 7047
rect 7415 7013 7449 7047
rect 7483 7013 7517 7047
rect 7551 7013 7585 7047
rect 7619 7013 7653 7047
rect 7687 7013 7756 7047
rect 1364 7004 7756 7013
rect 25 6997 7756 7004
rect 7183 6957 7756 6997
rect 8184 7315 14614 7317
rect 14648 7315 14692 7349
rect 14726 7315 14770 7349
rect 14804 7315 14848 7349
rect 14882 7315 14926 7349
rect 14966 7319 15000 7353
rect 15034 7349 15068 7353
rect 15038 7319 15068 7349
rect 14960 7315 15004 7319
rect 15038 7315 15102 7319
rect 8184 7282 15102 7315
rect 8184 7248 8210 7282
rect 8244 7248 8279 7282
rect 8313 7248 8348 7282
rect 8382 7248 8417 7282
rect 8451 7248 8486 7282
rect 8520 7248 8555 7282
rect 8589 7248 8624 7282
rect 8658 7248 8693 7282
rect 8727 7248 8762 7282
rect 8796 7248 8831 7282
rect 8865 7248 8900 7282
rect 8934 7248 8969 7282
rect 9003 7248 9038 7282
rect 9072 7248 9107 7282
rect 9141 7248 9176 7282
rect 9210 7248 9245 7282
rect 9279 7248 9314 7282
rect 9348 7248 9383 7282
rect 9417 7248 9452 7282
rect 9486 7248 9521 7282
rect 9555 7248 9590 7282
rect 9624 7248 9659 7282
rect 9693 7248 9728 7282
rect 9762 7248 9797 7282
rect 9831 7248 9866 7282
rect 9900 7248 9935 7282
rect 9969 7248 10004 7282
rect 10038 7248 10073 7282
rect 10107 7248 10142 7282
rect 10176 7248 10211 7282
rect 10245 7248 10280 7282
rect 10314 7248 10349 7282
rect 10383 7248 10418 7282
rect 10452 7248 10487 7282
rect 10521 7248 10556 7282
rect 10590 7248 10625 7282
rect 10659 7248 10694 7282
rect 10728 7248 10763 7282
rect 10797 7248 10832 7282
rect 10866 7248 10901 7282
rect 10935 7248 10970 7282
rect 11004 7248 11039 7282
rect 11073 7248 11108 7282
rect 11142 7248 11177 7282
rect 11211 7248 11246 7282
rect 11280 7248 11315 7282
rect 11349 7248 11384 7282
rect 11418 7248 11453 7282
rect 11487 7248 11522 7282
rect 11556 7248 11591 7282
rect 11625 7248 11660 7282
rect 11694 7248 11729 7282
rect 11763 7248 11798 7282
rect 11832 7248 11867 7282
rect 11901 7248 11936 7282
rect 11970 7248 12005 7282
rect 12039 7248 12074 7282
rect 12108 7248 12143 7282
rect 12177 7248 12212 7282
rect 12246 7248 12280 7282
rect 12314 7248 12348 7282
rect 12382 7248 12416 7282
rect 12450 7248 12484 7282
rect 12518 7248 12552 7282
rect 12586 7248 12620 7282
rect 12654 7248 12688 7282
rect 12722 7248 12756 7282
rect 12790 7248 12824 7282
rect 12858 7248 12892 7282
rect 12926 7248 12960 7282
rect 12994 7248 13028 7282
rect 13062 7248 13096 7282
rect 13130 7248 13164 7282
rect 13198 7248 13232 7282
rect 13266 7248 13300 7282
rect 13334 7248 13368 7282
rect 13402 7248 13436 7282
rect 13470 7248 13504 7282
rect 13538 7248 13572 7282
rect 13606 7248 13640 7282
rect 13674 7248 13708 7282
rect 13742 7248 13776 7282
rect 13810 7248 13844 7282
rect 13878 7248 13912 7282
rect 13946 7248 13980 7282
rect 14014 7248 14048 7282
rect 14082 7248 14116 7282
rect 14150 7248 14184 7282
rect 14218 7248 14252 7282
rect 14286 7248 14320 7282
rect 14354 7248 14388 7282
rect 14422 7248 14456 7282
rect 14490 7248 14524 7282
rect 14558 7248 14592 7282
rect 14626 7274 14660 7282
rect 14694 7274 14728 7282
rect 14648 7248 14660 7274
rect 14726 7248 14728 7274
rect 14762 7274 14796 7282
rect 14830 7274 14864 7282
rect 14898 7281 15102 7282
rect 14898 7274 14932 7281
rect 14762 7248 14770 7274
rect 14830 7248 14848 7274
rect 14898 7248 14926 7274
rect 8184 7240 14614 7248
rect 14648 7240 14692 7248
rect 14726 7240 14770 7248
rect 14804 7240 14848 7248
rect 14882 7240 14926 7248
rect 14966 7247 15000 7281
rect 15034 7274 15068 7281
rect 15038 7247 15068 7274
rect 14960 7240 15004 7247
rect 15038 7240 15102 7247
rect 8184 7210 15102 7240
rect 8184 7176 8210 7210
rect 8244 7176 8279 7210
rect 8313 7176 8348 7210
rect 8382 7176 8417 7210
rect 8451 7176 8486 7210
rect 8520 7176 8555 7210
rect 8589 7176 8624 7210
rect 8658 7176 8693 7210
rect 8727 7176 8762 7210
rect 8796 7176 8831 7210
rect 8865 7176 8900 7210
rect 8934 7176 8969 7210
rect 9003 7176 9038 7210
rect 9072 7176 9107 7210
rect 9141 7176 9176 7210
rect 9210 7176 9245 7210
rect 9279 7176 9314 7210
rect 9348 7176 9383 7210
rect 9417 7176 9452 7210
rect 9486 7176 9521 7210
rect 9555 7176 9590 7210
rect 9624 7176 9659 7210
rect 9693 7176 9728 7210
rect 9762 7176 9797 7210
rect 9831 7176 9866 7210
rect 9900 7176 9935 7210
rect 9969 7176 10004 7210
rect 10038 7176 10073 7210
rect 10107 7176 10142 7210
rect 10176 7176 10211 7210
rect 10245 7176 10280 7210
rect 10314 7176 10349 7210
rect 10383 7176 10418 7210
rect 10452 7176 10487 7210
rect 10521 7176 10556 7210
rect 10590 7176 10625 7210
rect 10659 7176 10694 7210
rect 10728 7176 10763 7210
rect 10797 7176 10832 7210
rect 10866 7176 10901 7210
rect 10935 7176 10970 7210
rect 11004 7176 11039 7210
rect 11073 7176 11108 7210
rect 11142 7176 11177 7210
rect 11211 7176 11246 7210
rect 11280 7176 11315 7210
rect 11349 7176 11384 7210
rect 11418 7176 11453 7210
rect 11487 7176 11522 7210
rect 11556 7176 11591 7210
rect 11625 7176 11660 7210
rect 11694 7176 11729 7210
rect 11763 7176 11798 7210
rect 11832 7176 11867 7210
rect 11901 7176 11936 7210
rect 11970 7176 12005 7210
rect 12039 7176 12074 7210
rect 12108 7176 12143 7210
rect 12177 7176 12212 7210
rect 12246 7176 12280 7210
rect 12314 7176 12348 7210
rect 12382 7176 12416 7210
rect 12450 7176 12484 7210
rect 12518 7176 12552 7210
rect 12586 7176 12620 7210
rect 12654 7176 12688 7210
rect 12722 7176 12756 7210
rect 12790 7176 12824 7210
rect 12858 7176 12892 7210
rect 12926 7176 12960 7210
rect 12994 7176 13028 7210
rect 13062 7176 13096 7210
rect 13130 7176 13164 7210
rect 13198 7176 13232 7210
rect 13266 7176 13300 7210
rect 13334 7176 13368 7210
rect 13402 7176 13436 7210
rect 13470 7176 13504 7210
rect 13538 7176 13572 7210
rect 13606 7176 13640 7210
rect 13674 7176 13708 7210
rect 13742 7176 13776 7210
rect 13810 7176 13844 7210
rect 13878 7176 13912 7210
rect 13946 7176 13980 7210
rect 14014 7176 14048 7210
rect 14082 7176 14116 7210
rect 14150 7176 14184 7210
rect 14218 7176 14252 7210
rect 14286 7176 14320 7210
rect 14354 7176 14388 7210
rect 14422 7176 14456 7210
rect 14490 7176 14524 7210
rect 14558 7176 14592 7210
rect 14626 7199 14660 7210
rect 14694 7199 14728 7210
rect 14648 7176 14660 7199
rect 14726 7176 14728 7199
rect 14762 7199 14796 7210
rect 14830 7199 14864 7210
rect 14898 7209 15102 7210
rect 14898 7199 14932 7209
rect 14762 7176 14770 7199
rect 14830 7176 14848 7199
rect 14898 7176 14926 7199
rect 8184 7165 14614 7176
rect 14648 7165 14692 7176
rect 14726 7165 14770 7176
rect 14804 7165 14848 7176
rect 14882 7165 14926 7176
rect 14966 7175 15000 7209
rect 15034 7199 15068 7209
rect 15038 7175 15068 7199
rect 14960 7165 15004 7175
rect 15038 7165 15102 7175
rect 8184 7138 15102 7165
rect 8184 7104 8210 7138
rect 8244 7104 8279 7138
rect 8313 7104 8348 7138
rect 8382 7104 8417 7138
rect 8451 7104 8486 7138
rect 8520 7104 8555 7138
rect 8589 7104 8624 7138
rect 8658 7104 8693 7138
rect 8727 7104 8762 7138
rect 8796 7104 8831 7138
rect 8865 7104 8900 7138
rect 8934 7104 8969 7138
rect 9003 7104 9038 7138
rect 9072 7104 9107 7138
rect 9141 7104 9176 7138
rect 9210 7104 9245 7138
rect 9279 7104 9314 7138
rect 9348 7104 9383 7138
rect 9417 7104 9452 7138
rect 9486 7104 9521 7138
rect 9555 7104 9590 7138
rect 9624 7104 9659 7138
rect 9693 7104 9728 7138
rect 9762 7104 9797 7138
rect 9831 7104 9866 7138
rect 9900 7104 9935 7138
rect 9969 7104 10004 7138
rect 10038 7104 10073 7138
rect 10107 7104 10142 7138
rect 10176 7104 10211 7138
rect 10245 7104 10280 7138
rect 10314 7104 10349 7138
rect 10383 7104 10418 7138
rect 10452 7104 10487 7138
rect 10521 7104 10556 7138
rect 10590 7104 10625 7138
rect 10659 7104 10694 7138
rect 10728 7104 10763 7138
rect 10797 7104 10832 7138
rect 10866 7104 10901 7138
rect 10935 7104 10970 7138
rect 11004 7104 11039 7138
rect 11073 7104 11108 7138
rect 11142 7104 11177 7138
rect 11211 7104 11246 7138
rect 11280 7104 11315 7138
rect 11349 7104 11384 7138
rect 11418 7104 11453 7138
rect 11487 7104 11522 7138
rect 11556 7104 11591 7138
rect 11625 7104 11660 7138
rect 11694 7104 11729 7138
rect 11763 7104 11798 7138
rect 11832 7104 11867 7138
rect 11901 7104 11936 7138
rect 11970 7104 12005 7138
rect 12039 7104 12074 7138
rect 12108 7104 12143 7138
rect 12177 7104 12212 7138
rect 12246 7104 12280 7138
rect 12314 7104 12348 7138
rect 12382 7104 12416 7138
rect 12450 7104 12484 7138
rect 12518 7104 12552 7138
rect 12586 7104 12620 7138
rect 12654 7104 12688 7138
rect 12722 7104 12756 7138
rect 12790 7104 12824 7138
rect 12858 7104 12892 7138
rect 12926 7104 12960 7138
rect 12994 7104 13028 7138
rect 13062 7104 13096 7138
rect 13130 7104 13164 7138
rect 13198 7104 13232 7138
rect 13266 7104 13300 7138
rect 13334 7104 13368 7138
rect 13402 7104 13436 7138
rect 13470 7104 13504 7138
rect 13538 7104 13572 7138
rect 13606 7104 13640 7138
rect 13674 7104 13708 7138
rect 13742 7104 13776 7138
rect 13810 7104 13844 7138
rect 13878 7104 13912 7138
rect 13946 7104 13980 7138
rect 14014 7104 14048 7138
rect 14082 7104 14116 7138
rect 14150 7104 14184 7138
rect 14218 7104 14252 7138
rect 14286 7104 14320 7138
rect 14354 7104 14388 7138
rect 14422 7104 14456 7138
rect 14490 7104 14524 7138
rect 14558 7104 14592 7138
rect 14626 7124 14660 7138
rect 14694 7124 14728 7138
rect 14648 7104 14660 7124
rect 14726 7104 14728 7124
rect 14762 7124 14796 7138
rect 14830 7124 14864 7138
rect 14898 7137 15102 7138
rect 14898 7124 14932 7137
rect 14762 7104 14770 7124
rect 14830 7104 14848 7124
rect 14898 7104 14926 7124
rect 8184 7090 14614 7104
rect 14648 7090 14692 7104
rect 14726 7090 14770 7104
rect 14804 7090 14848 7104
rect 14882 7090 14926 7104
rect 14966 7103 15000 7137
rect 15034 7124 15068 7137
rect 15038 7103 15068 7124
rect 14960 7090 15004 7103
rect 15038 7090 15102 7103
rect 8184 7066 15102 7090
rect 8184 7032 8210 7066
rect 8244 7032 8279 7066
rect 8313 7032 8348 7066
rect 8382 7032 8417 7066
rect 8451 7032 8486 7066
rect 8520 7032 8555 7066
rect 8589 7032 8624 7066
rect 8658 7032 8693 7066
rect 8727 7032 8762 7066
rect 8796 7032 8831 7066
rect 8865 7032 8900 7066
rect 8934 7032 8969 7066
rect 9003 7032 9038 7066
rect 9072 7032 9107 7066
rect 9141 7032 9176 7066
rect 9210 7032 9245 7066
rect 9279 7032 9314 7066
rect 9348 7032 9383 7066
rect 9417 7032 9452 7066
rect 9486 7032 9521 7066
rect 9555 7032 9590 7066
rect 9624 7032 9659 7066
rect 9693 7032 9728 7066
rect 9762 7032 9797 7066
rect 9831 7032 9866 7066
rect 9900 7032 9935 7066
rect 9969 7032 10004 7066
rect 10038 7032 10073 7066
rect 10107 7032 10142 7066
rect 10176 7032 10211 7066
rect 10245 7032 10280 7066
rect 10314 7032 10349 7066
rect 10383 7032 10418 7066
rect 10452 7032 10487 7066
rect 10521 7032 10556 7066
rect 10590 7032 10625 7066
rect 10659 7032 10694 7066
rect 10728 7032 10763 7066
rect 10797 7032 10832 7066
rect 10866 7032 10901 7066
rect 10935 7032 10970 7066
rect 11004 7032 11039 7066
rect 11073 7032 11108 7066
rect 11142 7032 11177 7066
rect 11211 7032 11246 7066
rect 11280 7032 11315 7066
rect 11349 7032 11384 7066
rect 11418 7032 11453 7066
rect 11487 7032 11522 7066
rect 11556 7032 11591 7066
rect 11625 7032 11660 7066
rect 11694 7032 11729 7066
rect 11763 7032 11798 7066
rect 11832 7032 11867 7066
rect 11901 7032 11936 7066
rect 11970 7032 12005 7066
rect 12039 7032 12074 7066
rect 12108 7032 12143 7066
rect 12177 7032 12212 7066
rect 12246 7032 12280 7066
rect 12314 7032 12348 7066
rect 12382 7032 12416 7066
rect 12450 7032 12484 7066
rect 12518 7032 12552 7066
rect 12586 7032 12620 7066
rect 12654 7032 12688 7066
rect 12722 7032 12756 7066
rect 12790 7032 12824 7066
rect 12858 7032 12892 7066
rect 12926 7032 12960 7066
rect 12994 7032 13028 7066
rect 13062 7032 13096 7066
rect 13130 7032 13164 7066
rect 13198 7032 13232 7066
rect 13266 7032 13300 7066
rect 13334 7032 13368 7066
rect 13402 7032 13436 7066
rect 13470 7032 13504 7066
rect 13538 7032 13572 7066
rect 13606 7032 13640 7066
rect 13674 7032 13708 7066
rect 13742 7032 13776 7066
rect 13810 7032 13844 7066
rect 13878 7032 13912 7066
rect 13946 7032 13980 7066
rect 14014 7032 14048 7066
rect 14082 7032 14116 7066
rect 14150 7032 14184 7066
rect 14218 7032 14252 7066
rect 14286 7032 14320 7066
rect 14354 7032 14388 7066
rect 14422 7032 14456 7066
rect 14490 7032 14524 7066
rect 14558 7032 14592 7066
rect 14626 7032 14660 7066
rect 14694 7032 14728 7066
rect 14762 7032 14796 7066
rect 14830 7032 14864 7066
rect 14898 7065 15102 7066
rect 14898 7032 14932 7065
rect 8184 7031 14932 7032
rect 14966 7031 15000 7065
rect 15034 7031 15068 7065
rect 8184 6997 15102 7031
rect 8184 6957 8488 6997
rect 44 6809 68 6843
rect 102 6809 137 6843
rect 171 6809 206 6843
rect 240 6809 275 6843
rect 309 6809 344 6843
rect 378 6809 413 6843
rect 447 6809 482 6843
rect 516 6809 551 6843
rect 585 6809 620 6843
rect 654 6809 689 6843
rect 723 6809 758 6843
rect 792 6809 827 6843
rect 861 6809 896 6843
rect 930 6809 965 6843
rect 999 6809 1034 6843
rect 1068 6809 1103 6843
rect 1137 6809 1172 6843
rect 1206 6809 1241 6843
rect 1275 6809 1310 6843
rect 1344 6809 1379 6843
rect 1413 6809 1448 6843
rect 1482 6809 1517 6843
rect 1551 6809 1586 6843
rect 1620 6809 1655 6843
rect 1689 6809 1724 6843
rect 1758 6809 1793 6843
rect 1827 6809 1862 6843
rect 1896 6809 1931 6843
rect 1965 6809 2000 6843
rect 2034 6809 2069 6843
rect 2103 6809 2138 6843
rect 2172 6809 2207 6843
rect 2241 6809 2276 6843
rect 2310 6809 2345 6843
rect 2379 6809 2414 6843
rect 2448 6809 2483 6843
rect 2517 6809 2552 6843
rect 2586 6809 2621 6843
rect 2655 6809 2690 6843
rect 2724 6809 2759 6843
rect 2793 6809 2828 6843
rect 2862 6809 2897 6843
rect 2931 6809 2966 6843
rect 3000 6809 3035 6843
rect 3069 6809 3104 6843
rect 3138 6809 3173 6843
rect 3207 6809 3242 6843
rect 3276 6809 3310 6843
rect 3344 6809 3378 6843
rect 3412 6809 3446 6843
rect 3480 6809 3514 6843
rect 3548 6809 3582 6843
rect 3616 6809 3650 6843
rect 3684 6809 3718 6843
rect 3752 6809 3786 6843
rect 3820 6809 3854 6843
rect 3888 6809 3922 6843
rect 3956 6809 3990 6843
rect 4024 6809 4058 6843
rect 4092 6809 4126 6843
rect 4160 6809 4194 6843
rect 4228 6809 4262 6843
rect 4296 6809 4330 6843
rect 4364 6809 4398 6843
rect 4432 6809 4466 6843
rect 4500 6809 4534 6843
rect 4568 6809 4602 6843
rect 4636 6809 4670 6843
rect 4704 6809 4738 6843
rect 4772 6809 4806 6843
rect 4840 6809 4874 6843
rect 4908 6809 4942 6843
rect 4976 6809 5010 6843
rect 5044 6809 5078 6843
rect 5112 6809 5146 6843
rect 5180 6809 5214 6843
rect 5248 6809 5282 6843
rect 5316 6809 5350 6843
rect 5384 6809 5418 6843
rect 5452 6809 5486 6843
rect 5520 6809 5554 6843
rect 5588 6809 5622 6843
rect 5656 6809 5690 6843
rect 5724 6809 5758 6843
rect 5792 6809 5826 6843
rect 5860 6809 5894 6843
rect 5928 6809 5962 6843
rect 5996 6809 6030 6843
rect 6064 6809 6098 6843
rect 6132 6809 6166 6843
rect 6200 6809 6234 6843
rect 6268 6809 6302 6843
rect 6336 6809 6370 6843
rect 6404 6809 6438 6843
rect 6472 6809 6506 6843
rect 6540 6809 6574 6843
rect 6608 6809 6642 6843
rect 6676 6809 6710 6843
rect 6744 6809 6778 6843
rect 6812 6809 6846 6843
rect 6880 6809 6914 6843
rect 6948 6809 6982 6843
rect 7016 6809 7050 6843
rect 7084 6809 7108 6843
rect 44 6756 7108 6809
rect 44 6722 68 6756
rect 102 6722 137 6756
rect 171 6722 206 6756
rect 240 6722 275 6756
rect 309 6722 344 6756
rect 378 6722 413 6756
rect 447 6722 482 6756
rect 516 6722 551 6756
rect 585 6722 620 6756
rect 654 6722 689 6756
rect 723 6722 758 6756
rect 792 6722 827 6756
rect 861 6722 896 6756
rect 930 6722 965 6756
rect 999 6722 1034 6756
rect 1068 6722 1103 6756
rect 1137 6722 1172 6756
rect 1206 6722 1241 6756
rect 1275 6722 1310 6756
rect 1344 6722 1379 6756
rect 1413 6722 1448 6756
rect 1482 6722 1517 6756
rect 1551 6722 1586 6756
rect 1620 6722 1655 6756
rect 1689 6722 1724 6756
rect 1758 6722 1793 6756
rect 1827 6722 1862 6756
rect 1896 6722 1931 6756
rect 1965 6722 2000 6756
rect 2034 6722 2069 6756
rect 2103 6722 2138 6756
rect 2172 6722 2207 6756
rect 2241 6722 2276 6756
rect 2310 6722 2345 6756
rect 2379 6722 2414 6756
rect 2448 6722 2483 6756
rect 2517 6722 2552 6756
rect 2586 6722 2621 6756
rect 2655 6722 2690 6756
rect 2724 6722 2759 6756
rect 2793 6722 2828 6756
rect 2862 6722 2897 6756
rect 2931 6722 2966 6756
rect 3000 6722 3035 6756
rect 3069 6722 3104 6756
rect 3138 6722 3173 6756
rect 3207 6722 3242 6756
rect 3276 6722 3310 6756
rect 3344 6722 3378 6756
rect 3412 6722 3446 6756
rect 3480 6722 3514 6756
rect 3548 6722 3582 6756
rect 3616 6722 3650 6756
rect 3684 6722 3718 6756
rect 3752 6722 3786 6756
rect 3820 6722 3854 6756
rect 3888 6722 3922 6756
rect 3956 6722 3990 6756
rect 4024 6722 4058 6756
rect 4092 6722 4126 6756
rect 4160 6722 4194 6756
rect 4228 6722 4262 6756
rect 4296 6722 4330 6756
rect 4364 6722 4398 6756
rect 4432 6722 4466 6756
rect 4500 6722 4534 6756
rect 4568 6722 4602 6756
rect 4636 6722 4670 6756
rect 4704 6722 4738 6756
rect 4772 6722 4806 6756
rect 4840 6722 4874 6756
rect 4908 6722 4942 6756
rect 4976 6722 5010 6756
rect 5044 6722 5078 6756
rect 5112 6722 5146 6756
rect 5180 6722 5214 6756
rect 5248 6722 5282 6756
rect 5316 6722 5350 6756
rect 5384 6722 5418 6756
rect 5452 6722 5486 6756
rect 5520 6722 5554 6756
rect 5588 6722 5622 6756
rect 5656 6722 5690 6756
rect 5724 6722 5758 6756
rect 5792 6722 5826 6756
rect 5860 6722 5894 6756
rect 5928 6722 5962 6756
rect 5996 6722 6030 6756
rect 6064 6722 6098 6756
rect 6132 6722 6166 6756
rect 6200 6722 6234 6756
rect 6268 6722 6302 6756
rect 6336 6722 6370 6756
rect 6404 6722 6438 6756
rect 6472 6722 6506 6756
rect 6540 6722 6574 6756
rect 6608 6722 6642 6756
rect 6676 6722 6710 6756
rect 6744 6722 6778 6756
rect 6812 6722 6846 6756
rect 6880 6722 6914 6756
rect 6948 6722 6982 6756
rect 7016 6722 7050 6756
rect 7084 6722 7108 6756
rect 7183 6739 8488 6957
rect 12493 6809 12517 6843
rect 12551 6809 12586 6843
rect 12620 6809 12655 6843
rect 12689 6809 12724 6843
rect 12758 6809 12793 6843
rect 12827 6809 12862 6843
rect 12896 6809 12931 6843
rect 12965 6809 13000 6843
rect 13034 6809 13069 6843
rect 13103 6809 13138 6843
rect 13172 6809 13207 6843
rect 13241 6809 13276 6843
rect 13310 6809 13345 6843
rect 13379 6809 13414 6843
rect 13448 6809 13483 6843
rect 13517 6809 13552 6843
rect 13586 6809 13621 6843
rect 13655 6809 13690 6843
rect 13724 6809 13759 6843
rect 13793 6809 13828 6843
rect 13862 6809 13897 6843
rect 13931 6809 13966 6843
rect 14000 6809 14035 6843
rect 14069 6809 14104 6843
rect 14138 6809 14173 6843
rect 14207 6809 14242 6843
rect 14276 6809 14311 6843
rect 14345 6809 14380 6843
rect 14414 6809 14449 6843
rect 14483 6809 14518 6843
rect 14552 6809 14587 6843
rect 14621 6809 14655 6843
rect 14689 6809 14723 6843
rect 14757 6809 14791 6843
rect 14825 6809 14859 6843
rect 14893 6825 15117 6843
rect 14893 6809 15068 6825
rect 12493 6805 15068 6809
rect 12493 6771 14932 6805
rect 14966 6771 15000 6805
rect 15034 6771 15068 6805
rect 15102 6771 15117 6825
rect 12493 6756 15117 6771
rect 44 6669 7108 6722
rect 44 6635 68 6669
rect 102 6635 137 6669
rect 171 6635 206 6669
rect 240 6635 275 6669
rect 309 6635 344 6669
rect 378 6635 413 6669
rect 447 6635 482 6669
rect 516 6635 551 6669
rect 585 6635 620 6669
rect 654 6635 689 6669
rect 723 6635 758 6669
rect 792 6635 827 6669
rect 861 6635 896 6669
rect 930 6635 965 6669
rect 999 6635 1034 6669
rect 1068 6635 1103 6669
rect 1137 6635 1172 6669
rect 1206 6635 1241 6669
rect 1275 6635 1310 6669
rect 1344 6635 1379 6669
rect 1413 6635 1448 6669
rect 1482 6635 1517 6669
rect 1551 6635 1586 6669
rect 1620 6635 1655 6669
rect 1689 6635 1724 6669
rect 1758 6635 1793 6669
rect 1827 6635 1862 6669
rect 1896 6635 1931 6669
rect 1965 6635 2000 6669
rect 2034 6635 2069 6669
rect 2103 6635 2138 6669
rect 2172 6635 2207 6669
rect 2241 6635 2276 6669
rect 2310 6635 2345 6669
rect 2379 6635 2414 6669
rect 2448 6635 2483 6669
rect 2517 6635 2552 6669
rect 2586 6635 2621 6669
rect 2655 6635 2690 6669
rect 2724 6635 2759 6669
rect 2793 6635 2828 6669
rect 2862 6635 2897 6669
rect 2931 6635 2966 6669
rect 3000 6635 3035 6669
rect 3069 6635 3104 6669
rect 3138 6635 3173 6669
rect 3207 6635 3242 6669
rect 3276 6635 3310 6669
rect 3344 6635 3378 6669
rect 3412 6635 3446 6669
rect 3480 6635 3514 6669
rect 3548 6635 3582 6669
rect 3616 6635 3650 6669
rect 3684 6635 3718 6669
rect 3752 6635 3786 6669
rect 3820 6635 3854 6669
rect 3888 6635 3922 6669
rect 3956 6635 3990 6669
rect 4024 6635 4058 6669
rect 4092 6635 4126 6669
rect 4160 6635 4194 6669
rect 4228 6635 4262 6669
rect 4296 6635 4330 6669
rect 4364 6635 4398 6669
rect 4432 6635 4466 6669
rect 4500 6635 4534 6669
rect 4568 6635 4602 6669
rect 4636 6635 4670 6669
rect 4704 6635 4738 6669
rect 4772 6635 4806 6669
rect 4840 6635 4874 6669
rect 4908 6635 4942 6669
rect 4976 6635 5010 6669
rect 5044 6635 5078 6669
rect 5112 6635 5146 6669
rect 5180 6635 5214 6669
rect 5248 6635 5282 6669
rect 5316 6635 5350 6669
rect 5384 6635 5418 6669
rect 5452 6635 5486 6669
rect 5520 6635 5554 6669
rect 5588 6635 5622 6669
rect 5656 6635 5690 6669
rect 5724 6635 5758 6669
rect 5792 6635 5826 6669
rect 5860 6635 5894 6669
rect 5928 6635 5962 6669
rect 5996 6635 6030 6669
rect 6064 6635 6098 6669
rect 6132 6635 6166 6669
rect 6200 6635 6234 6669
rect 6268 6635 6302 6669
rect 6336 6635 6370 6669
rect 6404 6635 6438 6669
rect 6472 6635 6506 6669
rect 6540 6635 6574 6669
rect 6608 6635 6642 6669
rect 6676 6635 6710 6669
rect 6744 6635 6778 6669
rect 6812 6635 6846 6669
rect 6880 6635 6914 6669
rect 6948 6635 6982 6669
rect 7016 6635 7050 6669
rect 7084 6635 7108 6669
rect 12493 6722 12517 6756
rect 12551 6722 12586 6756
rect 12620 6722 12655 6756
rect 12689 6722 12724 6756
rect 12758 6722 12793 6756
rect 12827 6722 12862 6756
rect 12896 6722 12931 6756
rect 12965 6722 13000 6756
rect 13034 6722 13069 6756
rect 13103 6722 13138 6756
rect 13172 6722 13207 6756
rect 13241 6722 13276 6756
rect 13310 6722 13345 6756
rect 13379 6722 13414 6756
rect 13448 6722 13483 6756
rect 13517 6722 13552 6756
rect 13586 6722 13621 6756
rect 13655 6722 13690 6756
rect 13724 6722 13759 6756
rect 13793 6722 13828 6756
rect 13862 6722 13897 6756
rect 13931 6722 13966 6756
rect 14000 6722 14035 6756
rect 14069 6722 14104 6756
rect 14138 6722 14173 6756
rect 14207 6722 14242 6756
rect 14276 6722 14311 6756
rect 14345 6722 14380 6756
rect 14414 6722 14449 6756
rect 14483 6722 14518 6756
rect 14552 6722 14587 6756
rect 14621 6722 14655 6756
rect 14689 6722 14723 6756
rect 14757 6722 14791 6756
rect 14825 6722 14859 6756
rect 14893 6753 15117 6756
rect 14893 6731 15068 6753
rect 14893 6722 14932 6731
rect 12493 6697 14932 6722
rect 14966 6697 15000 6731
rect 15034 6697 15068 6731
rect 15102 6697 15117 6753
rect 12493 6681 15117 6697
rect 12493 6669 15068 6681
rect 12493 6635 12517 6669
rect 12551 6635 12586 6669
rect 12620 6635 12655 6669
rect 12689 6635 12724 6669
rect 12758 6635 12793 6669
rect 12827 6635 12862 6669
rect 12896 6635 12931 6669
rect 12965 6635 13000 6669
rect 13034 6635 13069 6669
rect 13103 6635 13138 6669
rect 13172 6635 13207 6669
rect 13241 6635 13276 6669
rect 13310 6635 13345 6669
rect 13379 6635 13414 6669
rect 13448 6635 13483 6669
rect 13517 6635 13552 6669
rect 13586 6635 13621 6669
rect 13655 6635 13690 6669
rect 13724 6635 13759 6669
rect 13793 6635 13828 6669
rect 13862 6635 13897 6669
rect 13931 6635 13966 6669
rect 14000 6635 14035 6669
rect 14069 6635 14104 6669
rect 14138 6635 14173 6669
rect 14207 6635 14242 6669
rect 14276 6635 14311 6669
rect 14345 6635 14380 6669
rect 14414 6635 14449 6669
rect 14483 6635 14518 6669
rect 14552 6635 14587 6669
rect 14621 6635 14655 6669
rect 14689 6635 14723 6669
rect 14757 6635 14791 6669
rect 14825 6635 14859 6669
rect 14893 6657 15068 6669
rect 14893 6635 14932 6657
rect 44 6623 14932 6635
rect 14966 6623 15000 6657
rect 15034 6623 15068 6657
rect 15102 6623 15117 6681
rect 44 6609 15117 6623
rect 44 6583 15068 6609
rect 44 6582 14932 6583
rect 44 6548 68 6582
rect 102 6548 137 6582
rect 171 6548 206 6582
rect 240 6548 275 6582
rect 309 6548 344 6582
rect 378 6548 413 6582
rect 447 6548 482 6582
rect 516 6548 551 6582
rect 585 6548 620 6582
rect 654 6548 689 6582
rect 723 6548 758 6582
rect 792 6548 827 6582
rect 861 6548 896 6582
rect 930 6548 965 6582
rect 999 6548 1034 6582
rect 1068 6548 1103 6582
rect 1137 6548 1172 6582
rect 1206 6548 1241 6582
rect 1275 6548 1310 6582
rect 1344 6548 1379 6582
rect 1413 6548 1448 6582
rect 1482 6548 1517 6582
rect 1551 6548 1586 6582
rect 1620 6548 1655 6582
rect 1689 6548 1724 6582
rect 1758 6548 1793 6582
rect 1827 6548 1862 6582
rect 1896 6548 1931 6582
rect 1965 6548 2000 6582
rect 2034 6548 2069 6582
rect 2103 6548 2138 6582
rect 2172 6548 2207 6582
rect 2241 6548 2276 6582
rect 2310 6548 2345 6582
rect 2379 6548 2414 6582
rect 2448 6548 2483 6582
rect 2517 6548 2551 6582
rect 2585 6548 2619 6582
rect 2653 6548 2687 6582
rect 2721 6548 2755 6582
rect 2789 6548 2823 6582
rect 2857 6548 2891 6582
rect 2925 6548 2959 6582
rect 2993 6548 3027 6582
rect 3061 6548 3095 6582
rect 3129 6548 3163 6582
rect 3197 6548 3231 6582
rect 3265 6548 3299 6582
rect 3333 6548 3367 6582
rect 3401 6548 3435 6582
rect 3469 6548 3503 6582
rect 3537 6548 3571 6582
rect 3605 6548 3639 6582
rect 3673 6548 3707 6582
rect 3741 6548 3775 6582
rect 3809 6548 3843 6582
rect 3877 6548 3911 6582
rect 3945 6548 3979 6582
rect 4013 6548 4047 6582
rect 4081 6548 4115 6582
rect 4149 6548 4183 6582
rect 4217 6548 4251 6582
rect 4285 6548 4319 6582
rect 4353 6548 4387 6582
rect 4421 6548 4455 6582
rect 4489 6548 4523 6582
rect 4557 6548 4591 6582
rect 4625 6548 4659 6582
rect 4693 6548 4727 6582
rect 4761 6548 4795 6582
rect 4829 6548 4863 6582
rect 4897 6548 4931 6582
rect 4965 6548 4999 6582
rect 5033 6548 5067 6582
rect 5101 6548 5135 6582
rect 5169 6548 5203 6582
rect 5237 6548 5271 6582
rect 5305 6548 5339 6582
rect 5373 6548 5407 6582
rect 5441 6548 5475 6582
rect 5509 6548 5543 6582
rect 5577 6548 5611 6582
rect 5645 6548 5679 6582
rect 5713 6548 5747 6582
rect 5781 6548 5815 6582
rect 5849 6548 5883 6582
rect 5917 6548 5951 6582
rect 5985 6548 6019 6582
rect 6053 6548 6087 6582
rect 6121 6548 6155 6582
rect 6189 6548 6223 6582
rect 6257 6548 6291 6582
rect 6325 6548 6359 6582
rect 6393 6548 6427 6582
rect 6461 6548 6495 6582
rect 6529 6548 6563 6582
rect 6597 6548 6631 6582
rect 6665 6548 6699 6582
rect 6733 6548 6767 6582
rect 6801 6548 6835 6582
rect 6869 6548 6903 6582
rect 6937 6548 6971 6582
rect 7005 6548 7039 6582
rect 7073 6548 7107 6582
rect 7141 6548 7175 6582
rect 7209 6548 7243 6582
rect 7277 6548 7311 6582
rect 7345 6548 7379 6582
rect 7413 6548 7447 6582
rect 7481 6548 7515 6582
rect 7549 6548 7583 6582
rect 7617 6548 7651 6582
rect 7685 6548 7719 6582
rect 7753 6548 7787 6582
rect 7821 6548 7855 6582
rect 7889 6548 7923 6582
rect 7957 6548 7991 6582
rect 8025 6548 8059 6582
rect 8093 6548 8127 6582
rect 8161 6548 8195 6582
rect 8229 6548 8263 6582
rect 8297 6548 8331 6582
rect 8365 6548 8399 6582
rect 8433 6548 8467 6582
rect 8501 6548 8535 6582
rect 8569 6548 8603 6582
rect 8637 6548 8671 6582
rect 8705 6548 8739 6582
rect 8773 6548 8807 6582
rect 8841 6548 8875 6582
rect 8909 6548 8943 6582
rect 8977 6548 9011 6582
rect 9045 6548 9079 6582
rect 9113 6548 9147 6582
rect 9181 6548 9215 6582
rect 9249 6548 9283 6582
rect 9317 6548 9351 6582
rect 9385 6548 9419 6582
rect 9453 6548 9487 6582
rect 9521 6548 9555 6582
rect 9589 6548 9623 6582
rect 9657 6548 9691 6582
rect 9725 6548 9759 6582
rect 9793 6548 9827 6582
rect 9861 6548 9895 6582
rect 9929 6548 9963 6582
rect 9997 6548 10031 6582
rect 10065 6548 10099 6582
rect 10133 6548 10167 6582
rect 10201 6548 10235 6582
rect 10269 6548 10303 6582
rect 10337 6548 10371 6582
rect 10405 6548 10439 6582
rect 10473 6548 10507 6582
rect 10541 6548 10575 6582
rect 10609 6548 10643 6582
rect 10677 6548 10711 6582
rect 10745 6548 10779 6582
rect 10813 6548 10847 6582
rect 10881 6548 10915 6582
rect 10949 6548 10983 6582
rect 11017 6548 11051 6582
rect 11085 6548 11119 6582
rect 11153 6548 11187 6582
rect 11221 6548 11255 6582
rect 11289 6548 11323 6582
rect 11357 6548 11391 6582
rect 11425 6548 11459 6582
rect 11493 6548 11527 6582
rect 11561 6548 11595 6582
rect 11629 6548 11663 6582
rect 11697 6548 11731 6582
rect 11765 6548 11799 6582
rect 11833 6548 11867 6582
rect 11901 6548 11935 6582
rect 11969 6548 12003 6582
rect 12037 6548 12071 6582
rect 12105 6548 12139 6582
rect 12173 6548 12207 6582
rect 12241 6548 12275 6582
rect 12309 6548 12343 6582
rect 12377 6548 12411 6582
rect 12445 6548 12479 6582
rect 12513 6548 12547 6582
rect 12581 6548 12615 6582
rect 12649 6548 12683 6582
rect 12717 6548 12751 6582
rect 12785 6548 12819 6582
rect 12853 6548 12887 6582
rect 12921 6548 12955 6582
rect 12989 6548 13023 6582
rect 13057 6548 13091 6582
rect 13125 6548 13159 6582
rect 13193 6548 13227 6582
rect 13261 6548 13295 6582
rect 13329 6548 13363 6582
rect 13397 6548 13431 6582
rect 13465 6548 13499 6582
rect 13533 6548 13567 6582
rect 13601 6548 13635 6582
rect 13669 6548 13703 6582
rect 13737 6548 13771 6582
rect 13805 6548 13839 6582
rect 13873 6548 13907 6582
rect 13941 6548 13975 6582
rect 14009 6548 14043 6582
rect 14077 6548 14111 6582
rect 14145 6548 14179 6582
rect 14213 6548 14247 6582
rect 14281 6548 14315 6582
rect 14349 6548 14383 6582
rect 14417 6548 14451 6582
rect 14485 6548 14519 6582
rect 14553 6548 14587 6582
rect 14621 6548 14655 6582
rect 14689 6548 14723 6582
rect 14757 6548 14791 6582
rect 14825 6548 14859 6582
rect 14893 6549 14932 6582
rect 14966 6549 15000 6583
rect 15034 6549 15068 6583
rect 15102 6549 15117 6609
rect 14893 6548 15117 6549
rect 44 6537 15117 6548
rect 44 6509 15068 6537
rect 44 6508 14932 6509
rect 44 6474 68 6508
rect 102 6474 137 6508
rect 171 6474 206 6508
rect 240 6474 275 6508
rect 309 6474 344 6508
rect 378 6474 413 6508
rect 447 6474 482 6508
rect 516 6474 551 6508
rect 585 6474 620 6508
rect 654 6474 689 6508
rect 723 6474 758 6508
rect 792 6474 827 6508
rect 861 6474 896 6508
rect 930 6474 965 6508
rect 999 6474 1034 6508
rect 1068 6474 1103 6508
rect 1137 6474 1172 6508
rect 1206 6474 1241 6508
rect 1275 6474 1310 6508
rect 1344 6474 1379 6508
rect 1413 6474 1448 6508
rect 1482 6474 1517 6508
rect 1551 6474 1586 6508
rect 1620 6474 1655 6508
rect 1689 6474 1724 6508
rect 1758 6474 1793 6508
rect 1827 6474 1862 6508
rect 1896 6474 1931 6508
rect 1965 6474 2000 6508
rect 2034 6474 2069 6508
rect 2103 6474 2138 6508
rect 2172 6474 2207 6508
rect 2241 6474 2276 6508
rect 2310 6474 2345 6508
rect 2379 6474 2414 6508
rect 2448 6474 2483 6508
rect 2517 6474 2551 6508
rect 2585 6474 2619 6508
rect 2653 6474 2687 6508
rect 2721 6474 2755 6508
rect 2789 6474 2823 6508
rect 2857 6474 2891 6508
rect 2925 6474 2959 6508
rect 2993 6474 3027 6508
rect 3061 6474 3095 6508
rect 3129 6474 3163 6508
rect 3197 6474 3231 6508
rect 3265 6474 3299 6508
rect 3333 6474 3367 6508
rect 3401 6474 3435 6508
rect 3469 6474 3503 6508
rect 3537 6474 3571 6508
rect 3605 6474 3639 6508
rect 3673 6474 3707 6508
rect 3741 6474 3775 6508
rect 3809 6474 3843 6508
rect 3877 6474 3911 6508
rect 3945 6474 3979 6508
rect 4013 6474 4047 6508
rect 4081 6474 4115 6508
rect 4149 6474 4183 6508
rect 4217 6474 4251 6508
rect 4285 6474 4319 6508
rect 4353 6474 4387 6508
rect 4421 6474 4455 6508
rect 4489 6474 4523 6508
rect 4557 6474 4591 6508
rect 4625 6474 4659 6508
rect 4693 6474 4727 6508
rect 4761 6474 4795 6508
rect 4829 6474 4863 6508
rect 4897 6474 4931 6508
rect 4965 6474 4999 6508
rect 5033 6474 5067 6508
rect 5101 6474 5135 6508
rect 5169 6474 5203 6508
rect 5237 6474 5271 6508
rect 5305 6474 5339 6508
rect 5373 6474 5407 6508
rect 5441 6474 5475 6508
rect 5509 6474 5543 6508
rect 5577 6474 5611 6508
rect 5645 6474 5679 6508
rect 5713 6474 5747 6508
rect 5781 6474 5815 6508
rect 5849 6474 5883 6508
rect 5917 6474 5951 6508
rect 5985 6474 6019 6508
rect 6053 6474 6087 6508
rect 6121 6474 6155 6508
rect 6189 6474 6223 6508
rect 6257 6474 6291 6508
rect 6325 6474 6359 6508
rect 6393 6474 6427 6508
rect 6461 6474 6495 6508
rect 6529 6474 6563 6508
rect 6597 6474 6631 6508
rect 6665 6474 6699 6508
rect 6733 6474 6767 6508
rect 6801 6474 6835 6508
rect 6869 6474 6903 6508
rect 6937 6474 6971 6508
rect 7005 6474 7039 6508
rect 7073 6474 7107 6508
rect 7141 6474 7175 6508
rect 7209 6474 7243 6508
rect 7277 6474 7311 6508
rect 7345 6474 7379 6508
rect 7413 6474 7447 6508
rect 7481 6474 7515 6508
rect 7549 6474 7583 6508
rect 7617 6474 7651 6508
rect 7685 6474 7719 6508
rect 7753 6474 7787 6508
rect 7821 6474 7855 6508
rect 7889 6474 7923 6508
rect 7957 6474 7991 6508
rect 8025 6474 8059 6508
rect 8093 6474 8127 6508
rect 8161 6474 8195 6508
rect 8229 6474 8263 6508
rect 8297 6474 8331 6508
rect 8365 6474 8399 6508
rect 8433 6474 8467 6508
rect 8501 6474 8535 6508
rect 8569 6474 8603 6508
rect 8637 6474 8671 6508
rect 8705 6474 8739 6508
rect 8773 6474 8807 6508
rect 8841 6474 8875 6508
rect 8909 6474 8943 6508
rect 8977 6474 9011 6508
rect 9045 6474 9079 6508
rect 9113 6474 9147 6508
rect 9181 6474 9215 6508
rect 9249 6474 9283 6508
rect 9317 6474 9351 6508
rect 9385 6474 9419 6508
rect 9453 6474 9487 6508
rect 9521 6474 9555 6508
rect 9589 6474 9623 6508
rect 9657 6474 9691 6508
rect 9725 6474 9759 6508
rect 9793 6474 9827 6508
rect 9861 6474 9895 6508
rect 9929 6474 9963 6508
rect 9997 6474 10031 6508
rect 10065 6474 10099 6508
rect 10133 6474 10167 6508
rect 10201 6474 10235 6508
rect 10269 6474 10303 6508
rect 10337 6474 10371 6508
rect 10405 6474 10439 6508
rect 10473 6474 10507 6508
rect 10541 6474 10575 6508
rect 10609 6474 10643 6508
rect 10677 6474 10711 6508
rect 10745 6474 10779 6508
rect 10813 6474 10847 6508
rect 10881 6474 10915 6508
rect 10949 6474 10983 6508
rect 11017 6474 11051 6508
rect 11085 6474 11119 6508
rect 11153 6474 11187 6508
rect 11221 6474 11255 6508
rect 11289 6474 11323 6508
rect 11357 6474 11391 6508
rect 11425 6474 11459 6508
rect 11493 6474 11527 6508
rect 11561 6474 11595 6508
rect 11629 6474 11663 6508
rect 11697 6474 11731 6508
rect 11765 6474 11799 6508
rect 11833 6474 11867 6508
rect 11901 6474 11935 6508
rect 11969 6474 12003 6508
rect 12037 6474 12071 6508
rect 12105 6474 12139 6508
rect 12173 6474 12207 6508
rect 12241 6474 12275 6508
rect 12309 6474 12343 6508
rect 12377 6474 12411 6508
rect 12445 6474 12479 6508
rect 12513 6474 12547 6508
rect 12581 6474 12615 6508
rect 12649 6474 12683 6508
rect 12717 6474 12751 6508
rect 12785 6474 12819 6508
rect 12853 6474 12887 6508
rect 12921 6474 12955 6508
rect 12989 6474 13023 6508
rect 13057 6474 13091 6508
rect 13125 6474 13159 6508
rect 13193 6474 13227 6508
rect 13261 6474 13295 6508
rect 13329 6474 13363 6508
rect 13397 6474 13431 6508
rect 13465 6474 13499 6508
rect 13533 6474 13567 6508
rect 13601 6474 13635 6508
rect 13669 6474 13703 6508
rect 13737 6474 13771 6508
rect 13805 6474 13839 6508
rect 13873 6474 13907 6508
rect 13941 6474 13975 6508
rect 14009 6474 14043 6508
rect 14077 6474 14111 6508
rect 14145 6474 14179 6508
rect 14213 6474 14247 6508
rect 14281 6474 14315 6508
rect 14349 6474 14383 6508
rect 14417 6474 14451 6508
rect 14485 6474 14519 6508
rect 14553 6474 14587 6508
rect 14621 6474 14655 6508
rect 14689 6474 14723 6508
rect 14757 6474 14791 6508
rect 14825 6474 14859 6508
rect 14893 6475 14932 6508
rect 14966 6475 15000 6509
rect 15034 6475 15068 6509
rect 15102 6475 15117 6537
rect 14893 6474 15117 6475
rect 44 6465 15117 6474
rect 44 6439 15068 6465
rect 44 6400 68 6439
rect 102 6434 141 6439
rect 175 6434 214 6439
rect 248 6434 287 6439
rect 321 6434 360 6439
rect 394 6434 433 6439
rect 467 6434 506 6439
rect 540 6434 579 6439
rect 613 6434 652 6439
rect 686 6434 725 6439
rect 759 6434 798 6439
rect 832 6434 871 6439
rect 905 6434 944 6439
rect 978 6434 1017 6439
rect 1051 6434 1090 6439
rect 15020 6435 15068 6439
rect 102 6400 137 6434
rect 175 6405 206 6434
rect 248 6405 275 6434
rect 321 6405 344 6434
rect 394 6405 413 6434
rect 467 6405 482 6434
rect 540 6405 551 6434
rect 613 6405 620 6434
rect 686 6405 689 6434
rect 171 6400 206 6405
rect 240 6400 275 6405
rect 309 6400 344 6405
rect 378 6400 413 6405
rect 447 6400 482 6405
rect 516 6400 551 6405
rect 585 6400 620 6405
rect 654 6400 689 6405
rect 723 6405 725 6434
rect 792 6405 798 6434
rect 861 6405 871 6434
rect 930 6405 944 6434
rect 999 6405 1017 6434
rect 723 6400 758 6405
rect 792 6400 827 6405
rect 861 6400 896 6405
rect 930 6400 965 6405
rect 999 6400 1034 6405
rect 1068 6400 1090 6434
rect 15034 6401 15068 6435
rect 15102 6401 15117 6465
rect 44 6367 1090 6400
rect 44 6326 68 6367
rect 102 6360 141 6367
rect 175 6360 214 6367
rect 248 6360 287 6367
rect 321 6360 360 6367
rect 394 6360 433 6367
rect 467 6360 506 6367
rect 540 6360 579 6367
rect 613 6360 652 6367
rect 686 6360 725 6367
rect 759 6360 798 6367
rect 832 6360 871 6367
rect 905 6360 944 6367
rect 978 6360 1017 6367
rect 1051 6360 1090 6367
rect 15020 6393 15117 6401
rect 15020 6360 15068 6393
rect 102 6326 137 6360
rect 175 6333 206 6360
rect 248 6333 275 6360
rect 321 6333 344 6360
rect 394 6333 413 6360
rect 467 6333 482 6360
rect 540 6333 551 6360
rect 613 6333 620 6360
rect 686 6333 689 6360
rect 171 6326 206 6333
rect 240 6326 275 6333
rect 309 6326 344 6333
rect 378 6326 413 6333
rect 447 6326 482 6333
rect 516 6326 551 6333
rect 585 6326 620 6333
rect 654 6326 689 6333
rect 723 6333 725 6360
rect 792 6333 798 6360
rect 861 6333 871 6360
rect 930 6333 944 6360
rect 999 6333 1017 6360
rect 723 6326 758 6333
rect 792 6326 827 6333
rect 861 6326 896 6333
rect 930 6326 965 6333
rect 999 6326 1034 6333
rect 1068 6326 1090 6360
rect 15034 6326 15068 6360
rect 15102 6326 15117 6393
rect 44 6295 1090 6326
rect 44 6252 68 6295
rect 102 6286 141 6295
rect 175 6286 214 6295
rect 248 6286 287 6295
rect 321 6286 360 6295
rect 394 6286 433 6295
rect 467 6286 506 6295
rect 540 6286 579 6295
rect 613 6286 652 6295
rect 686 6286 725 6295
rect 759 6286 798 6295
rect 832 6286 871 6295
rect 905 6286 944 6295
rect 978 6286 1017 6295
rect 1051 6286 1090 6295
rect 15020 6321 15117 6326
rect 15020 6287 15068 6321
rect 15102 6287 15117 6321
rect 102 6252 137 6286
rect 175 6261 206 6286
rect 248 6261 275 6286
rect 321 6261 344 6286
rect 394 6261 413 6286
rect 467 6261 482 6286
rect 540 6261 551 6286
rect 613 6261 620 6286
rect 686 6261 689 6286
rect 171 6252 206 6261
rect 240 6252 275 6261
rect 309 6252 344 6261
rect 378 6252 413 6261
rect 447 6252 482 6261
rect 516 6252 551 6261
rect 585 6252 620 6261
rect 654 6252 689 6261
rect 723 6261 725 6286
rect 792 6261 798 6286
rect 861 6261 871 6286
rect 930 6261 944 6286
rect 999 6261 1017 6286
rect 723 6252 758 6261
rect 792 6252 827 6261
rect 861 6252 896 6261
rect 930 6252 965 6261
rect 999 6252 1034 6261
rect 1068 6252 1090 6286
rect 15020 6285 15117 6287
rect 44 6223 1090 6252
rect 15034 6251 15068 6285
rect 15102 6251 15117 6285
rect 44 6178 68 6223
rect 102 6212 141 6223
rect 175 6212 214 6223
rect 248 6212 287 6223
rect 321 6212 360 6223
rect 394 6212 433 6223
rect 467 6212 506 6223
rect 540 6212 579 6223
rect 613 6212 652 6223
rect 686 6212 725 6223
rect 759 6212 798 6223
rect 832 6212 871 6223
rect 905 6212 944 6223
rect 978 6212 1017 6223
rect 1051 6212 1090 6223
rect 15020 6249 15117 6251
rect 15020 6215 15068 6249
rect 15102 6215 15117 6249
rect 102 6178 137 6212
rect 175 6189 206 6212
rect 248 6189 275 6212
rect 321 6189 344 6212
rect 394 6189 413 6212
rect 467 6189 482 6212
rect 540 6189 551 6212
rect 613 6189 620 6212
rect 686 6189 689 6212
rect 171 6178 206 6189
rect 240 6178 275 6189
rect 309 6178 344 6189
rect 378 6178 413 6189
rect 447 6178 482 6189
rect 516 6178 551 6189
rect 585 6178 620 6189
rect 654 6178 689 6189
rect 723 6189 725 6212
rect 792 6189 798 6212
rect 861 6189 871 6212
rect 930 6189 944 6212
rect 999 6189 1017 6212
rect 723 6178 758 6189
rect 792 6178 827 6189
rect 861 6178 896 6189
rect 930 6178 965 6189
rect 999 6178 1034 6189
rect 1068 6178 1090 6212
rect 15020 6210 15117 6215
rect 44 6151 1090 6178
rect 15034 6176 15068 6210
rect 44 6104 68 6151
rect 102 6138 141 6151
rect 175 6138 214 6151
rect 248 6138 287 6151
rect 321 6138 360 6151
rect 394 6138 433 6151
rect 467 6138 506 6151
rect 540 6138 579 6151
rect 613 6138 652 6151
rect 686 6138 725 6151
rect 759 6138 798 6151
rect 832 6138 871 6151
rect 905 6138 944 6151
rect 978 6138 1017 6151
rect 1051 6138 1090 6151
rect 15020 6143 15068 6176
rect 15102 6143 15117 6210
rect 102 6104 137 6138
rect 175 6117 206 6138
rect 248 6117 275 6138
rect 321 6117 344 6138
rect 394 6117 413 6138
rect 467 6117 482 6138
rect 540 6117 551 6138
rect 613 6117 620 6138
rect 686 6117 689 6138
rect 171 6104 206 6117
rect 240 6104 275 6117
rect 309 6104 344 6117
rect 378 6104 413 6117
rect 447 6104 482 6117
rect 516 6104 551 6117
rect 585 6104 620 6117
rect 654 6104 689 6117
rect 723 6117 725 6138
rect 792 6117 798 6138
rect 861 6117 871 6138
rect 930 6117 944 6138
rect 999 6117 1017 6138
rect 1068 6117 1090 6138
rect 15020 6135 15117 6143
rect 723 6104 758 6117
rect 792 6104 827 6117
rect 861 6104 896 6117
rect 930 6104 965 6117
rect 999 6104 1034 6117
rect 1068 6104 1103 6117
rect 1137 6104 1172 6117
rect 1206 6104 1241 6117
rect 1275 6104 1310 6117
rect 1344 6104 1379 6117
rect 1413 6104 1448 6117
rect 1482 6104 1517 6117
rect 1551 6104 1586 6117
rect 1620 6104 1655 6117
rect 1689 6104 1724 6117
rect 1758 6104 1793 6117
rect 1827 6104 1862 6117
rect 1896 6104 1931 6117
rect 1965 6104 2000 6117
rect 2034 6104 2069 6117
rect 2103 6104 2138 6117
rect 2172 6104 2207 6117
rect 2241 6104 2276 6117
rect 2310 6104 2345 6117
rect 2379 6104 2414 6117
rect 2448 6104 2483 6117
rect 2517 6104 2551 6117
rect 2585 6104 2619 6117
rect 2653 6104 2687 6117
rect 2721 6104 2755 6117
rect 2789 6104 2823 6117
rect 2857 6104 2891 6117
rect 2925 6104 2959 6117
rect 2993 6104 3027 6117
rect 3061 6104 3095 6117
rect 3129 6104 3163 6117
rect 3197 6104 3231 6117
rect 3265 6104 3299 6117
rect 3333 6104 3367 6117
rect 3401 6104 3435 6117
rect 3469 6104 3503 6117
rect 3537 6104 3571 6117
rect 3605 6104 3639 6117
rect 3673 6104 3707 6117
rect 3741 6104 3775 6117
rect 3809 6104 3843 6117
rect 3877 6104 3911 6117
rect 3945 6104 3979 6117
rect 4013 6104 4047 6117
rect 4081 6104 4115 6117
rect 4149 6104 4183 6117
rect 4217 6104 4251 6117
rect 4285 6104 4319 6117
rect 4353 6104 4387 6117
rect 4421 6104 4455 6117
rect 4489 6104 4523 6117
rect 4557 6104 4591 6117
rect 4625 6104 4659 6117
rect 4693 6104 4727 6117
rect 4761 6104 4795 6117
rect 4829 6104 4863 6117
rect 4897 6104 4931 6117
rect 4965 6104 4999 6117
rect 5033 6104 5067 6117
rect 5101 6104 5135 6117
rect 5169 6104 5203 6117
rect 5237 6104 5271 6117
rect 5305 6104 5339 6117
rect 5373 6104 5407 6117
rect 5441 6104 5475 6117
rect 5509 6104 5543 6117
rect 5577 6104 5611 6117
rect 5645 6104 5679 6117
rect 5713 6104 5747 6117
rect 5781 6104 5815 6117
rect 5849 6104 5883 6117
rect 5917 6104 5951 6117
rect 5985 6104 6019 6117
rect 6053 6104 6087 6117
rect 6121 6104 6155 6117
rect 6189 6104 6223 6117
rect 6257 6104 6291 6117
rect 6325 6104 6359 6117
rect 6393 6104 6427 6117
rect 6461 6104 6495 6117
rect 6529 6104 6563 6117
rect 6597 6104 6631 6117
rect 6665 6104 6699 6117
rect 6733 6104 6767 6117
rect 6801 6104 6835 6117
rect 6869 6104 6903 6117
rect 6937 6104 6971 6117
rect 7005 6104 7039 6117
rect 7073 6104 7107 6117
rect 7141 6104 7175 6117
rect 7209 6104 7243 6117
rect 7277 6104 7311 6117
rect 7345 6104 7379 6117
rect 7413 6104 7447 6117
rect 7481 6104 7515 6117
rect 7549 6104 7583 6117
rect 7617 6104 7651 6117
rect 7685 6104 7719 6117
rect 7753 6104 7787 6117
rect 7821 6104 7855 6117
rect 7889 6104 7923 6117
rect 7957 6104 7991 6117
rect 8025 6104 8059 6117
rect 8093 6104 8127 6117
rect 8161 6104 8195 6117
rect 8229 6104 8263 6117
rect 8297 6104 8331 6117
rect 8365 6104 8399 6117
rect 8433 6104 8467 6117
rect 8501 6104 8535 6117
rect 8569 6104 8603 6117
rect 8637 6104 8671 6117
rect 8705 6104 8739 6117
rect 8773 6104 8807 6117
rect 8841 6104 8875 6117
rect 8909 6104 8943 6117
rect 8977 6104 9011 6117
rect 9045 6104 9079 6117
rect 9113 6104 9147 6117
rect 9181 6104 9215 6117
rect 9249 6104 9283 6117
rect 9317 6104 9351 6117
rect 9385 6104 9419 6117
rect 9453 6104 9487 6117
rect 9521 6104 9555 6117
rect 9589 6104 9623 6117
rect 9657 6104 9691 6117
rect 9725 6104 9759 6117
rect 9793 6104 9827 6117
rect 9861 6104 9895 6117
rect 9929 6104 9963 6117
rect 9997 6104 10031 6117
rect 10065 6104 10099 6117
rect 10133 6104 10167 6117
rect 10201 6104 10235 6117
rect 10269 6104 10303 6117
rect 10337 6104 10371 6117
rect 10405 6104 10439 6117
rect 10473 6104 10507 6117
rect 10541 6104 10575 6117
rect 10609 6104 10643 6117
rect 10677 6104 10711 6117
rect 10745 6104 10779 6117
rect 10813 6104 10847 6117
rect 10881 6104 10915 6117
rect 10949 6104 10983 6117
rect 11017 6104 11051 6117
rect 11085 6104 11119 6117
rect 11153 6104 11187 6117
rect 11221 6104 11255 6117
rect 11289 6104 11323 6117
rect 11357 6104 11391 6117
rect 11425 6104 11459 6117
rect 11493 6104 11527 6117
rect 11561 6104 11595 6117
rect 11629 6104 11663 6117
rect 11697 6104 11731 6117
rect 11765 6104 11799 6117
rect 11833 6104 11867 6117
rect 11901 6104 11935 6117
rect 11969 6104 12003 6117
rect 12037 6104 12071 6117
rect 12105 6104 12139 6117
rect 12173 6104 12207 6117
rect 12241 6104 12275 6117
rect 12309 6104 12343 6117
rect 12377 6104 12411 6117
rect 12445 6104 12479 6117
rect 12513 6104 12547 6117
rect 12581 6104 12615 6117
rect 12649 6104 12683 6117
rect 12717 6104 12751 6117
rect 12785 6104 12819 6117
rect 12853 6104 12887 6117
rect 12921 6104 12955 6117
rect 12989 6104 13023 6117
rect 13057 6104 13091 6117
rect 13125 6104 13159 6117
rect 13193 6104 13227 6117
rect 13261 6104 13295 6117
rect 13329 6104 13363 6117
rect 13397 6104 13431 6117
rect 13465 6104 13499 6117
rect 13533 6104 13567 6117
rect 13601 6104 13635 6117
rect 13669 6104 13703 6117
rect 13737 6104 13771 6117
rect 13805 6104 13839 6117
rect 13873 6104 13907 6117
rect 13941 6104 13975 6117
rect 14009 6104 14043 6117
rect 14077 6104 14111 6117
rect 14145 6104 14179 6117
rect 14213 6104 14247 6117
rect 14281 6104 14315 6117
rect 14349 6104 14383 6117
rect 14417 6104 14451 6117
rect 14485 6104 14519 6117
rect 14553 6104 14587 6117
rect 14621 6104 14655 6117
rect 14689 6104 14723 6117
rect 14757 6104 14791 6117
rect 14825 6104 14859 6117
rect 14893 6104 14932 6117
rect 44 6101 14932 6104
rect 14966 6101 15000 6117
rect 15034 6101 15068 6135
rect 44 6071 15068 6101
rect 15102 6071 15117 6135
rect 44 6060 15117 6071
rect 44 6051 14932 6060
rect 14917 6026 14932 6051
rect 14966 6026 15000 6060
rect 15034 6026 15068 6060
rect 14917 5999 15068 6026
rect 15102 5999 15117 6060
rect 14917 5988 15117 5999
rect 14977 5961 15117 5988
rect 14977 5954 15068 5961
rect 14977 4628 15000 5954
rect 15102 4628 15117 5961
rect 14977 4593 15117 4628
rect 14977 4559 15000 4593
rect 15034 4559 15068 4593
rect 15102 4559 15117 4593
rect 14977 4524 15117 4559
rect 14977 4490 15000 4524
rect 15034 4490 15068 4524
rect 14977 4487 15068 4490
rect 15102 4487 15117 4524
rect 14977 4455 15117 4487
rect 14977 4421 15000 4455
rect 15034 4421 15068 4455
rect 14977 4415 15068 4421
rect 15102 4415 15117 4455
rect 14977 4386 15117 4415
rect 14977 4352 15000 4386
rect 15034 4352 15068 4386
rect 14977 4343 15068 4352
rect 15102 4343 15117 4386
rect 14977 4317 15117 4343
rect 14977 4283 15000 4317
rect 15034 4283 15068 4317
rect 14977 4271 15068 4283
rect 15102 4271 15117 4317
rect 14977 4248 15117 4271
rect 14977 4214 15000 4248
rect 15034 4214 15068 4248
rect 14977 4199 15068 4214
rect 15102 4199 15117 4248
rect 14977 4179 15117 4199
rect 14977 4145 15000 4179
rect 15034 4145 15068 4179
rect 14977 4127 15068 4145
rect 15102 4127 15117 4179
rect 14977 4110 15117 4127
rect 14977 4076 15000 4110
rect 15034 4076 15068 4110
rect 14977 4055 15068 4076
rect 15102 4055 15117 4110
rect 14977 4041 15117 4055
rect 14977 4007 15000 4041
rect 15034 4007 15068 4041
rect 14977 3983 15068 4007
rect 15102 3983 15117 4041
rect 14977 3972 15117 3983
rect 14977 3938 15000 3972
rect 15034 3938 15068 3972
rect 14977 3911 15068 3938
rect 15102 3911 15117 3972
rect 14977 3903 15117 3911
rect 14977 3869 15000 3903
rect 15034 3869 15068 3903
rect 14977 3839 15068 3869
rect 15102 3839 15117 3903
rect 14977 3834 15117 3839
rect 14977 3800 15000 3834
rect 15034 3800 15068 3834
rect 14977 3767 15068 3800
rect 15102 3767 15117 3834
rect 14977 3765 15117 3767
rect 14977 3731 15000 3765
rect 15034 3731 15068 3765
rect 15102 3731 15117 3765
rect 14977 3729 15117 3731
rect 14977 3696 15068 3729
rect 14977 3662 15000 3696
rect 15034 3662 15068 3696
rect 15102 3662 15117 3729
rect 14977 3657 15117 3662
rect 14977 3627 15068 3657
rect 14977 3593 15000 3627
rect 15034 3593 15068 3627
rect 15102 3593 15117 3657
rect 14977 3585 15117 3593
rect 14977 3558 15068 3585
rect 14977 3524 15000 3558
rect 15034 3524 15068 3558
rect 15102 3524 15117 3585
rect 14977 3513 15117 3524
rect 14977 3489 15068 3513
rect 14977 3455 15000 3489
rect 15034 3455 15068 3489
rect 15102 3455 15117 3513
rect 14977 3441 15117 3455
rect 14977 3420 15068 3441
rect 14977 3386 15000 3420
rect 15034 3386 15068 3420
rect 15102 3386 15117 3441
rect 14977 3369 15117 3386
rect 14977 3351 15068 3369
rect 14977 3317 15000 3351
rect 15034 3317 15068 3351
rect 15102 3317 15117 3369
rect 14977 3297 15117 3317
rect 14977 3282 15068 3297
rect 14977 3248 15000 3282
rect 15034 3248 15068 3282
rect 15102 3248 15117 3297
rect 14977 3225 15117 3248
rect 14977 3213 15068 3225
rect 14977 3179 15000 3213
rect 15034 3179 15068 3213
rect 15102 3179 15117 3225
rect 14977 3153 15117 3179
rect 14977 3144 15068 3153
rect 14977 3110 15000 3144
rect 15034 3110 15068 3144
rect 15102 3110 15117 3153
rect 14977 3081 15117 3110
rect 14977 3075 15068 3081
rect 14977 3041 15000 3075
rect 15034 3041 15068 3075
rect 15102 3041 15117 3081
rect 14977 3009 15117 3041
rect 14977 3006 15068 3009
rect 14977 2972 15000 3006
rect 15034 2972 15068 3006
rect 15102 2972 15117 3009
rect 14977 2937 15117 2972
rect 14977 2903 15000 2937
rect 15034 2903 15068 2937
rect 15102 2903 15117 2937
rect 14977 2868 15117 2903
rect 14977 2834 15000 2868
rect 15034 2834 15068 2868
rect 14977 2831 15068 2834
rect 15102 2831 15117 2868
rect 14977 2799 15117 2831
rect 14977 2765 15000 2799
rect 15034 2765 15068 2799
rect 14977 2759 15068 2765
rect 15102 2759 15117 2799
rect 14977 2730 15117 2759
rect 14977 2696 15000 2730
rect 15034 2696 15068 2730
rect 14977 2687 15068 2696
rect 15102 2687 15117 2730
rect 14977 2661 15117 2687
rect 14977 2627 15000 2661
rect 15034 2627 15068 2661
rect 14977 2615 15068 2627
rect 15102 2615 15117 2661
rect 14977 2592 15117 2615
rect 14977 2558 15000 2592
rect 15034 2558 15068 2592
rect 14977 2543 15068 2558
rect 15102 2543 15117 2592
rect 14977 2523 15117 2543
rect 14977 2489 15000 2523
rect 15034 2489 15068 2523
rect 14977 2471 15068 2489
rect 15102 2471 15117 2523
rect 14977 2454 15117 2471
rect 14977 2420 15000 2454
rect 15034 2420 15068 2454
rect 14977 2399 15068 2420
rect 15102 2399 15117 2454
rect 14977 2385 15117 2399
rect 14977 2351 15000 2385
rect 15034 2351 15068 2385
rect 14977 2327 15068 2351
rect 15102 2327 15117 2385
rect 14977 2316 15117 2327
rect 14977 2282 15000 2316
rect 15034 2282 15068 2316
rect 14977 2255 15068 2282
rect 15102 2255 15117 2316
rect 14977 2247 15117 2255
rect 14977 2213 15000 2247
rect 15034 2213 15068 2247
rect 14977 2183 15068 2213
rect 15102 2183 15117 2247
rect 14977 2178 15117 2183
rect 14977 2144 15000 2178
rect 15034 2144 15068 2178
rect 14977 2111 15068 2144
rect 15102 2111 15117 2178
rect 14977 2109 15117 2111
rect 14977 2075 15000 2109
rect 15034 2075 15068 2109
rect 15102 2075 15117 2109
rect 14977 2073 15117 2075
rect 14977 2040 15068 2073
rect 14977 2006 15000 2040
rect 15034 2006 15068 2040
rect 15102 2006 15117 2073
rect 14977 2001 15117 2006
rect 14977 1971 15068 2001
rect 14977 1937 15000 1971
rect 15034 1937 15068 1971
rect 15102 1937 15117 2001
rect 14977 1929 15117 1937
rect 14977 1902 15068 1929
rect 14977 1868 15000 1902
rect 15034 1868 15068 1902
rect 15102 1868 15117 1929
rect 14977 1857 15117 1868
rect 14977 1833 15068 1857
rect 14977 1799 15000 1833
rect 15034 1799 15068 1833
rect 15102 1799 15117 1857
rect 14977 1785 15117 1799
rect 14977 1764 15068 1785
rect 14977 1730 15000 1764
rect 15034 1730 15068 1764
rect 15102 1730 15117 1785
rect 14977 1713 15117 1730
rect 14977 1695 15068 1713
rect 14977 1661 15000 1695
rect 15034 1661 15068 1695
rect 15102 1661 15117 1713
rect 14977 1641 15117 1661
rect 14977 1626 15068 1641
rect 14977 1592 15000 1626
rect 15034 1592 15068 1626
rect 15102 1592 15117 1641
rect 14977 1569 15117 1592
rect 14977 1557 15068 1569
rect 14977 1523 15000 1557
rect 15034 1523 15068 1557
rect 15102 1523 15117 1569
rect 14977 1497 15117 1523
rect 14977 1488 15068 1497
rect 14977 1454 15000 1488
rect 15034 1454 15068 1488
rect 15102 1454 15117 1497
rect 14977 1425 15117 1454
rect 14977 1419 15068 1425
rect 14977 1385 15000 1419
rect 15034 1385 15068 1419
rect 15102 1385 15117 1425
rect 310 1322 402 1368
rect 14977 1353 15117 1385
rect 14977 1350 15068 1353
rect 14977 1316 15000 1350
rect 15034 1316 15068 1350
rect 15102 1316 15117 1353
rect 7044 1282 14917 1288
rect 14977 1282 15117 1316
rect 68 1281 15117 1282
rect 68 1257 15068 1281
rect 68 1251 7068 1257
rect 7022 1223 7068 1251
rect 7102 1223 7137 1257
rect 7171 1223 7206 1257
rect 7240 1223 7275 1257
rect 7309 1223 7344 1257
rect 7378 1223 7413 1257
rect 7447 1223 7482 1257
rect 7516 1223 7551 1257
rect 7585 1223 7620 1257
rect 7654 1223 7689 1257
rect 7723 1223 7758 1257
rect 7792 1223 7827 1257
rect 7861 1223 7896 1257
rect 7930 1223 7965 1257
rect 7999 1223 8034 1257
rect 8068 1223 8103 1257
rect 8137 1223 8172 1257
rect 8206 1223 8241 1257
rect 8275 1223 8310 1257
rect 8344 1223 8379 1257
rect 8413 1223 8448 1257
rect 8482 1223 8517 1257
rect 8551 1223 8586 1257
rect 8620 1223 8655 1257
rect 8689 1223 8724 1257
rect 8758 1223 8793 1257
rect 8827 1223 8862 1257
rect 8896 1223 8931 1257
rect 8965 1223 9000 1257
rect 9034 1223 9069 1257
rect 9103 1223 9138 1257
rect 9172 1223 9207 1257
rect 9241 1223 9276 1257
rect 9310 1223 9345 1257
rect 9379 1223 9414 1257
rect 9448 1223 9483 1257
rect 9517 1223 9552 1257
rect 9586 1223 9621 1257
rect 9655 1223 9690 1257
rect 9724 1223 9759 1257
rect 7022 1217 9759 1223
rect 14893 1247 15068 1257
rect 15102 1247 15117 1281
rect 14893 1244 15117 1247
rect 14893 1217 14932 1244
rect 14966 1217 15000 1244
rect 7022 1189 7069 1217
rect 7103 1189 7142 1217
rect 7176 1189 7215 1217
rect 7249 1189 7288 1217
rect 7322 1189 7361 1217
rect 7395 1189 7434 1217
rect 7468 1189 7507 1217
rect 7541 1189 7580 1217
rect 7614 1189 7653 1217
rect 7687 1189 7726 1217
rect 7760 1189 7799 1217
rect 7833 1189 7872 1217
rect 7906 1189 7945 1217
rect 7979 1189 8018 1217
rect 8052 1189 8091 1217
rect 8125 1189 8164 1217
rect 8198 1189 8237 1217
rect 8271 1189 8310 1217
rect 8344 1189 8383 1217
rect 8417 1189 8456 1217
rect 8490 1189 8528 1217
rect 8562 1189 8600 1217
rect 8634 1189 8672 1217
rect 8706 1189 8744 1217
rect 8778 1189 8816 1217
rect 8850 1189 8888 1217
rect 8922 1189 8960 1217
rect 8994 1189 9032 1217
rect 9066 1189 9104 1217
rect 7022 1155 7068 1189
rect 7103 1183 7137 1189
rect 7176 1183 7206 1189
rect 7249 1183 7275 1189
rect 7322 1183 7344 1189
rect 7395 1183 7413 1189
rect 7468 1183 7482 1189
rect 7541 1183 7551 1189
rect 7614 1183 7620 1189
rect 7687 1183 7689 1189
rect 7102 1155 7137 1183
rect 7171 1155 7206 1183
rect 7240 1155 7275 1183
rect 7309 1155 7344 1183
rect 7378 1155 7413 1183
rect 7447 1155 7482 1183
rect 7516 1155 7551 1183
rect 7585 1155 7620 1183
rect 7654 1155 7689 1183
rect 7723 1183 7726 1189
rect 7792 1183 7799 1189
rect 7861 1183 7872 1189
rect 7930 1183 7945 1189
rect 7999 1183 8018 1189
rect 8068 1183 8091 1189
rect 8137 1183 8164 1189
rect 8206 1183 8237 1189
rect 7723 1155 7758 1183
rect 7792 1155 7827 1183
rect 7861 1155 7896 1183
rect 7930 1155 7965 1183
rect 7999 1155 8034 1183
rect 8068 1155 8103 1183
rect 8137 1155 8172 1183
rect 8206 1155 8241 1183
rect 8275 1155 8310 1189
rect 8344 1155 8379 1189
rect 8417 1183 8448 1189
rect 8490 1183 8517 1189
rect 8562 1183 8586 1189
rect 8634 1183 8655 1189
rect 8706 1183 8724 1189
rect 8778 1183 8793 1189
rect 8850 1183 8862 1189
rect 8922 1183 8931 1189
rect 8994 1183 9000 1189
rect 9066 1183 9069 1189
rect 8413 1155 8448 1183
rect 8482 1155 8517 1183
rect 8551 1155 8586 1183
rect 8620 1155 8655 1183
rect 8689 1155 8724 1183
rect 8758 1155 8793 1183
rect 8827 1155 8862 1183
rect 8896 1155 8931 1183
rect 8965 1155 9000 1183
rect 9034 1155 9069 1183
rect 9103 1183 9104 1189
rect 9138 1189 9176 1217
rect 9210 1189 9248 1217
rect 9282 1189 9320 1217
rect 9354 1189 9392 1217
rect 9426 1189 9464 1217
rect 9498 1189 9536 1217
rect 9570 1189 9608 1217
rect 9642 1189 9680 1217
rect 9714 1189 9752 1217
rect 9103 1155 9138 1183
rect 9172 1183 9176 1189
rect 9241 1183 9248 1189
rect 9310 1183 9320 1189
rect 9379 1183 9392 1189
rect 9448 1183 9464 1189
rect 9517 1183 9536 1189
rect 9586 1183 9608 1189
rect 9655 1183 9680 1189
rect 9724 1183 9752 1189
rect 14926 1210 14932 1217
rect 14998 1210 15000 1217
rect 15034 1210 15068 1244
rect 15102 1210 15117 1244
rect 14926 1183 14964 1210
rect 14998 1209 15117 1210
rect 14998 1183 15068 1209
rect 9172 1155 9207 1183
rect 9241 1155 9276 1183
rect 9310 1155 9345 1183
rect 9379 1155 9414 1183
rect 9448 1155 9483 1183
rect 9517 1155 9552 1183
rect 9586 1155 9621 1183
rect 9655 1155 9690 1183
rect 9724 1155 9759 1183
rect 7022 1139 9759 1155
rect 14893 1175 15068 1183
rect 15102 1175 15117 1209
rect 14893 1172 15117 1175
rect 14893 1139 14932 1172
rect 14966 1139 15000 1172
rect 7022 1121 7069 1139
rect 7103 1121 7142 1139
rect 7176 1121 7215 1139
rect 7249 1121 7288 1139
rect 7322 1121 7361 1139
rect 7395 1121 7434 1139
rect 7468 1121 7507 1139
rect 7541 1121 7580 1139
rect 7614 1121 7653 1139
rect 7687 1121 7726 1139
rect 7760 1121 7799 1139
rect 7833 1121 7872 1139
rect 7906 1121 7945 1139
rect 7979 1121 8018 1139
rect 8052 1121 8091 1139
rect 8125 1121 8164 1139
rect 8198 1121 8237 1139
rect 8271 1121 8310 1139
rect 8344 1121 8383 1139
rect 8417 1121 8456 1139
rect 8490 1121 8528 1139
rect 8562 1121 8600 1139
rect 8634 1121 8672 1139
rect 8706 1121 8744 1139
rect 8778 1121 8816 1139
rect 8850 1121 8888 1139
rect 8922 1121 8960 1139
rect 8994 1121 9032 1139
rect 9066 1121 9104 1139
rect 7022 1087 7068 1121
rect 7103 1105 7137 1121
rect 7176 1105 7206 1121
rect 7249 1105 7275 1121
rect 7322 1105 7344 1121
rect 7395 1105 7413 1121
rect 7468 1105 7482 1121
rect 7541 1105 7551 1121
rect 7614 1105 7620 1121
rect 7687 1105 7689 1121
rect 7102 1087 7137 1105
rect 7171 1087 7206 1105
rect 7240 1087 7275 1105
rect 7309 1087 7344 1105
rect 7378 1087 7413 1105
rect 7447 1087 7482 1105
rect 7516 1087 7551 1105
rect 7585 1087 7620 1105
rect 7654 1087 7689 1105
rect 7723 1105 7726 1121
rect 7792 1105 7799 1121
rect 7861 1105 7872 1121
rect 7930 1105 7945 1121
rect 7999 1105 8018 1121
rect 8068 1105 8091 1121
rect 8137 1105 8164 1121
rect 8206 1105 8237 1121
rect 7723 1087 7758 1105
rect 7792 1087 7827 1105
rect 7861 1087 7896 1105
rect 7930 1087 7965 1105
rect 7999 1087 8034 1105
rect 8068 1087 8103 1105
rect 8137 1087 8172 1105
rect 8206 1087 8241 1105
rect 8275 1087 8310 1121
rect 8344 1087 8379 1121
rect 8417 1105 8448 1121
rect 8490 1105 8517 1121
rect 8562 1105 8586 1121
rect 8634 1105 8655 1121
rect 8706 1105 8724 1121
rect 8778 1105 8793 1121
rect 8850 1105 8862 1121
rect 8922 1105 8931 1121
rect 8994 1105 9000 1121
rect 9066 1105 9069 1121
rect 8413 1087 8448 1105
rect 8482 1087 8517 1105
rect 8551 1087 8586 1105
rect 8620 1087 8655 1105
rect 8689 1087 8724 1105
rect 8758 1087 8793 1105
rect 8827 1087 8862 1105
rect 8896 1087 8931 1105
rect 8965 1087 9000 1105
rect 9034 1087 9069 1105
rect 9103 1105 9104 1121
rect 9138 1121 9176 1139
rect 9210 1121 9248 1139
rect 9282 1121 9320 1139
rect 9354 1121 9392 1139
rect 9426 1121 9464 1139
rect 9498 1121 9536 1139
rect 9570 1121 9608 1139
rect 9642 1121 9680 1139
rect 9714 1121 9752 1139
rect 9103 1087 9138 1105
rect 9172 1105 9176 1121
rect 9241 1105 9248 1121
rect 9310 1105 9320 1121
rect 9379 1105 9392 1121
rect 9448 1105 9464 1121
rect 9517 1105 9536 1121
rect 9586 1105 9608 1121
rect 9655 1105 9680 1121
rect 9724 1105 9752 1121
rect 14926 1138 14932 1139
rect 14998 1138 15000 1139
rect 15034 1138 15068 1172
rect 15102 1138 15117 1172
rect 14926 1105 14964 1138
rect 14998 1137 15117 1138
rect 14998 1105 15068 1137
rect 9172 1087 9207 1105
rect 9241 1087 9276 1105
rect 9310 1087 9345 1105
rect 9379 1087 9414 1105
rect 9448 1087 9483 1105
rect 9517 1087 9552 1105
rect 9586 1087 9621 1105
rect 9655 1087 9690 1105
rect 9724 1087 9759 1105
rect 7022 1061 9759 1087
rect 14893 1103 15068 1105
rect 15102 1103 15117 1137
rect 14893 1100 15117 1103
rect 14893 1066 14932 1100
rect 14966 1066 15000 1100
rect 15034 1066 15068 1100
rect 15102 1066 15117 1100
rect 14893 1065 15117 1066
rect 14893 1061 15068 1065
rect 7022 1053 7069 1061
rect 7103 1053 7142 1061
rect 7176 1053 7215 1061
rect 7249 1053 7288 1061
rect 7322 1053 7361 1061
rect 7395 1053 7434 1061
rect 7468 1053 7507 1061
rect 7541 1053 7580 1061
rect 7614 1053 7653 1061
rect 7687 1053 7726 1061
rect 7760 1053 7799 1061
rect 7833 1053 7872 1061
rect 7906 1053 7945 1061
rect 7979 1053 8018 1061
rect 8052 1053 8091 1061
rect 8125 1053 8164 1061
rect 8198 1053 8237 1061
rect 8271 1053 8310 1061
rect 8344 1053 8383 1061
rect 8417 1053 8456 1061
rect 8490 1053 8528 1061
rect 8562 1053 8600 1061
rect 8634 1053 8672 1061
rect 8706 1053 8744 1061
rect 8778 1053 8816 1061
rect 8850 1053 8888 1061
rect 8922 1053 8960 1061
rect 8994 1053 9032 1061
rect 9066 1053 9104 1061
rect 7022 1019 7068 1053
rect 7103 1027 7137 1053
rect 7176 1027 7206 1053
rect 7249 1027 7275 1053
rect 7322 1027 7344 1053
rect 7395 1027 7413 1053
rect 7468 1027 7482 1053
rect 7541 1027 7551 1053
rect 7614 1027 7620 1053
rect 7687 1027 7689 1053
rect 7102 1019 7137 1027
rect 7171 1019 7206 1027
rect 7240 1019 7275 1027
rect 7309 1019 7344 1027
rect 7378 1019 7413 1027
rect 7447 1019 7482 1027
rect 7516 1019 7551 1027
rect 7585 1019 7620 1027
rect 7654 1019 7689 1027
rect 7723 1027 7726 1053
rect 7792 1027 7799 1053
rect 7861 1027 7872 1053
rect 7930 1027 7945 1053
rect 7999 1027 8018 1053
rect 8068 1027 8091 1053
rect 8137 1027 8164 1053
rect 8206 1027 8237 1053
rect 7723 1019 7758 1027
rect 7792 1019 7827 1027
rect 7861 1019 7896 1027
rect 7930 1019 7965 1027
rect 7999 1019 8034 1027
rect 8068 1019 8103 1027
rect 8137 1019 8172 1027
rect 8206 1019 8241 1027
rect 8275 1019 8310 1053
rect 8344 1019 8379 1053
rect 8417 1027 8448 1053
rect 8490 1027 8517 1053
rect 8562 1027 8586 1053
rect 8634 1027 8655 1053
rect 8706 1027 8724 1053
rect 8778 1027 8793 1053
rect 8850 1027 8862 1053
rect 8922 1027 8931 1053
rect 8994 1027 9000 1053
rect 9066 1027 9069 1053
rect 8413 1019 8448 1027
rect 8482 1019 8517 1027
rect 8551 1019 8586 1027
rect 8620 1019 8655 1027
rect 8689 1019 8724 1027
rect 8758 1019 8793 1027
rect 8827 1019 8862 1027
rect 8896 1019 8931 1027
rect 8965 1019 9000 1027
rect 9034 1019 9069 1027
rect 9103 1027 9104 1053
rect 9138 1053 9176 1061
rect 9210 1053 9248 1061
rect 9282 1053 9320 1061
rect 9354 1053 9392 1061
rect 9426 1053 9464 1061
rect 9498 1053 9536 1061
rect 9570 1053 9608 1061
rect 9642 1053 9680 1061
rect 9714 1053 9752 1061
rect 9103 1019 9138 1027
rect 9172 1027 9176 1053
rect 9241 1027 9248 1053
rect 9310 1027 9320 1053
rect 9379 1027 9392 1053
rect 9448 1027 9464 1053
rect 9517 1027 9536 1053
rect 9586 1027 9608 1053
rect 9655 1027 9680 1053
rect 9724 1027 9752 1053
rect 14926 1028 14964 1061
rect 14998 1031 15068 1061
rect 15102 1031 15117 1065
rect 14998 1028 15117 1031
rect 14926 1027 14932 1028
rect 14998 1027 15000 1028
rect 9172 1019 9207 1027
rect 9241 1019 9276 1027
rect 9310 1019 9345 1027
rect 9379 1019 9414 1027
rect 9448 1019 9483 1027
rect 9517 1019 9552 1027
rect 9586 1019 9621 1027
rect 9655 1019 9690 1027
rect 9724 1019 9759 1027
rect 14893 1019 14932 1027
rect 7022 994 14932 1019
rect 14966 994 15000 1027
rect 15034 994 15068 1028
rect 15102 994 15117 1028
rect 7022 993 15117 994
rect 7022 989 15068 993
rect 7022 988 14576 989
rect 7022 947 7754 988
rect 7022 913 7067 947
rect 7101 918 7137 947
rect 7101 913 7104 918
rect 7171 913 7207 947
rect 7241 913 7277 947
rect 7311 913 7347 947
rect 7381 913 7417 947
rect 7451 913 7487 947
rect 7521 913 7557 947
rect 7591 913 7627 947
rect 7661 913 7696 947
rect 7730 913 7754 947
rect 7022 884 7104 913
rect 7138 884 7754 913
rect 7022 875 7754 884
rect 7022 841 7067 875
rect 7101 841 7137 875
rect 7171 841 7207 875
rect 7241 841 7277 875
rect 7311 841 7347 875
rect 7381 841 7417 875
rect 7451 841 7487 875
rect 7521 841 7557 875
rect 7591 841 7627 875
rect 7661 841 7696 875
rect 7730 841 7754 875
rect 7022 803 7754 841
rect 7022 769 7067 803
rect 7101 769 7137 803
rect 7171 769 7207 803
rect 7241 769 7277 803
rect 7311 769 7347 803
rect 7381 769 7417 803
rect 7451 769 7487 803
rect 7521 769 7557 803
rect 7591 769 7627 803
rect 7661 769 7696 803
rect 7730 769 7754 803
rect 7022 731 7754 769
rect 7022 697 7067 731
rect 7101 697 7137 731
rect 7171 697 7207 731
rect 7241 697 7277 731
rect 7311 697 7347 731
rect 7381 697 7417 731
rect 7451 697 7487 731
rect 7521 697 7557 731
rect 7591 697 7627 731
rect 7661 697 7696 731
rect 7730 697 7754 731
rect 7022 659 7754 697
rect 7022 625 7067 659
rect 7101 625 7137 659
rect 7171 625 7207 659
rect 7241 625 7277 659
rect 7311 625 7347 659
rect 7381 625 7417 659
rect 7451 625 7487 659
rect 7521 625 7557 659
rect 7591 625 7627 659
rect 7661 625 7696 659
rect 7730 625 7754 659
rect 7022 587 7754 625
rect 7022 553 7067 587
rect 7101 553 7137 587
rect 7171 553 7207 587
rect 7241 553 7277 587
rect 7311 553 7347 587
rect 7381 553 7417 587
rect 7451 553 7487 587
rect 7521 553 7557 587
rect 7591 553 7627 587
rect 7661 553 7696 587
rect 7730 553 7754 587
rect 7022 515 7754 553
rect 7022 481 7067 515
rect 7101 481 7137 515
rect 7171 481 7207 515
rect 7241 481 7277 515
rect 7311 481 7347 515
rect 7381 481 7417 515
rect 7451 481 7487 515
rect 7521 481 7557 515
rect 7591 481 7627 515
rect 7661 481 7696 515
rect 7730 481 7754 515
rect 7022 443 7754 481
rect 7022 409 7067 443
rect 7101 409 7137 443
rect 7171 409 7207 443
rect 7241 409 7277 443
rect 7311 409 7347 443
rect 7381 409 7417 443
rect 7451 409 7487 443
rect 7521 409 7557 443
rect 7591 409 7627 443
rect 7661 409 7696 443
rect 7730 409 7754 443
rect 7022 369 7754 409
rect 9687 955 14576 988
rect 14610 955 14654 989
rect 14688 955 14732 989
rect 14766 955 14810 989
rect 14844 955 14888 989
rect 14922 956 14966 989
rect 14922 955 14932 956
rect 9687 947 11680 955
rect 9687 913 9711 947
rect 9745 913 9781 947
rect 9815 923 9851 947
rect 9885 923 9921 947
rect 9955 923 9991 947
rect 10025 923 10061 947
rect 9830 913 9851 923
rect 9906 913 9921 923
rect 9982 913 9991 923
rect 10058 913 10061 923
rect 10095 923 10131 947
rect 10165 923 10201 947
rect 10235 923 10271 947
rect 10305 923 10341 947
rect 10375 923 10411 947
rect 10445 923 10481 947
rect 10095 913 10100 923
rect 10165 913 10176 923
rect 10235 913 10251 923
rect 10305 913 10326 923
rect 10375 913 10401 923
rect 10445 913 10476 923
rect 10515 913 10551 947
rect 10585 913 10621 947
rect 10655 923 10691 947
rect 10725 923 10761 947
rect 10795 923 10831 947
rect 10865 923 10901 947
rect 10935 923 10971 947
rect 11005 923 11041 947
rect 10660 913 10691 923
rect 10735 913 10761 923
rect 10810 913 10831 923
rect 10885 913 10901 923
rect 10960 913 10971 923
rect 11035 913 11041 923
rect 11075 923 11111 947
rect 11075 913 11076 923
rect 9687 889 9796 913
rect 9830 889 9872 913
rect 9906 889 9948 913
rect 9982 889 10024 913
rect 10058 889 10100 913
rect 10134 889 10176 913
rect 10210 889 10251 913
rect 10285 889 10326 913
rect 10360 889 10401 913
rect 10435 889 10476 913
rect 10510 889 10551 913
rect 10585 889 10626 913
rect 10660 889 10701 913
rect 10735 889 10776 913
rect 10810 889 10851 913
rect 10885 889 10926 913
rect 10960 889 11001 913
rect 11035 889 11076 913
rect 11110 913 11111 923
rect 11145 923 11181 947
rect 11215 923 11251 947
rect 11285 923 11321 947
rect 11145 913 11151 923
rect 11215 913 11226 923
rect 11285 913 11301 923
rect 11355 913 11391 947
rect 11425 913 11460 947
rect 11494 913 11529 947
rect 11563 913 11598 947
rect 11632 921 11680 947
rect 11714 921 11750 955
rect 11784 921 11820 955
rect 11854 921 11890 955
rect 11924 921 11960 955
rect 11994 921 12030 955
rect 12064 921 12099 955
rect 12133 921 12168 955
rect 12202 921 12237 955
rect 12271 921 12306 955
rect 12340 921 12375 955
rect 12409 921 12444 955
rect 12478 921 12513 955
rect 12547 921 12582 955
rect 12616 921 12651 955
rect 12685 921 12720 955
rect 12754 921 12789 955
rect 12823 921 12858 955
rect 12892 921 12927 955
rect 12961 921 12996 955
rect 13030 921 13065 955
rect 13099 921 13134 955
rect 13168 921 13203 955
rect 13237 921 13272 955
rect 13306 921 13341 955
rect 13375 921 13410 955
rect 13444 921 13479 955
rect 13513 921 13548 955
rect 13582 921 13617 955
rect 13651 921 13686 955
rect 13720 921 13755 955
rect 13789 921 13824 955
rect 13858 921 13893 955
rect 13927 921 13962 955
rect 13996 921 14031 955
rect 14065 921 14100 955
rect 14134 921 14169 955
rect 14203 921 14238 955
rect 14272 921 14307 955
rect 14341 921 14376 955
rect 14410 921 14445 955
rect 14479 921 14514 955
rect 14548 921 14583 955
rect 14617 921 14652 955
rect 14686 921 14721 955
rect 14755 921 14790 955
rect 14824 921 14859 955
rect 14893 922 14932 955
rect 15000 959 15068 989
rect 15102 959 15117 993
rect 15000 956 15117 959
rect 14966 922 15000 955
rect 15034 922 15068 956
rect 15102 922 15117 956
rect 14893 921 15117 922
rect 11632 916 15068 921
rect 11632 913 14576 916
rect 11110 889 11151 913
rect 11185 889 11226 913
rect 11260 889 11301 913
rect 11335 889 14576 913
rect 9687 882 14576 889
rect 14610 882 14654 916
rect 14688 882 14732 916
rect 14766 882 14810 916
rect 14844 882 14888 916
rect 14922 884 14966 916
rect 14922 882 14932 884
rect 9687 875 14932 882
rect 9687 841 9711 875
rect 9745 841 9781 875
rect 9815 841 9851 875
rect 9885 841 9921 875
rect 9955 841 9991 875
rect 10025 841 10061 875
rect 10095 841 10131 875
rect 10165 841 10201 875
rect 10235 841 10271 875
rect 10305 841 10341 875
rect 10375 841 10411 875
rect 10445 841 10481 875
rect 10515 841 10551 875
rect 10585 841 10621 875
rect 10655 841 10691 875
rect 10725 841 10761 875
rect 10795 841 10831 875
rect 10865 841 10901 875
rect 10935 841 10971 875
rect 11005 841 11041 875
rect 11075 841 11111 875
rect 11145 841 11181 875
rect 11215 841 11251 875
rect 11285 841 11321 875
rect 11355 841 11391 875
rect 11425 841 11460 875
rect 11494 841 11529 875
rect 11563 841 11598 875
rect 11632 841 11680 875
rect 11714 841 11750 875
rect 11784 841 11820 875
rect 11854 841 11890 875
rect 11924 841 11960 875
rect 11994 841 12030 875
rect 12064 841 12099 875
rect 12133 841 12168 875
rect 12202 841 12237 875
rect 12271 841 12306 875
rect 12340 841 12375 875
rect 12409 841 12444 875
rect 12478 841 12513 875
rect 12547 841 12582 875
rect 12616 841 12651 875
rect 12685 841 12720 875
rect 12754 841 12789 875
rect 12823 841 12858 875
rect 12892 841 12927 875
rect 12961 841 12996 875
rect 13030 841 13065 875
rect 13099 841 13134 875
rect 13168 841 13203 875
rect 13237 841 13272 875
rect 13306 841 13341 875
rect 13375 841 13410 875
rect 13444 841 13479 875
rect 13513 841 13548 875
rect 13582 841 13617 875
rect 13651 841 13686 875
rect 13720 841 13755 875
rect 13789 841 13824 875
rect 13858 841 13893 875
rect 13927 841 13962 875
rect 13996 841 14031 875
rect 14065 841 14100 875
rect 14134 841 14169 875
rect 14203 841 14238 875
rect 14272 841 14307 875
rect 14341 841 14376 875
rect 14410 841 14445 875
rect 14479 841 14514 875
rect 14548 843 14583 875
rect 14548 841 14576 843
rect 14617 841 14652 875
rect 14686 843 14721 875
rect 14755 843 14790 875
rect 14824 843 14859 875
rect 14893 850 14932 875
rect 15000 887 15068 916
rect 15102 887 15117 921
rect 15000 884 15117 887
rect 14966 850 15000 882
rect 15034 850 15068 884
rect 15102 850 15117 884
rect 14893 849 15117 850
rect 14893 843 15068 849
rect 14688 841 14721 843
rect 14766 841 14790 843
rect 14844 841 14859 843
rect 9687 839 14576 841
rect 9687 805 9796 839
rect 9830 805 9872 839
rect 9906 805 9948 839
rect 9982 805 10024 839
rect 10058 805 10100 839
rect 10134 805 10176 839
rect 10210 805 10251 839
rect 10285 805 10326 839
rect 10360 805 10401 839
rect 10435 805 10476 839
rect 10510 805 10551 839
rect 10585 805 10626 839
rect 10660 805 10701 839
rect 10735 805 10776 839
rect 10810 805 10851 839
rect 10885 805 10926 839
rect 10960 805 11001 839
rect 11035 805 11076 839
rect 11110 805 11151 839
rect 11185 805 11226 839
rect 11260 805 11301 839
rect 11335 809 14576 839
rect 14610 809 14654 841
rect 14688 809 14732 841
rect 14766 809 14810 841
rect 14844 809 14888 841
rect 14922 812 14966 843
rect 14922 809 14932 812
rect 11335 805 14932 809
rect 9687 803 14932 805
rect 9687 769 9711 803
rect 9745 769 9781 803
rect 9815 769 9851 803
rect 9885 769 9921 803
rect 9955 769 9991 803
rect 10025 769 10061 803
rect 10095 769 10131 803
rect 10165 769 10201 803
rect 10235 769 10271 803
rect 10305 769 10341 803
rect 10375 769 10411 803
rect 10445 769 10481 803
rect 10515 769 10551 803
rect 10585 769 10621 803
rect 10655 769 10691 803
rect 10725 769 10761 803
rect 10795 769 10831 803
rect 10865 769 10901 803
rect 10935 769 10971 803
rect 11005 769 11041 803
rect 11075 769 11111 803
rect 11145 769 11181 803
rect 11215 769 11251 803
rect 11285 769 11321 803
rect 11355 769 11391 803
rect 11425 769 11460 803
rect 11494 769 11529 803
rect 11563 769 11598 803
rect 11632 795 14932 803
rect 11632 769 11680 795
rect 9687 761 11680 769
rect 11714 761 11750 795
rect 11784 761 11820 795
rect 11854 761 11890 795
rect 11924 761 11960 795
rect 11994 761 12030 795
rect 12064 761 12099 795
rect 12133 761 12168 795
rect 12202 761 12237 795
rect 12271 761 12306 795
rect 12340 761 12375 795
rect 12409 761 12444 795
rect 12478 761 12513 795
rect 12547 761 12582 795
rect 12616 761 12651 795
rect 12685 761 12720 795
rect 12754 761 12789 795
rect 12823 761 12858 795
rect 12892 761 12927 795
rect 12961 761 12996 795
rect 13030 761 13065 795
rect 13099 761 13134 795
rect 13168 761 13203 795
rect 13237 761 13272 795
rect 13306 761 13341 795
rect 13375 761 13410 795
rect 13444 761 13479 795
rect 13513 761 13548 795
rect 13582 761 13617 795
rect 13651 761 13686 795
rect 13720 761 13755 795
rect 13789 761 13824 795
rect 13858 761 13893 795
rect 13927 761 13962 795
rect 13996 761 14031 795
rect 14065 761 14100 795
rect 14134 761 14169 795
rect 14203 761 14238 795
rect 14272 761 14307 795
rect 14341 761 14376 795
rect 14410 761 14445 795
rect 14479 761 14514 795
rect 14548 770 14583 795
rect 14548 761 14576 770
rect 14617 761 14652 795
rect 14686 770 14721 795
rect 14755 770 14790 795
rect 14824 770 14859 795
rect 14893 778 14932 795
rect 15000 815 15068 843
rect 15102 815 15117 849
rect 15000 812 15117 815
rect 14966 778 15000 809
rect 15034 778 15068 812
rect 15102 778 15117 812
rect 14893 777 15117 778
rect 14893 770 15068 777
rect 14688 761 14721 770
rect 14766 761 14790 770
rect 14844 761 14859 770
rect 9687 755 14576 761
rect 9687 731 9796 755
rect 9830 731 9872 755
rect 9906 731 9948 755
rect 9982 731 10024 755
rect 10058 731 10100 755
rect 10134 731 10176 755
rect 10210 731 10251 755
rect 10285 731 10326 755
rect 10360 731 10401 755
rect 10435 731 10476 755
rect 10510 731 10551 755
rect 10585 731 10626 755
rect 10660 731 10701 755
rect 10735 731 10776 755
rect 10810 731 10851 755
rect 10885 731 10926 755
rect 10960 731 11001 755
rect 11035 731 11076 755
rect 9687 697 9711 731
rect 9745 697 9781 731
rect 9830 721 9851 731
rect 9906 721 9921 731
rect 9982 721 9991 731
rect 10058 721 10061 731
rect 9815 697 9851 721
rect 9885 697 9921 721
rect 9955 697 9991 721
rect 10025 697 10061 721
rect 10095 721 10100 731
rect 10165 721 10176 731
rect 10235 721 10251 731
rect 10305 721 10326 731
rect 10375 721 10401 731
rect 10445 721 10476 731
rect 10095 697 10131 721
rect 10165 697 10201 721
rect 10235 697 10271 721
rect 10305 697 10341 721
rect 10375 697 10411 721
rect 10445 697 10481 721
rect 10515 697 10551 731
rect 10585 697 10621 731
rect 10660 721 10691 731
rect 10735 721 10761 731
rect 10810 721 10831 731
rect 10885 721 10901 731
rect 10960 721 10971 731
rect 11035 721 11041 731
rect 10655 697 10691 721
rect 10725 697 10761 721
rect 10795 697 10831 721
rect 10865 697 10901 721
rect 10935 697 10971 721
rect 11005 697 11041 721
rect 11075 721 11076 731
rect 11110 731 11151 755
rect 11185 731 11226 755
rect 11260 731 11301 755
rect 11335 736 14576 755
rect 14610 736 14654 761
rect 14688 736 14732 761
rect 14766 736 14810 761
rect 14844 736 14888 761
rect 14922 740 14966 770
rect 14922 736 14932 740
rect 11335 731 14932 736
rect 11110 721 11111 731
rect 11075 697 11111 721
rect 11145 721 11151 731
rect 11215 721 11226 731
rect 11285 721 11301 731
rect 11145 697 11181 721
rect 11215 697 11251 721
rect 11285 697 11321 721
rect 11355 697 11391 731
rect 11425 697 11460 731
rect 11494 697 11529 731
rect 11563 697 11598 731
rect 11632 728 14932 731
rect 11632 697 11656 728
rect 9687 671 11656 697
rect 9687 659 9796 671
rect 9830 659 9872 671
rect 9906 659 9948 671
rect 9982 659 10024 671
rect 10058 659 10100 671
rect 10134 659 10176 671
rect 10210 659 10251 671
rect 10285 659 10326 671
rect 10360 659 10401 671
rect 10435 659 10476 671
rect 10510 659 10551 671
rect 10585 659 10626 671
rect 10660 659 10701 671
rect 10735 659 10776 671
rect 10810 659 10851 671
rect 10885 659 10926 671
rect 10960 659 11001 671
rect 11035 659 11076 671
rect 9687 625 9711 659
rect 9745 625 9781 659
rect 9830 637 9851 659
rect 9906 637 9921 659
rect 9982 637 9991 659
rect 10058 637 10061 659
rect 9815 625 9851 637
rect 9885 625 9921 637
rect 9955 625 9991 637
rect 10025 625 10061 637
rect 10095 637 10100 659
rect 10165 637 10176 659
rect 10235 637 10251 659
rect 10305 637 10326 659
rect 10375 637 10401 659
rect 10445 637 10476 659
rect 10095 625 10131 637
rect 10165 625 10201 637
rect 10235 625 10271 637
rect 10305 625 10341 637
rect 10375 625 10411 637
rect 10445 625 10481 637
rect 10515 625 10551 659
rect 10585 625 10621 659
rect 10660 637 10691 659
rect 10735 637 10761 659
rect 10810 637 10831 659
rect 10885 637 10901 659
rect 10960 637 10971 659
rect 11035 637 11041 659
rect 10655 625 10691 637
rect 10725 625 10761 637
rect 10795 625 10831 637
rect 10865 625 10901 637
rect 10935 625 10971 637
rect 11005 625 11041 637
rect 11075 637 11076 659
rect 11110 659 11151 671
rect 11185 659 11226 671
rect 11260 659 11301 671
rect 11335 659 11656 671
rect 11110 637 11111 659
rect 11075 625 11111 637
rect 11145 637 11151 659
rect 11215 637 11226 659
rect 11285 637 11301 659
rect 11145 625 11181 637
rect 11215 625 11251 637
rect 11285 625 11321 637
rect 11355 625 11391 659
rect 11425 625 11460 659
rect 11494 625 11529 659
rect 11563 625 11598 659
rect 11632 625 11656 659
rect 9687 587 11656 625
rect 9687 553 9711 587
rect 9745 553 9781 587
rect 9830 553 9851 587
rect 9906 553 9921 587
rect 9982 553 9991 587
rect 10058 553 10061 587
rect 10095 553 10100 587
rect 10165 553 10176 587
rect 10235 553 10251 587
rect 10305 553 10326 587
rect 10375 553 10401 587
rect 10445 553 10476 587
rect 10515 553 10551 587
rect 10585 553 10621 587
rect 10660 553 10691 587
rect 10735 553 10761 587
rect 10810 553 10831 587
rect 10885 553 10901 587
rect 10960 553 10971 587
rect 11035 553 11041 587
rect 11075 553 11076 587
rect 11110 553 11111 587
rect 11145 553 11151 587
rect 11215 553 11226 587
rect 11285 553 11301 587
rect 11355 553 11391 587
rect 11425 553 11460 587
rect 11494 553 11529 587
rect 11563 553 11598 587
rect 11632 553 11656 587
rect 9687 515 11656 553
rect 9687 481 9711 515
rect 9745 481 9781 515
rect 9815 503 9851 515
rect 9885 503 9921 515
rect 9955 503 9991 515
rect 10025 503 10061 515
rect 9830 481 9851 503
rect 9906 481 9921 503
rect 9982 481 9991 503
rect 10058 481 10061 503
rect 10095 503 10131 515
rect 10165 503 10201 515
rect 10235 503 10271 515
rect 10305 503 10341 515
rect 10375 503 10411 515
rect 10445 503 10481 515
rect 10095 481 10100 503
rect 10165 481 10176 503
rect 10235 481 10251 503
rect 10305 481 10326 503
rect 10375 481 10401 503
rect 10445 481 10476 503
rect 10515 481 10551 515
rect 10585 481 10621 515
rect 10655 503 10691 515
rect 10725 503 10761 515
rect 10795 503 10831 515
rect 10865 503 10901 515
rect 10935 503 10971 515
rect 11005 503 11041 515
rect 10660 481 10691 503
rect 10735 481 10761 503
rect 10810 481 10831 503
rect 10885 481 10901 503
rect 10960 481 10971 503
rect 11035 481 11041 503
rect 11075 503 11111 515
rect 11075 481 11076 503
rect 9687 469 9796 481
rect 9830 469 9872 481
rect 9906 469 9948 481
rect 9982 469 10024 481
rect 10058 469 10100 481
rect 10134 469 10176 481
rect 10210 469 10251 481
rect 10285 469 10326 481
rect 10360 469 10401 481
rect 10435 469 10476 481
rect 10510 469 10551 481
rect 10585 469 10626 481
rect 10660 469 10701 481
rect 10735 469 10776 481
rect 10810 469 10851 481
rect 10885 469 10926 481
rect 10960 469 11001 481
rect 11035 469 11076 481
rect 11110 481 11111 503
rect 11145 503 11181 515
rect 11215 503 11251 515
rect 11285 503 11321 515
rect 11145 481 11151 503
rect 11215 481 11226 503
rect 11285 481 11301 503
rect 11355 481 11391 515
rect 11425 481 11460 515
rect 11494 481 11529 515
rect 11563 481 11598 515
rect 11632 481 11656 515
rect 11110 469 11151 481
rect 11185 469 11226 481
rect 11260 469 11301 481
rect 11335 469 11656 481
rect 9687 443 11656 469
rect 9687 409 9711 443
rect 9745 409 9781 443
rect 9815 409 9851 443
rect 9885 409 9921 443
rect 9955 409 9991 443
rect 10025 409 10061 443
rect 10095 409 10131 443
rect 10165 409 10201 443
rect 10235 409 10271 443
rect 10305 409 10341 443
rect 10375 409 10411 443
rect 10445 409 10481 443
rect 10515 409 10551 443
rect 10585 409 10621 443
rect 10655 409 10691 443
rect 10725 409 10761 443
rect 10795 409 10831 443
rect 10865 409 10901 443
rect 10935 409 10971 443
rect 11005 409 11041 443
rect 11075 409 11111 443
rect 11145 409 11181 443
rect 11215 409 11251 443
rect 11285 409 11321 443
rect 11355 409 11391 443
rect 11425 409 11460 443
rect 11494 409 11529 443
rect 11563 409 11598 443
rect 11632 409 11656 443
rect 9687 369 11656 409
rect 14465 706 14932 728
rect 15000 743 15068 770
rect 15102 743 15117 777
rect 15000 740 15117 743
rect 14966 706 15000 736
rect 15034 706 15068 740
rect 15102 706 15117 740
rect 14465 705 15117 706
rect 14465 697 15068 705
rect 14465 695 14576 697
rect 14610 695 14654 697
rect 14688 695 14732 697
rect 14499 661 14543 695
rect 14610 663 14621 695
rect 14688 663 14698 695
rect 14577 661 14621 663
rect 14655 661 14698 663
rect 14766 695 14810 697
rect 14766 663 14775 695
rect 14732 661 14775 663
rect 14809 663 14810 695
rect 14844 695 14888 697
rect 14844 663 14852 695
rect 14809 661 14852 663
rect 14886 663 14888 695
rect 14922 668 14966 697
rect 14922 663 14932 668
rect 14886 661 14932 663
rect 14465 634 14932 661
rect 15000 671 15068 697
rect 15102 671 15117 705
rect 15000 668 15117 671
rect 14966 634 15000 663
rect 15034 634 15068 668
rect 15102 634 15117 668
rect 14465 633 15117 634
rect 14465 623 15068 633
rect 14465 609 14576 623
rect 14610 609 14654 623
rect 14688 609 14732 623
rect 14499 575 14543 609
rect 14610 589 14621 609
rect 14688 589 14698 609
rect 14577 575 14621 589
rect 14655 575 14698 589
rect 14766 609 14810 623
rect 14766 589 14775 609
rect 14732 575 14775 589
rect 14809 589 14810 609
rect 14844 609 14888 623
rect 14844 589 14852 609
rect 14809 575 14852 589
rect 14886 589 14888 609
rect 14922 596 14966 623
rect 14922 589 14932 596
rect 14886 575 14932 589
rect 14465 562 14932 575
rect 15000 599 15068 623
rect 15102 599 15117 633
rect 15000 596 15117 599
rect 14966 562 15000 589
rect 15034 562 15068 596
rect 15102 562 15117 596
rect 14465 561 15117 562
rect 14465 549 15068 561
rect 14465 523 14576 549
rect 14610 523 14654 549
rect 14688 523 14732 549
rect 14499 489 14543 523
rect 14610 515 14621 523
rect 14688 515 14698 523
rect 14577 489 14621 515
rect 14655 489 14698 515
rect 14766 523 14810 549
rect 14766 515 14775 523
rect 14732 489 14775 515
rect 14809 515 14810 523
rect 14844 523 14888 549
rect 14844 515 14852 523
rect 14809 489 14852 515
rect 14886 515 14888 523
rect 14922 524 14966 549
rect 14922 515 14932 524
rect 14886 490 14932 515
rect 15000 527 15068 549
rect 15102 527 15117 561
rect 15000 524 15117 527
rect 14966 490 15000 515
rect 15034 490 15068 524
rect 15102 490 15117 524
rect 14886 489 15117 490
rect 14465 475 15068 489
rect 14465 441 14576 475
rect 14610 441 14654 475
rect 14688 441 14732 475
rect 14766 441 14810 475
rect 14844 441 14888 475
rect 14922 452 14966 475
rect 14922 441 14932 452
rect 14465 437 14932 441
rect 14499 403 14543 437
rect 14577 403 14621 437
rect 14655 403 14698 437
rect 14732 403 14775 437
rect 14809 403 14852 437
rect 14886 418 14932 437
rect 15000 455 15068 475
rect 15102 455 15117 489
rect 15000 452 15117 455
rect 14966 418 15000 441
rect 15034 418 15068 452
rect 15102 418 15117 452
rect 14886 417 15117 418
rect 14886 403 15068 417
rect 14465 390 15068 403
rect 14465 369 14657 390
rect 7022 367 14657 369
rect 14691 367 14735 390
rect 14769 367 14813 390
rect 14847 367 14891 390
rect 14925 380 14969 390
rect 15003 383 15068 390
rect 15102 383 15117 417
rect 15003 380 15117 383
rect 7022 333 7056 367
rect 7090 333 7125 367
rect 7159 333 7194 367
rect 7228 333 7263 367
rect 7297 333 7332 367
rect 7366 333 7401 367
rect 7435 333 7470 367
rect 7504 333 7539 367
rect 7573 333 7608 367
rect 7642 333 7677 367
rect 7711 333 7746 367
rect 7780 333 7815 367
rect 7849 333 7884 367
rect 7918 333 7953 367
rect 7987 333 8022 367
rect 8056 333 8091 367
rect 8125 333 8160 367
rect 8194 333 8229 367
rect 8263 333 8298 367
rect 8332 333 8367 367
rect 8401 333 8436 367
rect 8470 333 8505 367
rect 8539 333 8574 367
rect 8608 333 8643 367
rect 8677 333 8712 367
rect 8746 333 8781 367
rect 8815 333 8850 367
rect 8884 333 8919 367
rect 8953 333 8988 367
rect 9022 333 9057 367
rect 9091 333 9126 367
rect 9160 333 9195 367
rect 9229 333 9264 367
rect 9298 333 9333 367
rect 9367 333 9402 367
rect 9436 333 9471 367
rect 9505 333 9540 367
rect 9574 333 9609 367
rect 9643 333 9678 367
rect 9712 333 9747 367
rect 9781 333 9816 367
rect 9850 333 9885 367
rect 9919 333 9954 367
rect 9988 333 10023 367
rect 10057 333 10092 367
rect 10126 333 10161 367
rect 10195 333 10230 367
rect 10264 333 10299 367
rect 10333 333 10368 367
rect 10402 333 10437 367
rect 10471 333 10506 367
rect 10540 333 10575 367
rect 10609 333 10643 367
rect 10677 333 10711 367
rect 10745 333 10779 367
rect 10813 333 10847 367
rect 10881 333 10915 367
rect 10949 333 10983 367
rect 11017 333 11051 367
rect 11085 333 11119 367
rect 11153 333 11187 367
rect 11221 333 11255 367
rect 11289 333 11323 367
rect 11357 333 11391 367
rect 11425 333 11459 367
rect 11493 333 11527 367
rect 11561 333 11595 367
rect 11629 333 11663 367
rect 11697 333 11731 367
rect 11765 333 11799 367
rect 11833 333 11867 367
rect 11901 333 11935 367
rect 11969 333 12003 367
rect 12037 333 12071 367
rect 12105 333 12139 367
rect 12173 333 12207 367
rect 12241 333 12275 367
rect 12309 333 12343 367
rect 12377 333 12411 367
rect 12445 333 12479 367
rect 12513 333 12547 367
rect 12581 333 12615 367
rect 12649 333 12683 367
rect 12717 333 12751 367
rect 12785 333 12819 367
rect 12853 333 12887 367
rect 12921 333 12955 367
rect 12989 333 13023 367
rect 13057 333 13091 367
rect 13125 333 13159 367
rect 13193 333 13227 367
rect 13261 333 13295 367
rect 13329 333 13363 367
rect 13397 333 13431 367
rect 13465 333 13499 367
rect 13533 333 13567 367
rect 13601 333 13635 367
rect 13669 333 13703 367
rect 13737 333 13771 367
rect 13805 333 13839 367
rect 13873 333 13907 367
rect 13941 333 13975 367
rect 14009 333 14043 367
rect 14077 333 14111 367
rect 14145 333 14179 367
rect 14213 333 14247 367
rect 14281 333 14315 367
rect 14349 333 14383 367
rect 14417 333 14451 367
rect 14485 333 14519 367
rect 14553 333 14587 367
rect 14621 333 14655 367
rect 14691 356 14723 367
rect 14769 356 14791 367
rect 14847 356 14859 367
rect 14925 356 14932 380
rect 14689 333 14723 356
rect 14757 333 14791 356
rect 14825 333 14859 356
rect 14893 346 14932 356
rect 14966 356 14969 380
rect 14966 346 15000 356
rect 15034 346 15068 380
rect 15102 346 15117 380
rect 14893 345 15117 346
rect 14893 333 15068 345
rect 7022 312 15068 333
rect 7022 289 14657 312
rect 14691 289 14735 312
rect 14769 289 14813 312
rect 14847 289 14891 312
rect 14925 308 14969 312
rect 15003 311 15068 312
rect 15102 311 15117 345
rect 15003 308 15117 311
rect 7022 255 7056 289
rect 7090 255 7125 289
rect 7159 255 7194 289
rect 7228 255 7263 289
rect 7297 255 7332 289
rect 7366 255 7401 289
rect 7435 255 7470 289
rect 7504 255 7539 289
rect 7573 255 7608 289
rect 7642 255 7677 289
rect 7711 255 7746 289
rect 7780 255 7815 289
rect 7849 255 7884 289
rect 7918 255 7953 289
rect 7987 255 8022 289
rect 8056 255 8091 289
rect 8125 255 8160 289
rect 8194 255 8229 289
rect 8263 255 8298 289
rect 8332 255 8367 289
rect 8401 255 8436 289
rect 8470 255 8505 289
rect 8539 255 8574 289
rect 8608 255 8643 289
rect 8677 255 8712 289
rect 8746 255 8781 289
rect 8815 255 8850 289
rect 8884 255 8919 289
rect 8953 255 8988 289
rect 9022 255 9057 289
rect 9091 255 9126 289
rect 9160 255 9195 289
rect 9229 255 9264 289
rect 9298 255 9333 289
rect 9367 255 9402 289
rect 9436 255 9471 289
rect 9505 255 9540 289
rect 9574 255 9609 289
rect 9643 255 9678 289
rect 9712 255 9747 289
rect 9781 255 9816 289
rect 9850 255 9885 289
rect 9919 255 9954 289
rect 9988 255 10023 289
rect 10057 255 10092 289
rect 10126 255 10161 289
rect 10195 255 10230 289
rect 10264 255 10299 289
rect 10333 255 10368 289
rect 10402 255 10437 289
rect 10471 255 10506 289
rect 10540 255 10575 289
rect 10609 255 10643 289
rect 10677 255 10711 289
rect 10745 255 10779 289
rect 10813 255 10847 289
rect 10881 255 10915 289
rect 10949 255 10983 289
rect 11017 255 11051 289
rect 11085 255 11119 289
rect 11153 255 11187 289
rect 11221 255 11255 289
rect 11289 255 11323 289
rect 11357 255 11391 289
rect 11425 255 11459 289
rect 11493 255 11527 289
rect 11561 255 11595 289
rect 11629 255 11663 289
rect 11697 255 11731 289
rect 11765 255 11799 289
rect 11833 255 11867 289
rect 11901 255 11935 289
rect 11969 255 12003 289
rect 12037 255 12071 289
rect 12105 255 12139 289
rect 12173 255 12207 289
rect 12241 255 12275 289
rect 12309 255 12343 289
rect 12377 255 12411 289
rect 12445 255 12479 289
rect 12513 255 12547 289
rect 12581 255 12615 289
rect 12649 255 12683 289
rect 12717 255 12751 289
rect 12785 255 12819 289
rect 12853 255 12887 289
rect 12921 255 12955 289
rect 12989 255 13023 289
rect 13057 255 13091 289
rect 13125 255 13159 289
rect 13193 255 13227 289
rect 13261 255 13295 289
rect 13329 255 13363 289
rect 13397 255 13431 289
rect 13465 255 13499 289
rect 13533 255 13567 289
rect 13601 255 13635 289
rect 13669 255 13703 289
rect 13737 255 13771 289
rect 13805 255 13839 289
rect 13873 255 13907 289
rect 13941 255 13975 289
rect 14009 255 14043 289
rect 14077 255 14111 289
rect 14145 255 14179 289
rect 14213 255 14247 289
rect 14281 255 14315 289
rect 14349 255 14383 289
rect 14417 255 14451 289
rect 14485 255 14519 289
rect 14553 255 14587 289
rect 14621 255 14655 289
rect 14691 278 14723 289
rect 14769 278 14791 289
rect 14847 278 14859 289
rect 14925 278 14932 308
rect 14689 255 14723 278
rect 14757 255 14791 278
rect 14825 255 14859 278
rect 14893 274 14932 278
rect 14966 278 14969 308
rect 14966 274 15000 278
rect 15034 274 15068 308
rect 15102 274 15117 308
rect 14893 272 15117 274
rect 14893 255 15068 272
rect 7022 238 15068 255
rect 15102 238 15117 272
rect 7022 236 15117 238
rect 7022 234 14932 236
rect 7022 211 14657 234
rect 14691 211 14735 234
rect 14769 211 14813 234
rect 14847 211 14891 234
rect 7022 177 7056 211
rect 7090 177 7125 211
rect 7159 177 7194 211
rect 7228 177 7263 211
rect 7297 177 7332 211
rect 7366 177 7401 211
rect 7435 177 7470 211
rect 7504 177 7539 211
rect 7573 177 7608 211
rect 7642 177 7677 211
rect 7711 177 7746 211
rect 7780 177 7815 211
rect 7849 177 7884 211
rect 7918 177 7953 211
rect 7987 177 8022 211
rect 8056 177 8091 211
rect 8125 177 8160 211
rect 8194 177 8229 211
rect 8263 177 8298 211
rect 8332 177 8367 211
rect 8401 177 8436 211
rect 8470 177 8505 211
rect 8539 177 8574 211
rect 8608 177 8643 211
rect 8677 177 8712 211
rect 8746 177 8781 211
rect 8815 177 8850 211
rect 8884 177 8919 211
rect 8953 177 8988 211
rect 9022 177 9057 211
rect 9091 177 9126 211
rect 9160 177 9195 211
rect 9229 177 9264 211
rect 9298 177 9333 211
rect 9367 177 9402 211
rect 9436 177 9471 211
rect 9505 177 9540 211
rect 9574 177 9609 211
rect 9643 177 9678 211
rect 9712 177 9747 211
rect 9781 177 9816 211
rect 9850 177 9885 211
rect 9919 177 9954 211
rect 9988 177 10023 211
rect 10057 177 10092 211
rect 10126 177 10161 211
rect 10195 177 10230 211
rect 10264 177 10299 211
rect 10333 177 10368 211
rect 10402 177 10437 211
rect 10471 177 10506 211
rect 10540 177 10575 211
rect 10609 177 10643 211
rect 10677 177 10711 211
rect 10745 177 10779 211
rect 10813 177 10847 211
rect 10881 177 10915 211
rect 10949 177 10983 211
rect 11017 177 11051 211
rect 11085 177 11119 211
rect 11153 177 11187 211
rect 11221 177 11255 211
rect 11289 177 11323 211
rect 11357 177 11391 211
rect 11425 177 11459 211
rect 11493 177 11527 211
rect 11561 177 11595 211
rect 11629 177 11663 211
rect 11697 177 11731 211
rect 11765 177 11799 211
rect 11833 177 11867 211
rect 11901 177 11935 211
rect 11969 177 12003 211
rect 12037 177 12071 211
rect 12105 177 12139 211
rect 12173 177 12207 211
rect 12241 177 12275 211
rect 12309 177 12343 211
rect 12377 177 12411 211
rect 12445 177 12479 211
rect 12513 177 12547 211
rect 12581 177 12615 211
rect 12649 177 12683 211
rect 12717 177 12751 211
rect 12785 177 12819 211
rect 12853 177 12887 211
rect 12921 177 12955 211
rect 12989 177 13023 211
rect 13057 177 13091 211
rect 13125 177 13159 211
rect 13193 177 13227 211
rect 13261 177 13295 211
rect 13329 177 13363 211
rect 13397 177 13431 211
rect 13465 177 13499 211
rect 13533 177 13567 211
rect 13601 177 13635 211
rect 13669 177 13703 211
rect 13737 177 13771 211
rect 13805 177 13839 211
rect 13873 177 13907 211
rect 13941 177 13975 211
rect 14009 177 14043 211
rect 14077 177 14111 211
rect 14145 177 14179 211
rect 14213 177 14247 211
rect 14281 177 14315 211
rect 14349 177 14383 211
rect 14417 177 14451 211
rect 14485 177 14519 211
rect 14553 177 14587 211
rect 14621 177 14655 211
rect 14691 200 14723 211
rect 14769 200 14791 211
rect 14847 200 14859 211
rect 14925 202 14932 234
rect 14966 234 15000 236
rect 14966 202 14969 234
rect 15034 202 15068 236
rect 15102 202 15117 236
rect 14925 200 14969 202
rect 15003 200 15117 202
rect 14689 177 14723 200
rect 14757 177 14791 200
rect 14825 177 14859 200
rect 14893 199 15117 200
rect 14893 177 15068 199
rect 7022 165 15068 177
rect 15102 165 15117 199
rect 7022 164 15117 165
rect 7022 156 14932 164
rect 7022 133 14657 156
rect 14691 133 14735 156
rect 14769 133 14813 156
rect 14847 133 14891 156
rect 7022 99 7056 133
rect 7090 99 7125 133
rect 7159 99 7194 133
rect 7228 99 7263 133
rect 7297 99 7332 133
rect 7366 99 7401 133
rect 7435 99 7470 133
rect 7504 99 7539 133
rect 7573 99 7608 133
rect 7642 99 7677 133
rect 7711 99 7746 133
rect 7780 99 7815 133
rect 7849 99 7884 133
rect 7918 99 7953 133
rect 7987 99 8022 133
rect 8056 99 8091 133
rect 8125 99 8160 133
rect 8194 99 8229 133
rect 8263 99 8298 133
rect 8332 99 8367 133
rect 8401 99 8436 133
rect 8470 99 8505 133
rect 8539 99 8574 133
rect 8608 99 8643 133
rect 8677 99 8712 133
rect 8746 99 8781 133
rect 8815 99 8850 133
rect 8884 99 8919 133
rect 8953 99 8988 133
rect 9022 99 9057 133
rect 9091 99 9126 133
rect 9160 99 9195 133
rect 9229 99 9264 133
rect 9298 99 9333 133
rect 9367 99 9402 133
rect 9436 99 9471 133
rect 9505 99 9540 133
rect 9574 99 9609 133
rect 9643 99 9678 133
rect 9712 99 9747 133
rect 9781 99 9816 133
rect 9850 99 9885 133
rect 9919 99 9954 133
rect 9988 99 10023 133
rect 10057 99 10092 133
rect 10126 99 10161 133
rect 10195 99 10230 133
rect 10264 99 10299 133
rect 10333 99 10368 133
rect 10402 99 10437 133
rect 10471 99 10506 133
rect 10540 99 10575 133
rect 10609 99 10643 133
rect 10677 99 10711 133
rect 10745 99 10779 133
rect 10813 99 10847 133
rect 10881 99 10915 133
rect 10949 99 10983 133
rect 11017 99 11051 133
rect 11085 99 11119 133
rect 11153 99 11187 133
rect 11221 99 11255 133
rect 11289 99 11323 133
rect 11357 99 11391 133
rect 11425 99 11459 133
rect 11493 99 11527 133
rect 11561 99 11595 133
rect 11629 99 11663 133
rect 11697 99 11731 133
rect 11765 99 11799 133
rect 11833 99 11867 133
rect 11901 99 11935 133
rect 11969 99 12003 133
rect 12037 99 12071 133
rect 12105 99 12139 133
rect 12173 99 12207 133
rect 12241 99 12275 133
rect 12309 99 12343 133
rect 12377 99 12411 133
rect 12445 99 12479 133
rect 12513 99 12547 133
rect 12581 99 12615 133
rect 12649 99 12683 133
rect 12717 99 12751 133
rect 12785 99 12819 133
rect 12853 99 12887 133
rect 12921 99 12955 133
rect 12989 99 13023 133
rect 13057 99 13091 133
rect 13125 99 13159 133
rect 13193 99 13227 133
rect 13261 99 13295 133
rect 13329 99 13363 133
rect 13397 99 13431 133
rect 13465 99 13499 133
rect 13533 99 13567 133
rect 13601 99 13635 133
rect 13669 99 13703 133
rect 13737 99 13771 133
rect 13805 99 13839 133
rect 13873 99 13907 133
rect 13941 99 13975 133
rect 14009 99 14043 133
rect 14077 99 14111 133
rect 14145 99 14179 133
rect 14213 99 14247 133
rect 14281 99 14315 133
rect 14349 99 14383 133
rect 14417 99 14451 133
rect 14485 99 14519 133
rect 14553 99 14587 133
rect 14621 99 14655 133
rect 14691 122 14723 133
rect 14769 122 14791 133
rect 14847 122 14859 133
rect 14925 130 14932 156
rect 14966 156 15000 164
rect 14966 130 14969 156
rect 15034 130 15068 164
rect 15102 130 15117 164
rect 14925 122 14969 130
rect 15003 126 15117 130
rect 15003 122 15068 126
rect 14689 99 14723 122
rect 14757 99 14791 122
rect 14825 99 14859 122
rect 14893 99 15068 122
rect 7022 92 15068 99
rect 15102 92 15117 126
rect 7022 91 15117 92
rect 7022 77 14932 91
rect 7022 55 14657 77
rect 14691 55 14735 77
rect 14769 55 14813 77
rect 14847 55 14891 77
rect 14925 57 14932 77
rect 14966 77 15000 91
rect 14966 57 14969 77
rect 15034 57 15068 91
rect 15102 57 15117 91
rect 7022 21 7056 55
rect 7090 21 7125 55
rect 7159 21 7194 55
rect 7228 21 7263 55
rect 7297 21 7332 55
rect 7366 21 7401 55
rect 7435 21 7470 55
rect 7504 21 7539 55
rect 7573 21 7608 55
rect 7642 21 7677 55
rect 7711 21 7746 55
rect 7780 21 7815 55
rect 7849 21 7884 55
rect 7918 21 7953 55
rect 7987 21 8022 55
rect 8056 21 8091 55
rect 8125 21 8160 55
rect 8194 21 8229 55
rect 8263 21 8298 55
rect 8332 21 8367 55
rect 8401 21 8436 55
rect 8470 21 8505 55
rect 8539 21 8574 55
rect 8608 21 8643 55
rect 8677 21 8712 55
rect 8746 21 8781 55
rect 8815 21 8850 55
rect 8884 21 8919 55
rect 8953 21 8988 55
rect 9022 21 9057 55
rect 9091 21 9126 55
rect 9160 21 9195 55
rect 9229 21 9264 55
rect 9298 21 9333 55
rect 9367 21 9402 55
rect 9436 21 9471 55
rect 9505 21 9540 55
rect 9574 21 9609 55
rect 9643 21 9678 55
rect 9712 21 9747 55
rect 9781 21 9816 55
rect 9850 21 9885 55
rect 9919 21 9954 55
rect 9988 21 10023 55
rect 10057 21 10092 55
rect 10126 21 10161 55
rect 10195 21 10230 55
rect 10264 21 10299 55
rect 10333 21 10368 55
rect 10402 21 10437 55
rect 10471 21 10506 55
rect 10540 21 10575 55
rect 10609 21 10643 55
rect 10677 21 10711 55
rect 10745 21 10779 55
rect 10813 21 10847 55
rect 10881 21 10915 55
rect 10949 21 10983 55
rect 11017 21 11051 55
rect 11085 21 11119 55
rect 11153 21 11187 55
rect 11221 21 11255 55
rect 11289 21 11323 55
rect 11357 21 11391 55
rect 11425 21 11459 55
rect 11493 21 11527 55
rect 11561 21 11595 55
rect 11629 21 11663 55
rect 11697 21 11731 55
rect 11765 21 11799 55
rect 11833 21 11867 55
rect 11901 21 11935 55
rect 11969 21 12003 55
rect 12037 21 12071 55
rect 12105 21 12139 55
rect 12173 21 12207 55
rect 12241 21 12275 55
rect 12309 21 12343 55
rect 12377 21 12411 55
rect 12445 21 12479 55
rect 12513 21 12547 55
rect 12581 21 12615 55
rect 12649 21 12683 55
rect 12717 21 12751 55
rect 12785 21 12819 55
rect 12853 21 12887 55
rect 12921 21 12955 55
rect 12989 21 13023 55
rect 13057 21 13091 55
rect 13125 21 13159 55
rect 13193 21 13227 55
rect 13261 21 13295 55
rect 13329 21 13363 55
rect 13397 21 13431 55
rect 13465 21 13499 55
rect 13533 21 13567 55
rect 13601 21 13635 55
rect 13669 21 13703 55
rect 13737 21 13771 55
rect 13805 21 13839 55
rect 13873 21 13907 55
rect 13941 21 13975 55
rect 14009 21 14043 55
rect 14077 21 14111 55
rect 14145 21 14179 55
rect 14213 21 14247 55
rect 14281 21 14315 55
rect 14349 21 14383 55
rect 14417 21 14451 55
rect 14485 21 14519 55
rect 14553 21 14587 55
rect 14621 21 14655 55
rect 14691 43 14723 55
rect 14769 43 14791 55
rect 14847 43 14859 55
rect 14925 43 14969 57
rect 15003 53 15117 57
rect 15003 43 15068 53
rect 14689 21 14723 43
rect 14757 21 14791 43
rect 14825 21 14859 43
rect 14893 21 15068 43
rect 7022 19 15068 21
rect 15102 19 15117 53
rect 5884 -9229 5918 -9191
<< viali >>
rect -484 9510 -482 9514
rect -482 9510 -450 9514
rect -411 9510 -378 9514
rect -378 9510 -377 9514
rect -338 9510 -309 9514
rect -309 9510 -304 9514
rect -265 9510 -240 9514
rect -240 9510 -231 9514
rect -192 9510 -171 9514
rect -171 9510 -158 9514
rect -119 9510 -102 9514
rect -102 9510 -85 9514
rect -484 9480 -450 9510
rect -411 9480 -377 9510
rect -338 9480 -304 9510
rect -265 9480 -231 9510
rect -192 9480 -158 9510
rect -119 9480 -85 9510
rect -46 9480 -33 9514
rect -33 9480 -12 9514
rect 27 9480 61 9514
rect 100 9480 134 9514
rect 173 9480 207 9514
rect 246 9480 280 9514
rect 319 9480 353 9514
rect 392 9480 426 9514
rect 465 9480 499 9514
rect 538 9480 572 9514
rect 611 9480 645 9514
rect 684 9480 718 9514
rect 757 9480 791 9514
rect 830 9480 864 9514
rect 903 9480 937 9514
rect 976 9480 1010 9514
rect 1049 9480 1083 9514
rect 1122 9480 1156 9514
rect 1195 9480 1229 9514
rect 1268 9480 1302 9514
rect 1341 9480 1375 9514
rect 1414 9480 1448 9514
rect 1487 9480 1521 9514
rect 1559 9480 1593 9514
rect 1631 9480 1665 9514
rect 1703 9480 1737 9514
rect 1775 9480 1809 9514
rect 1847 9480 1881 9514
rect 1919 9480 1953 9514
rect 1991 9480 2025 9514
rect 2063 9480 2097 9514
rect 2135 9480 2169 9514
rect 2207 9480 2241 9514
rect 2279 9480 2313 9514
rect 2351 9480 2385 9514
rect 2423 9480 2457 9514
rect 2495 9480 2529 9514
rect 2567 9480 2601 9514
rect 2639 9480 2673 9514
rect 2711 9480 2745 9514
rect 2783 9480 2817 9514
rect 2855 9480 2889 9514
rect 2927 9480 2961 9514
rect 2999 9480 3033 9514
rect 3071 9480 3105 9514
rect 3143 9480 3177 9514
rect 3215 9480 3249 9514
rect 3287 9480 3321 9514
rect 3359 9480 3393 9514
rect 3431 9480 3465 9514
rect 3503 9480 3537 9514
rect 3575 9480 3609 9514
rect 3647 9480 3681 9514
rect 3719 9480 3753 9514
rect 3791 9480 3825 9514
rect 3863 9480 3897 9514
rect 3935 9480 3969 9514
rect 4007 9480 4041 9514
rect 4079 9480 4113 9514
rect 4151 9480 4185 9514
rect 4223 9480 4257 9514
rect 4295 9480 4329 9514
rect 4367 9480 4401 9514
rect 4439 9480 4473 9514
rect 4511 9480 4545 9514
rect 4583 9480 4617 9514
rect 4655 9480 4689 9514
rect 4727 9480 4761 9514
rect 4799 9480 4833 9514
rect 4871 9480 4905 9514
rect 4943 9480 4977 9514
rect 5015 9480 5049 9514
rect 5087 9480 5121 9514
rect 5159 9480 5193 9514
rect 5231 9480 5265 9514
rect 5303 9480 5337 9514
rect 5375 9480 5409 9514
rect 5447 9480 5481 9514
rect 5519 9480 5553 9514
rect 5591 9480 5625 9514
rect 5663 9480 5697 9514
rect 5735 9480 5769 9514
rect 5807 9480 5841 9514
rect 5879 9480 5913 9514
rect 5951 9480 5985 9514
rect 6023 9480 6057 9514
rect 6095 9480 6129 9514
rect 6167 9480 6201 9514
rect 6239 9480 6273 9514
rect 6311 9480 6345 9514
rect 6383 9480 6417 9514
rect 6455 9480 6489 9514
rect 6527 9480 6561 9514
rect 6599 9480 6633 9514
rect 6671 9480 6705 9514
rect 6743 9480 6777 9514
rect 6815 9480 6849 9514
rect 6887 9480 6921 9514
rect 6959 9480 6993 9514
rect 7031 9480 7065 9514
rect 7103 9480 7137 9514
rect 7175 9480 7209 9514
rect 7247 9480 7281 9514
rect 7319 9480 7353 9514
rect 7391 9480 7425 9514
rect 7463 9480 7497 9514
rect 7535 9480 7569 9514
rect 7607 9480 7641 9514
rect 7679 9480 7713 9514
rect 7751 9480 7785 9514
rect 7823 9480 7857 9514
rect 7895 9480 7929 9514
rect 7967 9480 8001 9514
rect 8039 9480 8073 9514
rect 8111 9480 8145 9514
rect 8183 9480 8217 9514
rect 8255 9480 8289 9514
rect 8327 9480 8361 9514
rect 8399 9480 8433 9514
rect 8471 9480 8505 9514
rect 8543 9480 8577 9514
rect 8615 9480 8649 9514
rect 8687 9480 8721 9514
rect 8759 9480 8793 9514
rect 8831 9480 8865 9514
rect 8903 9480 8937 9514
rect 8975 9480 9009 9514
rect 9047 9480 9081 9514
rect 9119 9480 9153 9514
rect 9191 9480 9225 9514
rect 9263 9480 9297 9514
rect 9335 9480 9369 9514
rect 9407 9480 9441 9514
rect 9479 9480 9513 9514
rect 9551 9480 9585 9514
rect 9623 9480 9657 9514
rect 9695 9480 9729 9514
rect 9767 9480 9801 9514
rect 9839 9480 9873 9514
rect 9911 9480 9945 9514
rect 9983 9480 10017 9514
rect 10055 9480 10089 9514
rect 10127 9480 10161 9514
rect 10199 9480 10233 9514
rect 10271 9480 10305 9514
rect 10343 9480 10377 9514
rect 10415 9480 10449 9514
rect 10487 9480 10521 9514
rect 10559 9480 10593 9514
rect 10631 9480 10665 9514
rect 10703 9480 10737 9514
rect 10775 9480 10809 9514
rect 10847 9480 10881 9514
rect 10919 9480 10953 9514
rect 10991 9480 11025 9514
rect 11063 9480 11097 9514
rect 11135 9480 11169 9514
rect 11207 9480 11241 9514
rect 11279 9480 11313 9514
rect 11351 9480 11385 9514
rect 11423 9480 11457 9514
rect 11495 9480 11529 9514
rect 11567 9480 11601 9514
rect 11639 9480 11673 9514
rect 11711 9480 11745 9514
rect 11783 9480 11817 9514
rect 11855 9480 11889 9514
rect 11927 9480 11961 9514
rect 11999 9480 12033 9514
rect 12071 9480 12105 9514
rect 12143 9480 12177 9514
rect 12215 9480 12249 9514
rect 12287 9480 12321 9514
rect 12359 9480 12393 9514
rect 12431 9480 12465 9514
rect 12503 9480 12537 9514
rect 12575 9480 12609 9514
rect 12647 9480 12681 9514
rect 12719 9480 12753 9514
rect 12791 9480 12825 9514
rect 12863 9480 12897 9514
rect 12935 9480 12969 9514
rect 13007 9480 13041 9514
rect 13079 9480 13113 9514
rect 13151 9480 13185 9514
rect 13223 9480 13257 9514
rect 13295 9480 13329 9514
rect 13367 9480 13401 9514
rect 13439 9480 13473 9514
rect 13511 9480 13545 9514
rect 13583 9480 13617 9514
rect 13655 9480 13689 9514
rect 13727 9480 13761 9514
rect 13799 9480 13833 9514
rect -484 9408 -450 9428
rect -411 9408 -377 9428
rect -338 9408 -304 9428
rect -265 9408 -231 9428
rect -192 9408 -158 9428
rect -119 9408 -85 9428
rect -484 9394 -482 9408
rect -482 9394 -450 9408
rect -411 9394 -378 9408
rect -378 9394 -377 9408
rect -338 9394 -309 9408
rect -309 9394 -304 9408
rect -265 9394 -240 9408
rect -240 9394 -231 9408
rect -192 9394 -171 9408
rect -171 9394 -158 9408
rect -119 9394 -102 9408
rect -102 9394 -85 9408
rect -46 9394 -33 9428
rect -33 9394 -12 9428
rect 27 9394 61 9428
rect 100 9394 134 9428
rect 173 9394 207 9428
rect 246 9394 280 9428
rect 319 9394 353 9428
rect 392 9394 426 9428
rect 465 9394 499 9428
rect 538 9394 572 9428
rect 611 9394 645 9428
rect 684 9394 718 9428
rect 757 9394 791 9428
rect 830 9394 864 9428
rect 903 9394 937 9428
rect 976 9394 1010 9428
rect 1049 9394 1083 9428
rect 1122 9394 1156 9428
rect 1195 9394 1229 9428
rect 1268 9394 1302 9428
rect 1341 9394 1375 9428
rect 1414 9394 1448 9428
rect 1487 9394 1521 9428
rect 1559 9394 1593 9428
rect 1631 9394 1665 9428
rect 1703 9394 1737 9428
rect 1775 9394 1809 9428
rect 1847 9394 1881 9428
rect 1919 9394 1953 9428
rect 1991 9394 2025 9428
rect 2063 9394 2097 9428
rect 2135 9394 2169 9428
rect 2207 9394 2241 9428
rect 2279 9394 2313 9428
rect 2351 9394 2385 9428
rect 2423 9394 2457 9428
rect 2495 9394 2529 9428
rect 2567 9394 2601 9428
rect 2639 9394 2673 9428
rect 2711 9394 2745 9428
rect 2783 9394 2817 9428
rect 2855 9394 2889 9428
rect 2927 9394 2961 9428
rect 2999 9394 3033 9428
rect 3071 9394 3105 9428
rect 3143 9394 3177 9428
rect 3215 9394 3249 9428
rect 3287 9394 3321 9428
rect 3359 9394 3393 9428
rect 3431 9394 3465 9428
rect 3503 9394 3537 9428
rect 3575 9394 3609 9428
rect 3647 9394 3681 9428
rect 3719 9394 3753 9428
rect 3791 9394 3825 9428
rect 3863 9394 3897 9428
rect 3935 9394 3969 9428
rect 4007 9394 4041 9428
rect 4079 9394 4113 9428
rect 4151 9394 4185 9428
rect 4223 9394 4257 9428
rect 4295 9394 4329 9428
rect 4367 9394 4401 9428
rect 4439 9394 4473 9428
rect 4511 9394 4545 9428
rect 4583 9394 4617 9428
rect 4655 9394 4689 9428
rect 4727 9394 4761 9428
rect 4799 9394 4833 9428
rect 4871 9394 4905 9428
rect 4943 9394 4977 9428
rect 5015 9394 5049 9428
rect 5087 9394 5121 9428
rect 5159 9394 5193 9428
rect 5231 9394 5265 9428
rect 5303 9394 5337 9428
rect 5375 9394 5409 9428
rect 5447 9394 5481 9428
rect 5519 9394 5553 9428
rect 5591 9394 5625 9428
rect 5663 9394 5697 9428
rect 5735 9394 5769 9428
rect 5807 9394 5841 9428
rect 5879 9394 5913 9428
rect 5951 9394 5985 9428
rect 6023 9394 6057 9428
rect 6095 9394 6129 9428
rect 6167 9394 6201 9428
rect 6239 9394 6273 9428
rect 6311 9394 6345 9428
rect 6383 9394 6417 9428
rect 6455 9394 6489 9428
rect 6527 9394 6561 9428
rect 6599 9394 6633 9428
rect 6671 9394 6705 9428
rect 6743 9394 6777 9428
rect 6815 9394 6849 9428
rect 6887 9394 6921 9428
rect 6959 9394 6993 9428
rect 7031 9394 7065 9428
rect 7103 9394 7137 9428
rect 7175 9394 7209 9428
rect 7247 9394 7281 9428
rect 7319 9394 7353 9428
rect 7391 9394 7425 9428
rect 7463 9394 7497 9428
rect 7535 9394 7569 9428
rect 7607 9394 7641 9428
rect 7679 9394 7713 9428
rect 7751 9394 7785 9428
rect 7823 9394 7857 9428
rect 7895 9394 7929 9428
rect 7967 9394 8001 9428
rect 8039 9394 8073 9428
rect 8111 9394 8145 9428
rect 8183 9394 8217 9428
rect 8255 9394 8289 9428
rect 8327 9394 8361 9428
rect 8399 9394 8433 9428
rect 8471 9394 8505 9428
rect 8543 9394 8577 9428
rect 8615 9394 8649 9428
rect 8687 9394 8721 9428
rect 8759 9394 8793 9428
rect 8831 9394 8865 9428
rect 8903 9394 8937 9428
rect 8975 9394 9009 9428
rect 9047 9394 9081 9428
rect 9119 9394 9153 9428
rect 9191 9394 9225 9428
rect 9263 9394 9297 9428
rect 9335 9394 9369 9428
rect 9407 9394 9441 9428
rect 9479 9394 9513 9428
rect 9551 9394 9585 9428
rect 9623 9394 9657 9428
rect 9695 9394 9729 9428
rect 9767 9394 9801 9428
rect 9839 9394 9873 9428
rect 9911 9394 9945 9428
rect 9983 9394 10017 9428
rect 10055 9394 10089 9428
rect 10127 9394 10161 9428
rect 10199 9394 10233 9428
rect 10271 9394 10305 9428
rect 10343 9394 10377 9428
rect 10415 9394 10449 9428
rect 10487 9394 10521 9428
rect 10559 9394 10593 9428
rect 10631 9394 10665 9428
rect 10703 9394 10737 9428
rect 10775 9394 10809 9428
rect 10847 9394 10881 9428
rect 10919 9394 10953 9428
rect 10991 9394 11025 9428
rect 11063 9394 11097 9428
rect 11135 9394 11169 9428
rect 11207 9394 11241 9428
rect 11279 9394 11313 9428
rect 11351 9394 11385 9428
rect 11423 9394 11457 9428
rect 11495 9394 11529 9428
rect 11567 9394 11601 9428
rect 11639 9394 11673 9428
rect 11711 9394 11745 9428
rect 11783 9394 11817 9428
rect 11855 9394 11889 9428
rect 11927 9394 11961 9428
rect 11999 9394 12033 9428
rect 12071 9394 12105 9428
rect 12143 9394 12177 9428
rect 12215 9394 12249 9428
rect 12287 9394 12321 9428
rect 12359 9394 12393 9428
rect 12431 9394 12465 9428
rect 12503 9394 12537 9428
rect 12575 9394 12609 9428
rect 12647 9394 12681 9428
rect 12719 9394 12753 9428
rect 12791 9394 12825 9428
rect 12863 9394 12897 9428
rect 12935 9394 12969 9428
rect 13007 9394 13041 9428
rect 13079 9394 13113 9428
rect 13151 9394 13185 9428
rect 13223 9394 13257 9428
rect 13295 9394 13329 9428
rect 13367 9394 13401 9428
rect 13439 9394 13473 9428
rect 13511 9394 13545 9428
rect 13583 9394 13617 9428
rect 13655 9394 13689 9428
rect 13727 9394 13761 9428
rect 13799 9394 13833 9428
rect -484 9340 -450 9342
rect -411 9340 -377 9342
rect -338 9340 -304 9342
rect -265 9340 -231 9342
rect -192 9340 -158 9342
rect -119 9340 -85 9342
rect -484 9308 -482 9340
rect -482 9308 -450 9340
rect -411 9308 -378 9340
rect -378 9308 -377 9340
rect -338 9308 -309 9340
rect -309 9308 -304 9340
rect -265 9308 -240 9340
rect -240 9308 -231 9340
rect -192 9308 -171 9340
rect -171 9308 -158 9340
rect -119 9308 -102 9340
rect -102 9308 -85 9340
rect -46 9308 -33 9342
rect -33 9308 -12 9342
rect 27 9308 61 9342
rect 100 9308 134 9342
rect 173 9308 207 9342
rect 246 9308 280 9342
rect 319 9308 353 9342
rect 392 9308 426 9342
rect 465 9308 499 9342
rect 538 9308 572 9342
rect 611 9308 645 9342
rect 684 9308 718 9342
rect 757 9308 791 9342
rect 830 9308 864 9342
rect 903 9308 937 9342
rect 976 9308 1010 9342
rect 1049 9308 1083 9342
rect 1122 9308 1156 9342
rect 1195 9308 1229 9342
rect 1268 9308 1302 9342
rect 1341 9308 1375 9342
rect 1414 9308 1448 9342
rect 1487 9308 1521 9342
rect 1559 9308 1593 9342
rect 1631 9308 1665 9342
rect 1703 9308 1737 9342
rect 1775 9308 1809 9342
rect 1847 9308 1881 9342
rect 1919 9308 1953 9342
rect 1991 9308 2025 9342
rect 2063 9308 2097 9342
rect 2135 9308 2169 9342
rect 2207 9308 2241 9342
rect 2279 9308 2313 9342
rect 2351 9308 2385 9342
rect 2423 9308 2457 9342
rect 2495 9308 2529 9342
rect 2567 9308 2601 9342
rect 2639 9308 2673 9342
rect 2711 9308 2745 9342
rect 2783 9308 2817 9342
rect 2855 9308 2889 9342
rect 2927 9308 2961 9342
rect 2999 9308 3033 9342
rect 3071 9308 3105 9342
rect 3143 9308 3177 9342
rect 3215 9308 3249 9342
rect 3287 9308 3321 9342
rect 3359 9308 3393 9342
rect 3431 9308 3465 9342
rect 3503 9308 3537 9342
rect 3575 9308 3609 9342
rect 3647 9308 3681 9342
rect 3719 9308 3753 9342
rect 3791 9308 3825 9342
rect 3863 9308 3897 9342
rect 3935 9308 3969 9342
rect 4007 9308 4041 9342
rect 4079 9308 4113 9342
rect 4151 9308 4185 9342
rect 4223 9308 4257 9342
rect 4295 9308 4329 9342
rect 4367 9308 4401 9342
rect 4439 9308 4473 9342
rect 4511 9308 4545 9342
rect 4583 9308 4617 9342
rect 4655 9308 4689 9342
rect 4727 9308 4761 9342
rect 4799 9308 4833 9342
rect 4871 9308 4905 9342
rect 4943 9308 4977 9342
rect 5015 9308 5049 9342
rect 5087 9308 5121 9342
rect 5159 9308 5193 9342
rect 5231 9308 5265 9342
rect 5303 9308 5337 9342
rect 5375 9308 5409 9342
rect 5447 9308 5481 9342
rect 5519 9308 5553 9342
rect 5591 9308 5625 9342
rect 5663 9308 5697 9342
rect 5735 9308 5769 9342
rect 5807 9308 5841 9342
rect 5879 9308 5913 9342
rect 5951 9308 5985 9342
rect 6023 9308 6057 9342
rect 6095 9308 6129 9342
rect 6167 9308 6201 9342
rect 6239 9308 6273 9342
rect 6311 9308 6345 9342
rect 6383 9308 6417 9342
rect 6455 9308 6489 9342
rect 6527 9308 6561 9342
rect 6599 9308 6633 9342
rect 6671 9308 6705 9342
rect 6743 9308 6777 9342
rect 6815 9308 6849 9342
rect 6887 9308 6921 9342
rect 6959 9308 6993 9342
rect 7031 9308 7065 9342
rect 7103 9308 7137 9342
rect 7175 9308 7209 9342
rect 7247 9308 7281 9342
rect 7319 9308 7353 9342
rect 7391 9308 7425 9342
rect 7463 9308 7497 9342
rect 7535 9308 7569 9342
rect 7607 9308 7641 9342
rect 7679 9308 7713 9342
rect 7751 9308 7785 9342
rect 7823 9308 7857 9342
rect 7895 9308 7929 9342
rect 7967 9308 8001 9342
rect 8039 9308 8073 9342
rect 8111 9308 8145 9342
rect 8183 9308 8217 9342
rect 8255 9308 8289 9342
rect 8327 9308 8361 9342
rect 8399 9308 8433 9342
rect 8471 9308 8505 9342
rect 8543 9308 8577 9342
rect 8615 9308 8649 9342
rect 8687 9308 8721 9342
rect 8759 9308 8793 9342
rect 8831 9308 8865 9342
rect 8903 9308 8937 9342
rect 8975 9308 9009 9342
rect 9047 9308 9081 9342
rect 9119 9308 9153 9342
rect 9191 9308 9225 9342
rect 9263 9308 9297 9342
rect 9335 9308 9369 9342
rect 9407 9308 9441 9342
rect 9479 9308 9513 9342
rect 9551 9308 9585 9342
rect 9623 9308 9657 9342
rect 9695 9308 9729 9342
rect 9767 9308 9801 9342
rect 9839 9308 9873 9342
rect 9911 9308 9945 9342
rect 9983 9308 10017 9342
rect 10055 9308 10089 9342
rect 10127 9308 10161 9342
rect 10199 9308 10233 9342
rect 10271 9308 10305 9342
rect 10343 9308 10377 9342
rect 10415 9308 10449 9342
rect 10487 9308 10521 9342
rect 10559 9308 10593 9342
rect 10631 9308 10665 9342
rect 10703 9308 10737 9342
rect 10775 9308 10809 9342
rect 10847 9308 10881 9342
rect 10919 9308 10953 9342
rect 10991 9308 11025 9342
rect 11063 9308 11097 9342
rect 11135 9308 11169 9342
rect 11207 9308 11241 9342
rect 11279 9308 11313 9342
rect 11351 9308 11385 9342
rect 11423 9308 11457 9342
rect 11495 9308 11529 9342
rect 11567 9308 11601 9342
rect 11639 9308 11673 9342
rect 11711 9308 11745 9342
rect 11783 9308 11817 9342
rect 11855 9308 11889 9342
rect 11927 9308 11961 9342
rect 11999 9308 12033 9342
rect 12071 9308 12105 9342
rect 12143 9308 12177 9342
rect 12215 9308 12249 9342
rect 12287 9308 12321 9342
rect 12359 9308 12393 9342
rect 12431 9308 12465 9342
rect 12503 9308 12537 9342
rect 12575 9308 12609 9342
rect 12647 9308 12681 9342
rect 12719 9308 12753 9342
rect 12791 9308 12825 9342
rect 12863 9308 12897 9342
rect 12935 9308 12969 9342
rect 13007 9308 13041 9342
rect 13079 9308 13113 9342
rect 13151 9308 13185 9342
rect 13223 9308 13257 9342
rect 13295 9308 13329 9342
rect 13367 9308 13401 9342
rect 13439 9308 13473 9342
rect 13511 9308 13545 9342
rect 13583 9308 13617 9342
rect 13655 9308 13689 9342
rect 13727 9308 13761 9342
rect 13799 9308 13833 9342
rect -484 9238 -482 9256
rect -482 9238 -450 9256
rect -411 9238 -378 9256
rect -378 9238 -377 9256
rect -338 9238 -309 9256
rect -309 9238 -304 9256
rect -265 9238 -240 9256
rect -240 9238 -231 9256
rect -192 9238 -171 9256
rect -171 9238 -158 9256
rect -119 9238 -102 9256
rect -102 9238 -85 9256
rect -484 9222 -450 9238
rect -411 9222 -377 9238
rect -338 9222 -304 9238
rect -265 9222 -231 9238
rect -192 9222 -158 9238
rect -119 9222 -85 9238
rect -46 9222 -33 9256
rect -33 9222 -12 9256
rect 27 9222 61 9256
rect 100 9222 134 9256
rect 173 9222 207 9256
rect 246 9222 280 9256
rect 319 9222 353 9256
rect 392 9222 426 9256
rect 465 9222 499 9256
rect 538 9222 572 9256
rect 611 9222 645 9256
rect 684 9222 718 9256
rect 757 9222 791 9256
rect 830 9222 864 9256
rect 903 9222 937 9256
rect 976 9222 1010 9256
rect 1049 9222 1083 9256
rect 1122 9222 1156 9256
rect 1195 9222 1229 9256
rect 1268 9222 1302 9256
rect 1341 9222 1375 9256
rect 1414 9222 1448 9256
rect 1487 9222 1521 9256
rect 1559 9222 1593 9256
rect 1631 9222 1665 9256
rect 1703 9222 1737 9256
rect 1775 9222 1809 9256
rect 1847 9222 1881 9256
rect 1919 9222 1953 9256
rect 1991 9222 2025 9256
rect 2063 9222 2097 9256
rect 2135 9222 2169 9256
rect 2207 9222 2241 9256
rect 2279 9222 2313 9256
rect 2351 9222 2385 9256
rect 2423 9222 2457 9256
rect 2495 9222 2529 9256
rect 2567 9222 2601 9256
rect 2639 9222 2673 9256
rect 2711 9222 2745 9256
rect 2783 9222 2817 9256
rect 2855 9222 2889 9256
rect 2927 9222 2961 9256
rect 2999 9222 3033 9256
rect 3071 9222 3105 9256
rect 3143 9222 3177 9256
rect 3215 9222 3249 9256
rect 3287 9222 3321 9256
rect 3359 9222 3393 9256
rect 3431 9222 3465 9256
rect 3503 9222 3537 9256
rect 3575 9222 3609 9256
rect 3647 9222 3681 9256
rect 3719 9222 3753 9256
rect 3791 9222 3825 9256
rect 3863 9222 3897 9256
rect 3935 9222 3969 9256
rect 4007 9222 4041 9256
rect 4079 9222 4113 9256
rect 4151 9222 4185 9256
rect 4223 9222 4257 9256
rect 4295 9222 4329 9256
rect 4367 9222 4401 9256
rect 4439 9222 4473 9256
rect 4511 9222 4545 9256
rect 4583 9222 4617 9256
rect 4655 9222 4689 9256
rect 4727 9222 4761 9256
rect 4799 9222 4833 9256
rect 4871 9222 4905 9256
rect 4943 9222 4977 9256
rect 5015 9222 5049 9256
rect 5087 9222 5121 9256
rect 5159 9222 5193 9256
rect 5231 9222 5265 9256
rect 5303 9222 5337 9256
rect 5375 9222 5409 9256
rect 5447 9222 5481 9256
rect 5519 9222 5553 9256
rect 5591 9222 5625 9256
rect 5663 9222 5697 9256
rect 5735 9222 5769 9256
rect 5807 9222 5841 9256
rect 5879 9222 5913 9256
rect 5951 9222 5985 9256
rect 6023 9222 6057 9256
rect 6095 9222 6129 9256
rect 6167 9222 6201 9256
rect 6239 9222 6273 9256
rect 6311 9222 6345 9256
rect 6383 9222 6417 9256
rect 6455 9222 6489 9256
rect 6527 9222 6561 9256
rect 6599 9222 6633 9256
rect 6671 9222 6705 9256
rect 6743 9222 6777 9256
rect 6815 9222 6849 9256
rect 6887 9222 6921 9256
rect 6959 9222 6993 9256
rect 7031 9222 7065 9256
rect 7103 9222 7137 9256
rect 7175 9222 7209 9256
rect 7247 9222 7281 9256
rect 7319 9222 7353 9256
rect 7391 9222 7425 9256
rect 7463 9222 7497 9256
rect 7535 9222 7569 9256
rect 7607 9222 7641 9256
rect 7679 9222 7713 9256
rect 7751 9222 7785 9256
rect 7823 9222 7857 9256
rect 7895 9222 7929 9256
rect 7967 9222 8001 9256
rect 8039 9222 8073 9256
rect 8111 9222 8145 9256
rect 8183 9222 8217 9256
rect 8255 9222 8289 9256
rect 8327 9222 8361 9256
rect 8399 9222 8433 9256
rect 8471 9222 8505 9256
rect 8543 9222 8577 9256
rect 8615 9222 8649 9256
rect 8687 9222 8721 9256
rect 8759 9222 8793 9256
rect 8831 9222 8865 9256
rect 8903 9222 8937 9256
rect 8975 9222 9009 9256
rect 9047 9222 9081 9256
rect 9119 9222 9153 9256
rect 9191 9222 9225 9256
rect 9263 9222 9297 9256
rect 9335 9222 9369 9256
rect 9407 9222 9441 9256
rect 9479 9222 9513 9256
rect 9551 9222 9585 9256
rect 9623 9222 9657 9256
rect 9695 9222 9729 9256
rect 9767 9222 9801 9256
rect 9839 9222 9873 9256
rect 9911 9222 9945 9256
rect 9983 9222 10017 9256
rect 10055 9222 10089 9256
rect 10127 9222 10161 9256
rect 10199 9222 10233 9256
rect 10271 9222 10305 9256
rect 10343 9222 10377 9256
rect 10415 9222 10449 9256
rect 10487 9222 10521 9256
rect 10559 9222 10593 9256
rect 10631 9222 10665 9256
rect 10703 9222 10737 9256
rect 10775 9222 10809 9256
rect 10847 9222 10881 9256
rect 10919 9222 10953 9256
rect 10991 9222 11025 9256
rect 11063 9222 11097 9256
rect 11135 9222 11169 9256
rect 11207 9222 11241 9256
rect 11279 9222 11313 9256
rect 11351 9222 11385 9256
rect 11423 9222 11457 9256
rect 11495 9222 11529 9256
rect 11567 9222 11601 9256
rect 11639 9222 11673 9256
rect 11711 9222 11745 9256
rect 11783 9222 11817 9256
rect 11855 9222 11889 9256
rect 11927 9222 11961 9256
rect 11999 9222 12033 9256
rect 12071 9222 12105 9256
rect 12143 9222 12177 9256
rect 12215 9222 12249 9256
rect 12287 9222 12321 9256
rect 12359 9222 12393 9256
rect 12431 9222 12465 9256
rect 12503 9222 12537 9256
rect 12575 9222 12609 9256
rect 12647 9222 12681 9256
rect 12719 9222 12753 9256
rect 12791 9222 12825 9256
rect 12863 9222 12897 9256
rect 12935 9222 12969 9256
rect 13007 9222 13041 9256
rect 13079 9222 13113 9256
rect 13151 9222 13185 9256
rect 13223 9222 13257 9256
rect 13295 9222 13329 9256
rect 13367 9222 13401 9256
rect 13439 9222 13473 9256
rect 13511 9222 13545 9256
rect 13583 9222 13617 9256
rect 13655 9222 13689 9256
rect 13727 9222 13761 9256
rect 13799 9222 13833 9256
rect -484 9136 -450 9170
rect -411 9136 -377 9170
rect -338 9136 -304 9170
rect -265 9136 -231 9170
rect -192 9136 -158 9170
rect -119 9136 -85 9170
rect -46 9136 -33 9170
rect -33 9136 -12 9170
rect 27 9136 61 9170
rect 100 9136 134 9170
rect 173 9136 207 9170
rect 246 9136 280 9170
rect 319 9136 353 9170
rect 392 9136 426 9170
rect 465 9136 499 9170
rect 538 9136 572 9170
rect 611 9136 645 9170
rect 684 9136 718 9170
rect 757 9136 791 9170
rect 830 9136 864 9170
rect 903 9136 937 9170
rect 976 9136 1010 9170
rect 1049 9136 1083 9170
rect 1122 9136 1156 9170
rect 1195 9136 1229 9170
rect 1268 9136 1302 9170
rect 1341 9136 1375 9170
rect 1414 9136 1448 9170
rect 1487 9136 1521 9170
rect 1559 9136 1593 9170
rect 1631 9136 1665 9170
rect 1703 9136 1737 9170
rect 1775 9136 1809 9170
rect 1847 9136 1881 9170
rect 1919 9136 1953 9170
rect 1991 9136 2025 9170
rect 2063 9136 2097 9170
rect 2135 9136 2169 9170
rect 2207 9136 2241 9170
rect 2279 9136 2313 9170
rect 2351 9136 2385 9170
rect 2423 9136 2457 9170
rect 2495 9136 2529 9170
rect 2567 9136 2601 9170
rect 2639 9136 2673 9170
rect 2711 9136 2745 9170
rect 2783 9136 2817 9170
rect 2855 9136 2889 9170
rect 2927 9136 2961 9170
rect 2999 9136 3033 9170
rect 3071 9136 3105 9170
rect 3143 9136 3177 9170
rect 3215 9136 3249 9170
rect 3287 9136 3321 9170
rect 3359 9136 3393 9170
rect 3431 9136 3465 9170
rect 3503 9136 3537 9170
rect 3575 9136 3609 9170
rect 3647 9136 3681 9170
rect 3719 9136 3753 9170
rect 3791 9136 3825 9170
rect 3863 9136 3897 9170
rect 3935 9136 3969 9170
rect 4007 9136 4041 9170
rect 4079 9136 4113 9170
rect 4151 9136 4185 9170
rect 4223 9136 4257 9170
rect 4295 9136 4329 9170
rect 4367 9136 4401 9170
rect 4439 9136 4473 9170
rect 4511 9136 4545 9170
rect 4583 9136 4617 9170
rect 4655 9136 4689 9170
rect 4727 9136 4761 9170
rect 4799 9136 4833 9170
rect 4871 9136 4905 9170
rect 4943 9136 4977 9170
rect 5015 9136 5049 9170
rect 5087 9136 5121 9170
rect 5159 9136 5193 9170
rect 5231 9136 5265 9170
rect 5303 9136 5337 9170
rect 5375 9136 5409 9170
rect 5447 9136 5481 9170
rect 5519 9136 5553 9170
rect 5591 9136 5625 9170
rect 5663 9136 5697 9170
rect 5735 9136 5769 9170
rect 5807 9136 5841 9170
rect 5879 9136 5913 9170
rect 5951 9136 5985 9170
rect 6023 9136 6057 9170
rect 6095 9136 6129 9170
rect 6167 9136 6201 9170
rect 6239 9136 6273 9170
rect 6311 9136 6345 9170
rect 6383 9136 6417 9170
rect 6455 9136 6489 9170
rect 6527 9136 6561 9170
rect 6599 9136 6633 9170
rect 6671 9136 6705 9170
rect 6743 9136 6777 9170
rect 6815 9136 6849 9170
rect 6887 9136 6921 9170
rect 6959 9136 6993 9170
rect 7031 9136 7065 9170
rect 7103 9136 7137 9170
rect 7175 9136 7209 9170
rect 7247 9136 7281 9170
rect 7319 9136 7353 9170
rect 7391 9136 7425 9170
rect 7463 9136 7497 9170
rect 7535 9136 7569 9170
rect 7607 9136 7641 9170
rect 7679 9136 7713 9170
rect 7751 9136 7785 9170
rect 7823 9136 7857 9170
rect 7895 9136 7929 9170
rect 7967 9136 8001 9170
rect 8039 9136 8073 9170
rect 8111 9136 8145 9170
rect 8183 9136 8217 9170
rect 8255 9136 8289 9170
rect 8327 9136 8361 9170
rect 8399 9136 8433 9170
rect 8471 9136 8505 9170
rect 8543 9136 8577 9170
rect 8615 9136 8649 9170
rect 8687 9136 8721 9170
rect 8759 9136 8793 9170
rect 8831 9136 8865 9170
rect 8903 9136 8937 9170
rect 8975 9136 9009 9170
rect 9047 9136 9081 9170
rect 9119 9136 9153 9170
rect 9191 9136 9225 9170
rect 9263 9136 9297 9170
rect 9335 9136 9369 9170
rect 9407 9136 9441 9170
rect 9479 9136 9513 9170
rect 9551 9136 9585 9170
rect 9623 9136 9657 9170
rect 9695 9136 9729 9170
rect 9767 9136 9801 9170
rect 9839 9136 9873 9170
rect 9911 9136 9945 9170
rect 9983 9136 10017 9170
rect 10055 9136 10089 9170
rect 10127 9136 10161 9170
rect 10199 9136 10233 9170
rect 10271 9136 10305 9170
rect 10343 9136 10377 9170
rect 10415 9136 10449 9170
rect 10487 9136 10521 9170
rect 10559 9136 10593 9170
rect 10631 9136 10665 9170
rect 10703 9136 10737 9170
rect 10775 9136 10809 9170
rect 10847 9136 10881 9170
rect 10919 9136 10953 9170
rect 10991 9136 11025 9170
rect 11063 9136 11097 9170
rect 11135 9136 11169 9170
rect 11207 9136 11241 9170
rect 11279 9136 11313 9170
rect 11351 9136 11385 9170
rect 11423 9136 11457 9170
rect 11495 9136 11529 9170
rect 11567 9136 11601 9170
rect 11639 9136 11673 9170
rect 11711 9136 11745 9170
rect 11783 9136 11817 9170
rect 11855 9136 11889 9170
rect 11927 9136 11961 9170
rect 11999 9136 12033 9170
rect 12071 9136 12105 9170
rect 12143 9136 12177 9170
rect 12215 9136 12249 9170
rect 12287 9136 12321 9170
rect 12359 9136 12393 9170
rect 12431 9136 12465 9170
rect 12503 9136 12537 9170
rect 12575 9136 12609 9170
rect 12647 9136 12681 9170
rect 12719 9136 12753 9170
rect 12791 9136 12825 9170
rect 12863 9136 12897 9170
rect 12935 9136 12969 9170
rect 13007 9136 13041 9170
rect 13079 9136 13113 9170
rect 13151 9136 13185 9170
rect 13223 9136 13257 9170
rect 13295 9136 13329 9170
rect 13367 9136 13401 9170
rect 13439 9136 13473 9170
rect 13511 9136 13545 9170
rect 13583 9136 13617 9170
rect 13655 9136 13689 9170
rect 13727 9136 13761 9170
rect 13799 9136 13833 9170
rect 248 8740 278 8753
rect 278 8740 282 8753
rect 322 8740 348 8753
rect 348 8740 356 8753
rect 396 8740 418 8753
rect 418 8740 430 8753
rect 470 8740 488 8753
rect 488 8740 504 8753
rect 544 8740 558 8753
rect 558 8740 578 8753
rect 618 8740 628 8753
rect 628 8740 652 8753
rect 691 8740 698 8753
rect 698 8740 725 8753
rect 764 8740 768 8753
rect 768 8740 798 8753
rect 837 8740 838 8753
rect 838 8740 871 8753
rect 912 8740 942 8760
rect 942 8740 946 8760
rect 984 8740 1012 8760
rect 1012 8740 1018 8760
rect 1056 8740 1082 8760
rect 1082 8740 1090 8760
rect 1128 8740 1152 8760
rect 1152 8740 1162 8760
rect 1200 8740 1222 8760
rect 1222 8740 1234 8760
rect 1272 8740 1292 8760
rect 1292 8740 1306 8760
rect 1344 8740 1362 8760
rect 1362 8740 1378 8760
rect 1416 8740 1432 8760
rect 1432 8740 1450 8760
rect 1488 8740 1501 8760
rect 1501 8740 1522 8760
rect 1560 8740 1570 8760
rect 1570 8740 1594 8760
rect 1632 8740 1639 8760
rect 1639 8740 1666 8760
rect 1704 8740 1708 8760
rect 1708 8740 1738 8760
rect 1776 8740 1777 8760
rect 1777 8740 1810 8760
rect 1849 8740 1881 8760
rect 1881 8740 1883 8760
rect 1922 8740 1950 8760
rect 1950 8740 1956 8760
rect 1995 8740 2019 8760
rect 2019 8740 2029 8760
rect 2068 8740 2088 8760
rect 2088 8740 2102 8760
rect 2141 8740 2157 8760
rect 2157 8740 2175 8760
rect 2227 8740 2260 8753
rect 2260 8740 2261 8753
rect 2306 8740 2329 8753
rect 2329 8740 2340 8753
rect 2385 8740 2398 8753
rect 2398 8740 2419 8753
rect 2464 8740 2467 8753
rect 2467 8740 2498 8753
rect 2543 8740 2571 8753
rect 2571 8740 2577 8753
rect 2621 8740 2640 8753
rect 2640 8740 2655 8753
rect 2699 8740 2709 8753
rect 2709 8740 2733 8753
rect 2777 8740 2778 8753
rect 2778 8740 2811 8753
rect 2855 8740 2881 8753
rect 2881 8740 2889 8753
rect 248 8719 282 8740
rect 322 8719 356 8740
rect 396 8719 430 8740
rect 470 8719 504 8740
rect 544 8719 578 8740
rect 618 8719 652 8740
rect 691 8719 725 8740
rect 764 8719 798 8740
rect 837 8719 871 8740
rect 912 8726 946 8740
rect 984 8726 1018 8740
rect 1056 8726 1090 8740
rect 1128 8726 1162 8740
rect 1200 8726 1234 8740
rect 1272 8726 1306 8740
rect 1344 8726 1378 8740
rect 1416 8726 1450 8740
rect 1488 8726 1522 8740
rect 1560 8726 1594 8740
rect 1632 8726 1666 8740
rect 1704 8726 1738 8740
rect 1776 8726 1810 8740
rect 1849 8726 1883 8740
rect 1922 8726 1956 8740
rect 1995 8726 2029 8740
rect 2068 8726 2102 8740
rect 2141 8726 2175 8740
rect 2227 8719 2261 8740
rect 2306 8719 2340 8740
rect 2385 8719 2419 8740
rect 2464 8719 2498 8740
rect 2543 8719 2577 8740
rect 2621 8719 2655 8740
rect 2699 8719 2733 8740
rect 2777 8719 2811 8740
rect 2855 8719 2889 8740
rect 2933 8736 2967 8753
rect 3011 8736 3036 8753
rect 3036 8736 3045 8753
rect 3477 8736 3479 8760
rect 3479 8736 3511 8760
rect 3550 8736 3581 8760
rect 3581 8736 3584 8760
rect 3623 8736 3649 8760
rect 3649 8736 3657 8760
rect 3696 8736 3717 8760
rect 3717 8736 3730 8760
rect 3769 8736 3785 8760
rect 3785 8736 3803 8760
rect 3842 8736 3853 8760
rect 3853 8736 3876 8760
rect 3915 8736 3921 8760
rect 3921 8736 3949 8760
rect 3988 8736 3989 8760
rect 3989 8736 4022 8760
rect 4061 8736 4091 8760
rect 4091 8736 4095 8760
rect 4134 8736 4159 8760
rect 4159 8736 4168 8760
rect 4207 8736 4227 8760
rect 4227 8736 4241 8760
rect 4280 8736 4295 8760
rect 4295 8736 4314 8760
rect 4353 8736 4363 8760
rect 4363 8736 4387 8760
rect 4426 8736 4431 8760
rect 4431 8736 4460 8760
rect 4499 8736 4533 8760
rect 4572 8736 4601 8760
rect 4601 8736 4606 8760
rect 4645 8736 4669 8760
rect 4669 8736 4679 8760
rect 4718 8736 4737 8760
rect 4737 8736 4752 8760
rect 4791 8736 4805 8760
rect 4805 8736 4825 8760
rect 4864 8736 4873 8760
rect 4873 8736 4898 8760
rect 4937 8736 4941 8760
rect 4941 8736 4971 8760
rect 5010 8736 5043 8760
rect 5043 8736 5044 8760
rect 5083 8736 5111 8760
rect 5111 8736 5117 8760
rect 5156 8736 5179 8760
rect 5179 8736 5190 8760
rect 5229 8736 5247 8760
rect 5247 8736 5263 8760
rect 5302 8736 5315 8760
rect 5315 8736 5336 8760
rect 5375 8736 5383 8760
rect 5383 8736 5409 8760
rect 5448 8736 5451 8760
rect 5451 8736 5482 8760
rect 5521 8736 5553 8760
rect 5553 8736 5555 8760
rect 5594 8736 5621 8760
rect 5621 8736 5628 8760
rect 5667 8736 5689 8760
rect 5689 8736 5701 8760
rect 5740 8736 5757 8760
rect 5757 8736 5774 8760
rect 5813 8736 5825 8760
rect 5825 8736 5847 8760
rect 5886 8736 5893 8760
rect 5893 8736 5920 8760
rect 5959 8736 5961 8760
rect 5961 8736 5993 8760
rect 6032 8736 6063 8760
rect 6063 8736 6066 8760
rect 6105 8736 6131 8760
rect 6131 8736 6139 8760
rect 6178 8736 6199 8760
rect 6199 8736 6212 8760
rect 6251 8736 6267 8760
rect 6267 8736 6285 8760
rect 6324 8736 6335 8760
rect 6335 8736 6358 8760
rect 6397 8736 6403 8760
rect 6403 8736 6431 8760
rect 6470 8736 6471 8760
rect 6471 8736 6504 8760
rect 6543 8736 6573 8760
rect 6573 8736 6577 8760
rect 6616 8736 6641 8760
rect 6641 8736 6650 8760
rect 6689 8736 6709 8760
rect 6709 8736 6723 8760
rect 6762 8736 6777 8760
rect 6777 8736 6796 8760
rect 6835 8736 6845 8760
rect 6845 8736 6869 8760
rect 6908 8736 6913 8760
rect 6913 8736 6942 8760
rect 2933 8719 2967 8736
rect 3011 8719 3045 8736
rect 3477 8726 3511 8736
rect 3550 8726 3584 8736
rect 3623 8726 3657 8736
rect 3696 8726 3730 8736
rect 3769 8726 3803 8736
rect 3842 8726 3876 8736
rect 3915 8726 3949 8736
rect 3988 8726 4022 8736
rect 4061 8726 4095 8736
rect 4134 8726 4168 8736
rect 4207 8726 4241 8736
rect 4280 8726 4314 8736
rect 4353 8726 4387 8736
rect 4426 8726 4460 8736
rect 4499 8726 4533 8736
rect 4572 8726 4606 8736
rect 4645 8726 4679 8736
rect 4718 8726 4752 8736
rect 4791 8726 4825 8736
rect 4864 8726 4898 8736
rect 4937 8726 4971 8736
rect 5010 8726 5044 8736
rect 5083 8726 5117 8736
rect 5156 8726 5190 8736
rect 5229 8726 5263 8736
rect 5302 8726 5336 8736
rect 5375 8726 5409 8736
rect 5448 8726 5482 8736
rect 5521 8726 5555 8736
rect 5594 8726 5628 8736
rect 5667 8726 5701 8736
rect 5740 8726 5774 8736
rect 5813 8726 5847 8736
rect 5886 8726 5920 8736
rect 5959 8726 5993 8736
rect 6032 8726 6066 8736
rect 6105 8726 6139 8736
rect 6178 8726 6212 8736
rect 6251 8726 6285 8736
rect 6324 8726 6358 8736
rect 6397 8726 6431 8736
rect 6470 8726 6504 8736
rect 6543 8726 6577 8736
rect 6616 8726 6650 8736
rect 6689 8726 6723 8736
rect 6762 8726 6796 8736
rect 6835 8726 6869 8736
rect 6908 8726 6942 8736
rect 6981 8726 7015 8760
rect 7054 8736 7083 8760
rect 7083 8736 7088 8760
rect 7127 8736 7151 8760
rect 7151 8736 7161 8760
rect 7200 8736 7219 8760
rect 7219 8736 7234 8760
rect 7273 8736 7287 8760
rect 7287 8736 7307 8760
rect 7346 8736 7355 8760
rect 7355 8736 7380 8760
rect 7419 8736 7423 8760
rect 7423 8736 7453 8760
rect 7492 8736 7525 8760
rect 7525 8736 7526 8760
rect 7565 8736 7593 8760
rect 7593 8736 7599 8760
rect 7638 8736 7661 8760
rect 7661 8736 7672 8760
rect 7711 8736 7729 8760
rect 7729 8736 7745 8760
rect 7784 8736 7797 8760
rect 7797 8736 7818 8760
rect 7857 8736 7865 8760
rect 7865 8736 7891 8760
rect 7930 8736 7933 8760
rect 7933 8736 7964 8760
rect 8003 8736 8035 8760
rect 8035 8736 8037 8760
rect 8075 8736 8103 8760
rect 8103 8736 8109 8760
rect 8147 8736 8171 8760
rect 8171 8736 8181 8760
rect 8219 8736 8239 8760
rect 8239 8736 8253 8760
rect 8291 8736 8307 8760
rect 8307 8736 8325 8760
rect 8363 8739 8393 8760
rect 8393 8739 8397 8760
rect 8435 8739 8462 8760
rect 8462 8739 8469 8760
rect 8507 8739 8531 8760
rect 8531 8739 8541 8760
rect 8579 8739 8600 8760
rect 8600 8739 8613 8760
rect 8651 8739 8669 8760
rect 8669 8739 8685 8760
rect 8723 8739 8738 8760
rect 8738 8739 8757 8760
rect 8795 8739 8807 8760
rect 8807 8739 8829 8760
rect 8867 8739 8876 8760
rect 8876 8739 8901 8760
rect 8939 8739 8945 8760
rect 8945 8739 8973 8760
rect 9011 8739 9014 8760
rect 9014 8739 9045 8760
rect 9083 8739 9117 8760
rect 9155 8739 9186 8760
rect 9186 8739 9189 8760
rect 9227 8739 9254 8760
rect 9254 8739 9261 8760
rect 9299 8739 9322 8760
rect 9322 8739 9333 8760
rect 9371 8739 9390 8760
rect 9390 8739 9405 8760
rect 9443 8739 9458 8760
rect 9458 8739 9477 8760
rect 9515 8739 9526 8760
rect 9526 8739 9549 8760
rect 9587 8739 9594 8760
rect 9594 8739 9621 8760
rect 9659 8739 9662 8760
rect 9662 8739 9693 8760
rect 9731 8739 9764 8760
rect 9764 8739 9765 8760
rect 9803 8739 9832 8760
rect 9832 8739 9837 8760
rect 9875 8739 9900 8760
rect 9900 8739 9909 8760
rect 9947 8739 9968 8760
rect 9968 8739 9981 8760
rect 10019 8739 10036 8760
rect 10036 8739 10053 8760
rect 10091 8739 10104 8760
rect 10104 8739 10125 8760
rect 10163 8739 10172 8760
rect 10172 8739 10197 8760
rect 10235 8739 10240 8760
rect 10240 8739 10269 8760
rect 10307 8739 10308 8760
rect 10308 8739 10341 8760
rect 10379 8739 10410 8760
rect 10410 8739 10413 8760
rect 10451 8739 10478 8760
rect 10478 8739 10485 8760
rect 10523 8739 10546 8760
rect 10546 8739 10557 8760
rect 10595 8739 10614 8760
rect 10614 8739 10629 8760
rect 10667 8739 10682 8760
rect 10682 8739 10701 8760
rect 10739 8739 10750 8760
rect 10750 8739 10773 8760
rect 10811 8739 10818 8760
rect 10818 8739 10845 8760
rect 10883 8739 10886 8760
rect 10886 8739 10917 8760
rect 10955 8739 10988 8760
rect 10988 8739 10989 8760
rect 11027 8739 11056 8760
rect 11056 8739 11061 8760
rect 11099 8739 11124 8760
rect 11124 8739 11133 8760
rect 11171 8739 11192 8760
rect 11192 8739 11205 8760
rect 11243 8739 11260 8760
rect 11260 8739 11277 8760
rect 11315 8739 11328 8760
rect 11328 8739 11349 8760
rect 11387 8739 11396 8760
rect 11396 8739 11421 8760
rect 11459 8739 11464 8760
rect 11464 8739 11493 8760
rect 11531 8739 11532 8760
rect 11532 8739 11565 8760
rect 11603 8739 11634 8760
rect 11634 8739 11637 8760
rect 11675 8739 11702 8760
rect 11702 8739 11709 8760
rect 11747 8739 11770 8760
rect 11770 8739 11781 8760
rect 11819 8739 11838 8760
rect 11838 8739 11853 8760
rect 11891 8739 11906 8760
rect 11906 8739 11925 8760
rect 11963 8739 11974 8760
rect 11974 8739 11997 8760
rect 12035 8739 12042 8760
rect 12042 8739 12069 8760
rect 12107 8739 12110 8760
rect 12110 8739 12141 8760
rect 12179 8739 12212 8760
rect 12212 8739 12213 8760
rect 12251 8739 12280 8760
rect 12280 8739 12285 8760
rect 12323 8739 12348 8760
rect 12348 8739 12357 8760
rect 12395 8739 12416 8760
rect 12416 8739 12429 8760
rect 12467 8739 12484 8760
rect 12484 8739 12501 8760
rect 12539 8739 12552 8760
rect 12552 8739 12573 8760
rect 12611 8739 12620 8760
rect 12620 8739 12645 8760
rect 12683 8739 12688 8760
rect 12688 8739 12717 8760
rect 12755 8739 12756 8760
rect 12756 8739 12789 8760
rect 12827 8739 12858 8760
rect 12858 8739 12861 8760
rect 12899 8739 12926 8760
rect 12926 8739 12933 8760
rect 12971 8739 12994 8760
rect 12994 8739 13005 8760
rect 13043 8739 13062 8760
rect 13062 8739 13077 8760
rect 13115 8739 13130 8760
rect 13130 8739 13149 8760
rect 13187 8739 13198 8760
rect 13198 8739 13221 8760
rect 13259 8739 13266 8760
rect 13266 8739 13293 8760
rect 13331 8739 13334 8760
rect 13334 8739 13365 8760
rect 13403 8739 13436 8760
rect 13436 8739 13437 8760
rect 13475 8739 13504 8760
rect 13504 8739 13509 8760
rect 13547 8739 13572 8760
rect 13572 8739 13581 8760
rect 13619 8739 13640 8760
rect 13640 8739 13653 8760
rect 13691 8739 13708 8760
rect 13708 8739 13725 8760
rect 13763 8739 13776 8760
rect 13776 8739 13797 8760
rect 13835 8739 13844 8760
rect 13844 8739 13869 8760
rect 13907 8739 13912 8760
rect 13912 8739 13941 8760
rect 13979 8739 13980 8760
rect 13980 8739 14013 8760
rect 14051 8739 14082 8760
rect 14082 8739 14085 8760
rect 14123 8739 14150 8760
rect 14150 8739 14157 8760
rect 14195 8739 14218 8760
rect 14218 8739 14229 8760
rect 14267 8739 14286 8760
rect 14286 8739 14301 8760
rect 14339 8739 14354 8760
rect 14354 8739 14373 8760
rect 14411 8739 14422 8760
rect 14422 8739 14445 8760
rect 14483 8739 14490 8760
rect 14490 8739 14517 8760
rect 14555 8739 14558 8760
rect 14558 8739 14589 8760
rect 14627 8739 14660 8760
rect 14660 8739 14661 8760
rect 14699 8739 14728 8760
rect 14728 8739 14733 8760
rect 14771 8739 14796 8760
rect 14796 8739 14805 8760
rect 14843 8739 14864 8760
rect 14864 8739 14877 8760
rect 7054 8726 7088 8736
rect 7127 8726 7161 8736
rect 7200 8726 7234 8736
rect 7273 8726 7307 8736
rect 7346 8726 7380 8736
rect 7419 8726 7453 8736
rect 7492 8726 7526 8736
rect 7565 8726 7599 8736
rect 7638 8726 7672 8736
rect 7711 8726 7745 8736
rect 7784 8726 7818 8736
rect 7857 8726 7891 8736
rect 7930 8726 7964 8736
rect 8003 8726 8037 8736
rect 8075 8726 8109 8736
rect 8147 8726 8181 8736
rect 8219 8726 8253 8736
rect 8291 8726 8325 8736
rect 8363 8726 8397 8739
rect 8435 8726 8469 8739
rect 8507 8726 8541 8739
rect 8579 8726 8613 8739
rect 8651 8726 8685 8739
rect 8723 8726 8757 8739
rect 8795 8726 8829 8739
rect 8867 8726 8901 8739
rect 8939 8726 8973 8739
rect 9011 8726 9045 8739
rect 9083 8726 9117 8739
rect 9155 8726 9189 8739
rect 9227 8726 9261 8739
rect 9299 8726 9333 8739
rect 9371 8726 9405 8739
rect 9443 8726 9477 8739
rect 9515 8726 9549 8739
rect 9587 8726 9621 8739
rect 9659 8726 9693 8739
rect 9731 8726 9765 8739
rect 9803 8726 9837 8739
rect 9875 8726 9909 8739
rect 9947 8726 9981 8739
rect 10019 8726 10053 8739
rect 10091 8726 10125 8739
rect 10163 8726 10197 8739
rect 10235 8726 10269 8739
rect 10307 8726 10341 8739
rect 10379 8726 10413 8739
rect 10451 8726 10485 8739
rect 10523 8726 10557 8739
rect 10595 8726 10629 8739
rect 10667 8726 10701 8739
rect 10739 8726 10773 8739
rect 10811 8726 10845 8739
rect 10883 8726 10917 8739
rect 10955 8726 10989 8739
rect 11027 8726 11061 8739
rect 11099 8726 11133 8739
rect 11171 8726 11205 8739
rect 11243 8726 11277 8739
rect 11315 8726 11349 8739
rect 11387 8726 11421 8739
rect 11459 8726 11493 8739
rect 11531 8726 11565 8739
rect 11603 8726 11637 8739
rect 11675 8726 11709 8739
rect 11747 8726 11781 8739
rect 11819 8726 11853 8739
rect 11891 8726 11925 8739
rect 11963 8726 11997 8739
rect 12035 8726 12069 8739
rect 12107 8726 12141 8739
rect 12179 8726 12213 8739
rect 12251 8726 12285 8739
rect 12323 8726 12357 8739
rect 12395 8726 12429 8739
rect 12467 8726 12501 8739
rect 12539 8726 12573 8739
rect 12611 8726 12645 8739
rect 12683 8726 12717 8739
rect 12755 8726 12789 8739
rect 12827 8726 12861 8739
rect 12899 8726 12933 8739
rect 12971 8726 13005 8739
rect 13043 8726 13077 8739
rect 13115 8726 13149 8739
rect 13187 8726 13221 8739
rect 13259 8726 13293 8739
rect 13331 8726 13365 8739
rect 13403 8726 13437 8739
rect 13475 8726 13509 8739
rect 13547 8726 13581 8739
rect 13619 8726 13653 8739
rect 13691 8726 13725 8739
rect 13763 8726 13797 8739
rect 13835 8726 13869 8739
rect 13907 8726 13941 8739
rect 13979 8726 14013 8739
rect 14051 8726 14085 8739
rect 14123 8726 14157 8739
rect 14195 8726 14229 8739
rect 14267 8726 14301 8739
rect 14339 8726 14373 8739
rect 14411 8726 14445 8739
rect 14483 8726 14517 8739
rect 14555 8726 14589 8739
rect 14627 8726 14661 8739
rect 14699 8726 14733 8739
rect 14771 8726 14805 8739
rect 14843 8726 14877 8739
rect 912 8626 946 8636
rect 984 8626 1018 8636
rect 1056 8626 1090 8636
rect 1128 8626 1162 8636
rect 1200 8626 1234 8636
rect 1272 8626 1306 8636
rect 1344 8626 1378 8636
rect 1416 8626 1450 8636
rect 1488 8626 1522 8636
rect 1560 8626 1594 8636
rect 1632 8626 1666 8636
rect 1704 8626 1738 8636
rect 1776 8626 1810 8636
rect 1849 8626 1883 8636
rect 1922 8626 1956 8636
rect 1995 8626 2029 8636
rect 2068 8626 2102 8636
rect 2141 8626 2175 8636
rect 3477 8630 3511 8636
rect 3550 8630 3584 8636
rect 3623 8630 3657 8636
rect 3696 8630 3730 8636
rect 3769 8630 3803 8636
rect 3842 8630 3876 8636
rect 3915 8630 3949 8636
rect 3988 8630 4022 8636
rect 4061 8630 4095 8636
rect 4134 8630 4168 8636
rect 4207 8630 4241 8636
rect 4280 8630 4314 8636
rect 4353 8630 4387 8636
rect 4426 8630 4460 8636
rect 4499 8630 4533 8636
rect 4572 8630 4606 8636
rect 4645 8630 4679 8636
rect 4718 8630 4752 8636
rect 4791 8630 4825 8636
rect 4864 8630 4898 8636
rect 4937 8630 4971 8636
rect 5010 8630 5044 8636
rect 5083 8630 5117 8636
rect 5156 8630 5190 8636
rect 5229 8630 5263 8636
rect 5302 8630 5336 8636
rect 5375 8630 5409 8636
rect 5448 8630 5482 8636
rect 5521 8630 5555 8636
rect 5594 8630 5628 8636
rect 5667 8630 5701 8636
rect 5740 8630 5774 8636
rect 5813 8630 5847 8636
rect 5886 8630 5920 8636
rect 5959 8630 5993 8636
rect 6032 8630 6066 8636
rect 6105 8630 6139 8636
rect 6178 8630 6212 8636
rect 6251 8630 6285 8636
rect 6324 8630 6358 8636
rect 6397 8630 6431 8636
rect 6470 8630 6504 8636
rect 6543 8630 6577 8636
rect 6616 8630 6650 8636
rect 6689 8630 6723 8636
rect 6762 8630 6796 8636
rect 6835 8630 6869 8636
rect 6908 8630 6942 8636
rect 912 8602 942 8626
rect 942 8602 946 8626
rect 984 8602 1012 8626
rect 1012 8602 1018 8626
rect 1056 8602 1082 8626
rect 1082 8602 1090 8626
rect 1128 8602 1152 8626
rect 1152 8602 1162 8626
rect 1200 8602 1222 8626
rect 1222 8602 1234 8626
rect 1272 8602 1292 8626
rect 1292 8602 1306 8626
rect 1344 8602 1362 8626
rect 1362 8602 1378 8626
rect 1416 8602 1432 8626
rect 1432 8602 1450 8626
rect 1488 8602 1501 8626
rect 1501 8602 1522 8626
rect 1560 8602 1570 8626
rect 1570 8602 1594 8626
rect 1632 8602 1639 8626
rect 1639 8602 1666 8626
rect 1704 8602 1708 8626
rect 1708 8602 1738 8626
rect 1776 8602 1777 8626
rect 1777 8602 1810 8626
rect 1849 8602 1881 8626
rect 1881 8602 1883 8626
rect 1922 8602 1950 8626
rect 1950 8602 1956 8626
rect 1995 8602 2019 8626
rect 2019 8602 2029 8626
rect 2068 8602 2088 8626
rect 2088 8602 2102 8626
rect 2141 8602 2157 8626
rect 2157 8602 2175 8626
rect 3477 8602 3479 8630
rect 3479 8602 3511 8630
rect 3550 8602 3581 8630
rect 3581 8602 3584 8630
rect 3623 8602 3649 8630
rect 3649 8602 3657 8630
rect 3696 8602 3717 8630
rect 3717 8602 3730 8630
rect 3769 8602 3785 8630
rect 3785 8602 3803 8630
rect 3842 8602 3853 8630
rect 3853 8602 3876 8630
rect 3915 8602 3921 8630
rect 3921 8602 3949 8630
rect 3988 8602 3989 8630
rect 3989 8602 4022 8630
rect 4061 8602 4091 8630
rect 4091 8602 4095 8630
rect 4134 8602 4159 8630
rect 4159 8602 4168 8630
rect 4207 8602 4227 8630
rect 4227 8602 4241 8630
rect 4280 8602 4295 8630
rect 4295 8602 4314 8630
rect 4353 8602 4363 8630
rect 4363 8602 4387 8630
rect 4426 8602 4431 8630
rect 4431 8602 4460 8630
rect 4499 8602 4533 8630
rect 4572 8602 4601 8630
rect 4601 8602 4606 8630
rect 4645 8602 4669 8630
rect 4669 8602 4679 8630
rect 4718 8602 4737 8630
rect 4737 8602 4752 8630
rect 4791 8602 4805 8630
rect 4805 8602 4825 8630
rect 4864 8602 4873 8630
rect 4873 8602 4898 8630
rect 4937 8602 4941 8630
rect 4941 8602 4971 8630
rect 5010 8602 5043 8630
rect 5043 8602 5044 8630
rect 5083 8602 5111 8630
rect 5111 8602 5117 8630
rect 5156 8602 5179 8630
rect 5179 8602 5190 8630
rect 5229 8602 5247 8630
rect 5247 8602 5263 8630
rect 5302 8602 5315 8630
rect 5315 8602 5336 8630
rect 5375 8602 5383 8630
rect 5383 8602 5409 8630
rect 5448 8602 5451 8630
rect 5451 8602 5482 8630
rect 5521 8602 5553 8630
rect 5553 8602 5555 8630
rect 5594 8602 5621 8630
rect 5621 8602 5628 8630
rect 5667 8602 5689 8630
rect 5689 8602 5701 8630
rect 5740 8602 5757 8630
rect 5757 8602 5774 8630
rect 5813 8602 5825 8630
rect 5825 8602 5847 8630
rect 5886 8602 5893 8630
rect 5893 8602 5920 8630
rect 5959 8602 5961 8630
rect 5961 8602 5993 8630
rect 6032 8602 6063 8630
rect 6063 8602 6066 8630
rect 6105 8602 6131 8630
rect 6131 8602 6139 8630
rect 6178 8602 6199 8630
rect 6199 8602 6212 8630
rect 6251 8602 6267 8630
rect 6267 8602 6285 8630
rect 6324 8602 6335 8630
rect 6335 8602 6358 8630
rect 6397 8602 6403 8630
rect 6403 8602 6431 8630
rect 6470 8602 6471 8630
rect 6471 8602 6504 8630
rect 6543 8602 6573 8630
rect 6573 8602 6577 8630
rect 6616 8602 6641 8630
rect 6641 8602 6650 8630
rect 6689 8602 6709 8630
rect 6709 8602 6723 8630
rect 6762 8602 6777 8630
rect 6777 8602 6796 8630
rect 6835 8602 6845 8630
rect 6845 8602 6869 8630
rect 6908 8602 6913 8630
rect 6913 8602 6942 8630
rect 6981 8602 7015 8636
rect 7054 8630 7088 8636
rect 7127 8630 7161 8636
rect 7200 8630 7234 8636
rect 7273 8630 7307 8636
rect 7346 8630 7380 8636
rect 7419 8630 7453 8636
rect 7492 8630 7526 8636
rect 7565 8630 7599 8636
rect 7638 8630 7672 8636
rect 7711 8630 7745 8636
rect 7784 8630 7818 8636
rect 7857 8630 7891 8636
rect 7930 8630 7964 8636
rect 8003 8630 8037 8636
rect 8075 8630 8109 8636
rect 8147 8630 8181 8636
rect 8219 8630 8253 8636
rect 8291 8630 8325 8636
rect 7054 8602 7083 8630
rect 7083 8602 7088 8630
rect 7127 8602 7151 8630
rect 7151 8602 7161 8630
rect 7200 8602 7219 8630
rect 7219 8602 7234 8630
rect 7273 8602 7287 8630
rect 7287 8602 7307 8630
rect 7346 8602 7355 8630
rect 7355 8602 7380 8630
rect 7419 8602 7423 8630
rect 7423 8602 7453 8630
rect 7492 8602 7525 8630
rect 7525 8602 7526 8630
rect 7565 8602 7593 8630
rect 7593 8602 7599 8630
rect 7638 8602 7661 8630
rect 7661 8602 7672 8630
rect 7711 8602 7729 8630
rect 7729 8602 7745 8630
rect 7784 8602 7797 8630
rect 7797 8602 7818 8630
rect 7857 8602 7865 8630
rect 7865 8602 7891 8630
rect 7930 8602 7933 8630
rect 7933 8602 7964 8630
rect 8003 8602 8035 8630
rect 8035 8602 8037 8630
rect 8075 8602 8103 8630
rect 8103 8602 8109 8630
rect 8147 8602 8171 8630
rect 8171 8602 8181 8630
rect 8219 8602 8239 8630
rect 8239 8602 8253 8630
rect 8291 8602 8307 8630
rect 8307 8602 8325 8630
rect 8363 8613 8397 8636
rect 8435 8613 8469 8636
rect 8507 8613 8541 8636
rect 8579 8613 8613 8636
rect 8651 8613 8685 8636
rect 8723 8613 8757 8636
rect 8795 8613 8829 8636
rect 8867 8613 8901 8636
rect 8939 8613 8973 8636
rect 9011 8613 9045 8636
rect 9083 8613 9117 8636
rect 9155 8613 9189 8636
rect 9227 8613 9261 8636
rect 9299 8613 9333 8636
rect 9371 8613 9405 8636
rect 9443 8613 9477 8636
rect 9515 8613 9549 8636
rect 9587 8613 9621 8636
rect 9659 8613 9693 8636
rect 9731 8613 9765 8636
rect 9803 8613 9837 8636
rect 9875 8613 9909 8636
rect 9947 8613 9981 8636
rect 10019 8613 10053 8636
rect 10091 8613 10125 8636
rect 10163 8613 10197 8636
rect 10235 8613 10269 8636
rect 10307 8613 10341 8636
rect 10379 8613 10413 8636
rect 10451 8613 10485 8636
rect 10523 8613 10557 8636
rect 10595 8613 10629 8636
rect 10667 8613 10701 8636
rect 10739 8613 10773 8636
rect 10811 8613 10845 8636
rect 10883 8613 10917 8636
rect 10955 8613 10989 8636
rect 11027 8613 11061 8636
rect 11099 8613 11133 8636
rect 11171 8613 11205 8636
rect 11243 8613 11277 8636
rect 11315 8613 11349 8636
rect 11387 8613 11421 8636
rect 11459 8613 11493 8636
rect 11531 8613 11565 8636
rect 11603 8613 11637 8636
rect 11675 8613 11709 8636
rect 11747 8613 11781 8636
rect 11819 8613 11853 8636
rect 11891 8613 11925 8636
rect 11963 8613 11997 8636
rect 12035 8613 12069 8636
rect 12107 8613 12141 8636
rect 12179 8613 12213 8636
rect 12251 8613 12285 8636
rect 12323 8613 12357 8636
rect 12395 8613 12429 8636
rect 12467 8613 12501 8636
rect 12539 8613 12573 8636
rect 12611 8613 12645 8636
rect 12683 8613 12717 8636
rect 12755 8613 12789 8636
rect 12827 8613 12861 8636
rect 12899 8613 12933 8636
rect 12971 8613 13005 8636
rect 13043 8613 13077 8636
rect 13115 8613 13149 8636
rect 13187 8613 13221 8636
rect 13259 8613 13293 8636
rect 13331 8613 13365 8636
rect 13403 8613 13437 8636
rect 13475 8613 13509 8636
rect 13547 8613 13581 8636
rect 13619 8613 13653 8636
rect 13691 8613 13725 8636
rect 13763 8613 13797 8636
rect 13835 8613 13869 8636
rect 13907 8613 13941 8636
rect 13979 8613 14013 8636
rect 14051 8613 14085 8636
rect 14123 8613 14157 8636
rect 14195 8613 14229 8636
rect 14267 8613 14301 8636
rect 14339 8613 14373 8636
rect 14411 8613 14445 8636
rect 14483 8613 14517 8636
rect 14555 8613 14589 8636
rect 14627 8613 14661 8636
rect 14699 8613 14733 8636
rect 14771 8613 14805 8636
rect 14843 8613 14877 8636
rect 8363 8602 8393 8613
rect 8393 8602 8397 8613
rect 8435 8602 8462 8613
rect 8462 8602 8469 8613
rect 8507 8602 8531 8613
rect 8531 8602 8541 8613
rect 8579 8602 8600 8613
rect 8600 8602 8613 8613
rect 8651 8602 8669 8613
rect 8669 8602 8685 8613
rect 8723 8602 8738 8613
rect 8738 8602 8757 8613
rect 8795 8602 8807 8613
rect 8807 8602 8829 8613
rect 8867 8602 8876 8613
rect 8876 8602 8901 8613
rect 8939 8602 8945 8613
rect 8945 8602 8973 8613
rect 9011 8602 9014 8613
rect 9014 8602 9045 8613
rect 9083 8602 9117 8613
rect 9155 8602 9186 8613
rect 9186 8602 9189 8613
rect 9227 8602 9254 8613
rect 9254 8602 9261 8613
rect 9299 8602 9322 8613
rect 9322 8602 9333 8613
rect 9371 8602 9390 8613
rect 9390 8602 9405 8613
rect 9443 8602 9458 8613
rect 9458 8602 9477 8613
rect 9515 8602 9526 8613
rect 9526 8602 9549 8613
rect 9587 8602 9594 8613
rect 9594 8602 9621 8613
rect 9659 8602 9662 8613
rect 9662 8602 9693 8613
rect 9731 8602 9764 8613
rect 9764 8602 9765 8613
rect 9803 8602 9832 8613
rect 9832 8602 9837 8613
rect 9875 8602 9900 8613
rect 9900 8602 9909 8613
rect 9947 8602 9968 8613
rect 9968 8602 9981 8613
rect 10019 8602 10036 8613
rect 10036 8602 10053 8613
rect 10091 8602 10104 8613
rect 10104 8602 10125 8613
rect 10163 8602 10172 8613
rect 10172 8602 10197 8613
rect 10235 8602 10240 8613
rect 10240 8602 10269 8613
rect 10307 8602 10308 8613
rect 10308 8602 10341 8613
rect 10379 8602 10410 8613
rect 10410 8602 10413 8613
rect 10451 8602 10478 8613
rect 10478 8602 10485 8613
rect 10523 8602 10546 8613
rect 10546 8602 10557 8613
rect 10595 8602 10614 8613
rect 10614 8602 10629 8613
rect 10667 8602 10682 8613
rect 10682 8602 10701 8613
rect 10739 8602 10750 8613
rect 10750 8602 10773 8613
rect 10811 8602 10818 8613
rect 10818 8602 10845 8613
rect 10883 8602 10886 8613
rect 10886 8602 10917 8613
rect 10955 8602 10988 8613
rect 10988 8602 10989 8613
rect 11027 8602 11056 8613
rect 11056 8602 11061 8613
rect 11099 8602 11124 8613
rect 11124 8602 11133 8613
rect 11171 8602 11192 8613
rect 11192 8602 11205 8613
rect 11243 8602 11260 8613
rect 11260 8602 11277 8613
rect 11315 8602 11328 8613
rect 11328 8602 11349 8613
rect 11387 8602 11396 8613
rect 11396 8602 11421 8613
rect 11459 8602 11464 8613
rect 11464 8602 11493 8613
rect 11531 8602 11532 8613
rect 11532 8602 11565 8613
rect 11603 8602 11634 8613
rect 11634 8602 11637 8613
rect 11675 8602 11702 8613
rect 11702 8602 11709 8613
rect 11747 8602 11770 8613
rect 11770 8602 11781 8613
rect 11819 8602 11838 8613
rect 11838 8602 11853 8613
rect 11891 8602 11906 8613
rect 11906 8602 11925 8613
rect 11963 8602 11974 8613
rect 11974 8602 11997 8613
rect 12035 8602 12042 8613
rect 12042 8602 12069 8613
rect 12107 8602 12110 8613
rect 12110 8602 12141 8613
rect 12179 8602 12212 8613
rect 12212 8602 12213 8613
rect 12251 8602 12280 8613
rect 12280 8602 12285 8613
rect 12323 8602 12348 8613
rect 12348 8602 12357 8613
rect 12395 8602 12416 8613
rect 12416 8602 12429 8613
rect 12467 8602 12484 8613
rect 12484 8602 12501 8613
rect 12539 8602 12552 8613
rect 12552 8602 12573 8613
rect 12611 8602 12620 8613
rect 12620 8602 12645 8613
rect 12683 8602 12688 8613
rect 12688 8602 12717 8613
rect 12755 8602 12756 8613
rect 12756 8602 12789 8613
rect 12827 8602 12858 8613
rect 12858 8602 12861 8613
rect 12899 8602 12926 8613
rect 12926 8602 12933 8613
rect 12971 8602 12994 8613
rect 12994 8602 13005 8613
rect 13043 8602 13062 8613
rect 13062 8602 13077 8613
rect 13115 8602 13130 8613
rect 13130 8602 13149 8613
rect 13187 8602 13198 8613
rect 13198 8602 13221 8613
rect 13259 8602 13266 8613
rect 13266 8602 13293 8613
rect 13331 8602 13334 8613
rect 13334 8602 13365 8613
rect 13403 8602 13436 8613
rect 13436 8602 13437 8613
rect 13475 8602 13504 8613
rect 13504 8602 13509 8613
rect 13547 8602 13572 8613
rect 13572 8602 13581 8613
rect 13619 8602 13640 8613
rect 13640 8602 13653 8613
rect 13691 8602 13708 8613
rect 13708 8602 13725 8613
rect 13763 8602 13776 8613
rect 13776 8602 13797 8613
rect 13835 8602 13844 8613
rect 13844 8602 13869 8613
rect 13907 8602 13912 8613
rect 13912 8602 13941 8613
rect 13979 8602 13980 8613
rect 13980 8602 14013 8613
rect 14051 8602 14082 8613
rect 14082 8602 14085 8613
rect 14123 8602 14150 8613
rect 14150 8602 14157 8613
rect 14195 8602 14218 8613
rect 14218 8602 14229 8613
rect 14267 8602 14286 8613
rect 14286 8602 14301 8613
rect 14339 8602 14354 8613
rect 14354 8602 14373 8613
rect 14411 8602 14422 8613
rect 14422 8602 14445 8613
rect 14483 8602 14490 8613
rect 14490 8602 14517 8613
rect 14555 8602 14558 8613
rect 14558 8602 14589 8613
rect 14627 8602 14660 8613
rect 14660 8602 14661 8613
rect 14699 8602 14728 8613
rect 14728 8602 14733 8613
rect 14771 8602 14796 8613
rect 14796 8602 14805 8613
rect 14843 8602 14864 8613
rect 14864 8602 14877 8613
rect 13992 8533 14026 8546
rect 14076 8533 14110 8546
rect 13992 8512 14014 8533
rect 14014 8512 14026 8533
rect 14076 8512 14082 8533
rect 14082 8512 14110 8533
rect 14185 8499 14218 8512
rect 14218 8499 14219 8512
rect 14257 8499 14286 8512
rect 14286 8499 14291 8512
rect 14329 8499 14354 8512
rect 14354 8499 14363 8512
rect 14401 8499 14422 8512
rect 14422 8499 14435 8512
rect 14473 8499 14490 8512
rect 14490 8499 14507 8512
rect 14185 8478 14219 8499
rect 14257 8478 14291 8499
rect 14329 8478 14363 8499
rect 14401 8478 14435 8499
rect 14473 8478 14507 8499
rect 13992 8453 14026 8474
rect 14076 8453 14110 8474
rect 14614 8453 14648 8462
rect 14692 8453 14726 8462
rect 14770 8453 14804 8462
rect 14848 8453 14882 8462
rect 13992 8440 14014 8453
rect 14014 8440 14026 8453
rect 14076 8440 14082 8453
rect 14082 8440 14110 8453
rect 14185 8419 14218 8435
rect 14218 8419 14219 8435
rect 14257 8419 14286 8435
rect 14286 8419 14291 8435
rect 14329 8419 14354 8435
rect 14354 8419 14363 8435
rect 14401 8419 14422 8435
rect 14422 8419 14435 8435
rect 14473 8419 14490 8435
rect 14490 8419 14507 8435
rect 14614 8428 14626 8453
rect 14626 8428 14648 8453
rect 14692 8428 14694 8453
rect 14694 8428 14726 8453
rect 14770 8428 14796 8453
rect 14796 8428 14804 8453
rect 14848 8428 14864 8453
rect 14864 8428 14882 8453
rect 14926 8433 14960 8462
rect 15004 8433 15038 8462
rect 14926 8428 14932 8433
rect 14932 8428 14960 8433
rect 14185 8401 14219 8419
rect 14257 8401 14291 8419
rect 14329 8401 14363 8419
rect 14401 8401 14435 8419
rect 14473 8401 14507 8419
rect 13992 8367 14026 8401
rect 14076 8367 14110 8401
rect 15004 8428 15034 8433
rect 15034 8428 15038 8433
rect 14185 8357 14219 8358
rect 14257 8357 14291 8358
rect 14329 8357 14363 8358
rect 14401 8357 14435 8358
rect 14473 8357 14507 8358
rect 14614 8357 14648 8388
rect 14692 8357 14726 8388
rect 14770 8357 14804 8388
rect 14848 8357 14882 8388
rect 14926 8361 14960 8388
rect 15004 8361 15038 8388
rect 14185 8324 14198 8357
rect 14198 8324 14219 8357
rect 14257 8324 14268 8357
rect 14268 8324 14291 8357
rect 14329 8324 14338 8357
rect 14338 8324 14363 8357
rect 14401 8324 14408 8357
rect 14408 8324 14435 8357
rect 14473 8324 14478 8357
rect 14478 8324 14507 8357
rect 14614 8354 14618 8357
rect 14618 8354 14648 8357
rect 14692 8354 14724 8357
rect 14724 8354 14726 8357
rect 14770 8354 14794 8357
rect 14794 8354 14804 8357
rect 14848 8354 14864 8357
rect 14864 8354 14882 8357
rect 14926 8354 14932 8361
rect 14932 8354 14960 8361
rect 15004 8354 15034 8361
rect 15034 8354 15038 8361
rect 14614 8283 14648 8314
rect 14692 8283 14726 8314
rect 14770 8283 14804 8314
rect 14848 8283 14882 8314
rect 14926 8289 14960 8314
rect 15004 8289 15038 8314
rect 8509 8239 8615 8254
rect 8509 7933 8510 8239
rect 8510 7933 8612 8239
rect 8612 7933 8615 8239
rect 8509 7932 8615 7933
rect 9596 8239 9630 8247
rect 9678 8239 9712 8247
rect 9596 8213 9612 8239
rect 9612 8213 9630 8239
rect 9678 8213 9712 8239
rect 9596 8110 9612 8144
rect 9612 8110 9630 8144
rect 9678 8110 9712 8144
rect 9596 8007 9612 8041
rect 9612 8007 9630 8041
rect 9678 8007 9712 8041
rect 10314 8239 10348 8247
rect 10396 8239 10430 8247
rect 10314 8213 10348 8239
rect 10396 8213 10416 8239
rect 10416 8213 10430 8239
rect 10314 8110 10348 8144
rect 10396 8110 10416 8144
rect 10416 8110 10430 8144
rect 10314 8007 10348 8041
rect 10396 8007 10416 8041
rect 10416 8007 10430 8041
rect 10804 8239 10838 8254
rect 10898 8239 10932 8254
rect 10804 8220 10816 8239
rect 10816 8220 10838 8239
rect 10898 8220 10918 8239
rect 10918 8220 10932 8239
rect 10804 8145 10816 8179
rect 10816 8145 10838 8179
rect 10898 8145 10918 8179
rect 10918 8145 10932 8179
rect 10804 8070 10816 8104
rect 10816 8070 10838 8104
rect 10898 8070 10918 8104
rect 10918 8070 10932 8104
rect 10804 7994 10816 8028
rect 10816 7994 10838 8028
rect 10898 7994 10918 8028
rect 10918 7994 10932 8028
rect 10804 7933 10816 7952
rect 10816 7933 10838 7952
rect 10898 7933 10918 7952
rect 10918 7933 10932 7952
rect 10804 7918 10838 7933
rect 10898 7918 10932 7933
rect 14185 8249 14198 8280
rect 14198 8249 14219 8280
rect 14257 8249 14268 8280
rect 14268 8249 14291 8280
rect 14329 8249 14338 8280
rect 14338 8249 14363 8280
rect 14401 8249 14408 8280
rect 14408 8249 14435 8280
rect 14473 8249 14478 8280
rect 14478 8249 14507 8280
rect 14614 8280 14618 8283
rect 14618 8280 14648 8283
rect 14692 8280 14724 8283
rect 14724 8280 14726 8283
rect 14770 8280 14794 8283
rect 14794 8280 14804 8283
rect 14848 8280 14864 8283
rect 14864 8280 14882 8283
rect 14926 8280 14932 8289
rect 14932 8280 14960 8289
rect 15004 8280 15034 8289
rect 15034 8280 15038 8289
rect 14185 8246 14219 8249
rect 14257 8246 14291 8249
rect 14329 8246 14363 8249
rect 14401 8246 14435 8249
rect 14473 8246 14507 8249
rect 14614 8209 14648 8240
rect 14692 8209 14726 8240
rect 14770 8209 14804 8240
rect 14848 8209 14882 8240
rect 14926 8217 14960 8240
rect 15004 8217 15038 8240
rect 14185 8175 14198 8202
rect 14198 8175 14219 8202
rect 14257 8175 14268 8202
rect 14268 8175 14291 8202
rect 14329 8175 14338 8202
rect 14338 8175 14363 8202
rect 14401 8175 14408 8202
rect 14408 8175 14435 8202
rect 14473 8175 14478 8202
rect 14478 8175 14507 8202
rect 14614 8206 14618 8209
rect 14618 8206 14648 8209
rect 14692 8206 14724 8209
rect 14724 8206 14726 8209
rect 14770 8206 14794 8209
rect 14794 8206 14804 8209
rect 14848 8206 14864 8209
rect 14864 8206 14882 8209
rect 14926 8206 14932 8217
rect 14932 8206 14960 8217
rect 15004 8206 15034 8217
rect 15034 8206 15038 8217
rect 14185 8168 14219 8175
rect 14257 8168 14291 8175
rect 14329 8168 14363 8175
rect 14401 8168 14435 8175
rect 14473 8168 14507 8175
rect 14614 8135 14648 8166
rect 14692 8135 14726 8166
rect 14770 8135 14804 8166
rect 14848 8135 14882 8166
rect 14926 8145 14960 8166
rect 15004 8145 15038 8166
rect 14431 8101 14444 8115
rect 14444 8101 14465 8115
rect 14511 8101 14514 8115
rect 14514 8101 14545 8115
rect 14614 8132 14618 8135
rect 14618 8132 14648 8135
rect 14692 8132 14724 8135
rect 14724 8132 14726 8135
rect 14770 8132 14794 8135
rect 14794 8132 14804 8135
rect 14848 8132 14864 8135
rect 14864 8132 14882 8135
rect 14926 8132 14932 8145
rect 14932 8132 14960 8145
rect 15004 8132 15034 8145
rect 15034 8132 15038 8145
rect 14431 8081 14465 8101
rect 14511 8081 14545 8101
rect 14614 8061 14648 8092
rect 14692 8061 14726 8092
rect 14770 8061 14804 8092
rect 14848 8061 14882 8092
rect 14926 8073 14960 8092
rect 15004 8073 15038 8092
rect 14431 8027 14444 8033
rect 14444 8027 14465 8033
rect 14511 8027 14514 8033
rect 14514 8027 14545 8033
rect 14614 8058 14618 8061
rect 14618 8058 14648 8061
rect 14692 8058 14724 8061
rect 14724 8058 14726 8061
rect 14770 8058 14794 8061
rect 14794 8058 14804 8061
rect 14848 8058 14864 8061
rect 14864 8058 14882 8061
rect 14926 8058 14932 8073
rect 14932 8058 14960 8073
rect 15004 8058 15034 8073
rect 15034 8058 15038 8073
rect 14431 7999 14465 8027
rect 14511 7999 14545 8027
rect 14614 7987 14648 8018
rect 14692 7987 14726 8018
rect 14770 7987 14804 8018
rect 14848 7987 14882 8018
rect 14926 8001 14960 8018
rect 15004 8001 15038 8018
rect 14614 7984 14618 7987
rect 14618 7984 14648 7987
rect 14692 7984 14724 7987
rect 14724 7984 14726 7987
rect 14770 7984 14794 7987
rect 14794 7984 14804 7987
rect 14848 7984 14864 7987
rect 14864 7984 14882 7987
rect 14926 7984 14932 8001
rect 14932 7984 14960 8001
rect 15004 7984 15034 8001
rect 15034 7984 15038 8001
rect 14431 7916 14465 7950
rect 14511 7916 14545 7950
rect 14614 7913 14648 7944
rect 14692 7913 14726 7944
rect 14770 7913 14804 7944
rect 14848 7913 14882 7944
rect 14926 7929 14960 7944
rect 15004 7929 15038 7944
rect 14614 7910 14618 7913
rect 14618 7910 14648 7913
rect 14692 7910 14724 7913
rect 14724 7910 14726 7913
rect 14770 7910 14794 7913
rect 14794 7910 14804 7913
rect 14848 7910 14864 7913
rect 14864 7910 14882 7913
rect 14926 7910 14932 7929
rect 14932 7910 14960 7929
rect 15004 7910 15034 7929
rect 15034 7910 15038 7929
rect 14614 7839 14648 7870
rect 14692 7839 14726 7870
rect 14770 7839 14804 7870
rect 14848 7839 14882 7870
rect 14926 7857 14960 7870
rect 15004 7857 15038 7870
rect 14614 7836 14618 7839
rect 14618 7836 14648 7839
rect 14692 7836 14724 7839
rect 14724 7836 14726 7839
rect 14770 7836 14794 7839
rect 14794 7836 14804 7839
rect 14848 7836 14864 7839
rect 14864 7836 14882 7839
rect 14926 7836 14932 7857
rect 14932 7836 14960 7857
rect 15004 7836 15034 7857
rect 15034 7836 15038 7857
rect 14614 7762 14648 7796
rect 14692 7762 14726 7796
rect 14770 7762 14804 7796
rect 14848 7762 14882 7796
rect 14926 7785 14960 7796
rect 15004 7785 15038 7796
rect 14926 7762 14932 7785
rect 14932 7762 14960 7785
rect 15004 7762 15034 7785
rect 15034 7762 15038 7785
rect 14614 7715 14626 7722
rect 14626 7715 14648 7722
rect 14692 7715 14694 7722
rect 14694 7715 14726 7722
rect 14770 7715 14796 7722
rect 14796 7715 14804 7722
rect 14848 7715 14864 7722
rect 14864 7715 14882 7722
rect 14614 7688 14648 7715
rect 14692 7688 14726 7715
rect 14770 7688 14804 7715
rect 14848 7688 14882 7715
rect 14926 7713 14960 7722
rect 15004 7713 15038 7722
rect 14926 7688 14932 7713
rect 14932 7688 14960 7713
rect 15004 7688 15034 7713
rect 15034 7688 15038 7713
rect 14614 7640 14648 7648
rect 14692 7640 14726 7648
rect 14770 7640 14804 7648
rect 14848 7640 14882 7648
rect 14926 7641 14960 7648
rect 15004 7641 15038 7648
rect 14614 7614 14626 7640
rect 14626 7614 14648 7640
rect 14692 7614 14694 7640
rect 14694 7614 14726 7640
rect 14770 7614 14796 7640
rect 14796 7614 14804 7640
rect 14848 7614 14864 7640
rect 14864 7614 14882 7640
rect 14926 7614 14932 7641
rect 14932 7614 14960 7641
rect 15004 7614 15034 7641
rect 15034 7614 15038 7641
rect 14614 7556 14648 7574
rect 14692 7556 14726 7574
rect 14770 7556 14804 7574
rect 14848 7556 14882 7574
rect 14926 7569 14960 7574
rect 15004 7569 15038 7574
rect 14614 7540 14626 7556
rect 14626 7540 14648 7556
rect 14692 7540 14694 7556
rect 14694 7540 14726 7556
rect 14770 7540 14796 7556
rect 14796 7540 14804 7556
rect 14848 7540 14864 7556
rect 14864 7540 14882 7556
rect 14926 7540 14932 7569
rect 14932 7540 14960 7569
rect 15004 7540 15034 7569
rect 15034 7540 15038 7569
rect 14614 7472 14648 7499
rect 14692 7472 14726 7499
rect 14770 7472 14804 7499
rect 14848 7472 14882 7499
rect 14926 7497 14960 7499
rect 15004 7497 15038 7499
rect 14614 7465 14626 7472
rect 14626 7465 14648 7472
rect 14692 7465 14694 7472
rect 14694 7465 14726 7472
rect 14770 7465 14796 7472
rect 14796 7465 14804 7472
rect 14848 7465 14864 7472
rect 14864 7465 14882 7472
rect 14926 7465 14932 7497
rect 14932 7465 14960 7497
rect 15004 7465 15034 7497
rect 15034 7465 15038 7497
rect 14614 7390 14648 7424
rect 14692 7390 14726 7424
rect 14770 7390 14804 7424
rect 14848 7390 14882 7424
rect 14926 7391 14932 7424
rect 14932 7391 14960 7424
rect 15004 7391 15034 7424
rect 15034 7391 15038 7424
rect 14926 7390 14960 7391
rect 15004 7390 15038 7391
rect 57 7354 91 7374
rect 132 7354 166 7374
rect 207 7354 241 7374
rect 282 7354 316 7374
rect 357 7354 391 7374
rect 432 7354 466 7374
rect 507 7354 541 7374
rect 582 7354 616 7374
rect 657 7354 691 7374
rect 732 7354 766 7374
rect 807 7354 841 7374
rect 882 7354 916 7374
rect 957 7354 991 7374
rect 1032 7354 1066 7374
rect 1107 7354 1141 7374
rect 1182 7354 1216 7374
rect 1256 7354 1290 7374
rect 1330 7354 1364 7374
rect 57 7340 68 7354
rect 68 7340 91 7354
rect 132 7340 137 7354
rect 137 7340 166 7354
rect 207 7340 240 7354
rect 240 7340 241 7354
rect 282 7340 309 7354
rect 309 7340 316 7354
rect 357 7340 378 7354
rect 378 7340 391 7354
rect 432 7340 447 7354
rect 447 7340 466 7354
rect 507 7340 516 7354
rect 516 7340 541 7354
rect 582 7340 585 7354
rect 585 7340 616 7354
rect 657 7340 689 7354
rect 689 7340 691 7354
rect 732 7340 758 7354
rect 758 7340 766 7354
rect 807 7340 827 7354
rect 827 7340 841 7354
rect 882 7340 896 7354
rect 896 7340 916 7354
rect 957 7340 965 7354
rect 965 7340 991 7354
rect 1032 7340 1033 7354
rect 1033 7340 1066 7354
rect 1107 7340 1135 7354
rect 1135 7340 1141 7354
rect 1182 7340 1203 7354
rect 1203 7340 1216 7354
rect 1256 7340 1271 7354
rect 1271 7340 1290 7354
rect 1330 7340 1339 7354
rect 1339 7340 1364 7354
rect 57 7282 91 7290
rect 132 7282 166 7290
rect 207 7282 241 7290
rect 282 7282 316 7290
rect 357 7282 391 7290
rect 432 7282 466 7290
rect 507 7282 541 7290
rect 582 7282 616 7290
rect 657 7282 691 7290
rect 732 7282 766 7290
rect 807 7282 841 7290
rect 882 7282 916 7290
rect 957 7282 991 7290
rect 1032 7282 1066 7290
rect 1107 7282 1141 7290
rect 1182 7282 1216 7290
rect 1256 7282 1290 7290
rect 1330 7282 1364 7290
rect 57 7256 68 7282
rect 68 7256 91 7282
rect 132 7256 137 7282
rect 137 7256 166 7282
rect 207 7256 240 7282
rect 240 7256 241 7282
rect 282 7256 309 7282
rect 309 7256 316 7282
rect 357 7256 378 7282
rect 378 7256 391 7282
rect 432 7256 447 7282
rect 447 7256 466 7282
rect 507 7256 516 7282
rect 516 7256 541 7282
rect 582 7256 585 7282
rect 585 7256 616 7282
rect 657 7256 689 7282
rect 689 7256 691 7282
rect 732 7256 758 7282
rect 758 7256 766 7282
rect 807 7256 827 7282
rect 827 7256 841 7282
rect 882 7256 896 7282
rect 896 7256 916 7282
rect 957 7256 965 7282
rect 965 7256 991 7282
rect 1032 7256 1033 7282
rect 1033 7256 1066 7282
rect 1107 7256 1135 7282
rect 1135 7256 1141 7282
rect 1182 7256 1203 7282
rect 1203 7256 1216 7282
rect 1256 7256 1271 7282
rect 1271 7256 1290 7282
rect 1330 7256 1339 7282
rect 1339 7256 1364 7282
rect 1431 7210 1465 7220
rect 1504 7210 1538 7220
rect 1577 7210 1611 7220
rect 1650 7210 1684 7220
rect 1723 7210 1757 7220
rect 1796 7210 1830 7220
rect 1869 7210 1903 7220
rect 1942 7210 1976 7220
rect 2015 7210 2049 7220
rect 2088 7210 2122 7220
rect 2161 7210 2195 7220
rect 2234 7210 2268 7220
rect 2307 7210 2341 7220
rect 2380 7210 2414 7220
rect 2453 7210 2487 7220
rect 2526 7210 2560 7220
rect 2599 7210 2633 7220
rect 2672 7210 2706 7220
rect 57 7176 68 7206
rect 68 7176 91 7206
rect 132 7176 137 7206
rect 137 7176 166 7206
rect 207 7176 240 7206
rect 240 7176 241 7206
rect 282 7176 309 7206
rect 309 7176 316 7206
rect 357 7176 378 7206
rect 378 7176 391 7206
rect 432 7176 447 7206
rect 447 7176 466 7206
rect 507 7176 516 7206
rect 516 7176 541 7206
rect 582 7176 585 7206
rect 585 7176 616 7206
rect 657 7176 689 7206
rect 689 7176 691 7206
rect 732 7176 758 7206
rect 758 7176 766 7206
rect 807 7176 827 7206
rect 827 7176 841 7206
rect 882 7176 896 7206
rect 896 7176 916 7206
rect 957 7176 965 7206
rect 965 7176 991 7206
rect 1032 7176 1033 7206
rect 1033 7176 1066 7206
rect 1107 7176 1135 7206
rect 1135 7176 1141 7206
rect 1182 7176 1203 7206
rect 1203 7176 1216 7206
rect 1256 7176 1271 7206
rect 1271 7176 1290 7206
rect 1330 7176 1339 7206
rect 1339 7176 1364 7206
rect 1431 7186 1441 7210
rect 1441 7186 1465 7210
rect 1504 7186 1509 7210
rect 1509 7186 1538 7210
rect 1577 7186 1611 7210
rect 1650 7186 1679 7210
rect 1679 7186 1684 7210
rect 1723 7186 1747 7210
rect 1747 7186 1757 7210
rect 1796 7186 1815 7210
rect 1815 7186 1830 7210
rect 1869 7186 1883 7210
rect 1883 7186 1903 7210
rect 1942 7186 1951 7210
rect 1951 7186 1976 7210
rect 2015 7186 2019 7210
rect 2019 7186 2049 7210
rect 2088 7186 2121 7210
rect 2121 7186 2122 7210
rect 2161 7186 2189 7210
rect 2189 7186 2195 7210
rect 2234 7186 2257 7210
rect 2257 7186 2268 7210
rect 2307 7186 2325 7210
rect 2325 7186 2341 7210
rect 2380 7186 2393 7210
rect 2393 7186 2414 7210
rect 2453 7186 2461 7210
rect 2461 7186 2487 7210
rect 2526 7186 2529 7210
rect 2529 7186 2560 7210
rect 2599 7186 2631 7210
rect 2631 7186 2633 7210
rect 2672 7186 2699 7210
rect 2699 7186 2706 7210
rect 2745 7186 2779 7220
rect 2818 7186 2852 7220
rect 2891 7186 2925 7220
rect 2964 7186 2998 7220
rect 3037 7186 3071 7220
rect 3110 7186 3144 7220
rect 3183 7186 3217 7220
rect 3256 7186 3290 7220
rect 3329 7186 3363 7220
rect 3402 7186 3436 7220
rect 3475 7186 3509 7220
rect 3548 7186 3582 7220
rect 3621 7186 3655 7220
rect 3694 7186 3728 7220
rect 3767 7186 3801 7220
rect 3840 7186 3874 7220
rect 3913 7186 3947 7220
rect 3986 7186 4020 7220
rect 4059 7186 4093 7220
rect 4132 7186 4166 7220
rect 4205 7186 4239 7220
rect 4278 7186 4312 7220
rect 4351 7186 4385 7220
rect 4424 7186 4458 7220
rect 4497 7186 4531 7220
rect 4570 7186 4604 7220
rect 4643 7186 4677 7220
rect 4716 7186 4750 7220
rect 4789 7186 4823 7220
rect 4862 7186 4896 7220
rect 4935 7186 4969 7220
rect 5008 7186 5042 7220
rect 5081 7186 5115 7220
rect 5154 7186 5188 7220
rect 5227 7186 5261 7220
rect 5300 7186 5334 7220
rect 5373 7186 5407 7220
rect 5446 7186 5480 7220
rect 5519 7186 5553 7220
rect 5592 7186 5626 7220
rect 5665 7186 5699 7220
rect 5738 7186 5772 7220
rect 5811 7186 5845 7220
rect 5884 7186 5918 7220
rect 5957 7186 5991 7220
rect 6030 7186 6064 7220
rect 6103 7186 6137 7220
rect 6176 7186 6210 7220
rect 6249 7186 6283 7220
rect 6322 7186 6356 7220
rect 6395 7186 6429 7220
rect 6468 7186 6502 7220
rect 6540 7186 6574 7220
rect 6612 7186 6646 7220
rect 6684 7186 6718 7220
rect 6756 7186 6790 7220
rect 6828 7186 6862 7220
rect 6900 7186 6934 7220
rect 6972 7186 7006 7220
rect 7044 7186 7078 7220
rect 7116 7186 7150 7220
rect 57 7172 91 7176
rect 132 7172 166 7176
rect 207 7172 241 7176
rect 282 7172 316 7176
rect 357 7172 391 7176
rect 432 7172 466 7176
rect 507 7172 541 7176
rect 582 7172 616 7176
rect 657 7172 691 7176
rect 732 7172 766 7176
rect 807 7172 841 7176
rect 882 7172 916 7176
rect 957 7172 991 7176
rect 1032 7172 1066 7176
rect 1107 7172 1141 7176
rect 1182 7172 1216 7176
rect 1256 7172 1290 7176
rect 1330 7172 1364 7176
rect 57 7104 68 7122
rect 68 7104 91 7122
rect 132 7104 137 7122
rect 137 7104 166 7122
rect 207 7104 240 7122
rect 240 7104 241 7122
rect 282 7104 309 7122
rect 309 7104 316 7122
rect 357 7104 378 7122
rect 378 7104 391 7122
rect 432 7104 447 7122
rect 447 7104 466 7122
rect 507 7104 516 7122
rect 516 7104 541 7122
rect 582 7104 585 7122
rect 585 7104 616 7122
rect 657 7104 689 7122
rect 689 7104 691 7122
rect 732 7104 758 7122
rect 758 7104 766 7122
rect 807 7104 827 7122
rect 827 7104 841 7122
rect 882 7104 896 7122
rect 896 7104 916 7122
rect 957 7104 965 7122
rect 965 7104 991 7122
rect 1032 7104 1033 7122
rect 1033 7104 1066 7122
rect 1107 7104 1135 7122
rect 1135 7104 1141 7122
rect 1182 7104 1203 7122
rect 1203 7104 1216 7122
rect 1256 7104 1271 7122
rect 1271 7104 1290 7122
rect 1330 7104 1339 7122
rect 1339 7104 1364 7122
rect 57 7088 91 7104
rect 132 7088 166 7104
rect 207 7088 241 7104
rect 282 7088 316 7104
rect 357 7088 391 7104
rect 432 7088 466 7104
rect 507 7088 541 7104
rect 582 7088 616 7104
rect 657 7088 691 7104
rect 732 7088 766 7104
rect 807 7088 841 7104
rect 882 7088 916 7104
rect 957 7088 991 7104
rect 1032 7088 1066 7104
rect 1107 7088 1141 7104
rect 1182 7088 1216 7104
rect 1256 7088 1290 7104
rect 1330 7088 1364 7104
rect 57 7032 68 7038
rect 68 7032 91 7038
rect 132 7032 137 7038
rect 137 7032 166 7038
rect 207 7032 240 7038
rect 240 7032 241 7038
rect 282 7032 309 7038
rect 309 7032 316 7038
rect 357 7032 378 7038
rect 378 7032 391 7038
rect 432 7032 447 7038
rect 447 7032 466 7038
rect 507 7032 516 7038
rect 516 7032 541 7038
rect 582 7032 585 7038
rect 585 7032 616 7038
rect 657 7032 689 7038
rect 689 7032 691 7038
rect 732 7032 758 7038
rect 758 7032 766 7038
rect 807 7032 827 7038
rect 827 7032 841 7038
rect 882 7032 896 7038
rect 896 7032 916 7038
rect 957 7032 965 7038
rect 965 7032 991 7038
rect 1032 7032 1033 7038
rect 1033 7032 1066 7038
rect 1107 7032 1135 7038
rect 1135 7032 1141 7038
rect 1182 7032 1203 7038
rect 1203 7032 1216 7038
rect 1256 7032 1271 7038
rect 1271 7032 1290 7038
rect 1330 7032 1339 7038
rect 1339 7032 1364 7038
rect 57 7004 91 7032
rect 132 7004 166 7032
rect 207 7004 241 7032
rect 282 7004 316 7032
rect 357 7004 391 7032
rect 432 7004 466 7032
rect 507 7004 541 7032
rect 582 7004 616 7032
rect 657 7004 691 7032
rect 732 7004 766 7032
rect 807 7004 841 7032
rect 882 7004 916 7032
rect 957 7004 991 7032
rect 1032 7004 1066 7032
rect 1107 7004 1141 7032
rect 1182 7004 1216 7032
rect 1256 7004 1290 7032
rect 1330 7004 1364 7032
rect 14614 7315 14648 7349
rect 14692 7315 14726 7349
rect 14770 7315 14804 7349
rect 14848 7315 14882 7349
rect 14926 7319 14932 7349
rect 14932 7319 14960 7349
rect 15004 7319 15034 7349
rect 15034 7319 15038 7349
rect 14926 7315 14960 7319
rect 15004 7315 15038 7319
rect 14614 7248 14626 7274
rect 14626 7248 14648 7274
rect 14692 7248 14694 7274
rect 14694 7248 14726 7274
rect 14770 7248 14796 7274
rect 14796 7248 14804 7274
rect 14848 7248 14864 7274
rect 14864 7248 14882 7274
rect 14614 7240 14648 7248
rect 14692 7240 14726 7248
rect 14770 7240 14804 7248
rect 14848 7240 14882 7248
rect 14926 7247 14932 7274
rect 14932 7247 14960 7274
rect 15004 7247 15034 7274
rect 15034 7247 15038 7274
rect 14926 7240 14960 7247
rect 15004 7240 15038 7247
rect 14614 7176 14626 7199
rect 14626 7176 14648 7199
rect 14692 7176 14694 7199
rect 14694 7176 14726 7199
rect 14770 7176 14796 7199
rect 14796 7176 14804 7199
rect 14848 7176 14864 7199
rect 14864 7176 14882 7199
rect 14614 7165 14648 7176
rect 14692 7165 14726 7176
rect 14770 7165 14804 7176
rect 14848 7165 14882 7176
rect 14926 7175 14932 7199
rect 14932 7175 14960 7199
rect 15004 7175 15034 7199
rect 15034 7175 15038 7199
rect 14926 7165 14960 7175
rect 15004 7165 15038 7175
rect 14614 7104 14626 7124
rect 14626 7104 14648 7124
rect 14692 7104 14694 7124
rect 14694 7104 14726 7124
rect 14770 7104 14796 7124
rect 14796 7104 14804 7124
rect 14848 7104 14864 7124
rect 14864 7104 14882 7124
rect 14614 7090 14648 7104
rect 14692 7090 14726 7104
rect 14770 7090 14804 7104
rect 14848 7090 14882 7104
rect 14926 7103 14932 7124
rect 14932 7103 14960 7124
rect 15004 7103 15034 7124
rect 15034 7103 15038 7124
rect 14926 7090 14960 7103
rect 15004 7090 15038 7103
rect 15068 6805 15102 6825
rect 15068 6791 15102 6805
rect 15068 6731 15102 6753
rect 15068 6719 15102 6731
rect 15068 6657 15102 6681
rect 15068 6647 15102 6657
rect 15068 6583 15102 6609
rect 15068 6575 15102 6583
rect 15068 6509 15102 6537
rect 15068 6503 15102 6509
rect 68 6434 102 6439
rect 141 6434 175 6439
rect 214 6434 248 6439
rect 287 6434 321 6439
rect 360 6434 394 6439
rect 433 6434 467 6439
rect 506 6434 540 6439
rect 579 6434 613 6439
rect 652 6434 686 6439
rect 725 6434 759 6439
rect 798 6434 832 6439
rect 871 6434 905 6439
rect 944 6434 978 6439
rect 1017 6434 1051 6439
rect 1090 6435 15020 6439
rect 15068 6435 15102 6465
rect 1090 6434 14932 6435
rect 68 6405 102 6434
rect 141 6405 171 6434
rect 171 6405 175 6434
rect 214 6405 240 6434
rect 240 6405 248 6434
rect 287 6405 309 6434
rect 309 6405 321 6434
rect 360 6405 378 6434
rect 378 6405 394 6434
rect 433 6405 447 6434
rect 447 6405 467 6434
rect 506 6405 516 6434
rect 516 6405 540 6434
rect 579 6405 585 6434
rect 585 6405 613 6434
rect 652 6405 654 6434
rect 654 6405 686 6434
rect 725 6405 758 6434
rect 758 6405 759 6434
rect 798 6405 827 6434
rect 827 6405 832 6434
rect 871 6405 896 6434
rect 896 6405 905 6434
rect 944 6405 965 6434
rect 965 6405 978 6434
rect 1017 6405 1034 6434
rect 1034 6405 1051 6434
rect 1090 6400 1103 6434
rect 1103 6400 1137 6434
rect 1137 6400 1172 6434
rect 1172 6400 1206 6434
rect 1206 6400 1241 6434
rect 1241 6400 1275 6434
rect 1275 6400 1310 6434
rect 1310 6400 1344 6434
rect 1344 6400 1379 6434
rect 1379 6400 1413 6434
rect 1413 6400 1448 6434
rect 1448 6400 1482 6434
rect 1482 6400 1517 6434
rect 1517 6400 1551 6434
rect 1551 6400 1586 6434
rect 1586 6400 1620 6434
rect 1620 6400 1655 6434
rect 1655 6400 1689 6434
rect 1689 6400 1724 6434
rect 1724 6400 1758 6434
rect 1758 6400 1793 6434
rect 1793 6400 1827 6434
rect 1827 6400 1862 6434
rect 1862 6400 1896 6434
rect 1896 6400 1931 6434
rect 1931 6400 1965 6434
rect 1965 6400 2000 6434
rect 2000 6400 2034 6434
rect 2034 6400 2069 6434
rect 2069 6400 2103 6434
rect 2103 6400 2138 6434
rect 2138 6400 2172 6434
rect 2172 6400 2207 6434
rect 2207 6400 2241 6434
rect 2241 6400 2276 6434
rect 2276 6400 2310 6434
rect 2310 6400 2345 6434
rect 2345 6400 2379 6434
rect 2379 6400 2414 6434
rect 2414 6400 2448 6434
rect 2448 6400 2483 6434
rect 2483 6400 2517 6434
rect 2517 6400 2551 6434
rect 2551 6400 2585 6434
rect 2585 6400 2619 6434
rect 2619 6400 2653 6434
rect 2653 6400 2687 6434
rect 2687 6400 2721 6434
rect 2721 6400 2755 6434
rect 2755 6400 2789 6434
rect 2789 6400 2823 6434
rect 2823 6400 2857 6434
rect 2857 6400 2891 6434
rect 2891 6400 2925 6434
rect 2925 6400 2959 6434
rect 2959 6400 2993 6434
rect 2993 6400 3027 6434
rect 3027 6400 3061 6434
rect 3061 6400 3095 6434
rect 3095 6400 3129 6434
rect 3129 6400 3163 6434
rect 3163 6400 3197 6434
rect 3197 6400 3231 6434
rect 3231 6400 3265 6434
rect 3265 6400 3299 6434
rect 3299 6400 3333 6434
rect 3333 6400 3367 6434
rect 3367 6400 3401 6434
rect 3401 6400 3435 6434
rect 3435 6400 3469 6434
rect 3469 6400 3503 6434
rect 3503 6400 3537 6434
rect 3537 6400 3571 6434
rect 3571 6400 3605 6434
rect 3605 6400 3639 6434
rect 3639 6400 3673 6434
rect 3673 6400 3707 6434
rect 3707 6400 3741 6434
rect 3741 6400 3775 6434
rect 3775 6400 3809 6434
rect 3809 6400 3843 6434
rect 3843 6400 3877 6434
rect 3877 6400 3911 6434
rect 3911 6400 3945 6434
rect 3945 6400 3979 6434
rect 3979 6400 4013 6434
rect 4013 6400 4047 6434
rect 4047 6400 4081 6434
rect 4081 6400 4115 6434
rect 4115 6400 4149 6434
rect 4149 6400 4183 6434
rect 4183 6400 4217 6434
rect 4217 6400 4251 6434
rect 4251 6400 4285 6434
rect 4285 6400 4319 6434
rect 4319 6400 4353 6434
rect 4353 6400 4387 6434
rect 4387 6400 4421 6434
rect 4421 6400 4455 6434
rect 4455 6400 4489 6434
rect 4489 6400 4523 6434
rect 4523 6400 4557 6434
rect 4557 6400 4591 6434
rect 4591 6400 4625 6434
rect 4625 6400 4659 6434
rect 4659 6400 4693 6434
rect 4693 6400 4727 6434
rect 4727 6400 4761 6434
rect 4761 6400 4795 6434
rect 4795 6400 4829 6434
rect 4829 6400 4863 6434
rect 4863 6400 4897 6434
rect 4897 6400 4931 6434
rect 4931 6400 4965 6434
rect 4965 6400 4999 6434
rect 4999 6400 5033 6434
rect 5033 6400 5067 6434
rect 5067 6400 5101 6434
rect 5101 6400 5135 6434
rect 5135 6400 5169 6434
rect 5169 6400 5203 6434
rect 5203 6400 5237 6434
rect 5237 6400 5271 6434
rect 5271 6400 5305 6434
rect 5305 6400 5339 6434
rect 5339 6400 5373 6434
rect 5373 6400 5407 6434
rect 5407 6400 5441 6434
rect 5441 6400 5475 6434
rect 5475 6400 5509 6434
rect 5509 6400 5543 6434
rect 5543 6400 5577 6434
rect 5577 6400 5611 6434
rect 5611 6400 5645 6434
rect 5645 6400 5679 6434
rect 5679 6400 5713 6434
rect 5713 6400 5747 6434
rect 5747 6400 5781 6434
rect 5781 6400 5815 6434
rect 5815 6400 5849 6434
rect 5849 6400 5883 6434
rect 5883 6400 5917 6434
rect 5917 6400 5951 6434
rect 5951 6400 5985 6434
rect 5985 6400 6019 6434
rect 6019 6400 6053 6434
rect 6053 6400 6087 6434
rect 6087 6400 6121 6434
rect 6121 6400 6155 6434
rect 6155 6400 6189 6434
rect 6189 6400 6223 6434
rect 6223 6400 6257 6434
rect 6257 6400 6291 6434
rect 6291 6400 6325 6434
rect 6325 6400 6359 6434
rect 6359 6400 6393 6434
rect 6393 6400 6427 6434
rect 6427 6400 6461 6434
rect 6461 6400 6495 6434
rect 6495 6400 6529 6434
rect 6529 6400 6563 6434
rect 6563 6400 6597 6434
rect 6597 6400 6631 6434
rect 6631 6400 6665 6434
rect 6665 6400 6699 6434
rect 6699 6400 6733 6434
rect 6733 6400 6767 6434
rect 6767 6400 6801 6434
rect 6801 6400 6835 6434
rect 6835 6400 6869 6434
rect 6869 6400 6903 6434
rect 6903 6400 6937 6434
rect 6937 6400 6971 6434
rect 6971 6400 7005 6434
rect 7005 6400 7039 6434
rect 7039 6400 7073 6434
rect 7073 6400 7107 6434
rect 7107 6400 7141 6434
rect 7141 6400 7175 6434
rect 7175 6400 7209 6434
rect 7209 6400 7243 6434
rect 7243 6400 7277 6434
rect 7277 6400 7311 6434
rect 7311 6400 7345 6434
rect 7345 6400 7379 6434
rect 7379 6400 7413 6434
rect 7413 6400 7447 6434
rect 7447 6400 7481 6434
rect 7481 6400 7515 6434
rect 7515 6400 7549 6434
rect 7549 6400 7583 6434
rect 7583 6400 7617 6434
rect 7617 6400 7651 6434
rect 7651 6400 7685 6434
rect 7685 6400 7719 6434
rect 7719 6400 7753 6434
rect 7753 6400 7787 6434
rect 7787 6400 7821 6434
rect 7821 6400 7855 6434
rect 7855 6400 7889 6434
rect 7889 6400 7923 6434
rect 7923 6400 7957 6434
rect 7957 6400 7991 6434
rect 7991 6400 8025 6434
rect 8025 6400 8059 6434
rect 8059 6400 8093 6434
rect 8093 6400 8127 6434
rect 8127 6400 8161 6434
rect 8161 6400 8195 6434
rect 8195 6400 8229 6434
rect 8229 6400 8263 6434
rect 8263 6400 8297 6434
rect 8297 6400 8331 6434
rect 8331 6400 8365 6434
rect 8365 6400 8399 6434
rect 8399 6400 8433 6434
rect 8433 6400 8467 6434
rect 8467 6400 8501 6434
rect 8501 6400 8535 6434
rect 8535 6400 8569 6434
rect 8569 6400 8603 6434
rect 8603 6400 8637 6434
rect 8637 6400 8671 6434
rect 8671 6400 8705 6434
rect 8705 6400 8739 6434
rect 8739 6400 8773 6434
rect 8773 6400 8807 6434
rect 8807 6400 8841 6434
rect 8841 6400 8875 6434
rect 8875 6400 8909 6434
rect 8909 6400 8943 6434
rect 8943 6400 8977 6434
rect 8977 6400 9011 6434
rect 9011 6400 9045 6434
rect 9045 6400 9079 6434
rect 9079 6400 9113 6434
rect 9113 6400 9147 6434
rect 9147 6400 9181 6434
rect 9181 6400 9215 6434
rect 9215 6400 9249 6434
rect 9249 6400 9283 6434
rect 9283 6400 9317 6434
rect 9317 6400 9351 6434
rect 9351 6400 9385 6434
rect 9385 6400 9419 6434
rect 9419 6400 9453 6434
rect 9453 6400 9487 6434
rect 9487 6400 9521 6434
rect 9521 6400 9555 6434
rect 9555 6400 9589 6434
rect 9589 6400 9623 6434
rect 9623 6400 9657 6434
rect 9657 6400 9691 6434
rect 9691 6400 9725 6434
rect 9725 6400 9759 6434
rect 9759 6400 9793 6434
rect 9793 6400 9827 6434
rect 9827 6400 9861 6434
rect 9861 6400 9895 6434
rect 9895 6400 9929 6434
rect 9929 6400 9963 6434
rect 9963 6400 9997 6434
rect 9997 6400 10031 6434
rect 10031 6400 10065 6434
rect 10065 6400 10099 6434
rect 10099 6400 10133 6434
rect 10133 6400 10167 6434
rect 10167 6400 10201 6434
rect 10201 6400 10235 6434
rect 10235 6400 10269 6434
rect 10269 6400 10303 6434
rect 10303 6400 10337 6434
rect 10337 6400 10371 6434
rect 10371 6400 10405 6434
rect 10405 6400 10439 6434
rect 10439 6400 10473 6434
rect 10473 6400 10507 6434
rect 10507 6400 10541 6434
rect 10541 6400 10575 6434
rect 10575 6400 10609 6434
rect 10609 6400 10643 6434
rect 10643 6400 10677 6434
rect 10677 6400 10711 6434
rect 10711 6400 10745 6434
rect 10745 6400 10779 6434
rect 10779 6400 10813 6434
rect 10813 6400 10847 6434
rect 10847 6400 10881 6434
rect 10881 6400 10915 6434
rect 10915 6400 10949 6434
rect 10949 6400 10983 6434
rect 10983 6400 11017 6434
rect 11017 6400 11051 6434
rect 11051 6400 11085 6434
rect 11085 6400 11119 6434
rect 11119 6400 11153 6434
rect 11153 6400 11187 6434
rect 11187 6400 11221 6434
rect 11221 6400 11255 6434
rect 11255 6400 11289 6434
rect 11289 6400 11323 6434
rect 11323 6400 11357 6434
rect 11357 6400 11391 6434
rect 11391 6400 11425 6434
rect 11425 6400 11459 6434
rect 11459 6400 11493 6434
rect 11493 6400 11527 6434
rect 11527 6400 11561 6434
rect 11561 6400 11595 6434
rect 11595 6400 11629 6434
rect 11629 6400 11663 6434
rect 11663 6400 11697 6434
rect 11697 6400 11731 6434
rect 11731 6400 11765 6434
rect 11765 6400 11799 6434
rect 11799 6400 11833 6434
rect 11833 6400 11867 6434
rect 11867 6400 11901 6434
rect 11901 6400 11935 6434
rect 11935 6400 11969 6434
rect 11969 6400 12003 6434
rect 12003 6400 12037 6434
rect 12037 6400 12071 6434
rect 12071 6400 12105 6434
rect 12105 6400 12139 6434
rect 12139 6400 12173 6434
rect 12173 6400 12207 6434
rect 12207 6400 12241 6434
rect 12241 6400 12275 6434
rect 12275 6400 12309 6434
rect 12309 6400 12343 6434
rect 12343 6400 12377 6434
rect 12377 6400 12411 6434
rect 12411 6400 12445 6434
rect 12445 6400 12479 6434
rect 12479 6400 12513 6434
rect 12513 6400 12547 6434
rect 12547 6400 12581 6434
rect 12581 6400 12615 6434
rect 12615 6400 12649 6434
rect 12649 6400 12683 6434
rect 12683 6400 12717 6434
rect 12717 6400 12751 6434
rect 12751 6400 12785 6434
rect 12785 6400 12819 6434
rect 12819 6400 12853 6434
rect 12853 6400 12887 6434
rect 12887 6400 12921 6434
rect 12921 6400 12955 6434
rect 12955 6400 12989 6434
rect 12989 6400 13023 6434
rect 13023 6400 13057 6434
rect 13057 6400 13091 6434
rect 13091 6400 13125 6434
rect 13125 6400 13159 6434
rect 13159 6400 13193 6434
rect 13193 6400 13227 6434
rect 13227 6400 13261 6434
rect 13261 6400 13295 6434
rect 13295 6400 13329 6434
rect 13329 6400 13363 6434
rect 13363 6400 13397 6434
rect 13397 6400 13431 6434
rect 13431 6400 13465 6434
rect 13465 6400 13499 6434
rect 13499 6400 13533 6434
rect 13533 6400 13567 6434
rect 13567 6400 13601 6434
rect 13601 6400 13635 6434
rect 13635 6400 13669 6434
rect 13669 6400 13703 6434
rect 13703 6400 13737 6434
rect 13737 6400 13771 6434
rect 13771 6400 13805 6434
rect 13805 6400 13839 6434
rect 13839 6400 13873 6434
rect 13873 6400 13907 6434
rect 13907 6400 13941 6434
rect 13941 6400 13975 6434
rect 13975 6400 14009 6434
rect 14009 6400 14043 6434
rect 14043 6400 14077 6434
rect 14077 6400 14111 6434
rect 14111 6400 14145 6434
rect 14145 6400 14179 6434
rect 14179 6400 14213 6434
rect 14213 6400 14247 6434
rect 14247 6400 14281 6434
rect 14281 6400 14315 6434
rect 14315 6400 14349 6434
rect 14349 6400 14383 6434
rect 14383 6400 14417 6434
rect 14417 6400 14451 6434
rect 14451 6400 14485 6434
rect 14485 6400 14519 6434
rect 14519 6400 14553 6434
rect 14553 6400 14587 6434
rect 14587 6400 14621 6434
rect 14621 6400 14655 6434
rect 14655 6400 14689 6434
rect 14689 6400 14723 6434
rect 14723 6400 14757 6434
rect 14757 6400 14791 6434
rect 14791 6400 14825 6434
rect 14825 6400 14859 6434
rect 14859 6400 14893 6434
rect 14893 6401 14932 6434
rect 14932 6401 14966 6435
rect 14966 6401 15000 6435
rect 15000 6401 15020 6435
rect 15068 6431 15102 6435
rect 14893 6400 15020 6401
rect 68 6360 102 6367
rect 141 6360 175 6367
rect 214 6360 248 6367
rect 287 6360 321 6367
rect 360 6360 394 6367
rect 433 6360 467 6367
rect 506 6360 540 6367
rect 579 6360 613 6367
rect 652 6360 686 6367
rect 725 6360 759 6367
rect 798 6360 832 6367
rect 871 6360 905 6367
rect 944 6360 978 6367
rect 1017 6360 1051 6367
rect 1090 6360 15020 6400
rect 15068 6360 15102 6393
rect 68 6333 102 6360
rect 141 6333 171 6360
rect 171 6333 175 6360
rect 214 6333 240 6360
rect 240 6333 248 6360
rect 287 6333 309 6360
rect 309 6333 321 6360
rect 360 6333 378 6360
rect 378 6333 394 6360
rect 433 6333 447 6360
rect 447 6333 467 6360
rect 506 6333 516 6360
rect 516 6333 540 6360
rect 579 6333 585 6360
rect 585 6333 613 6360
rect 652 6333 654 6360
rect 654 6333 686 6360
rect 725 6333 758 6360
rect 758 6333 759 6360
rect 798 6333 827 6360
rect 827 6333 832 6360
rect 871 6333 896 6360
rect 896 6333 905 6360
rect 944 6333 965 6360
rect 965 6333 978 6360
rect 1017 6333 1034 6360
rect 1034 6333 1051 6360
rect 1090 6326 1103 6360
rect 1103 6326 1137 6360
rect 1137 6326 1172 6360
rect 1172 6326 1206 6360
rect 1206 6326 1241 6360
rect 1241 6326 1275 6360
rect 1275 6326 1310 6360
rect 1310 6326 1344 6360
rect 1344 6326 1379 6360
rect 1379 6326 1413 6360
rect 1413 6326 1448 6360
rect 1448 6326 1482 6360
rect 1482 6326 1517 6360
rect 1517 6326 1551 6360
rect 1551 6326 1586 6360
rect 1586 6326 1620 6360
rect 1620 6326 1655 6360
rect 1655 6326 1689 6360
rect 1689 6326 1724 6360
rect 1724 6326 1758 6360
rect 1758 6326 1793 6360
rect 1793 6326 1827 6360
rect 1827 6326 1862 6360
rect 1862 6326 1896 6360
rect 1896 6326 1931 6360
rect 1931 6326 1965 6360
rect 1965 6326 2000 6360
rect 2000 6326 2034 6360
rect 2034 6326 2069 6360
rect 2069 6326 2103 6360
rect 2103 6326 2138 6360
rect 2138 6326 2172 6360
rect 2172 6326 2207 6360
rect 2207 6326 2241 6360
rect 2241 6326 2276 6360
rect 2276 6326 2310 6360
rect 2310 6326 2345 6360
rect 2345 6326 2379 6360
rect 2379 6326 2414 6360
rect 2414 6326 2448 6360
rect 2448 6326 2483 6360
rect 2483 6326 2517 6360
rect 2517 6326 2551 6360
rect 2551 6326 2585 6360
rect 2585 6326 2619 6360
rect 2619 6326 2653 6360
rect 2653 6326 2687 6360
rect 2687 6326 2721 6360
rect 2721 6326 2755 6360
rect 2755 6326 2789 6360
rect 2789 6326 2823 6360
rect 2823 6326 2857 6360
rect 2857 6326 2891 6360
rect 2891 6326 2925 6360
rect 2925 6326 2959 6360
rect 2959 6326 2993 6360
rect 2993 6326 3027 6360
rect 3027 6326 3061 6360
rect 3061 6326 3095 6360
rect 3095 6326 3129 6360
rect 3129 6326 3163 6360
rect 3163 6326 3197 6360
rect 3197 6326 3231 6360
rect 3231 6326 3265 6360
rect 3265 6326 3299 6360
rect 3299 6326 3333 6360
rect 3333 6326 3367 6360
rect 3367 6326 3401 6360
rect 3401 6326 3435 6360
rect 3435 6326 3469 6360
rect 3469 6326 3503 6360
rect 3503 6326 3537 6360
rect 3537 6326 3571 6360
rect 3571 6326 3605 6360
rect 3605 6326 3639 6360
rect 3639 6326 3673 6360
rect 3673 6326 3707 6360
rect 3707 6326 3741 6360
rect 3741 6326 3775 6360
rect 3775 6326 3809 6360
rect 3809 6326 3843 6360
rect 3843 6326 3877 6360
rect 3877 6326 3911 6360
rect 3911 6326 3945 6360
rect 3945 6326 3979 6360
rect 3979 6326 4013 6360
rect 4013 6326 4047 6360
rect 4047 6326 4081 6360
rect 4081 6326 4115 6360
rect 4115 6326 4149 6360
rect 4149 6326 4183 6360
rect 4183 6326 4217 6360
rect 4217 6326 4251 6360
rect 4251 6326 4285 6360
rect 4285 6326 4319 6360
rect 4319 6326 4353 6360
rect 4353 6326 4387 6360
rect 4387 6326 4421 6360
rect 4421 6326 4455 6360
rect 4455 6326 4489 6360
rect 4489 6326 4523 6360
rect 4523 6326 4557 6360
rect 4557 6326 4591 6360
rect 4591 6326 4625 6360
rect 4625 6326 4659 6360
rect 4659 6326 4693 6360
rect 4693 6326 4727 6360
rect 4727 6326 4761 6360
rect 4761 6326 4795 6360
rect 4795 6326 4829 6360
rect 4829 6326 4863 6360
rect 4863 6326 4897 6360
rect 4897 6326 4931 6360
rect 4931 6326 4965 6360
rect 4965 6326 4999 6360
rect 4999 6326 5033 6360
rect 5033 6326 5067 6360
rect 5067 6326 5101 6360
rect 5101 6326 5135 6360
rect 5135 6326 5169 6360
rect 5169 6326 5203 6360
rect 5203 6326 5237 6360
rect 5237 6326 5271 6360
rect 5271 6326 5305 6360
rect 5305 6326 5339 6360
rect 5339 6326 5373 6360
rect 5373 6326 5407 6360
rect 5407 6326 5441 6360
rect 5441 6326 5475 6360
rect 5475 6326 5509 6360
rect 5509 6326 5543 6360
rect 5543 6326 5577 6360
rect 5577 6326 5611 6360
rect 5611 6326 5645 6360
rect 5645 6326 5679 6360
rect 5679 6326 5713 6360
rect 5713 6326 5747 6360
rect 5747 6326 5781 6360
rect 5781 6326 5815 6360
rect 5815 6326 5849 6360
rect 5849 6326 5883 6360
rect 5883 6326 5917 6360
rect 5917 6326 5951 6360
rect 5951 6326 5985 6360
rect 5985 6326 6019 6360
rect 6019 6326 6053 6360
rect 6053 6326 6087 6360
rect 6087 6326 6121 6360
rect 6121 6326 6155 6360
rect 6155 6326 6189 6360
rect 6189 6326 6223 6360
rect 6223 6326 6257 6360
rect 6257 6326 6291 6360
rect 6291 6326 6325 6360
rect 6325 6326 6359 6360
rect 6359 6326 6393 6360
rect 6393 6326 6427 6360
rect 6427 6326 6461 6360
rect 6461 6326 6495 6360
rect 6495 6326 6529 6360
rect 6529 6326 6563 6360
rect 6563 6326 6597 6360
rect 6597 6326 6631 6360
rect 6631 6326 6665 6360
rect 6665 6326 6699 6360
rect 6699 6326 6733 6360
rect 6733 6326 6767 6360
rect 6767 6326 6801 6360
rect 6801 6326 6835 6360
rect 6835 6326 6869 6360
rect 6869 6326 6903 6360
rect 6903 6326 6937 6360
rect 6937 6326 6971 6360
rect 6971 6326 7005 6360
rect 7005 6326 7039 6360
rect 7039 6326 7073 6360
rect 7073 6326 7107 6360
rect 7107 6326 7141 6360
rect 7141 6326 7175 6360
rect 7175 6326 7209 6360
rect 7209 6326 7243 6360
rect 7243 6326 7277 6360
rect 7277 6326 7311 6360
rect 7311 6326 7345 6360
rect 7345 6326 7379 6360
rect 7379 6326 7413 6360
rect 7413 6326 7447 6360
rect 7447 6326 7481 6360
rect 7481 6326 7515 6360
rect 7515 6326 7549 6360
rect 7549 6326 7583 6360
rect 7583 6326 7617 6360
rect 7617 6326 7651 6360
rect 7651 6326 7685 6360
rect 7685 6326 7719 6360
rect 7719 6326 7753 6360
rect 7753 6326 7787 6360
rect 7787 6326 7821 6360
rect 7821 6326 7855 6360
rect 7855 6326 7889 6360
rect 7889 6326 7923 6360
rect 7923 6326 7957 6360
rect 7957 6326 7991 6360
rect 7991 6326 8025 6360
rect 8025 6326 8059 6360
rect 8059 6326 8093 6360
rect 8093 6326 8127 6360
rect 8127 6326 8161 6360
rect 8161 6326 8195 6360
rect 8195 6326 8229 6360
rect 8229 6326 8263 6360
rect 8263 6326 8297 6360
rect 8297 6326 8331 6360
rect 8331 6326 8365 6360
rect 8365 6326 8399 6360
rect 8399 6326 8433 6360
rect 8433 6326 8467 6360
rect 8467 6326 8501 6360
rect 8501 6326 8535 6360
rect 8535 6326 8569 6360
rect 8569 6326 8603 6360
rect 8603 6326 8637 6360
rect 8637 6326 8671 6360
rect 8671 6326 8705 6360
rect 8705 6326 8739 6360
rect 8739 6326 8773 6360
rect 8773 6326 8807 6360
rect 8807 6326 8841 6360
rect 8841 6326 8875 6360
rect 8875 6326 8909 6360
rect 8909 6326 8943 6360
rect 8943 6326 8977 6360
rect 8977 6326 9011 6360
rect 9011 6326 9045 6360
rect 9045 6326 9079 6360
rect 9079 6326 9113 6360
rect 9113 6326 9147 6360
rect 9147 6326 9181 6360
rect 9181 6326 9215 6360
rect 9215 6326 9249 6360
rect 9249 6326 9283 6360
rect 9283 6326 9317 6360
rect 9317 6326 9351 6360
rect 9351 6326 9385 6360
rect 9385 6326 9419 6360
rect 9419 6326 9453 6360
rect 9453 6326 9487 6360
rect 9487 6326 9521 6360
rect 9521 6326 9555 6360
rect 9555 6326 9589 6360
rect 9589 6326 9623 6360
rect 9623 6326 9657 6360
rect 9657 6326 9691 6360
rect 9691 6326 9725 6360
rect 9725 6326 9759 6360
rect 9759 6326 9793 6360
rect 9793 6326 9827 6360
rect 9827 6326 9861 6360
rect 9861 6326 9895 6360
rect 9895 6326 9929 6360
rect 9929 6326 9963 6360
rect 9963 6326 9997 6360
rect 9997 6326 10031 6360
rect 10031 6326 10065 6360
rect 10065 6326 10099 6360
rect 10099 6326 10133 6360
rect 10133 6326 10167 6360
rect 10167 6326 10201 6360
rect 10201 6326 10235 6360
rect 10235 6326 10269 6360
rect 10269 6326 10303 6360
rect 10303 6326 10337 6360
rect 10337 6326 10371 6360
rect 10371 6326 10405 6360
rect 10405 6326 10439 6360
rect 10439 6326 10473 6360
rect 10473 6326 10507 6360
rect 10507 6326 10541 6360
rect 10541 6326 10575 6360
rect 10575 6326 10609 6360
rect 10609 6326 10643 6360
rect 10643 6326 10677 6360
rect 10677 6326 10711 6360
rect 10711 6326 10745 6360
rect 10745 6326 10779 6360
rect 10779 6326 10813 6360
rect 10813 6326 10847 6360
rect 10847 6326 10881 6360
rect 10881 6326 10915 6360
rect 10915 6326 10949 6360
rect 10949 6326 10983 6360
rect 10983 6326 11017 6360
rect 11017 6326 11051 6360
rect 11051 6326 11085 6360
rect 11085 6326 11119 6360
rect 11119 6326 11153 6360
rect 11153 6326 11187 6360
rect 11187 6326 11221 6360
rect 11221 6326 11255 6360
rect 11255 6326 11289 6360
rect 11289 6326 11323 6360
rect 11323 6326 11357 6360
rect 11357 6326 11391 6360
rect 11391 6326 11425 6360
rect 11425 6326 11459 6360
rect 11459 6326 11493 6360
rect 11493 6326 11527 6360
rect 11527 6326 11561 6360
rect 11561 6326 11595 6360
rect 11595 6326 11629 6360
rect 11629 6326 11663 6360
rect 11663 6326 11697 6360
rect 11697 6326 11731 6360
rect 11731 6326 11765 6360
rect 11765 6326 11799 6360
rect 11799 6326 11833 6360
rect 11833 6326 11867 6360
rect 11867 6326 11901 6360
rect 11901 6326 11935 6360
rect 11935 6326 11969 6360
rect 11969 6326 12003 6360
rect 12003 6326 12037 6360
rect 12037 6326 12071 6360
rect 12071 6326 12105 6360
rect 12105 6326 12139 6360
rect 12139 6326 12173 6360
rect 12173 6326 12207 6360
rect 12207 6326 12241 6360
rect 12241 6326 12275 6360
rect 12275 6326 12309 6360
rect 12309 6326 12343 6360
rect 12343 6326 12377 6360
rect 12377 6326 12411 6360
rect 12411 6326 12445 6360
rect 12445 6326 12479 6360
rect 12479 6326 12513 6360
rect 12513 6326 12547 6360
rect 12547 6326 12581 6360
rect 12581 6326 12615 6360
rect 12615 6326 12649 6360
rect 12649 6326 12683 6360
rect 12683 6326 12717 6360
rect 12717 6326 12751 6360
rect 12751 6326 12785 6360
rect 12785 6326 12819 6360
rect 12819 6326 12853 6360
rect 12853 6326 12887 6360
rect 12887 6326 12921 6360
rect 12921 6326 12955 6360
rect 12955 6326 12989 6360
rect 12989 6326 13023 6360
rect 13023 6326 13057 6360
rect 13057 6326 13091 6360
rect 13091 6326 13125 6360
rect 13125 6326 13159 6360
rect 13159 6326 13193 6360
rect 13193 6326 13227 6360
rect 13227 6326 13261 6360
rect 13261 6326 13295 6360
rect 13295 6326 13329 6360
rect 13329 6326 13363 6360
rect 13363 6326 13397 6360
rect 13397 6326 13431 6360
rect 13431 6326 13465 6360
rect 13465 6326 13499 6360
rect 13499 6326 13533 6360
rect 13533 6326 13567 6360
rect 13567 6326 13601 6360
rect 13601 6326 13635 6360
rect 13635 6326 13669 6360
rect 13669 6326 13703 6360
rect 13703 6326 13737 6360
rect 13737 6326 13771 6360
rect 13771 6326 13805 6360
rect 13805 6326 13839 6360
rect 13839 6326 13873 6360
rect 13873 6326 13907 6360
rect 13907 6326 13941 6360
rect 13941 6326 13975 6360
rect 13975 6326 14009 6360
rect 14009 6326 14043 6360
rect 14043 6326 14077 6360
rect 14077 6326 14111 6360
rect 14111 6326 14145 6360
rect 14145 6326 14179 6360
rect 14179 6326 14213 6360
rect 14213 6326 14247 6360
rect 14247 6326 14281 6360
rect 14281 6326 14315 6360
rect 14315 6326 14349 6360
rect 14349 6326 14383 6360
rect 14383 6326 14417 6360
rect 14417 6326 14451 6360
rect 14451 6326 14485 6360
rect 14485 6326 14519 6360
rect 14519 6326 14553 6360
rect 14553 6326 14587 6360
rect 14587 6326 14621 6360
rect 14621 6326 14655 6360
rect 14655 6326 14689 6360
rect 14689 6326 14723 6360
rect 14723 6326 14757 6360
rect 14757 6326 14791 6360
rect 14791 6326 14825 6360
rect 14825 6326 14859 6360
rect 14859 6326 14893 6360
rect 14893 6326 14932 6360
rect 14932 6326 14966 6360
rect 14966 6326 15000 6360
rect 15000 6326 15020 6360
rect 15068 6359 15102 6360
rect 68 6286 102 6295
rect 141 6286 175 6295
rect 214 6286 248 6295
rect 287 6286 321 6295
rect 360 6286 394 6295
rect 433 6286 467 6295
rect 506 6286 540 6295
rect 579 6286 613 6295
rect 652 6286 686 6295
rect 725 6286 759 6295
rect 798 6286 832 6295
rect 871 6286 905 6295
rect 944 6286 978 6295
rect 1017 6286 1051 6295
rect 1090 6286 15020 6326
rect 15068 6287 15102 6321
rect 68 6261 102 6286
rect 141 6261 171 6286
rect 171 6261 175 6286
rect 214 6261 240 6286
rect 240 6261 248 6286
rect 287 6261 309 6286
rect 309 6261 321 6286
rect 360 6261 378 6286
rect 378 6261 394 6286
rect 433 6261 447 6286
rect 447 6261 467 6286
rect 506 6261 516 6286
rect 516 6261 540 6286
rect 579 6261 585 6286
rect 585 6261 613 6286
rect 652 6261 654 6286
rect 654 6261 686 6286
rect 725 6261 758 6286
rect 758 6261 759 6286
rect 798 6261 827 6286
rect 827 6261 832 6286
rect 871 6261 896 6286
rect 896 6261 905 6286
rect 944 6261 965 6286
rect 965 6261 978 6286
rect 1017 6261 1034 6286
rect 1034 6261 1051 6286
rect 1090 6252 1103 6286
rect 1103 6252 1137 6286
rect 1137 6252 1172 6286
rect 1172 6252 1206 6286
rect 1206 6252 1241 6286
rect 1241 6252 1275 6286
rect 1275 6252 1310 6286
rect 1310 6252 1344 6286
rect 1344 6252 1379 6286
rect 1379 6252 1413 6286
rect 1413 6252 1448 6286
rect 1448 6252 1482 6286
rect 1482 6252 1517 6286
rect 1517 6252 1551 6286
rect 1551 6252 1586 6286
rect 1586 6252 1620 6286
rect 1620 6252 1655 6286
rect 1655 6252 1689 6286
rect 1689 6252 1724 6286
rect 1724 6252 1758 6286
rect 1758 6252 1793 6286
rect 1793 6252 1827 6286
rect 1827 6252 1862 6286
rect 1862 6252 1896 6286
rect 1896 6252 1931 6286
rect 1931 6252 1965 6286
rect 1965 6252 2000 6286
rect 2000 6252 2034 6286
rect 2034 6252 2069 6286
rect 2069 6252 2103 6286
rect 2103 6252 2138 6286
rect 2138 6252 2172 6286
rect 2172 6252 2207 6286
rect 2207 6252 2241 6286
rect 2241 6252 2276 6286
rect 2276 6252 2310 6286
rect 2310 6252 2345 6286
rect 2345 6252 2379 6286
rect 2379 6252 2414 6286
rect 2414 6252 2448 6286
rect 2448 6252 2483 6286
rect 2483 6252 2517 6286
rect 2517 6252 2551 6286
rect 2551 6252 2585 6286
rect 2585 6252 2619 6286
rect 2619 6252 2653 6286
rect 2653 6252 2687 6286
rect 2687 6252 2721 6286
rect 2721 6252 2755 6286
rect 2755 6252 2789 6286
rect 2789 6252 2823 6286
rect 2823 6252 2857 6286
rect 2857 6252 2891 6286
rect 2891 6252 2925 6286
rect 2925 6252 2959 6286
rect 2959 6252 2993 6286
rect 2993 6252 3027 6286
rect 3027 6252 3061 6286
rect 3061 6252 3095 6286
rect 3095 6252 3129 6286
rect 3129 6252 3163 6286
rect 3163 6252 3197 6286
rect 3197 6252 3231 6286
rect 3231 6252 3265 6286
rect 3265 6252 3299 6286
rect 3299 6252 3333 6286
rect 3333 6252 3367 6286
rect 3367 6252 3401 6286
rect 3401 6252 3435 6286
rect 3435 6252 3469 6286
rect 3469 6252 3503 6286
rect 3503 6252 3537 6286
rect 3537 6252 3571 6286
rect 3571 6252 3605 6286
rect 3605 6252 3639 6286
rect 3639 6252 3673 6286
rect 3673 6252 3707 6286
rect 3707 6252 3741 6286
rect 3741 6252 3775 6286
rect 3775 6252 3809 6286
rect 3809 6252 3843 6286
rect 3843 6252 3877 6286
rect 3877 6252 3911 6286
rect 3911 6252 3945 6286
rect 3945 6252 3979 6286
rect 3979 6252 4013 6286
rect 4013 6252 4047 6286
rect 4047 6252 4081 6286
rect 4081 6252 4115 6286
rect 4115 6252 4149 6286
rect 4149 6252 4183 6286
rect 4183 6252 4217 6286
rect 4217 6252 4251 6286
rect 4251 6252 4285 6286
rect 4285 6252 4319 6286
rect 4319 6252 4353 6286
rect 4353 6252 4387 6286
rect 4387 6252 4421 6286
rect 4421 6252 4455 6286
rect 4455 6252 4489 6286
rect 4489 6252 4523 6286
rect 4523 6252 4557 6286
rect 4557 6252 4591 6286
rect 4591 6252 4625 6286
rect 4625 6252 4659 6286
rect 4659 6252 4693 6286
rect 4693 6252 4727 6286
rect 4727 6252 4761 6286
rect 4761 6252 4795 6286
rect 4795 6252 4829 6286
rect 4829 6252 4863 6286
rect 4863 6252 4897 6286
rect 4897 6252 4931 6286
rect 4931 6252 4965 6286
rect 4965 6252 4999 6286
rect 4999 6252 5033 6286
rect 5033 6252 5067 6286
rect 5067 6252 5101 6286
rect 5101 6252 5135 6286
rect 5135 6252 5169 6286
rect 5169 6252 5203 6286
rect 5203 6252 5237 6286
rect 5237 6252 5271 6286
rect 5271 6252 5305 6286
rect 5305 6252 5339 6286
rect 5339 6252 5373 6286
rect 5373 6252 5407 6286
rect 5407 6252 5441 6286
rect 5441 6252 5475 6286
rect 5475 6252 5509 6286
rect 5509 6252 5543 6286
rect 5543 6252 5577 6286
rect 5577 6252 5611 6286
rect 5611 6252 5645 6286
rect 5645 6252 5679 6286
rect 5679 6252 5713 6286
rect 5713 6252 5747 6286
rect 5747 6252 5781 6286
rect 5781 6252 5815 6286
rect 5815 6252 5849 6286
rect 5849 6252 5883 6286
rect 5883 6252 5917 6286
rect 5917 6252 5951 6286
rect 5951 6252 5985 6286
rect 5985 6252 6019 6286
rect 6019 6252 6053 6286
rect 6053 6252 6087 6286
rect 6087 6252 6121 6286
rect 6121 6252 6155 6286
rect 6155 6252 6189 6286
rect 6189 6252 6223 6286
rect 6223 6252 6257 6286
rect 6257 6252 6291 6286
rect 6291 6252 6325 6286
rect 6325 6252 6359 6286
rect 6359 6252 6393 6286
rect 6393 6252 6427 6286
rect 6427 6252 6461 6286
rect 6461 6252 6495 6286
rect 6495 6252 6529 6286
rect 6529 6252 6563 6286
rect 6563 6252 6597 6286
rect 6597 6252 6631 6286
rect 6631 6252 6665 6286
rect 6665 6252 6699 6286
rect 6699 6252 6733 6286
rect 6733 6252 6767 6286
rect 6767 6252 6801 6286
rect 6801 6252 6835 6286
rect 6835 6252 6869 6286
rect 6869 6252 6903 6286
rect 6903 6252 6937 6286
rect 6937 6252 6971 6286
rect 6971 6252 7005 6286
rect 7005 6252 7039 6286
rect 7039 6252 7073 6286
rect 7073 6252 7107 6286
rect 7107 6252 7141 6286
rect 7141 6252 7175 6286
rect 7175 6252 7209 6286
rect 7209 6252 7243 6286
rect 7243 6252 7277 6286
rect 7277 6252 7311 6286
rect 7311 6252 7345 6286
rect 7345 6252 7379 6286
rect 7379 6252 7413 6286
rect 7413 6252 7447 6286
rect 7447 6252 7481 6286
rect 7481 6252 7515 6286
rect 7515 6252 7549 6286
rect 7549 6252 7583 6286
rect 7583 6252 7617 6286
rect 7617 6252 7651 6286
rect 7651 6252 7685 6286
rect 7685 6252 7719 6286
rect 7719 6252 7753 6286
rect 7753 6252 7787 6286
rect 7787 6252 7821 6286
rect 7821 6252 7855 6286
rect 7855 6252 7889 6286
rect 7889 6252 7923 6286
rect 7923 6252 7957 6286
rect 7957 6252 7991 6286
rect 7991 6252 8025 6286
rect 8025 6252 8059 6286
rect 8059 6252 8093 6286
rect 8093 6252 8127 6286
rect 8127 6252 8161 6286
rect 8161 6252 8195 6286
rect 8195 6252 8229 6286
rect 8229 6252 8263 6286
rect 8263 6252 8297 6286
rect 8297 6252 8331 6286
rect 8331 6252 8365 6286
rect 8365 6252 8399 6286
rect 8399 6252 8433 6286
rect 8433 6252 8467 6286
rect 8467 6252 8501 6286
rect 8501 6252 8535 6286
rect 8535 6252 8569 6286
rect 8569 6252 8603 6286
rect 8603 6252 8637 6286
rect 8637 6252 8671 6286
rect 8671 6252 8705 6286
rect 8705 6252 8739 6286
rect 8739 6252 8773 6286
rect 8773 6252 8807 6286
rect 8807 6252 8841 6286
rect 8841 6252 8875 6286
rect 8875 6252 8909 6286
rect 8909 6252 8943 6286
rect 8943 6252 8977 6286
rect 8977 6252 9011 6286
rect 9011 6252 9045 6286
rect 9045 6252 9079 6286
rect 9079 6252 9113 6286
rect 9113 6252 9147 6286
rect 9147 6252 9181 6286
rect 9181 6252 9215 6286
rect 9215 6252 9249 6286
rect 9249 6252 9283 6286
rect 9283 6252 9317 6286
rect 9317 6252 9351 6286
rect 9351 6252 9385 6286
rect 9385 6252 9419 6286
rect 9419 6252 9453 6286
rect 9453 6252 9487 6286
rect 9487 6252 9521 6286
rect 9521 6252 9555 6286
rect 9555 6252 9589 6286
rect 9589 6252 9623 6286
rect 9623 6252 9657 6286
rect 9657 6252 9691 6286
rect 9691 6252 9725 6286
rect 9725 6252 9759 6286
rect 9759 6252 9793 6286
rect 9793 6252 9827 6286
rect 9827 6252 9861 6286
rect 9861 6252 9895 6286
rect 9895 6252 9929 6286
rect 9929 6252 9963 6286
rect 9963 6252 9997 6286
rect 9997 6252 10031 6286
rect 10031 6252 10065 6286
rect 10065 6252 10099 6286
rect 10099 6252 10133 6286
rect 10133 6252 10167 6286
rect 10167 6252 10201 6286
rect 10201 6252 10235 6286
rect 10235 6252 10269 6286
rect 10269 6252 10303 6286
rect 10303 6252 10337 6286
rect 10337 6252 10371 6286
rect 10371 6252 10405 6286
rect 10405 6252 10439 6286
rect 10439 6252 10473 6286
rect 10473 6252 10507 6286
rect 10507 6252 10541 6286
rect 10541 6252 10575 6286
rect 10575 6252 10609 6286
rect 10609 6252 10643 6286
rect 10643 6252 10677 6286
rect 10677 6252 10711 6286
rect 10711 6252 10745 6286
rect 10745 6252 10779 6286
rect 10779 6252 10813 6286
rect 10813 6252 10847 6286
rect 10847 6252 10881 6286
rect 10881 6252 10915 6286
rect 10915 6252 10949 6286
rect 10949 6252 10983 6286
rect 10983 6252 11017 6286
rect 11017 6252 11051 6286
rect 11051 6252 11085 6286
rect 11085 6252 11119 6286
rect 11119 6252 11153 6286
rect 11153 6252 11187 6286
rect 11187 6252 11221 6286
rect 11221 6252 11255 6286
rect 11255 6252 11289 6286
rect 11289 6252 11323 6286
rect 11323 6252 11357 6286
rect 11357 6252 11391 6286
rect 11391 6252 11425 6286
rect 11425 6252 11459 6286
rect 11459 6252 11493 6286
rect 11493 6252 11527 6286
rect 11527 6252 11561 6286
rect 11561 6252 11595 6286
rect 11595 6252 11629 6286
rect 11629 6252 11663 6286
rect 11663 6252 11697 6286
rect 11697 6252 11731 6286
rect 11731 6252 11765 6286
rect 11765 6252 11799 6286
rect 11799 6252 11833 6286
rect 11833 6252 11867 6286
rect 11867 6252 11901 6286
rect 11901 6252 11935 6286
rect 11935 6252 11969 6286
rect 11969 6252 12003 6286
rect 12003 6252 12037 6286
rect 12037 6252 12071 6286
rect 12071 6252 12105 6286
rect 12105 6252 12139 6286
rect 12139 6252 12173 6286
rect 12173 6252 12207 6286
rect 12207 6252 12241 6286
rect 12241 6252 12275 6286
rect 12275 6252 12309 6286
rect 12309 6252 12343 6286
rect 12343 6252 12377 6286
rect 12377 6252 12411 6286
rect 12411 6252 12445 6286
rect 12445 6252 12479 6286
rect 12479 6252 12513 6286
rect 12513 6252 12547 6286
rect 12547 6252 12581 6286
rect 12581 6252 12615 6286
rect 12615 6252 12649 6286
rect 12649 6252 12683 6286
rect 12683 6252 12717 6286
rect 12717 6252 12751 6286
rect 12751 6252 12785 6286
rect 12785 6252 12819 6286
rect 12819 6252 12853 6286
rect 12853 6252 12887 6286
rect 12887 6252 12921 6286
rect 12921 6252 12955 6286
rect 12955 6252 12989 6286
rect 12989 6252 13023 6286
rect 13023 6252 13057 6286
rect 13057 6252 13091 6286
rect 13091 6252 13125 6286
rect 13125 6252 13159 6286
rect 13159 6252 13193 6286
rect 13193 6252 13227 6286
rect 13227 6252 13261 6286
rect 13261 6252 13295 6286
rect 13295 6252 13329 6286
rect 13329 6252 13363 6286
rect 13363 6252 13397 6286
rect 13397 6252 13431 6286
rect 13431 6252 13465 6286
rect 13465 6252 13499 6286
rect 13499 6252 13533 6286
rect 13533 6252 13567 6286
rect 13567 6252 13601 6286
rect 13601 6252 13635 6286
rect 13635 6252 13669 6286
rect 13669 6252 13703 6286
rect 13703 6252 13737 6286
rect 13737 6252 13771 6286
rect 13771 6252 13805 6286
rect 13805 6252 13839 6286
rect 13839 6252 13873 6286
rect 13873 6252 13907 6286
rect 13907 6252 13941 6286
rect 13941 6252 13975 6286
rect 13975 6252 14009 6286
rect 14009 6252 14043 6286
rect 14043 6252 14077 6286
rect 14077 6252 14111 6286
rect 14111 6252 14145 6286
rect 14145 6252 14179 6286
rect 14179 6252 14213 6286
rect 14213 6252 14247 6286
rect 14247 6252 14281 6286
rect 14281 6252 14315 6286
rect 14315 6252 14349 6286
rect 14349 6252 14383 6286
rect 14383 6252 14417 6286
rect 14417 6252 14451 6286
rect 14451 6252 14485 6286
rect 14485 6252 14519 6286
rect 14519 6252 14553 6286
rect 14553 6252 14587 6286
rect 14587 6252 14621 6286
rect 14621 6252 14655 6286
rect 14655 6252 14689 6286
rect 14689 6252 14723 6286
rect 14723 6252 14757 6286
rect 14757 6252 14791 6286
rect 14791 6252 14825 6286
rect 14825 6252 14859 6286
rect 14859 6252 14893 6286
rect 14893 6285 15020 6286
rect 14893 6252 14932 6285
rect 1090 6251 14932 6252
rect 14932 6251 14966 6285
rect 14966 6251 15000 6285
rect 15000 6251 15020 6285
rect 68 6212 102 6223
rect 141 6212 175 6223
rect 214 6212 248 6223
rect 287 6212 321 6223
rect 360 6212 394 6223
rect 433 6212 467 6223
rect 506 6212 540 6223
rect 579 6212 613 6223
rect 652 6212 686 6223
rect 725 6212 759 6223
rect 798 6212 832 6223
rect 871 6212 905 6223
rect 944 6212 978 6223
rect 1017 6212 1051 6223
rect 1090 6212 15020 6251
rect 15068 6215 15102 6249
rect 68 6189 102 6212
rect 141 6189 171 6212
rect 171 6189 175 6212
rect 214 6189 240 6212
rect 240 6189 248 6212
rect 287 6189 309 6212
rect 309 6189 321 6212
rect 360 6189 378 6212
rect 378 6189 394 6212
rect 433 6189 447 6212
rect 447 6189 467 6212
rect 506 6189 516 6212
rect 516 6189 540 6212
rect 579 6189 585 6212
rect 585 6189 613 6212
rect 652 6189 654 6212
rect 654 6189 686 6212
rect 725 6189 758 6212
rect 758 6189 759 6212
rect 798 6189 827 6212
rect 827 6189 832 6212
rect 871 6189 896 6212
rect 896 6189 905 6212
rect 944 6189 965 6212
rect 965 6189 978 6212
rect 1017 6189 1034 6212
rect 1034 6189 1051 6212
rect 1090 6178 1103 6212
rect 1103 6178 1137 6212
rect 1137 6178 1172 6212
rect 1172 6178 1206 6212
rect 1206 6178 1241 6212
rect 1241 6178 1275 6212
rect 1275 6178 1310 6212
rect 1310 6178 1344 6212
rect 1344 6178 1379 6212
rect 1379 6178 1413 6212
rect 1413 6178 1448 6212
rect 1448 6178 1482 6212
rect 1482 6178 1517 6212
rect 1517 6178 1551 6212
rect 1551 6178 1586 6212
rect 1586 6178 1620 6212
rect 1620 6178 1655 6212
rect 1655 6178 1689 6212
rect 1689 6178 1724 6212
rect 1724 6178 1758 6212
rect 1758 6178 1793 6212
rect 1793 6178 1827 6212
rect 1827 6178 1862 6212
rect 1862 6178 1896 6212
rect 1896 6178 1931 6212
rect 1931 6178 1965 6212
rect 1965 6178 2000 6212
rect 2000 6178 2034 6212
rect 2034 6178 2069 6212
rect 2069 6178 2103 6212
rect 2103 6178 2138 6212
rect 2138 6178 2172 6212
rect 2172 6178 2207 6212
rect 2207 6178 2241 6212
rect 2241 6178 2276 6212
rect 2276 6178 2310 6212
rect 2310 6178 2345 6212
rect 2345 6178 2379 6212
rect 2379 6178 2414 6212
rect 2414 6178 2448 6212
rect 2448 6178 2483 6212
rect 2483 6178 2517 6212
rect 2517 6178 2551 6212
rect 2551 6178 2585 6212
rect 2585 6178 2619 6212
rect 2619 6178 2653 6212
rect 2653 6178 2687 6212
rect 2687 6178 2721 6212
rect 2721 6178 2755 6212
rect 2755 6178 2789 6212
rect 2789 6178 2823 6212
rect 2823 6178 2857 6212
rect 2857 6178 2891 6212
rect 2891 6178 2925 6212
rect 2925 6178 2959 6212
rect 2959 6178 2993 6212
rect 2993 6178 3027 6212
rect 3027 6178 3061 6212
rect 3061 6178 3095 6212
rect 3095 6178 3129 6212
rect 3129 6178 3163 6212
rect 3163 6178 3197 6212
rect 3197 6178 3231 6212
rect 3231 6178 3265 6212
rect 3265 6178 3299 6212
rect 3299 6178 3333 6212
rect 3333 6178 3367 6212
rect 3367 6178 3401 6212
rect 3401 6178 3435 6212
rect 3435 6178 3469 6212
rect 3469 6178 3503 6212
rect 3503 6178 3537 6212
rect 3537 6178 3571 6212
rect 3571 6178 3605 6212
rect 3605 6178 3639 6212
rect 3639 6178 3673 6212
rect 3673 6178 3707 6212
rect 3707 6178 3741 6212
rect 3741 6178 3775 6212
rect 3775 6178 3809 6212
rect 3809 6178 3843 6212
rect 3843 6178 3877 6212
rect 3877 6178 3911 6212
rect 3911 6178 3945 6212
rect 3945 6178 3979 6212
rect 3979 6178 4013 6212
rect 4013 6178 4047 6212
rect 4047 6178 4081 6212
rect 4081 6178 4115 6212
rect 4115 6178 4149 6212
rect 4149 6178 4183 6212
rect 4183 6178 4217 6212
rect 4217 6178 4251 6212
rect 4251 6178 4285 6212
rect 4285 6178 4319 6212
rect 4319 6178 4353 6212
rect 4353 6178 4387 6212
rect 4387 6178 4421 6212
rect 4421 6178 4455 6212
rect 4455 6178 4489 6212
rect 4489 6178 4523 6212
rect 4523 6178 4557 6212
rect 4557 6178 4591 6212
rect 4591 6178 4625 6212
rect 4625 6178 4659 6212
rect 4659 6178 4693 6212
rect 4693 6178 4727 6212
rect 4727 6178 4761 6212
rect 4761 6178 4795 6212
rect 4795 6178 4829 6212
rect 4829 6178 4863 6212
rect 4863 6178 4897 6212
rect 4897 6178 4931 6212
rect 4931 6178 4965 6212
rect 4965 6178 4999 6212
rect 4999 6178 5033 6212
rect 5033 6178 5067 6212
rect 5067 6178 5101 6212
rect 5101 6178 5135 6212
rect 5135 6178 5169 6212
rect 5169 6178 5203 6212
rect 5203 6178 5237 6212
rect 5237 6178 5271 6212
rect 5271 6178 5305 6212
rect 5305 6178 5339 6212
rect 5339 6178 5373 6212
rect 5373 6178 5407 6212
rect 5407 6178 5441 6212
rect 5441 6178 5475 6212
rect 5475 6178 5509 6212
rect 5509 6178 5543 6212
rect 5543 6178 5577 6212
rect 5577 6178 5611 6212
rect 5611 6178 5645 6212
rect 5645 6178 5679 6212
rect 5679 6178 5713 6212
rect 5713 6178 5747 6212
rect 5747 6178 5781 6212
rect 5781 6178 5815 6212
rect 5815 6178 5849 6212
rect 5849 6178 5883 6212
rect 5883 6178 5917 6212
rect 5917 6178 5951 6212
rect 5951 6178 5985 6212
rect 5985 6178 6019 6212
rect 6019 6178 6053 6212
rect 6053 6178 6087 6212
rect 6087 6178 6121 6212
rect 6121 6178 6155 6212
rect 6155 6178 6189 6212
rect 6189 6178 6223 6212
rect 6223 6178 6257 6212
rect 6257 6178 6291 6212
rect 6291 6178 6325 6212
rect 6325 6178 6359 6212
rect 6359 6178 6393 6212
rect 6393 6178 6427 6212
rect 6427 6178 6461 6212
rect 6461 6178 6495 6212
rect 6495 6178 6529 6212
rect 6529 6178 6563 6212
rect 6563 6178 6597 6212
rect 6597 6178 6631 6212
rect 6631 6178 6665 6212
rect 6665 6178 6699 6212
rect 6699 6178 6733 6212
rect 6733 6178 6767 6212
rect 6767 6178 6801 6212
rect 6801 6178 6835 6212
rect 6835 6178 6869 6212
rect 6869 6178 6903 6212
rect 6903 6178 6937 6212
rect 6937 6178 6971 6212
rect 6971 6178 7005 6212
rect 7005 6178 7039 6212
rect 7039 6178 7073 6212
rect 7073 6178 7107 6212
rect 7107 6178 7141 6212
rect 7141 6178 7175 6212
rect 7175 6178 7209 6212
rect 7209 6178 7243 6212
rect 7243 6178 7277 6212
rect 7277 6178 7311 6212
rect 7311 6178 7345 6212
rect 7345 6178 7379 6212
rect 7379 6178 7413 6212
rect 7413 6178 7447 6212
rect 7447 6178 7481 6212
rect 7481 6178 7515 6212
rect 7515 6178 7549 6212
rect 7549 6178 7583 6212
rect 7583 6178 7617 6212
rect 7617 6178 7651 6212
rect 7651 6178 7685 6212
rect 7685 6178 7719 6212
rect 7719 6178 7753 6212
rect 7753 6178 7787 6212
rect 7787 6178 7821 6212
rect 7821 6178 7855 6212
rect 7855 6178 7889 6212
rect 7889 6178 7923 6212
rect 7923 6178 7957 6212
rect 7957 6178 7991 6212
rect 7991 6178 8025 6212
rect 8025 6178 8059 6212
rect 8059 6178 8093 6212
rect 8093 6178 8127 6212
rect 8127 6178 8161 6212
rect 8161 6178 8195 6212
rect 8195 6178 8229 6212
rect 8229 6178 8263 6212
rect 8263 6178 8297 6212
rect 8297 6178 8331 6212
rect 8331 6178 8365 6212
rect 8365 6178 8399 6212
rect 8399 6178 8433 6212
rect 8433 6178 8467 6212
rect 8467 6178 8501 6212
rect 8501 6178 8535 6212
rect 8535 6178 8569 6212
rect 8569 6178 8603 6212
rect 8603 6178 8637 6212
rect 8637 6178 8671 6212
rect 8671 6178 8705 6212
rect 8705 6178 8739 6212
rect 8739 6178 8773 6212
rect 8773 6178 8807 6212
rect 8807 6178 8841 6212
rect 8841 6178 8875 6212
rect 8875 6178 8909 6212
rect 8909 6178 8943 6212
rect 8943 6178 8977 6212
rect 8977 6178 9011 6212
rect 9011 6178 9045 6212
rect 9045 6178 9079 6212
rect 9079 6178 9113 6212
rect 9113 6178 9147 6212
rect 9147 6178 9181 6212
rect 9181 6178 9215 6212
rect 9215 6178 9249 6212
rect 9249 6178 9283 6212
rect 9283 6178 9317 6212
rect 9317 6178 9351 6212
rect 9351 6178 9385 6212
rect 9385 6178 9419 6212
rect 9419 6178 9453 6212
rect 9453 6178 9487 6212
rect 9487 6178 9521 6212
rect 9521 6178 9555 6212
rect 9555 6178 9589 6212
rect 9589 6178 9623 6212
rect 9623 6178 9657 6212
rect 9657 6178 9691 6212
rect 9691 6178 9725 6212
rect 9725 6178 9759 6212
rect 9759 6178 9793 6212
rect 9793 6178 9827 6212
rect 9827 6178 9861 6212
rect 9861 6178 9895 6212
rect 9895 6178 9929 6212
rect 9929 6178 9963 6212
rect 9963 6178 9997 6212
rect 9997 6178 10031 6212
rect 10031 6178 10065 6212
rect 10065 6178 10099 6212
rect 10099 6178 10133 6212
rect 10133 6178 10167 6212
rect 10167 6178 10201 6212
rect 10201 6178 10235 6212
rect 10235 6178 10269 6212
rect 10269 6178 10303 6212
rect 10303 6178 10337 6212
rect 10337 6178 10371 6212
rect 10371 6178 10405 6212
rect 10405 6178 10439 6212
rect 10439 6178 10473 6212
rect 10473 6178 10507 6212
rect 10507 6178 10541 6212
rect 10541 6178 10575 6212
rect 10575 6178 10609 6212
rect 10609 6178 10643 6212
rect 10643 6178 10677 6212
rect 10677 6178 10711 6212
rect 10711 6178 10745 6212
rect 10745 6178 10779 6212
rect 10779 6178 10813 6212
rect 10813 6178 10847 6212
rect 10847 6178 10881 6212
rect 10881 6178 10915 6212
rect 10915 6178 10949 6212
rect 10949 6178 10983 6212
rect 10983 6178 11017 6212
rect 11017 6178 11051 6212
rect 11051 6178 11085 6212
rect 11085 6178 11119 6212
rect 11119 6178 11153 6212
rect 11153 6178 11187 6212
rect 11187 6178 11221 6212
rect 11221 6178 11255 6212
rect 11255 6178 11289 6212
rect 11289 6178 11323 6212
rect 11323 6178 11357 6212
rect 11357 6178 11391 6212
rect 11391 6178 11425 6212
rect 11425 6178 11459 6212
rect 11459 6178 11493 6212
rect 11493 6178 11527 6212
rect 11527 6178 11561 6212
rect 11561 6178 11595 6212
rect 11595 6178 11629 6212
rect 11629 6178 11663 6212
rect 11663 6178 11697 6212
rect 11697 6178 11731 6212
rect 11731 6178 11765 6212
rect 11765 6178 11799 6212
rect 11799 6178 11833 6212
rect 11833 6178 11867 6212
rect 11867 6178 11901 6212
rect 11901 6178 11935 6212
rect 11935 6178 11969 6212
rect 11969 6178 12003 6212
rect 12003 6178 12037 6212
rect 12037 6178 12071 6212
rect 12071 6178 12105 6212
rect 12105 6178 12139 6212
rect 12139 6178 12173 6212
rect 12173 6178 12207 6212
rect 12207 6178 12241 6212
rect 12241 6178 12275 6212
rect 12275 6178 12309 6212
rect 12309 6178 12343 6212
rect 12343 6178 12377 6212
rect 12377 6178 12411 6212
rect 12411 6178 12445 6212
rect 12445 6178 12479 6212
rect 12479 6178 12513 6212
rect 12513 6178 12547 6212
rect 12547 6178 12581 6212
rect 12581 6178 12615 6212
rect 12615 6178 12649 6212
rect 12649 6178 12683 6212
rect 12683 6178 12717 6212
rect 12717 6178 12751 6212
rect 12751 6178 12785 6212
rect 12785 6178 12819 6212
rect 12819 6178 12853 6212
rect 12853 6178 12887 6212
rect 12887 6178 12921 6212
rect 12921 6178 12955 6212
rect 12955 6178 12989 6212
rect 12989 6178 13023 6212
rect 13023 6178 13057 6212
rect 13057 6178 13091 6212
rect 13091 6178 13125 6212
rect 13125 6178 13159 6212
rect 13159 6178 13193 6212
rect 13193 6178 13227 6212
rect 13227 6178 13261 6212
rect 13261 6178 13295 6212
rect 13295 6178 13329 6212
rect 13329 6178 13363 6212
rect 13363 6178 13397 6212
rect 13397 6178 13431 6212
rect 13431 6178 13465 6212
rect 13465 6178 13499 6212
rect 13499 6178 13533 6212
rect 13533 6178 13567 6212
rect 13567 6178 13601 6212
rect 13601 6178 13635 6212
rect 13635 6178 13669 6212
rect 13669 6178 13703 6212
rect 13703 6178 13737 6212
rect 13737 6178 13771 6212
rect 13771 6178 13805 6212
rect 13805 6178 13839 6212
rect 13839 6178 13873 6212
rect 13873 6178 13907 6212
rect 13907 6178 13941 6212
rect 13941 6178 13975 6212
rect 13975 6178 14009 6212
rect 14009 6178 14043 6212
rect 14043 6178 14077 6212
rect 14077 6178 14111 6212
rect 14111 6178 14145 6212
rect 14145 6178 14179 6212
rect 14179 6178 14213 6212
rect 14213 6178 14247 6212
rect 14247 6178 14281 6212
rect 14281 6178 14315 6212
rect 14315 6178 14349 6212
rect 14349 6178 14383 6212
rect 14383 6178 14417 6212
rect 14417 6178 14451 6212
rect 14451 6178 14485 6212
rect 14485 6178 14519 6212
rect 14519 6178 14553 6212
rect 14553 6178 14587 6212
rect 14587 6178 14621 6212
rect 14621 6178 14655 6212
rect 14655 6178 14689 6212
rect 14689 6178 14723 6212
rect 14723 6178 14757 6212
rect 14757 6178 14791 6212
rect 14791 6178 14825 6212
rect 14825 6178 14859 6212
rect 14859 6178 14893 6212
rect 14893 6210 15020 6212
rect 14893 6178 14932 6210
rect 1090 6176 14932 6178
rect 14932 6176 14966 6210
rect 14966 6176 15000 6210
rect 15000 6176 15020 6210
rect 15068 6176 15102 6177
rect 68 6138 102 6151
rect 141 6138 175 6151
rect 214 6138 248 6151
rect 287 6138 321 6151
rect 360 6138 394 6151
rect 433 6138 467 6151
rect 506 6138 540 6151
rect 579 6138 613 6151
rect 652 6138 686 6151
rect 725 6138 759 6151
rect 798 6138 832 6151
rect 871 6138 905 6151
rect 944 6138 978 6151
rect 1017 6138 1051 6151
rect 1090 6138 15020 6176
rect 15068 6143 15102 6176
rect 68 6117 102 6138
rect 141 6117 171 6138
rect 171 6117 175 6138
rect 214 6117 240 6138
rect 240 6117 248 6138
rect 287 6117 309 6138
rect 309 6117 321 6138
rect 360 6117 378 6138
rect 378 6117 394 6138
rect 433 6117 447 6138
rect 447 6117 467 6138
rect 506 6117 516 6138
rect 516 6117 540 6138
rect 579 6117 585 6138
rect 585 6117 613 6138
rect 652 6117 654 6138
rect 654 6117 686 6138
rect 725 6117 758 6138
rect 758 6117 759 6138
rect 798 6117 827 6138
rect 827 6117 832 6138
rect 871 6117 896 6138
rect 896 6117 905 6138
rect 944 6117 965 6138
rect 965 6117 978 6138
rect 1017 6117 1034 6138
rect 1034 6117 1051 6138
rect 1090 6117 1103 6138
rect 1103 6117 1137 6138
rect 1137 6117 1172 6138
rect 1172 6117 1206 6138
rect 1206 6117 1241 6138
rect 1241 6117 1275 6138
rect 1275 6117 1310 6138
rect 1310 6117 1344 6138
rect 1344 6117 1379 6138
rect 1379 6117 1413 6138
rect 1413 6117 1448 6138
rect 1448 6117 1482 6138
rect 1482 6117 1517 6138
rect 1517 6117 1551 6138
rect 1551 6117 1586 6138
rect 1586 6117 1620 6138
rect 1620 6117 1655 6138
rect 1655 6117 1689 6138
rect 1689 6117 1724 6138
rect 1724 6117 1758 6138
rect 1758 6117 1793 6138
rect 1793 6117 1827 6138
rect 1827 6117 1862 6138
rect 1862 6117 1896 6138
rect 1896 6117 1931 6138
rect 1931 6117 1965 6138
rect 1965 6117 2000 6138
rect 2000 6117 2034 6138
rect 2034 6117 2069 6138
rect 2069 6117 2103 6138
rect 2103 6117 2138 6138
rect 2138 6117 2172 6138
rect 2172 6117 2207 6138
rect 2207 6117 2241 6138
rect 2241 6117 2276 6138
rect 2276 6117 2310 6138
rect 2310 6117 2345 6138
rect 2345 6117 2379 6138
rect 2379 6117 2414 6138
rect 2414 6117 2448 6138
rect 2448 6117 2483 6138
rect 2483 6117 2517 6138
rect 2517 6117 2551 6138
rect 2551 6117 2585 6138
rect 2585 6117 2619 6138
rect 2619 6117 2653 6138
rect 2653 6117 2687 6138
rect 2687 6117 2721 6138
rect 2721 6117 2755 6138
rect 2755 6117 2789 6138
rect 2789 6117 2823 6138
rect 2823 6117 2857 6138
rect 2857 6117 2891 6138
rect 2891 6117 2925 6138
rect 2925 6117 2959 6138
rect 2959 6117 2993 6138
rect 2993 6117 3027 6138
rect 3027 6117 3061 6138
rect 3061 6117 3095 6138
rect 3095 6117 3129 6138
rect 3129 6117 3163 6138
rect 3163 6117 3197 6138
rect 3197 6117 3231 6138
rect 3231 6117 3265 6138
rect 3265 6117 3299 6138
rect 3299 6117 3333 6138
rect 3333 6117 3367 6138
rect 3367 6117 3401 6138
rect 3401 6117 3435 6138
rect 3435 6117 3469 6138
rect 3469 6117 3503 6138
rect 3503 6117 3537 6138
rect 3537 6117 3571 6138
rect 3571 6117 3605 6138
rect 3605 6117 3639 6138
rect 3639 6117 3673 6138
rect 3673 6117 3707 6138
rect 3707 6117 3741 6138
rect 3741 6117 3775 6138
rect 3775 6117 3809 6138
rect 3809 6117 3843 6138
rect 3843 6117 3877 6138
rect 3877 6117 3911 6138
rect 3911 6117 3945 6138
rect 3945 6117 3979 6138
rect 3979 6117 4013 6138
rect 4013 6117 4047 6138
rect 4047 6117 4081 6138
rect 4081 6117 4115 6138
rect 4115 6117 4149 6138
rect 4149 6117 4183 6138
rect 4183 6117 4217 6138
rect 4217 6117 4251 6138
rect 4251 6117 4285 6138
rect 4285 6117 4319 6138
rect 4319 6117 4353 6138
rect 4353 6117 4387 6138
rect 4387 6117 4421 6138
rect 4421 6117 4455 6138
rect 4455 6117 4489 6138
rect 4489 6117 4523 6138
rect 4523 6117 4557 6138
rect 4557 6117 4591 6138
rect 4591 6117 4625 6138
rect 4625 6117 4659 6138
rect 4659 6117 4693 6138
rect 4693 6117 4727 6138
rect 4727 6117 4761 6138
rect 4761 6117 4795 6138
rect 4795 6117 4829 6138
rect 4829 6117 4863 6138
rect 4863 6117 4897 6138
rect 4897 6117 4931 6138
rect 4931 6117 4965 6138
rect 4965 6117 4999 6138
rect 4999 6117 5033 6138
rect 5033 6117 5067 6138
rect 5067 6117 5101 6138
rect 5101 6117 5135 6138
rect 5135 6117 5169 6138
rect 5169 6117 5203 6138
rect 5203 6117 5237 6138
rect 5237 6117 5271 6138
rect 5271 6117 5305 6138
rect 5305 6117 5339 6138
rect 5339 6117 5373 6138
rect 5373 6117 5407 6138
rect 5407 6117 5441 6138
rect 5441 6117 5475 6138
rect 5475 6117 5509 6138
rect 5509 6117 5543 6138
rect 5543 6117 5577 6138
rect 5577 6117 5611 6138
rect 5611 6117 5645 6138
rect 5645 6117 5679 6138
rect 5679 6117 5713 6138
rect 5713 6117 5747 6138
rect 5747 6117 5781 6138
rect 5781 6117 5815 6138
rect 5815 6117 5849 6138
rect 5849 6117 5883 6138
rect 5883 6117 5917 6138
rect 5917 6117 5951 6138
rect 5951 6117 5985 6138
rect 5985 6117 6019 6138
rect 6019 6117 6053 6138
rect 6053 6117 6087 6138
rect 6087 6117 6121 6138
rect 6121 6117 6155 6138
rect 6155 6117 6189 6138
rect 6189 6117 6223 6138
rect 6223 6117 6257 6138
rect 6257 6117 6291 6138
rect 6291 6117 6325 6138
rect 6325 6117 6359 6138
rect 6359 6117 6393 6138
rect 6393 6117 6427 6138
rect 6427 6117 6461 6138
rect 6461 6117 6495 6138
rect 6495 6117 6529 6138
rect 6529 6117 6563 6138
rect 6563 6117 6597 6138
rect 6597 6117 6631 6138
rect 6631 6117 6665 6138
rect 6665 6117 6699 6138
rect 6699 6117 6733 6138
rect 6733 6117 6767 6138
rect 6767 6117 6801 6138
rect 6801 6117 6835 6138
rect 6835 6117 6869 6138
rect 6869 6117 6903 6138
rect 6903 6117 6937 6138
rect 6937 6117 6971 6138
rect 6971 6117 7005 6138
rect 7005 6117 7039 6138
rect 7039 6117 7073 6138
rect 7073 6117 7107 6138
rect 7107 6117 7141 6138
rect 7141 6117 7175 6138
rect 7175 6117 7209 6138
rect 7209 6117 7243 6138
rect 7243 6117 7277 6138
rect 7277 6117 7311 6138
rect 7311 6117 7345 6138
rect 7345 6117 7379 6138
rect 7379 6117 7413 6138
rect 7413 6117 7447 6138
rect 7447 6117 7481 6138
rect 7481 6117 7515 6138
rect 7515 6117 7549 6138
rect 7549 6117 7583 6138
rect 7583 6117 7617 6138
rect 7617 6117 7651 6138
rect 7651 6117 7685 6138
rect 7685 6117 7719 6138
rect 7719 6117 7753 6138
rect 7753 6117 7787 6138
rect 7787 6117 7821 6138
rect 7821 6117 7855 6138
rect 7855 6117 7889 6138
rect 7889 6117 7923 6138
rect 7923 6117 7957 6138
rect 7957 6117 7991 6138
rect 7991 6117 8025 6138
rect 8025 6117 8059 6138
rect 8059 6117 8093 6138
rect 8093 6117 8127 6138
rect 8127 6117 8161 6138
rect 8161 6117 8195 6138
rect 8195 6117 8229 6138
rect 8229 6117 8263 6138
rect 8263 6117 8297 6138
rect 8297 6117 8331 6138
rect 8331 6117 8365 6138
rect 8365 6117 8399 6138
rect 8399 6117 8433 6138
rect 8433 6117 8467 6138
rect 8467 6117 8501 6138
rect 8501 6117 8535 6138
rect 8535 6117 8569 6138
rect 8569 6117 8603 6138
rect 8603 6117 8637 6138
rect 8637 6117 8671 6138
rect 8671 6117 8705 6138
rect 8705 6117 8739 6138
rect 8739 6117 8773 6138
rect 8773 6117 8807 6138
rect 8807 6117 8841 6138
rect 8841 6117 8875 6138
rect 8875 6117 8909 6138
rect 8909 6117 8943 6138
rect 8943 6117 8977 6138
rect 8977 6117 9011 6138
rect 9011 6117 9045 6138
rect 9045 6117 9079 6138
rect 9079 6117 9113 6138
rect 9113 6117 9147 6138
rect 9147 6117 9181 6138
rect 9181 6117 9215 6138
rect 9215 6117 9249 6138
rect 9249 6117 9283 6138
rect 9283 6117 9317 6138
rect 9317 6117 9351 6138
rect 9351 6117 9385 6138
rect 9385 6117 9419 6138
rect 9419 6117 9453 6138
rect 9453 6117 9487 6138
rect 9487 6117 9521 6138
rect 9521 6117 9555 6138
rect 9555 6117 9589 6138
rect 9589 6117 9623 6138
rect 9623 6117 9657 6138
rect 9657 6117 9691 6138
rect 9691 6117 9725 6138
rect 9725 6117 9759 6138
rect 9759 6117 9793 6138
rect 9793 6117 9827 6138
rect 9827 6117 9861 6138
rect 9861 6117 9895 6138
rect 9895 6117 9929 6138
rect 9929 6117 9963 6138
rect 9963 6117 9997 6138
rect 9997 6117 10031 6138
rect 10031 6117 10065 6138
rect 10065 6117 10099 6138
rect 10099 6117 10133 6138
rect 10133 6117 10167 6138
rect 10167 6117 10201 6138
rect 10201 6117 10235 6138
rect 10235 6117 10269 6138
rect 10269 6117 10303 6138
rect 10303 6117 10337 6138
rect 10337 6117 10371 6138
rect 10371 6117 10405 6138
rect 10405 6117 10439 6138
rect 10439 6117 10473 6138
rect 10473 6117 10507 6138
rect 10507 6117 10541 6138
rect 10541 6117 10575 6138
rect 10575 6117 10609 6138
rect 10609 6117 10643 6138
rect 10643 6117 10677 6138
rect 10677 6117 10711 6138
rect 10711 6117 10745 6138
rect 10745 6117 10779 6138
rect 10779 6117 10813 6138
rect 10813 6117 10847 6138
rect 10847 6117 10881 6138
rect 10881 6117 10915 6138
rect 10915 6117 10949 6138
rect 10949 6117 10983 6138
rect 10983 6117 11017 6138
rect 11017 6117 11051 6138
rect 11051 6117 11085 6138
rect 11085 6117 11119 6138
rect 11119 6117 11153 6138
rect 11153 6117 11187 6138
rect 11187 6117 11221 6138
rect 11221 6117 11255 6138
rect 11255 6117 11289 6138
rect 11289 6117 11323 6138
rect 11323 6117 11357 6138
rect 11357 6117 11391 6138
rect 11391 6117 11425 6138
rect 11425 6117 11459 6138
rect 11459 6117 11493 6138
rect 11493 6117 11527 6138
rect 11527 6117 11561 6138
rect 11561 6117 11595 6138
rect 11595 6117 11629 6138
rect 11629 6117 11663 6138
rect 11663 6117 11697 6138
rect 11697 6117 11731 6138
rect 11731 6117 11765 6138
rect 11765 6117 11799 6138
rect 11799 6117 11833 6138
rect 11833 6117 11867 6138
rect 11867 6117 11901 6138
rect 11901 6117 11935 6138
rect 11935 6117 11969 6138
rect 11969 6117 12003 6138
rect 12003 6117 12037 6138
rect 12037 6117 12071 6138
rect 12071 6117 12105 6138
rect 12105 6117 12139 6138
rect 12139 6117 12173 6138
rect 12173 6117 12207 6138
rect 12207 6117 12241 6138
rect 12241 6117 12275 6138
rect 12275 6117 12309 6138
rect 12309 6117 12343 6138
rect 12343 6117 12377 6138
rect 12377 6117 12411 6138
rect 12411 6117 12445 6138
rect 12445 6117 12479 6138
rect 12479 6117 12513 6138
rect 12513 6117 12547 6138
rect 12547 6117 12581 6138
rect 12581 6117 12615 6138
rect 12615 6117 12649 6138
rect 12649 6117 12683 6138
rect 12683 6117 12717 6138
rect 12717 6117 12751 6138
rect 12751 6117 12785 6138
rect 12785 6117 12819 6138
rect 12819 6117 12853 6138
rect 12853 6117 12887 6138
rect 12887 6117 12921 6138
rect 12921 6117 12955 6138
rect 12955 6117 12989 6138
rect 12989 6117 13023 6138
rect 13023 6117 13057 6138
rect 13057 6117 13091 6138
rect 13091 6117 13125 6138
rect 13125 6117 13159 6138
rect 13159 6117 13193 6138
rect 13193 6117 13227 6138
rect 13227 6117 13261 6138
rect 13261 6117 13295 6138
rect 13295 6117 13329 6138
rect 13329 6117 13363 6138
rect 13363 6117 13397 6138
rect 13397 6117 13431 6138
rect 13431 6117 13465 6138
rect 13465 6117 13499 6138
rect 13499 6117 13533 6138
rect 13533 6117 13567 6138
rect 13567 6117 13601 6138
rect 13601 6117 13635 6138
rect 13635 6117 13669 6138
rect 13669 6117 13703 6138
rect 13703 6117 13737 6138
rect 13737 6117 13771 6138
rect 13771 6117 13805 6138
rect 13805 6117 13839 6138
rect 13839 6117 13873 6138
rect 13873 6117 13907 6138
rect 13907 6117 13941 6138
rect 13941 6117 13975 6138
rect 13975 6117 14009 6138
rect 14009 6117 14043 6138
rect 14043 6117 14077 6138
rect 14077 6117 14111 6138
rect 14111 6117 14145 6138
rect 14145 6117 14179 6138
rect 14179 6117 14213 6138
rect 14213 6117 14247 6138
rect 14247 6117 14281 6138
rect 14281 6117 14315 6138
rect 14315 6117 14349 6138
rect 14349 6117 14383 6138
rect 14383 6117 14417 6138
rect 14417 6117 14451 6138
rect 14451 6117 14485 6138
rect 14485 6117 14519 6138
rect 14519 6117 14553 6138
rect 14553 6117 14587 6138
rect 14587 6117 14621 6138
rect 14621 6117 14655 6138
rect 14655 6117 14689 6138
rect 14689 6117 14723 6138
rect 14723 6117 14757 6138
rect 14757 6117 14791 6138
rect 14791 6117 14825 6138
rect 14825 6117 14859 6138
rect 14859 6117 14893 6138
rect 14893 6135 15020 6138
rect 14893 6117 14932 6135
rect 14932 6117 14966 6135
rect 14966 6117 15000 6135
rect 15000 6117 15020 6135
rect 15068 6101 15102 6105
rect 15068 6071 15102 6101
rect 15068 6026 15102 6033
rect 15068 5999 15102 6026
rect 15068 5954 15102 5961
rect 15068 5927 15102 5954
rect 15068 5855 15102 5889
rect 15068 5783 15102 5817
rect 15068 5711 15102 5745
rect 15068 5639 15102 5673
rect 15068 5567 15102 5601
rect 15068 5495 15102 5529
rect 15068 5423 15102 5457
rect 15068 5351 15102 5385
rect 15068 5279 15102 5313
rect 15068 5207 15102 5241
rect 15068 5135 15102 5169
rect 15068 5063 15102 5097
rect 15068 4991 15102 5025
rect 15068 4919 15102 4953
rect 15068 4847 15102 4881
rect 15068 4775 15102 4809
rect 15068 4703 15102 4737
rect 15068 4631 15102 4665
rect 15068 4559 15102 4593
rect 15068 4490 15102 4521
rect 15068 4487 15102 4490
rect 15068 4421 15102 4449
rect 15068 4415 15102 4421
rect 15068 4352 15102 4377
rect 15068 4343 15102 4352
rect 15068 4283 15102 4305
rect 15068 4271 15102 4283
rect 15068 4214 15102 4233
rect 15068 4199 15102 4214
rect 15068 4145 15102 4161
rect 15068 4127 15102 4145
rect 15068 4076 15102 4089
rect 15068 4055 15102 4076
rect 15068 4007 15102 4017
rect 15068 3983 15102 4007
rect 15068 3938 15102 3945
rect 15068 3911 15102 3938
rect 15068 3869 15102 3873
rect 15068 3839 15102 3869
rect 15068 3800 15102 3801
rect 15068 3767 15102 3800
rect 15068 3696 15102 3729
rect 15068 3695 15102 3696
rect 15068 3627 15102 3657
rect 15068 3623 15102 3627
rect 15068 3558 15102 3585
rect 15068 3551 15102 3558
rect 15068 3489 15102 3513
rect 15068 3479 15102 3489
rect 15068 3420 15102 3441
rect 15068 3407 15102 3420
rect 15068 3351 15102 3369
rect 15068 3335 15102 3351
rect 15068 3282 15102 3297
rect 15068 3263 15102 3282
rect 15068 3213 15102 3225
rect 15068 3191 15102 3213
rect 15068 3144 15102 3153
rect 15068 3119 15102 3144
rect 15068 3075 15102 3081
rect 15068 3047 15102 3075
rect 15068 3006 15102 3009
rect 15068 2975 15102 3006
rect 15068 2903 15102 2937
rect 15068 2834 15102 2865
rect 15068 2831 15102 2834
rect 15068 2765 15102 2793
rect 15068 2759 15102 2765
rect 15068 2696 15102 2721
rect 15068 2687 15102 2696
rect 15068 2627 15102 2649
rect 15068 2615 15102 2627
rect 15068 2558 15102 2577
rect 15068 2543 15102 2558
rect 15068 2489 15102 2505
rect 15068 2471 15102 2489
rect 15068 2420 15102 2433
rect 15068 2399 15102 2420
rect 15068 2351 15102 2361
rect 15068 2327 15102 2351
rect 15068 2282 15102 2289
rect 15068 2255 15102 2282
rect 15068 2213 15102 2217
rect 15068 2183 15102 2213
rect 15068 2144 15102 2145
rect 15068 2111 15102 2144
rect 15068 2040 15102 2073
rect 15068 2039 15102 2040
rect 15068 1971 15102 2001
rect 15068 1967 15102 1971
rect 15068 1902 15102 1929
rect 15068 1895 15102 1902
rect 15068 1833 15102 1857
rect 15068 1823 15102 1833
rect 15068 1764 15102 1785
rect 15068 1751 15102 1764
rect 15068 1695 15102 1713
rect 15068 1679 15102 1695
rect 15068 1626 15102 1641
rect 15068 1607 15102 1626
rect 15068 1557 15102 1569
rect 15068 1535 15102 1557
rect 15068 1488 15102 1497
rect 15068 1463 15102 1488
rect 15068 1419 15102 1425
rect 15068 1391 15102 1419
rect 15068 1350 15102 1353
rect 15068 1319 15102 1350
rect 15068 1247 15102 1281
rect 7069 1189 7103 1217
rect 7142 1189 7176 1217
rect 7215 1189 7249 1217
rect 7288 1189 7322 1217
rect 7361 1189 7395 1217
rect 7434 1189 7468 1217
rect 7507 1189 7541 1217
rect 7580 1189 7614 1217
rect 7653 1189 7687 1217
rect 7726 1189 7760 1217
rect 7799 1189 7833 1217
rect 7872 1189 7906 1217
rect 7945 1189 7979 1217
rect 8018 1189 8052 1217
rect 8091 1189 8125 1217
rect 8164 1189 8198 1217
rect 8237 1189 8271 1217
rect 8310 1189 8344 1217
rect 8383 1189 8417 1217
rect 8456 1189 8490 1217
rect 8528 1189 8562 1217
rect 8600 1189 8634 1217
rect 8672 1189 8706 1217
rect 8744 1189 8778 1217
rect 8816 1189 8850 1217
rect 8888 1189 8922 1217
rect 8960 1189 8994 1217
rect 9032 1189 9066 1217
rect 7069 1183 7102 1189
rect 7102 1183 7103 1189
rect 7142 1183 7171 1189
rect 7171 1183 7176 1189
rect 7215 1183 7240 1189
rect 7240 1183 7249 1189
rect 7288 1183 7309 1189
rect 7309 1183 7322 1189
rect 7361 1183 7378 1189
rect 7378 1183 7395 1189
rect 7434 1183 7447 1189
rect 7447 1183 7468 1189
rect 7507 1183 7516 1189
rect 7516 1183 7541 1189
rect 7580 1183 7585 1189
rect 7585 1183 7614 1189
rect 7653 1183 7654 1189
rect 7654 1183 7687 1189
rect 7726 1183 7758 1189
rect 7758 1183 7760 1189
rect 7799 1183 7827 1189
rect 7827 1183 7833 1189
rect 7872 1183 7896 1189
rect 7896 1183 7906 1189
rect 7945 1183 7965 1189
rect 7965 1183 7979 1189
rect 8018 1183 8034 1189
rect 8034 1183 8052 1189
rect 8091 1183 8103 1189
rect 8103 1183 8125 1189
rect 8164 1183 8172 1189
rect 8172 1183 8198 1189
rect 8237 1183 8241 1189
rect 8241 1183 8271 1189
rect 8310 1183 8344 1189
rect 8383 1183 8413 1189
rect 8413 1183 8417 1189
rect 8456 1183 8482 1189
rect 8482 1183 8490 1189
rect 8528 1183 8551 1189
rect 8551 1183 8562 1189
rect 8600 1183 8620 1189
rect 8620 1183 8634 1189
rect 8672 1183 8689 1189
rect 8689 1183 8706 1189
rect 8744 1183 8758 1189
rect 8758 1183 8778 1189
rect 8816 1183 8827 1189
rect 8827 1183 8850 1189
rect 8888 1183 8896 1189
rect 8896 1183 8922 1189
rect 8960 1183 8965 1189
rect 8965 1183 8994 1189
rect 9032 1183 9034 1189
rect 9034 1183 9066 1189
rect 9104 1183 9138 1217
rect 9176 1189 9210 1217
rect 9248 1189 9282 1217
rect 9320 1189 9354 1217
rect 9392 1189 9426 1217
rect 9464 1189 9498 1217
rect 9536 1189 9570 1217
rect 9608 1189 9642 1217
rect 9680 1189 9714 1217
rect 9176 1183 9207 1189
rect 9207 1183 9210 1189
rect 9248 1183 9276 1189
rect 9276 1183 9282 1189
rect 9320 1183 9345 1189
rect 9345 1183 9354 1189
rect 9392 1183 9414 1189
rect 9414 1183 9426 1189
rect 9464 1183 9483 1189
rect 9483 1183 9498 1189
rect 9536 1183 9552 1189
rect 9552 1183 9570 1189
rect 9608 1183 9621 1189
rect 9621 1183 9642 1189
rect 9680 1183 9690 1189
rect 9690 1183 9714 1189
rect 9752 1183 9759 1217
rect 9759 1183 9786 1217
rect 9824 1183 9858 1217
rect 9896 1183 9930 1217
rect 9968 1183 10002 1217
rect 10040 1183 10074 1217
rect 10112 1183 10146 1217
rect 10184 1183 10218 1217
rect 10256 1183 10290 1217
rect 10328 1183 10362 1217
rect 10400 1183 10434 1217
rect 10472 1183 10506 1217
rect 10544 1183 10578 1217
rect 10616 1183 10650 1217
rect 10688 1183 10722 1217
rect 10760 1183 10794 1217
rect 10832 1183 10866 1217
rect 10904 1183 10938 1217
rect 10976 1183 11010 1217
rect 11048 1183 11082 1217
rect 11120 1183 11154 1217
rect 11192 1183 11226 1217
rect 11264 1183 11298 1217
rect 11336 1183 11370 1217
rect 11408 1183 11442 1217
rect 11480 1183 11514 1217
rect 11552 1183 11586 1217
rect 11624 1183 11658 1217
rect 11696 1183 11730 1217
rect 11768 1183 11802 1217
rect 11840 1183 11874 1217
rect 11912 1183 11946 1217
rect 11984 1183 12018 1217
rect 12056 1183 12090 1217
rect 12139 1183 12173 1217
rect 12212 1183 12246 1217
rect 12285 1183 12319 1217
rect 12358 1183 12392 1217
rect 12431 1183 12465 1217
rect 12504 1183 12538 1217
rect 12577 1183 12611 1217
rect 12650 1183 12684 1217
rect 12723 1183 12757 1217
rect 12796 1183 12830 1217
rect 12869 1183 12903 1217
rect 12942 1183 12976 1217
rect 13015 1183 13049 1217
rect 13088 1183 13122 1217
rect 13161 1183 13195 1217
rect 13234 1183 13268 1217
rect 13307 1183 13341 1217
rect 13380 1183 13414 1217
rect 13452 1183 13486 1217
rect 13524 1183 13558 1217
rect 13596 1183 13630 1217
rect 13668 1183 13702 1217
rect 13740 1183 13774 1217
rect 13812 1183 13846 1217
rect 13884 1183 13918 1217
rect 13956 1183 13990 1217
rect 14028 1183 14062 1217
rect 14100 1183 14134 1217
rect 14172 1183 14206 1217
rect 14244 1183 14278 1217
rect 14316 1183 14350 1217
rect 14388 1183 14422 1217
rect 14460 1183 14494 1217
rect 14532 1183 14566 1217
rect 14604 1183 14638 1217
rect 14676 1183 14710 1217
rect 14748 1183 14782 1217
rect 14820 1183 14854 1217
rect 14892 1183 14893 1217
rect 14893 1183 14926 1217
rect 14964 1210 14966 1217
rect 14966 1210 14998 1217
rect 14964 1183 14998 1210
rect 15068 1175 15102 1209
rect 7069 1121 7103 1139
rect 7142 1121 7176 1139
rect 7215 1121 7249 1139
rect 7288 1121 7322 1139
rect 7361 1121 7395 1139
rect 7434 1121 7468 1139
rect 7507 1121 7541 1139
rect 7580 1121 7614 1139
rect 7653 1121 7687 1139
rect 7726 1121 7760 1139
rect 7799 1121 7833 1139
rect 7872 1121 7906 1139
rect 7945 1121 7979 1139
rect 8018 1121 8052 1139
rect 8091 1121 8125 1139
rect 8164 1121 8198 1139
rect 8237 1121 8271 1139
rect 8310 1121 8344 1139
rect 8383 1121 8417 1139
rect 8456 1121 8490 1139
rect 8528 1121 8562 1139
rect 8600 1121 8634 1139
rect 8672 1121 8706 1139
rect 8744 1121 8778 1139
rect 8816 1121 8850 1139
rect 8888 1121 8922 1139
rect 8960 1121 8994 1139
rect 9032 1121 9066 1139
rect 7069 1105 7102 1121
rect 7102 1105 7103 1121
rect 7142 1105 7171 1121
rect 7171 1105 7176 1121
rect 7215 1105 7240 1121
rect 7240 1105 7249 1121
rect 7288 1105 7309 1121
rect 7309 1105 7322 1121
rect 7361 1105 7378 1121
rect 7378 1105 7395 1121
rect 7434 1105 7447 1121
rect 7447 1105 7468 1121
rect 7507 1105 7516 1121
rect 7516 1105 7541 1121
rect 7580 1105 7585 1121
rect 7585 1105 7614 1121
rect 7653 1105 7654 1121
rect 7654 1105 7687 1121
rect 7726 1105 7758 1121
rect 7758 1105 7760 1121
rect 7799 1105 7827 1121
rect 7827 1105 7833 1121
rect 7872 1105 7896 1121
rect 7896 1105 7906 1121
rect 7945 1105 7965 1121
rect 7965 1105 7979 1121
rect 8018 1105 8034 1121
rect 8034 1105 8052 1121
rect 8091 1105 8103 1121
rect 8103 1105 8125 1121
rect 8164 1105 8172 1121
rect 8172 1105 8198 1121
rect 8237 1105 8241 1121
rect 8241 1105 8271 1121
rect 8310 1105 8344 1121
rect 8383 1105 8413 1121
rect 8413 1105 8417 1121
rect 8456 1105 8482 1121
rect 8482 1105 8490 1121
rect 8528 1105 8551 1121
rect 8551 1105 8562 1121
rect 8600 1105 8620 1121
rect 8620 1105 8634 1121
rect 8672 1105 8689 1121
rect 8689 1105 8706 1121
rect 8744 1105 8758 1121
rect 8758 1105 8778 1121
rect 8816 1105 8827 1121
rect 8827 1105 8850 1121
rect 8888 1105 8896 1121
rect 8896 1105 8922 1121
rect 8960 1105 8965 1121
rect 8965 1105 8994 1121
rect 9032 1105 9034 1121
rect 9034 1105 9066 1121
rect 9104 1105 9138 1139
rect 9176 1121 9210 1139
rect 9248 1121 9282 1139
rect 9320 1121 9354 1139
rect 9392 1121 9426 1139
rect 9464 1121 9498 1139
rect 9536 1121 9570 1139
rect 9608 1121 9642 1139
rect 9680 1121 9714 1139
rect 9176 1105 9207 1121
rect 9207 1105 9210 1121
rect 9248 1105 9276 1121
rect 9276 1105 9282 1121
rect 9320 1105 9345 1121
rect 9345 1105 9354 1121
rect 9392 1105 9414 1121
rect 9414 1105 9426 1121
rect 9464 1105 9483 1121
rect 9483 1105 9498 1121
rect 9536 1105 9552 1121
rect 9552 1105 9570 1121
rect 9608 1105 9621 1121
rect 9621 1105 9642 1121
rect 9680 1105 9690 1121
rect 9690 1105 9714 1121
rect 9752 1105 9759 1139
rect 9759 1105 9786 1139
rect 9824 1105 9858 1139
rect 9896 1105 9930 1139
rect 9968 1105 10002 1139
rect 10040 1105 10074 1139
rect 10112 1105 10146 1139
rect 10184 1105 10218 1139
rect 10256 1105 10290 1139
rect 10328 1105 10362 1139
rect 10400 1105 10434 1139
rect 10472 1105 10506 1139
rect 10544 1105 10578 1139
rect 10616 1105 10650 1139
rect 10688 1105 10722 1139
rect 10760 1105 10794 1139
rect 10832 1105 10866 1139
rect 10904 1105 10938 1139
rect 10976 1105 11010 1139
rect 11048 1105 11082 1139
rect 11120 1105 11154 1139
rect 11192 1105 11226 1139
rect 11264 1105 11298 1139
rect 11336 1105 11370 1139
rect 11408 1105 11442 1139
rect 11480 1105 11514 1139
rect 11552 1105 11586 1139
rect 11624 1105 11658 1139
rect 11696 1105 11730 1139
rect 11768 1105 11802 1139
rect 11840 1105 11874 1139
rect 11912 1105 11946 1139
rect 11984 1105 12018 1139
rect 12056 1105 12090 1139
rect 12139 1105 12173 1139
rect 12212 1105 12246 1139
rect 12285 1105 12319 1139
rect 12358 1105 12392 1139
rect 12431 1105 12465 1139
rect 12504 1105 12538 1139
rect 12577 1105 12611 1139
rect 12650 1105 12684 1139
rect 12723 1105 12757 1139
rect 12796 1105 12830 1139
rect 12869 1105 12903 1139
rect 12942 1105 12976 1139
rect 13015 1105 13049 1139
rect 13088 1105 13122 1139
rect 13161 1105 13195 1139
rect 13234 1105 13268 1139
rect 13307 1105 13341 1139
rect 13380 1105 13414 1139
rect 13452 1105 13486 1139
rect 13524 1105 13558 1139
rect 13596 1105 13630 1139
rect 13668 1105 13702 1139
rect 13740 1105 13774 1139
rect 13812 1105 13846 1139
rect 13884 1105 13918 1139
rect 13956 1105 13990 1139
rect 14028 1105 14062 1139
rect 14100 1105 14134 1139
rect 14172 1105 14206 1139
rect 14244 1105 14278 1139
rect 14316 1105 14350 1139
rect 14388 1105 14422 1139
rect 14460 1105 14494 1139
rect 14532 1105 14566 1139
rect 14604 1105 14638 1139
rect 14676 1105 14710 1139
rect 14748 1105 14782 1139
rect 14820 1105 14854 1139
rect 14892 1105 14893 1139
rect 14893 1105 14926 1139
rect 14964 1138 14966 1139
rect 14966 1138 14998 1139
rect 14964 1105 14998 1138
rect 15068 1103 15102 1137
rect 7069 1053 7103 1061
rect 7142 1053 7176 1061
rect 7215 1053 7249 1061
rect 7288 1053 7322 1061
rect 7361 1053 7395 1061
rect 7434 1053 7468 1061
rect 7507 1053 7541 1061
rect 7580 1053 7614 1061
rect 7653 1053 7687 1061
rect 7726 1053 7760 1061
rect 7799 1053 7833 1061
rect 7872 1053 7906 1061
rect 7945 1053 7979 1061
rect 8018 1053 8052 1061
rect 8091 1053 8125 1061
rect 8164 1053 8198 1061
rect 8237 1053 8271 1061
rect 8310 1053 8344 1061
rect 8383 1053 8417 1061
rect 8456 1053 8490 1061
rect 8528 1053 8562 1061
rect 8600 1053 8634 1061
rect 8672 1053 8706 1061
rect 8744 1053 8778 1061
rect 8816 1053 8850 1061
rect 8888 1053 8922 1061
rect 8960 1053 8994 1061
rect 9032 1053 9066 1061
rect 7069 1027 7102 1053
rect 7102 1027 7103 1053
rect 7142 1027 7171 1053
rect 7171 1027 7176 1053
rect 7215 1027 7240 1053
rect 7240 1027 7249 1053
rect 7288 1027 7309 1053
rect 7309 1027 7322 1053
rect 7361 1027 7378 1053
rect 7378 1027 7395 1053
rect 7434 1027 7447 1053
rect 7447 1027 7468 1053
rect 7507 1027 7516 1053
rect 7516 1027 7541 1053
rect 7580 1027 7585 1053
rect 7585 1027 7614 1053
rect 7653 1027 7654 1053
rect 7654 1027 7687 1053
rect 7726 1027 7758 1053
rect 7758 1027 7760 1053
rect 7799 1027 7827 1053
rect 7827 1027 7833 1053
rect 7872 1027 7896 1053
rect 7896 1027 7906 1053
rect 7945 1027 7965 1053
rect 7965 1027 7979 1053
rect 8018 1027 8034 1053
rect 8034 1027 8052 1053
rect 8091 1027 8103 1053
rect 8103 1027 8125 1053
rect 8164 1027 8172 1053
rect 8172 1027 8198 1053
rect 8237 1027 8241 1053
rect 8241 1027 8271 1053
rect 8310 1027 8344 1053
rect 8383 1027 8413 1053
rect 8413 1027 8417 1053
rect 8456 1027 8482 1053
rect 8482 1027 8490 1053
rect 8528 1027 8551 1053
rect 8551 1027 8562 1053
rect 8600 1027 8620 1053
rect 8620 1027 8634 1053
rect 8672 1027 8689 1053
rect 8689 1027 8706 1053
rect 8744 1027 8758 1053
rect 8758 1027 8778 1053
rect 8816 1027 8827 1053
rect 8827 1027 8850 1053
rect 8888 1027 8896 1053
rect 8896 1027 8922 1053
rect 8960 1027 8965 1053
rect 8965 1027 8994 1053
rect 9032 1027 9034 1053
rect 9034 1027 9066 1053
rect 9104 1027 9138 1061
rect 9176 1053 9210 1061
rect 9248 1053 9282 1061
rect 9320 1053 9354 1061
rect 9392 1053 9426 1061
rect 9464 1053 9498 1061
rect 9536 1053 9570 1061
rect 9608 1053 9642 1061
rect 9680 1053 9714 1061
rect 9176 1027 9207 1053
rect 9207 1027 9210 1053
rect 9248 1027 9276 1053
rect 9276 1027 9282 1053
rect 9320 1027 9345 1053
rect 9345 1027 9354 1053
rect 9392 1027 9414 1053
rect 9414 1027 9426 1053
rect 9464 1027 9483 1053
rect 9483 1027 9498 1053
rect 9536 1027 9552 1053
rect 9552 1027 9570 1053
rect 9608 1027 9621 1053
rect 9621 1027 9642 1053
rect 9680 1027 9690 1053
rect 9690 1027 9714 1053
rect 9752 1027 9759 1061
rect 9759 1027 9786 1061
rect 9824 1027 9858 1061
rect 9896 1027 9930 1061
rect 9968 1027 10002 1061
rect 10040 1027 10074 1061
rect 10112 1027 10146 1061
rect 10184 1027 10218 1061
rect 10256 1027 10290 1061
rect 10328 1027 10362 1061
rect 10400 1027 10434 1061
rect 10472 1027 10506 1061
rect 10544 1027 10578 1061
rect 10616 1027 10650 1061
rect 10688 1027 10722 1061
rect 10760 1027 10794 1061
rect 10832 1027 10866 1061
rect 10904 1027 10938 1061
rect 10976 1027 11010 1061
rect 11048 1027 11082 1061
rect 11120 1027 11154 1061
rect 11192 1027 11226 1061
rect 11264 1027 11298 1061
rect 11336 1027 11370 1061
rect 11408 1027 11442 1061
rect 11480 1027 11514 1061
rect 11552 1027 11586 1061
rect 11624 1027 11658 1061
rect 11696 1027 11730 1061
rect 11768 1027 11802 1061
rect 11840 1027 11874 1061
rect 11912 1027 11946 1061
rect 11984 1027 12018 1061
rect 12056 1027 12090 1061
rect 12139 1027 12173 1061
rect 12212 1027 12246 1061
rect 12285 1027 12319 1061
rect 12358 1027 12392 1061
rect 12431 1027 12465 1061
rect 12504 1027 12538 1061
rect 12577 1027 12611 1061
rect 12650 1027 12684 1061
rect 12723 1027 12757 1061
rect 12796 1027 12830 1061
rect 12869 1027 12903 1061
rect 12942 1027 12976 1061
rect 13015 1027 13049 1061
rect 13088 1027 13122 1061
rect 13161 1027 13195 1061
rect 13234 1027 13268 1061
rect 13307 1027 13341 1061
rect 13380 1027 13414 1061
rect 13452 1027 13486 1061
rect 13524 1027 13558 1061
rect 13596 1027 13630 1061
rect 13668 1027 13702 1061
rect 13740 1027 13774 1061
rect 13812 1027 13846 1061
rect 13884 1027 13918 1061
rect 13956 1027 13990 1061
rect 14028 1027 14062 1061
rect 14100 1027 14134 1061
rect 14172 1027 14206 1061
rect 14244 1027 14278 1061
rect 14316 1027 14350 1061
rect 14388 1027 14422 1061
rect 14460 1027 14494 1061
rect 14532 1027 14566 1061
rect 14604 1027 14638 1061
rect 14676 1027 14710 1061
rect 14748 1027 14782 1061
rect 14820 1027 14854 1061
rect 14892 1027 14893 1061
rect 14893 1027 14926 1061
rect 14964 1028 14998 1061
rect 15068 1031 15102 1065
rect 14964 1027 14966 1028
rect 14966 1027 14998 1028
rect 7104 913 7137 918
rect 7137 913 7138 918
rect 7104 884 7138 913
rect 14576 955 14610 989
rect 14654 955 14688 989
rect 14732 955 14766 989
rect 14810 955 14844 989
rect 14888 955 14922 989
rect 9796 913 9815 923
rect 9815 913 9830 923
rect 9872 913 9885 923
rect 9885 913 9906 923
rect 9948 913 9955 923
rect 9955 913 9982 923
rect 10024 913 10025 923
rect 10025 913 10058 923
rect 10100 913 10131 923
rect 10131 913 10134 923
rect 10176 913 10201 923
rect 10201 913 10210 923
rect 10251 913 10271 923
rect 10271 913 10285 923
rect 10326 913 10341 923
rect 10341 913 10360 923
rect 10401 913 10411 923
rect 10411 913 10435 923
rect 10476 913 10481 923
rect 10481 913 10510 923
rect 10551 913 10585 923
rect 10626 913 10655 923
rect 10655 913 10660 923
rect 10701 913 10725 923
rect 10725 913 10735 923
rect 10776 913 10795 923
rect 10795 913 10810 923
rect 10851 913 10865 923
rect 10865 913 10885 923
rect 10926 913 10935 923
rect 10935 913 10960 923
rect 11001 913 11005 923
rect 11005 913 11035 923
rect 9796 889 9830 913
rect 9872 889 9906 913
rect 9948 889 9982 913
rect 10024 889 10058 913
rect 10100 889 10134 913
rect 10176 889 10210 913
rect 10251 889 10285 913
rect 10326 889 10360 913
rect 10401 889 10435 913
rect 10476 889 10510 913
rect 10551 889 10585 913
rect 10626 889 10660 913
rect 10701 889 10735 913
rect 10776 889 10810 913
rect 10851 889 10885 913
rect 10926 889 10960 913
rect 11001 889 11035 913
rect 11076 889 11110 923
rect 11151 913 11181 923
rect 11181 913 11185 923
rect 11226 913 11251 923
rect 11251 913 11260 923
rect 11301 913 11321 923
rect 11321 913 11335 923
rect 14966 955 15000 989
rect 15068 959 15102 993
rect 11151 889 11185 913
rect 11226 889 11260 913
rect 11301 889 11335 913
rect 14576 882 14610 916
rect 14654 882 14688 916
rect 14732 882 14766 916
rect 14810 882 14844 916
rect 14888 882 14922 916
rect 14576 841 14583 843
rect 14583 841 14610 843
rect 14966 882 15000 916
rect 15068 887 15102 921
rect 14654 841 14686 843
rect 14686 841 14688 843
rect 14732 841 14755 843
rect 14755 841 14766 843
rect 14810 841 14824 843
rect 14824 841 14844 843
rect 14888 841 14893 843
rect 14893 841 14922 843
rect 9796 805 9830 839
rect 9872 805 9906 839
rect 9948 805 9982 839
rect 10024 805 10058 839
rect 10100 805 10134 839
rect 10176 805 10210 839
rect 10251 805 10285 839
rect 10326 805 10360 839
rect 10401 805 10435 839
rect 10476 805 10510 839
rect 10551 805 10585 839
rect 10626 805 10660 839
rect 10701 805 10735 839
rect 10776 805 10810 839
rect 10851 805 10885 839
rect 10926 805 10960 839
rect 11001 805 11035 839
rect 11076 805 11110 839
rect 11151 805 11185 839
rect 11226 805 11260 839
rect 11301 805 11335 839
rect 14576 809 14610 841
rect 14654 809 14688 841
rect 14732 809 14766 841
rect 14810 809 14844 841
rect 14888 809 14922 841
rect 14576 761 14583 770
rect 14583 761 14610 770
rect 14966 809 15000 843
rect 15068 815 15102 849
rect 14654 761 14686 770
rect 14686 761 14688 770
rect 14732 761 14755 770
rect 14755 761 14766 770
rect 14810 761 14824 770
rect 14824 761 14844 770
rect 14888 761 14893 770
rect 14893 761 14922 770
rect 9796 731 9830 755
rect 9872 731 9906 755
rect 9948 731 9982 755
rect 10024 731 10058 755
rect 10100 731 10134 755
rect 10176 731 10210 755
rect 10251 731 10285 755
rect 10326 731 10360 755
rect 10401 731 10435 755
rect 10476 731 10510 755
rect 10551 731 10585 755
rect 10626 731 10660 755
rect 10701 731 10735 755
rect 10776 731 10810 755
rect 10851 731 10885 755
rect 10926 731 10960 755
rect 11001 731 11035 755
rect 9796 721 9815 731
rect 9815 721 9830 731
rect 9872 721 9885 731
rect 9885 721 9906 731
rect 9948 721 9955 731
rect 9955 721 9982 731
rect 10024 721 10025 731
rect 10025 721 10058 731
rect 10100 721 10131 731
rect 10131 721 10134 731
rect 10176 721 10201 731
rect 10201 721 10210 731
rect 10251 721 10271 731
rect 10271 721 10285 731
rect 10326 721 10341 731
rect 10341 721 10360 731
rect 10401 721 10411 731
rect 10411 721 10435 731
rect 10476 721 10481 731
rect 10481 721 10510 731
rect 10551 721 10585 731
rect 10626 721 10655 731
rect 10655 721 10660 731
rect 10701 721 10725 731
rect 10725 721 10735 731
rect 10776 721 10795 731
rect 10795 721 10810 731
rect 10851 721 10865 731
rect 10865 721 10885 731
rect 10926 721 10935 731
rect 10935 721 10960 731
rect 11001 721 11005 731
rect 11005 721 11035 731
rect 11076 721 11110 755
rect 11151 731 11185 755
rect 11226 731 11260 755
rect 11301 731 11335 755
rect 14576 736 14610 761
rect 14654 736 14688 761
rect 14732 736 14766 761
rect 14810 736 14844 761
rect 14888 736 14922 761
rect 11151 721 11181 731
rect 11181 721 11185 731
rect 11226 721 11251 731
rect 11251 721 11260 731
rect 11301 721 11321 731
rect 11321 721 11335 731
rect 9796 659 9830 671
rect 9872 659 9906 671
rect 9948 659 9982 671
rect 10024 659 10058 671
rect 10100 659 10134 671
rect 10176 659 10210 671
rect 10251 659 10285 671
rect 10326 659 10360 671
rect 10401 659 10435 671
rect 10476 659 10510 671
rect 10551 659 10585 671
rect 10626 659 10660 671
rect 10701 659 10735 671
rect 10776 659 10810 671
rect 10851 659 10885 671
rect 10926 659 10960 671
rect 11001 659 11035 671
rect 9796 637 9815 659
rect 9815 637 9830 659
rect 9872 637 9885 659
rect 9885 637 9906 659
rect 9948 637 9955 659
rect 9955 637 9982 659
rect 10024 637 10025 659
rect 10025 637 10058 659
rect 10100 637 10131 659
rect 10131 637 10134 659
rect 10176 637 10201 659
rect 10201 637 10210 659
rect 10251 637 10271 659
rect 10271 637 10285 659
rect 10326 637 10341 659
rect 10341 637 10360 659
rect 10401 637 10411 659
rect 10411 637 10435 659
rect 10476 637 10481 659
rect 10481 637 10510 659
rect 10551 637 10585 659
rect 10626 637 10655 659
rect 10655 637 10660 659
rect 10701 637 10725 659
rect 10725 637 10735 659
rect 10776 637 10795 659
rect 10795 637 10810 659
rect 10851 637 10865 659
rect 10865 637 10885 659
rect 10926 637 10935 659
rect 10935 637 10960 659
rect 11001 637 11005 659
rect 11005 637 11035 659
rect 11076 637 11110 671
rect 11151 659 11185 671
rect 11226 659 11260 671
rect 11301 659 11335 671
rect 11151 637 11181 659
rect 11181 637 11185 659
rect 11226 637 11251 659
rect 11251 637 11260 659
rect 11301 637 11321 659
rect 11321 637 11335 659
rect 9796 553 9815 587
rect 9815 553 9830 587
rect 9872 553 9885 587
rect 9885 553 9906 587
rect 9948 553 9955 587
rect 9955 553 9982 587
rect 10024 553 10025 587
rect 10025 553 10058 587
rect 10100 553 10131 587
rect 10131 553 10134 587
rect 10176 553 10201 587
rect 10201 553 10210 587
rect 10251 553 10271 587
rect 10271 553 10285 587
rect 10326 553 10341 587
rect 10341 553 10360 587
rect 10401 553 10411 587
rect 10411 553 10435 587
rect 10476 553 10481 587
rect 10481 553 10510 587
rect 10551 553 10585 587
rect 10626 553 10655 587
rect 10655 553 10660 587
rect 10701 553 10725 587
rect 10725 553 10735 587
rect 10776 553 10795 587
rect 10795 553 10810 587
rect 10851 553 10865 587
rect 10865 553 10885 587
rect 10926 553 10935 587
rect 10935 553 10960 587
rect 11001 553 11005 587
rect 11005 553 11035 587
rect 11076 553 11110 587
rect 11151 553 11181 587
rect 11181 553 11185 587
rect 11226 553 11251 587
rect 11251 553 11260 587
rect 11301 553 11321 587
rect 11321 553 11335 587
rect 9796 481 9815 503
rect 9815 481 9830 503
rect 9872 481 9885 503
rect 9885 481 9906 503
rect 9948 481 9955 503
rect 9955 481 9982 503
rect 10024 481 10025 503
rect 10025 481 10058 503
rect 10100 481 10131 503
rect 10131 481 10134 503
rect 10176 481 10201 503
rect 10201 481 10210 503
rect 10251 481 10271 503
rect 10271 481 10285 503
rect 10326 481 10341 503
rect 10341 481 10360 503
rect 10401 481 10411 503
rect 10411 481 10435 503
rect 10476 481 10481 503
rect 10481 481 10510 503
rect 10551 481 10585 503
rect 10626 481 10655 503
rect 10655 481 10660 503
rect 10701 481 10725 503
rect 10725 481 10735 503
rect 10776 481 10795 503
rect 10795 481 10810 503
rect 10851 481 10865 503
rect 10865 481 10885 503
rect 10926 481 10935 503
rect 10935 481 10960 503
rect 11001 481 11005 503
rect 11005 481 11035 503
rect 9796 469 9830 481
rect 9872 469 9906 481
rect 9948 469 9982 481
rect 10024 469 10058 481
rect 10100 469 10134 481
rect 10176 469 10210 481
rect 10251 469 10285 481
rect 10326 469 10360 481
rect 10401 469 10435 481
rect 10476 469 10510 481
rect 10551 469 10585 481
rect 10626 469 10660 481
rect 10701 469 10735 481
rect 10776 469 10810 481
rect 10851 469 10885 481
rect 10926 469 10960 481
rect 11001 469 11035 481
rect 11076 469 11110 503
rect 11151 481 11181 503
rect 11181 481 11185 503
rect 11226 481 11251 503
rect 11251 481 11260 503
rect 11301 481 11321 503
rect 11321 481 11335 503
rect 11151 469 11185 481
rect 11226 469 11260 481
rect 11301 469 11335 481
rect 14966 736 15000 770
rect 15068 743 15102 777
rect 14576 695 14610 697
rect 14654 695 14688 697
rect 14576 663 14577 695
rect 14577 663 14610 695
rect 14654 663 14655 695
rect 14655 663 14688 695
rect 14732 663 14766 697
rect 14810 663 14844 697
rect 14888 663 14922 697
rect 14966 663 15000 697
rect 15068 671 15102 705
rect 14576 609 14610 623
rect 14654 609 14688 623
rect 14576 589 14577 609
rect 14577 589 14610 609
rect 14654 589 14655 609
rect 14655 589 14688 609
rect 14732 589 14766 623
rect 14810 589 14844 623
rect 14888 589 14922 623
rect 14966 589 15000 623
rect 15068 599 15102 633
rect 14576 523 14610 549
rect 14654 523 14688 549
rect 14576 515 14577 523
rect 14577 515 14610 523
rect 14654 515 14655 523
rect 14655 515 14688 523
rect 14732 515 14766 549
rect 14810 515 14844 549
rect 14888 515 14922 549
rect 14966 515 15000 549
rect 15068 527 15102 561
rect 14576 441 14610 475
rect 14654 441 14688 475
rect 14732 441 14766 475
rect 14810 441 14844 475
rect 14888 441 14922 475
rect 14966 441 15000 475
rect 15068 455 15102 489
rect 14657 367 14691 390
rect 14735 367 14769 390
rect 14813 367 14847 390
rect 14891 367 14925 390
rect 14969 380 15003 390
rect 15068 383 15102 417
rect 14657 356 14689 367
rect 14689 356 14691 367
rect 14735 356 14757 367
rect 14757 356 14769 367
rect 14813 356 14825 367
rect 14825 356 14847 367
rect 14891 356 14893 367
rect 14893 356 14925 367
rect 14969 356 15000 380
rect 15000 356 15003 380
rect 14657 289 14691 312
rect 14735 289 14769 312
rect 14813 289 14847 312
rect 14891 289 14925 312
rect 14969 308 15003 312
rect 15068 311 15102 345
rect 14657 278 14689 289
rect 14689 278 14691 289
rect 14735 278 14757 289
rect 14757 278 14769 289
rect 14813 278 14825 289
rect 14825 278 14847 289
rect 14891 278 14893 289
rect 14893 278 14925 289
rect 14969 278 15000 308
rect 15000 278 15003 308
rect 15068 238 15102 272
rect 14657 211 14691 234
rect 14735 211 14769 234
rect 14813 211 14847 234
rect 14891 211 14925 234
rect 14657 200 14689 211
rect 14689 200 14691 211
rect 14735 200 14757 211
rect 14757 200 14769 211
rect 14813 200 14825 211
rect 14825 200 14847 211
rect 14891 200 14893 211
rect 14893 200 14925 211
rect 14969 202 15000 234
rect 15000 202 15003 234
rect 14969 200 15003 202
rect 15068 165 15102 199
rect 14657 133 14691 156
rect 14735 133 14769 156
rect 14813 133 14847 156
rect 14891 133 14925 156
rect 14657 122 14689 133
rect 14689 122 14691 133
rect 14735 122 14757 133
rect 14757 122 14769 133
rect 14813 122 14825 133
rect 14825 122 14847 133
rect 14891 122 14893 133
rect 14893 122 14925 133
rect 14969 130 15000 156
rect 15000 130 15003 156
rect 14969 122 15003 130
rect 15068 92 15102 126
rect 14657 55 14691 77
rect 14735 55 14769 77
rect 14813 55 14847 77
rect 14891 55 14925 77
rect 14969 57 15000 77
rect 15000 57 15003 77
rect 14657 43 14689 55
rect 14689 43 14691 55
rect 14735 43 14757 55
rect 14757 43 14769 55
rect 14813 43 14825 55
rect 14825 43 14847 55
rect 14891 43 14893 55
rect 14893 43 14925 55
rect 14969 43 15003 57
rect 15068 19 15102 53
rect 5884 -9191 5918 -9157
rect 5884 -9263 5918 -9229
<< metal1 >>
rect 359 16145 411 16151
rect 359 16081 411 16093
rect 359 16023 411 16029
rect 278 15989 330 15995
rect 278 15925 330 15937
rect 278 15867 330 15873
rect 535 10030 970 10031
rect 535 9978 541 10030
rect 593 9978 616 10030
rect 668 9978 690 10030
rect 742 9978 764 10030
rect 816 9978 838 10030
rect 890 9978 912 10030
rect 964 9978 970 10030
rect 535 9956 970 9978
rect 535 9904 541 9956
rect 593 9904 616 9956
rect 668 9904 690 9956
rect 742 9904 764 9956
rect 816 9904 838 9956
rect 890 9904 912 9956
rect 964 9904 970 9956
rect 535 9882 970 9904
rect 535 9830 541 9882
rect 593 9830 616 9882
rect 668 9830 690 9882
rect 742 9830 764 9882
rect 816 9830 838 9882
rect 890 9830 912 9882
rect 964 9830 970 9882
rect 535 9829 970 9830
tri 13999 9622 14206 9829 ne
rect -496 9514 13845 9521
rect -496 9480 -484 9514
rect -450 9480 -411 9514
rect -377 9480 -338 9514
rect -304 9480 -265 9514
rect -231 9480 -192 9514
rect -158 9480 -119 9514
rect -85 9480 -46 9514
rect -12 9480 27 9514
rect 61 9480 100 9514
rect 134 9480 173 9514
rect 207 9480 246 9514
rect 280 9480 319 9514
rect 353 9480 392 9514
rect 426 9480 465 9514
rect 499 9480 538 9514
rect 572 9480 611 9514
rect 645 9480 684 9514
rect 718 9480 757 9514
rect 791 9480 830 9514
rect 864 9480 903 9514
rect 937 9480 976 9514
rect 1010 9480 1049 9514
rect 1083 9480 1122 9514
rect 1156 9480 1195 9514
rect 1229 9480 1268 9514
rect 1302 9480 1341 9514
rect 1375 9480 1414 9514
rect 1448 9480 1487 9514
rect 1521 9480 1559 9514
rect 1593 9480 1631 9514
rect 1665 9480 1703 9514
rect 1737 9480 1775 9514
rect 1809 9480 1847 9514
rect 1881 9480 1919 9514
rect 1953 9480 1991 9514
rect 2025 9480 2063 9514
rect 2097 9480 2135 9514
rect 2169 9480 2207 9514
rect 2241 9480 2279 9514
rect 2313 9480 2351 9514
rect 2385 9480 2423 9514
rect 2457 9480 2495 9514
rect 2529 9480 2567 9514
rect 2601 9480 2639 9514
rect 2673 9480 2711 9514
rect 2745 9480 2783 9514
rect 2817 9480 2855 9514
rect 2889 9480 2927 9514
rect 2961 9480 2999 9514
rect 3033 9480 3071 9514
rect 3105 9480 3143 9514
rect 3177 9480 3215 9514
rect 3249 9480 3287 9514
rect 3321 9480 3359 9514
rect 3393 9480 3431 9514
rect 3465 9480 3503 9514
rect 3537 9480 3575 9514
rect 3609 9480 3647 9514
rect 3681 9480 3719 9514
rect 3753 9480 3791 9514
rect 3825 9480 3863 9514
rect 3897 9480 3935 9514
rect 3969 9480 4007 9514
rect 4041 9480 4079 9514
rect 4113 9480 4151 9514
rect 4185 9480 4223 9514
rect 4257 9480 4295 9514
rect 4329 9480 4367 9514
rect 4401 9480 4439 9514
rect 4473 9480 4511 9514
rect 4545 9480 4583 9514
rect 4617 9480 4655 9514
rect 4689 9480 4727 9514
rect 4761 9480 4799 9514
rect 4833 9480 4871 9514
rect 4905 9480 4943 9514
rect 4977 9480 5015 9514
rect 5049 9480 5087 9514
rect 5121 9480 5159 9514
rect 5193 9480 5231 9514
rect 5265 9480 5303 9514
rect 5337 9480 5375 9514
rect 5409 9480 5447 9514
rect 5481 9480 5519 9514
rect 5553 9480 5591 9514
rect 5625 9480 5663 9514
rect 5697 9480 5735 9514
rect 5769 9480 5807 9514
rect 5841 9480 5879 9514
rect 5913 9480 5951 9514
rect 5985 9480 6023 9514
rect 6057 9480 6095 9514
rect 6129 9480 6167 9514
rect 6201 9480 6239 9514
rect 6273 9480 6311 9514
rect 6345 9480 6383 9514
rect 6417 9480 6455 9514
rect 6489 9480 6527 9514
rect 6561 9480 6599 9514
rect 6633 9480 6671 9514
rect 6705 9480 6743 9514
rect 6777 9480 6815 9514
rect 6849 9480 6887 9514
rect 6921 9480 6959 9514
rect 6993 9480 7031 9514
rect 7065 9480 7103 9514
rect 7137 9480 7175 9514
rect 7209 9480 7247 9514
rect 7281 9480 7319 9514
rect 7353 9480 7391 9514
rect 7425 9480 7463 9514
rect 7497 9480 7535 9514
rect 7569 9480 7607 9514
rect 7641 9480 7679 9514
rect 7713 9480 7751 9514
rect 7785 9480 7823 9514
rect 7857 9480 7895 9514
rect 7929 9480 7967 9514
rect 8001 9480 8039 9514
rect 8073 9480 8111 9514
rect 8145 9480 8183 9514
rect 8217 9480 8255 9514
rect 8289 9480 8327 9514
rect 8361 9480 8399 9514
rect 8433 9480 8471 9514
rect 8505 9480 8543 9514
rect 8577 9480 8615 9514
rect 8649 9480 8687 9514
rect 8721 9480 8759 9514
rect 8793 9480 8831 9514
rect 8865 9480 8903 9514
rect 8937 9480 8975 9514
rect 9009 9480 9047 9514
rect 9081 9480 9119 9514
rect 9153 9480 9191 9514
rect 9225 9480 9263 9514
rect 9297 9480 9335 9514
rect 9369 9480 9407 9514
rect 9441 9480 9479 9514
rect 9513 9480 9551 9514
rect 9585 9480 9623 9514
rect 9657 9480 9695 9514
rect 9729 9480 9767 9514
rect 9801 9480 9839 9514
rect 9873 9480 9911 9514
rect 9945 9480 9983 9514
rect 10017 9480 10055 9514
rect 10089 9480 10127 9514
rect 10161 9480 10199 9514
rect 10233 9480 10271 9514
rect 10305 9480 10343 9514
rect 10377 9480 10415 9514
rect 10449 9480 10487 9514
rect 10521 9480 10559 9514
rect 10593 9480 10631 9514
rect 10665 9480 10703 9514
rect 10737 9480 10775 9514
rect 10809 9480 10847 9514
rect 10881 9480 10919 9514
rect 10953 9480 10991 9514
rect 11025 9480 11063 9514
rect 11097 9480 11135 9514
rect 11169 9480 11207 9514
rect 11241 9480 11279 9514
rect 11313 9480 11351 9514
rect 11385 9480 11423 9514
rect 11457 9480 11495 9514
rect 11529 9480 11567 9514
rect 11601 9480 11639 9514
rect 11673 9480 11711 9514
rect 11745 9480 11783 9514
rect 11817 9480 11855 9514
rect 11889 9480 11927 9514
rect 11961 9480 11999 9514
rect 12033 9480 12071 9514
rect 12105 9480 12143 9514
rect 12177 9480 12215 9514
rect 12249 9480 12287 9514
rect 12321 9480 12359 9514
rect 12393 9480 12431 9514
rect 12465 9480 12503 9514
rect 12537 9480 12575 9514
rect 12609 9480 12647 9514
rect 12681 9480 12719 9514
rect 12753 9480 12791 9514
rect 12825 9480 12863 9514
rect 12897 9480 12935 9514
rect 12969 9480 13007 9514
rect 13041 9480 13079 9514
rect 13113 9480 13151 9514
rect 13185 9480 13223 9514
rect 13257 9480 13295 9514
rect 13329 9480 13367 9514
rect 13401 9480 13439 9514
rect 13473 9480 13511 9514
rect 13545 9480 13583 9514
rect 13617 9480 13655 9514
rect 13689 9480 13727 9514
rect 13761 9480 13799 9514
rect 13833 9480 13845 9514
rect -496 9428 13845 9480
rect -496 9394 -484 9428
rect -450 9394 -411 9428
rect -377 9394 -338 9428
rect -304 9394 -265 9428
rect -231 9394 -192 9428
rect -158 9394 -119 9428
rect -85 9394 -46 9428
rect -12 9394 27 9428
rect 61 9394 100 9428
rect 134 9394 173 9428
rect 207 9394 246 9428
rect 280 9394 319 9428
rect 353 9394 392 9428
rect 426 9394 465 9428
rect 499 9394 538 9428
rect 572 9394 611 9428
rect 645 9394 684 9428
rect 718 9394 757 9428
rect 791 9394 830 9428
rect 864 9394 903 9428
rect 937 9394 976 9428
rect 1010 9394 1049 9428
rect 1083 9394 1122 9428
rect 1156 9394 1195 9428
rect 1229 9394 1268 9428
rect 1302 9394 1341 9428
rect 1375 9394 1414 9428
rect 1448 9394 1487 9428
rect 1521 9394 1559 9428
rect 1593 9394 1631 9428
rect 1665 9394 1703 9428
rect 1737 9394 1775 9428
rect 1809 9394 1847 9428
rect 1881 9394 1919 9428
rect 1953 9394 1991 9428
rect 2025 9394 2063 9428
rect 2097 9394 2135 9428
rect 2169 9394 2207 9428
rect 2241 9394 2279 9428
rect 2313 9394 2351 9428
rect 2385 9394 2423 9428
rect 2457 9394 2495 9428
rect 2529 9394 2567 9428
rect 2601 9394 2639 9428
rect 2673 9394 2711 9428
rect 2745 9394 2783 9428
rect 2817 9394 2855 9428
rect 2889 9394 2927 9428
rect 2961 9394 2999 9428
rect 3033 9394 3071 9428
rect 3105 9394 3143 9428
rect 3177 9394 3215 9428
rect 3249 9394 3287 9428
rect 3321 9394 3359 9428
rect 3393 9394 3431 9428
rect 3465 9394 3503 9428
rect 3537 9394 3575 9428
rect 3609 9394 3647 9428
rect 3681 9394 3719 9428
rect 3753 9394 3791 9428
rect 3825 9394 3863 9428
rect 3897 9394 3935 9428
rect 3969 9394 4007 9428
rect 4041 9394 4079 9428
rect 4113 9394 4151 9428
rect 4185 9394 4223 9428
rect 4257 9394 4295 9428
rect 4329 9394 4367 9428
rect 4401 9394 4439 9428
rect 4473 9394 4511 9428
rect 4545 9394 4583 9428
rect 4617 9394 4655 9428
rect 4689 9394 4727 9428
rect 4761 9394 4799 9428
rect 4833 9394 4871 9428
rect 4905 9394 4943 9428
rect 4977 9394 5015 9428
rect 5049 9394 5087 9428
rect 5121 9394 5159 9428
rect 5193 9394 5231 9428
rect 5265 9394 5303 9428
rect 5337 9394 5375 9428
rect 5409 9394 5447 9428
rect 5481 9394 5519 9428
rect 5553 9394 5591 9428
rect 5625 9394 5663 9428
rect 5697 9394 5735 9428
rect 5769 9394 5807 9428
rect 5841 9394 5879 9428
rect 5913 9394 5951 9428
rect 5985 9394 6023 9428
rect 6057 9394 6095 9428
rect 6129 9394 6167 9428
rect 6201 9394 6239 9428
rect 6273 9394 6311 9428
rect 6345 9394 6383 9428
rect 6417 9394 6455 9428
rect 6489 9394 6527 9428
rect 6561 9394 6599 9428
rect 6633 9394 6671 9428
rect 6705 9394 6743 9428
rect 6777 9394 6815 9428
rect 6849 9394 6887 9428
rect 6921 9394 6959 9428
rect 6993 9394 7031 9428
rect 7065 9394 7103 9428
rect 7137 9394 7175 9428
rect 7209 9394 7247 9428
rect 7281 9394 7319 9428
rect 7353 9394 7391 9428
rect 7425 9394 7463 9428
rect 7497 9394 7535 9428
rect 7569 9394 7607 9428
rect 7641 9394 7679 9428
rect 7713 9394 7751 9428
rect 7785 9394 7823 9428
rect 7857 9394 7895 9428
rect 7929 9394 7967 9428
rect 8001 9394 8039 9428
rect 8073 9394 8111 9428
rect 8145 9394 8183 9428
rect 8217 9394 8255 9428
rect 8289 9394 8327 9428
rect 8361 9394 8399 9428
rect 8433 9394 8471 9428
rect 8505 9394 8543 9428
rect 8577 9394 8615 9428
rect 8649 9394 8687 9428
rect 8721 9394 8759 9428
rect 8793 9394 8831 9428
rect 8865 9394 8903 9428
rect 8937 9394 8975 9428
rect 9009 9394 9047 9428
rect 9081 9394 9119 9428
rect 9153 9394 9191 9428
rect 9225 9394 9263 9428
rect 9297 9394 9335 9428
rect 9369 9394 9407 9428
rect 9441 9394 9479 9428
rect 9513 9394 9551 9428
rect 9585 9394 9623 9428
rect 9657 9394 9695 9428
rect 9729 9394 9767 9428
rect 9801 9394 9839 9428
rect 9873 9394 9911 9428
rect 9945 9394 9983 9428
rect 10017 9394 10055 9428
rect 10089 9394 10127 9428
rect 10161 9394 10199 9428
rect 10233 9394 10271 9428
rect 10305 9394 10343 9428
rect 10377 9394 10415 9428
rect 10449 9394 10487 9428
rect 10521 9394 10559 9428
rect 10593 9394 10631 9428
rect 10665 9394 10703 9428
rect 10737 9394 10775 9428
rect 10809 9394 10847 9428
rect 10881 9394 10919 9428
rect 10953 9394 10991 9428
rect 11025 9394 11063 9428
rect 11097 9394 11135 9428
rect 11169 9394 11207 9428
rect 11241 9394 11279 9428
rect 11313 9394 11351 9428
rect 11385 9394 11423 9428
rect 11457 9394 11495 9428
rect 11529 9394 11567 9428
rect 11601 9394 11639 9428
rect 11673 9394 11711 9428
rect 11745 9394 11783 9428
rect 11817 9394 11855 9428
rect 11889 9394 11927 9428
rect 11961 9394 11999 9428
rect 12033 9394 12071 9428
rect 12105 9394 12143 9428
rect 12177 9394 12215 9428
rect 12249 9394 12287 9428
rect 12321 9394 12359 9428
rect 12393 9394 12431 9428
rect 12465 9394 12503 9428
rect 12537 9394 12575 9428
rect 12609 9394 12647 9428
rect 12681 9394 12719 9428
rect 12753 9394 12791 9428
rect 12825 9394 12863 9428
rect 12897 9394 12935 9428
rect 12969 9394 13007 9428
rect 13041 9394 13079 9428
rect 13113 9394 13151 9428
rect 13185 9394 13223 9428
rect 13257 9394 13295 9428
rect 13329 9394 13367 9428
rect 13401 9394 13439 9428
rect 13473 9394 13511 9428
rect 13545 9394 13583 9428
rect 13617 9394 13655 9428
rect 13689 9394 13727 9428
rect 13761 9394 13799 9428
rect 13833 9394 13845 9428
rect -496 9359 13845 9394
rect -496 9342 12258 9359
rect 12310 9342 12335 9359
rect 12387 9342 12412 9359
rect 12464 9342 12488 9359
rect -496 9308 -484 9342
rect -450 9308 -411 9342
rect -377 9308 -338 9342
rect -304 9308 -265 9342
rect -231 9308 -192 9342
rect -158 9308 -119 9342
rect -85 9308 -46 9342
rect -12 9308 27 9342
rect 61 9308 100 9342
rect 134 9308 173 9342
rect 207 9308 246 9342
rect 280 9308 319 9342
rect 353 9308 392 9342
rect 426 9308 465 9342
rect 499 9308 538 9342
rect 572 9308 611 9342
rect 645 9308 684 9342
rect 718 9308 757 9342
rect 791 9308 830 9342
rect 864 9308 903 9342
rect 937 9308 976 9342
rect 1010 9308 1049 9342
rect 1083 9308 1122 9342
rect 1156 9308 1195 9342
rect 1229 9308 1268 9342
rect 1302 9308 1341 9342
rect 1375 9308 1414 9342
rect 1448 9308 1487 9342
rect 1521 9308 1559 9342
rect 1593 9308 1631 9342
rect 1665 9308 1703 9342
rect 1737 9308 1775 9342
rect 1809 9308 1847 9342
rect 1881 9308 1919 9342
rect 1953 9308 1991 9342
rect 2025 9308 2063 9342
rect 2097 9308 2135 9342
rect 2169 9308 2207 9342
rect 2241 9308 2279 9342
rect 2313 9308 2351 9342
rect 2385 9308 2423 9342
rect 2457 9308 2495 9342
rect 2529 9308 2567 9342
rect 2601 9308 2639 9342
rect 2673 9308 2711 9342
rect 2745 9308 2783 9342
rect 2817 9308 2855 9342
rect 2889 9308 2927 9342
rect 2961 9308 2999 9342
rect 3033 9308 3071 9342
rect 3105 9308 3143 9342
rect 3177 9308 3215 9342
rect 3249 9308 3287 9342
rect 3321 9308 3359 9342
rect 3393 9308 3431 9342
rect 3465 9308 3503 9342
rect 3537 9308 3575 9342
rect 3609 9308 3647 9342
rect 3681 9308 3719 9342
rect 3753 9308 3791 9342
rect 3825 9308 3863 9342
rect 3897 9308 3935 9342
rect 3969 9308 4007 9342
rect 4041 9308 4079 9342
rect 4113 9308 4151 9342
rect 4185 9308 4223 9342
rect 4257 9308 4295 9342
rect 4329 9308 4367 9342
rect 4401 9308 4439 9342
rect 4473 9308 4511 9342
rect 4545 9308 4583 9342
rect 4617 9308 4655 9342
rect 4689 9308 4727 9342
rect 4761 9308 4799 9342
rect 4833 9308 4871 9342
rect 4905 9308 4943 9342
rect 4977 9308 5015 9342
rect 5049 9308 5087 9342
rect 5121 9308 5159 9342
rect 5193 9308 5231 9342
rect 5265 9308 5303 9342
rect 5337 9308 5375 9342
rect 5409 9308 5447 9342
rect 5481 9308 5519 9342
rect 5553 9308 5591 9342
rect 5625 9308 5663 9342
rect 5697 9308 5735 9342
rect 5769 9308 5807 9342
rect 5841 9308 5879 9342
rect 5913 9308 5951 9342
rect 5985 9308 6023 9342
rect 6057 9308 6095 9342
rect 6129 9308 6167 9342
rect 6201 9308 6239 9342
rect 6273 9308 6311 9342
rect 6345 9308 6383 9342
rect 6417 9308 6455 9342
rect 6489 9308 6527 9342
rect 6561 9308 6599 9342
rect 6633 9308 6671 9342
rect 6705 9308 6743 9342
rect 6777 9308 6815 9342
rect 6849 9308 6887 9342
rect 6921 9308 6959 9342
rect 6993 9308 7031 9342
rect 7065 9308 7103 9342
rect 7137 9308 7175 9342
rect 7209 9308 7247 9342
rect 7281 9308 7319 9342
rect 7353 9308 7391 9342
rect 7425 9308 7463 9342
rect 7497 9308 7535 9342
rect 7569 9308 7607 9342
rect 7641 9308 7679 9342
rect 7713 9308 7751 9342
rect 7785 9308 7823 9342
rect 7857 9308 7895 9342
rect 7929 9308 7967 9342
rect 8001 9308 8039 9342
rect 8073 9308 8111 9342
rect 8145 9308 8183 9342
rect 8217 9308 8255 9342
rect 8289 9308 8327 9342
rect 8361 9308 8399 9342
rect 8433 9308 8471 9342
rect 8505 9308 8543 9342
rect 8577 9308 8615 9342
rect 8649 9308 8687 9342
rect 8721 9308 8759 9342
rect 8793 9308 8831 9342
rect 8865 9308 8903 9342
rect 8937 9308 8975 9342
rect 9009 9308 9047 9342
rect 9081 9308 9119 9342
rect 9153 9308 9191 9342
rect 9225 9308 9263 9342
rect 9297 9308 9335 9342
rect 9369 9308 9407 9342
rect 9441 9308 9479 9342
rect 9513 9308 9551 9342
rect 9585 9308 9623 9342
rect 9657 9308 9695 9342
rect 9729 9308 9767 9342
rect 9801 9308 9839 9342
rect 9873 9308 9911 9342
rect 9945 9308 9983 9342
rect 10017 9308 10055 9342
rect 10089 9308 10127 9342
rect 10161 9308 10199 9342
rect 10233 9308 10271 9342
rect 10305 9308 10343 9342
rect 10377 9308 10415 9342
rect 10449 9308 10487 9342
rect 10521 9308 10559 9342
rect 10593 9308 10631 9342
rect 10665 9308 10703 9342
rect 10737 9308 10775 9342
rect 10809 9308 10847 9342
rect 10881 9308 10919 9342
rect 10953 9308 10991 9342
rect 11025 9308 11063 9342
rect 11097 9308 11135 9342
rect 11169 9308 11207 9342
rect 11241 9308 11279 9342
rect 11313 9308 11351 9342
rect 11385 9308 11423 9342
rect 11457 9308 11495 9342
rect 11529 9308 11567 9342
rect 11601 9308 11639 9342
rect 11673 9308 11711 9342
rect 11745 9308 11783 9342
rect 11817 9308 11855 9342
rect 11889 9308 11927 9342
rect 11961 9308 11999 9342
rect 12033 9308 12071 9342
rect 12105 9308 12143 9342
rect 12177 9308 12215 9342
rect 12249 9308 12258 9342
rect 12321 9308 12335 9342
rect 12393 9308 12412 9342
rect 12465 9308 12488 9342
rect -496 9307 12258 9308
rect 12310 9307 12335 9308
rect 12387 9307 12412 9308
rect 12464 9307 12488 9308
rect 12540 9307 12564 9359
rect 12616 9342 13845 9359
rect 12616 9308 12647 9342
rect 12681 9308 12719 9342
rect 12753 9308 12791 9342
rect 12825 9308 12863 9342
rect 12897 9308 12935 9342
rect 12969 9308 13007 9342
rect 13041 9308 13079 9342
rect 13113 9308 13151 9342
rect 13185 9308 13223 9342
rect 13257 9308 13295 9342
rect 13329 9308 13367 9342
rect 13401 9308 13439 9342
rect 13473 9308 13511 9342
rect 13545 9308 13583 9342
rect 13617 9308 13655 9342
rect 13689 9308 13727 9342
rect 13761 9308 13799 9342
rect 13833 9308 13845 9342
rect 12616 9307 13845 9308
rect -496 9271 13845 9307
rect -496 9256 12258 9271
rect 12310 9256 12335 9271
rect 12387 9256 12412 9271
rect 12464 9256 12488 9271
rect -496 9222 -484 9256
rect -450 9222 -411 9256
rect -377 9222 -338 9256
rect -304 9222 -265 9256
rect -231 9222 -192 9256
rect -158 9222 -119 9256
rect -85 9222 -46 9256
rect -12 9222 27 9256
rect 61 9222 100 9256
rect 134 9222 173 9256
rect 207 9222 246 9256
rect 280 9222 319 9256
rect 353 9222 392 9256
rect 426 9222 465 9256
rect 499 9222 538 9256
rect 572 9222 611 9256
rect 645 9222 684 9256
rect 718 9222 757 9256
rect 791 9222 830 9256
rect 864 9222 903 9256
rect 937 9222 976 9256
rect 1010 9222 1049 9256
rect 1083 9222 1122 9256
rect 1156 9222 1195 9256
rect 1229 9222 1268 9256
rect 1302 9222 1341 9256
rect 1375 9222 1414 9256
rect 1448 9222 1487 9256
rect 1521 9222 1559 9256
rect 1593 9222 1631 9256
rect 1665 9222 1703 9256
rect 1737 9222 1775 9256
rect 1809 9222 1847 9256
rect 1881 9222 1919 9256
rect 1953 9222 1991 9256
rect 2025 9222 2063 9256
rect 2097 9222 2135 9256
rect 2169 9222 2207 9256
rect 2241 9222 2279 9256
rect 2313 9222 2351 9256
rect 2385 9222 2423 9256
rect 2457 9222 2495 9256
rect 2529 9222 2567 9256
rect 2601 9222 2639 9256
rect 2673 9222 2711 9256
rect 2745 9222 2783 9256
rect 2817 9222 2855 9256
rect 2889 9222 2927 9256
rect 2961 9222 2999 9256
rect 3033 9222 3071 9256
rect 3105 9222 3143 9256
rect 3177 9222 3215 9256
rect 3249 9222 3287 9256
rect 3321 9222 3359 9256
rect 3393 9222 3431 9256
rect 3465 9222 3503 9256
rect 3537 9222 3575 9256
rect 3609 9222 3647 9256
rect 3681 9222 3719 9256
rect 3753 9222 3791 9256
rect 3825 9222 3863 9256
rect 3897 9222 3935 9256
rect 3969 9222 4007 9256
rect 4041 9222 4079 9256
rect 4113 9222 4151 9256
rect 4185 9222 4223 9256
rect 4257 9222 4295 9256
rect 4329 9222 4367 9256
rect 4401 9222 4439 9256
rect 4473 9222 4511 9256
rect 4545 9222 4583 9256
rect 4617 9222 4655 9256
rect 4689 9222 4727 9256
rect 4761 9222 4799 9256
rect 4833 9222 4871 9256
rect 4905 9222 4943 9256
rect 4977 9222 5015 9256
rect 5049 9222 5087 9256
rect 5121 9222 5159 9256
rect 5193 9222 5231 9256
rect 5265 9222 5303 9256
rect 5337 9222 5375 9256
rect 5409 9222 5447 9256
rect 5481 9222 5519 9256
rect 5553 9222 5591 9256
rect 5625 9222 5663 9256
rect 5697 9222 5735 9256
rect 5769 9222 5807 9256
rect 5841 9222 5879 9256
rect 5913 9222 5951 9256
rect 5985 9222 6023 9256
rect 6057 9222 6095 9256
rect 6129 9222 6167 9256
rect 6201 9222 6239 9256
rect 6273 9222 6311 9256
rect 6345 9222 6383 9256
rect 6417 9222 6455 9256
rect 6489 9222 6527 9256
rect 6561 9222 6599 9256
rect 6633 9222 6671 9256
rect 6705 9222 6743 9256
rect 6777 9222 6815 9256
rect 6849 9222 6887 9256
rect 6921 9222 6959 9256
rect 6993 9222 7031 9256
rect 7065 9222 7103 9256
rect 7137 9222 7175 9256
rect 7209 9222 7247 9256
rect 7281 9222 7319 9256
rect 7353 9222 7391 9256
rect 7425 9222 7463 9256
rect 7497 9222 7535 9256
rect 7569 9222 7607 9256
rect 7641 9222 7679 9256
rect 7713 9222 7751 9256
rect 7785 9222 7823 9256
rect 7857 9222 7895 9256
rect 7929 9222 7967 9256
rect 8001 9222 8039 9256
rect 8073 9222 8111 9256
rect 8145 9222 8183 9256
rect 8217 9222 8255 9256
rect 8289 9222 8327 9256
rect 8361 9222 8399 9256
rect 8433 9222 8471 9256
rect 8505 9222 8543 9256
rect 8577 9222 8615 9256
rect 8649 9222 8687 9256
rect 8721 9222 8759 9256
rect 8793 9222 8831 9256
rect 8865 9222 8903 9256
rect 8937 9222 8975 9256
rect 9009 9222 9047 9256
rect 9081 9222 9119 9256
rect 9153 9222 9191 9256
rect 9225 9222 9263 9256
rect 9297 9222 9335 9256
rect 9369 9222 9407 9256
rect 9441 9222 9479 9256
rect 9513 9222 9551 9256
rect 9585 9222 9623 9256
rect 9657 9222 9695 9256
rect 9729 9222 9767 9256
rect 9801 9222 9839 9256
rect 9873 9222 9911 9256
rect 9945 9222 9983 9256
rect 10017 9222 10055 9256
rect 10089 9222 10127 9256
rect 10161 9222 10199 9256
rect 10233 9222 10271 9256
rect 10305 9222 10343 9256
rect 10377 9222 10415 9256
rect 10449 9222 10487 9256
rect 10521 9222 10559 9256
rect 10593 9222 10631 9256
rect 10665 9222 10703 9256
rect 10737 9222 10775 9256
rect 10809 9222 10847 9256
rect 10881 9222 10919 9256
rect 10953 9222 10991 9256
rect 11025 9222 11063 9256
rect 11097 9222 11135 9256
rect 11169 9222 11207 9256
rect 11241 9222 11279 9256
rect 11313 9222 11351 9256
rect 11385 9222 11423 9256
rect 11457 9222 11495 9256
rect 11529 9222 11567 9256
rect 11601 9222 11639 9256
rect 11673 9222 11711 9256
rect 11745 9222 11783 9256
rect 11817 9222 11855 9256
rect 11889 9222 11927 9256
rect 11961 9222 11999 9256
rect 12033 9222 12071 9256
rect 12105 9222 12143 9256
rect 12177 9222 12215 9256
rect 12249 9222 12258 9256
rect 12321 9222 12335 9256
rect 12393 9222 12412 9256
rect 12465 9222 12488 9256
rect -496 9219 12258 9222
rect 12310 9219 12335 9222
rect 12387 9219 12412 9222
rect 12464 9219 12488 9222
rect 12540 9219 12564 9271
rect 12616 9256 13845 9271
rect 12616 9222 12647 9256
rect 12681 9222 12719 9256
rect 12753 9222 12791 9256
rect 12825 9222 12863 9256
rect 12897 9222 12935 9256
rect 12969 9222 13007 9256
rect 13041 9222 13079 9256
rect 13113 9222 13151 9256
rect 13185 9222 13223 9256
rect 13257 9222 13295 9256
rect 13329 9222 13367 9256
rect 13401 9222 13439 9256
rect 13473 9222 13511 9256
rect 13545 9222 13583 9256
rect 13617 9222 13655 9256
rect 13689 9222 13727 9256
rect 13761 9222 13799 9256
rect 13833 9222 13845 9256
rect 12616 9219 13845 9222
rect -496 9183 13845 9219
rect -496 9170 12258 9183
rect 12310 9170 12335 9183
rect 12387 9170 12412 9183
rect 12464 9170 12488 9183
rect -496 9136 -484 9170
rect -450 9136 -411 9170
rect -377 9136 -338 9170
rect -304 9136 -265 9170
rect -231 9136 -192 9170
rect -158 9136 -119 9170
rect -85 9136 -46 9170
rect -12 9136 27 9170
rect 61 9136 100 9170
rect 134 9136 173 9170
rect 207 9136 246 9170
rect 280 9136 319 9170
rect 353 9136 392 9170
rect 426 9136 465 9170
rect 499 9136 538 9170
rect 572 9136 611 9170
rect 645 9136 684 9170
rect 718 9136 757 9170
rect 791 9136 830 9170
rect 864 9136 903 9170
rect 937 9136 976 9170
rect 1010 9136 1049 9170
rect 1083 9136 1122 9170
rect 1156 9136 1195 9170
rect 1229 9136 1268 9170
rect 1302 9136 1341 9170
rect 1375 9136 1414 9170
rect 1448 9136 1487 9170
rect 1521 9136 1559 9170
rect 1593 9136 1631 9170
rect 1665 9136 1703 9170
rect 1737 9136 1775 9170
rect 1809 9136 1847 9170
rect 1881 9136 1919 9170
rect 1953 9136 1991 9170
rect 2025 9136 2063 9170
rect 2097 9136 2135 9170
rect 2169 9136 2207 9170
rect 2241 9136 2279 9170
rect 2313 9136 2351 9170
rect 2385 9136 2423 9170
rect 2457 9136 2495 9170
rect 2529 9136 2567 9170
rect 2601 9136 2639 9170
rect 2673 9136 2711 9170
rect 2745 9136 2783 9170
rect 2817 9136 2855 9170
rect 2889 9136 2927 9170
rect 2961 9136 2999 9170
rect 3033 9136 3071 9170
rect 3105 9136 3143 9170
rect 3177 9136 3215 9170
rect 3249 9136 3287 9170
rect 3321 9136 3359 9170
rect 3393 9136 3431 9170
rect 3465 9136 3503 9170
rect 3537 9136 3575 9170
rect 3609 9136 3647 9170
rect 3681 9136 3719 9170
rect 3753 9136 3791 9170
rect 3825 9136 3863 9170
rect 3897 9136 3935 9170
rect 3969 9136 4007 9170
rect 4041 9136 4079 9170
rect 4113 9136 4151 9170
rect 4185 9136 4223 9170
rect 4257 9136 4295 9170
rect 4329 9136 4367 9170
rect 4401 9136 4439 9170
rect 4473 9136 4511 9170
rect 4545 9136 4583 9170
rect 4617 9136 4655 9170
rect 4689 9136 4727 9170
rect 4761 9136 4799 9170
rect 4833 9136 4871 9170
rect 4905 9136 4943 9170
rect 4977 9136 5015 9170
rect 5049 9136 5087 9170
rect 5121 9136 5159 9170
rect 5193 9136 5231 9170
rect 5265 9136 5303 9170
rect 5337 9136 5375 9170
rect 5409 9136 5447 9170
rect 5481 9136 5519 9170
rect 5553 9136 5591 9170
rect 5625 9136 5663 9170
rect 5697 9136 5735 9170
rect 5769 9136 5807 9170
rect 5841 9136 5879 9170
rect 5913 9136 5951 9170
rect 5985 9136 6023 9170
rect 6057 9136 6095 9170
rect 6129 9136 6167 9170
rect 6201 9136 6239 9170
rect 6273 9136 6311 9170
rect 6345 9136 6383 9170
rect 6417 9136 6455 9170
rect 6489 9136 6527 9170
rect 6561 9136 6599 9170
rect 6633 9136 6671 9170
rect 6705 9136 6743 9170
rect 6777 9136 6815 9170
rect 6849 9136 6887 9170
rect 6921 9136 6959 9170
rect 6993 9136 7031 9170
rect 7065 9136 7103 9170
rect 7137 9136 7175 9170
rect 7209 9136 7247 9170
rect 7281 9136 7319 9170
rect 7353 9136 7391 9170
rect 7425 9136 7463 9170
rect 7497 9136 7535 9170
rect 7569 9136 7607 9170
rect 7641 9136 7679 9170
rect 7713 9136 7751 9170
rect 7785 9136 7823 9170
rect 7857 9136 7895 9170
rect 7929 9136 7967 9170
rect 8001 9136 8039 9170
rect 8073 9136 8111 9170
rect 8145 9136 8183 9170
rect 8217 9136 8255 9170
rect 8289 9136 8327 9170
rect 8361 9136 8399 9170
rect 8433 9136 8471 9170
rect 8505 9136 8543 9170
rect 8577 9136 8615 9170
rect 8649 9136 8687 9170
rect 8721 9136 8759 9170
rect 8793 9136 8831 9170
rect 8865 9136 8903 9170
rect 8937 9136 8975 9170
rect 9009 9136 9047 9170
rect 9081 9136 9119 9170
rect 9153 9136 9191 9170
rect 9225 9136 9263 9170
rect 9297 9136 9335 9170
rect 9369 9136 9407 9170
rect 9441 9136 9479 9170
rect 9513 9136 9551 9170
rect 9585 9136 9623 9170
rect 9657 9136 9695 9170
rect 9729 9136 9767 9170
rect 9801 9136 9839 9170
rect 9873 9136 9911 9170
rect 9945 9136 9983 9170
rect 10017 9136 10055 9170
rect 10089 9136 10127 9170
rect 10161 9136 10199 9170
rect 10233 9136 10271 9170
rect 10305 9136 10343 9170
rect 10377 9136 10415 9170
rect 10449 9136 10487 9170
rect 10521 9136 10559 9170
rect 10593 9136 10631 9170
rect 10665 9136 10703 9170
rect 10737 9136 10775 9170
rect 10809 9136 10847 9170
rect 10881 9136 10919 9170
rect 10953 9136 10991 9170
rect 11025 9136 11063 9170
rect 11097 9136 11135 9170
rect 11169 9136 11207 9170
rect 11241 9136 11279 9170
rect 11313 9136 11351 9170
rect 11385 9136 11423 9170
rect 11457 9136 11495 9170
rect 11529 9136 11567 9170
rect 11601 9136 11639 9170
rect 11673 9136 11711 9170
rect 11745 9136 11783 9170
rect 11817 9136 11855 9170
rect 11889 9136 11927 9170
rect 11961 9136 11999 9170
rect 12033 9136 12071 9170
rect 12105 9136 12143 9170
rect 12177 9136 12215 9170
rect 12249 9136 12258 9170
rect 12321 9136 12335 9170
rect 12393 9136 12412 9170
rect 12465 9136 12488 9170
rect -496 9131 12258 9136
rect 12310 9131 12335 9136
rect 12387 9131 12412 9136
rect 12464 9131 12488 9136
rect 12540 9131 12564 9183
rect 12616 9170 13845 9183
rect 12616 9136 12647 9170
rect 12681 9136 12719 9170
rect 12753 9136 12791 9170
rect 12825 9136 12863 9170
rect 12897 9136 12935 9170
rect 12969 9136 13007 9170
rect 13041 9136 13079 9170
rect 13113 9136 13151 9170
rect 13185 9136 13223 9170
rect 13257 9136 13295 9170
rect 13329 9136 13367 9170
rect 13401 9136 13439 9170
rect 13473 9136 13511 9170
rect 13545 9136 13583 9170
rect 13617 9136 13655 9170
rect 13689 9136 13727 9170
rect 13761 9136 13799 9170
rect 13833 9136 13845 9170
rect 12616 9131 13845 9136
rect -496 9129 13845 9131
rect 14206 9460 15114 9829
rect 14206 9408 14240 9460
rect 14292 9408 14312 9460
rect 14364 9408 14384 9460
rect 14436 9408 14456 9460
rect 14508 9408 14528 9460
rect 14580 9408 14600 9460
rect 14652 9408 15114 9460
rect 14206 9395 15114 9408
rect 14206 9343 14240 9395
rect 14292 9343 14312 9395
rect 14364 9343 14384 9395
rect 14436 9343 14456 9395
rect 14508 9343 14528 9395
rect 14580 9343 14600 9395
rect 14652 9343 15114 9395
rect 14206 9330 15114 9343
rect 14206 9278 14240 9330
rect 14292 9278 14312 9330
rect 14364 9278 14384 9330
rect 14436 9278 14456 9330
rect 14508 9278 14528 9330
rect 14580 9278 14600 9330
rect 14652 9278 15114 9330
rect 14206 9265 15114 9278
rect 14206 9213 14240 9265
rect 14292 9213 14312 9265
rect 14364 9213 14384 9265
rect 14436 9213 14456 9265
rect 14508 9213 14528 9265
rect 14580 9213 14600 9265
rect 14652 9213 15114 9265
rect 14206 9200 15114 9213
rect 14206 9148 14240 9200
rect 14292 9148 14312 9200
rect 14364 9148 14384 9200
rect 14436 9148 14456 9200
rect 14508 9148 14528 9200
rect 14580 9148 14600 9200
rect 14652 9148 15114 9200
rect 14206 9135 15114 9148
rect 14206 9083 14240 9135
rect 14292 9083 14312 9135
rect 14364 9083 14384 9135
rect 14436 9083 14456 9135
rect 14508 9083 14528 9135
rect 14580 9083 14600 9135
rect 14652 9083 15114 9135
rect 14206 9070 15114 9083
rect 14206 9018 14240 9070
rect 14292 9018 14312 9070
rect 14364 9018 14384 9070
rect 14436 9018 14456 9070
rect 14508 9018 14528 9070
rect 14580 9018 14600 9070
rect 14652 9018 15114 9070
rect 14206 9005 15114 9018
tri 14031 8828 14206 9003 se
rect 14206 8953 14240 9005
rect 14292 8953 14312 9005
rect 14364 8953 14384 9005
rect 14436 8953 14456 9005
rect 14508 8953 14528 9005
rect 14580 8953 14600 9005
rect 14652 8953 15114 9005
rect 14206 8940 15114 8953
rect 14206 8888 14240 8940
rect 14292 8888 14312 8940
rect 14364 8888 14384 8940
rect 14436 8888 14456 8940
rect 14508 8888 14528 8940
rect 14580 8888 14600 8940
rect 14652 8888 15114 8940
rect 14206 8875 15114 8888
rect 14206 8828 14240 8875
rect 56 8827 14240 8828
rect 56 8775 541 8827
rect 593 8775 616 8827
rect 668 8775 690 8827
rect 742 8775 764 8827
rect 816 8775 838 8827
rect 890 8775 912 8827
rect 964 8823 14240 8827
rect 14292 8823 14312 8875
rect 14364 8823 14384 8875
rect 14436 8823 14456 8875
rect 14508 8823 14528 8875
rect 14580 8823 14600 8875
rect 14652 8823 15114 8875
rect 964 8810 15114 8823
rect 964 8775 14240 8810
rect 56 8760 14240 8775
rect 14292 8760 14312 8810
rect 14364 8760 14384 8810
rect 14436 8760 14456 8810
rect 14508 8760 14528 8810
rect 14580 8760 14600 8810
rect 14652 8760 15114 8810
rect 56 8753 912 8760
rect 56 8719 248 8753
rect 282 8719 322 8753
rect 356 8719 396 8753
rect 430 8719 470 8753
rect 504 8751 544 8753
rect 578 8751 618 8753
rect 652 8751 691 8753
rect 725 8751 764 8753
rect 798 8751 837 8753
rect 871 8751 912 8753
rect 946 8751 984 8760
rect 504 8719 541 8751
rect 56 8699 541 8719
rect 593 8699 616 8751
rect 668 8699 690 8751
rect 742 8699 764 8751
rect 816 8719 837 8751
rect 816 8699 838 8719
rect 890 8699 912 8751
rect 964 8726 984 8751
rect 1018 8726 1056 8760
rect 1090 8726 1128 8760
rect 1162 8726 1200 8760
rect 1234 8726 1272 8760
rect 1306 8726 1344 8760
rect 1378 8726 1416 8760
rect 1450 8726 1488 8760
rect 1522 8726 1560 8760
rect 1594 8726 1632 8760
rect 1666 8726 1704 8760
rect 1738 8726 1776 8760
rect 1810 8726 1849 8760
rect 1883 8726 1922 8760
rect 1956 8726 1995 8760
rect 2029 8726 2068 8760
rect 2102 8726 2141 8760
rect 2175 8753 3477 8760
rect 2175 8726 2227 8753
rect 964 8719 2227 8726
rect 2261 8719 2306 8753
rect 2340 8719 2385 8753
rect 2419 8719 2464 8753
rect 2498 8719 2543 8753
rect 2577 8719 2621 8753
rect 2655 8719 2699 8753
rect 2733 8719 2777 8753
rect 2811 8719 2855 8753
rect 2889 8719 2933 8753
rect 2967 8719 3011 8753
rect 3045 8726 3477 8753
rect 3511 8726 3550 8760
rect 3584 8726 3623 8760
rect 3657 8726 3696 8760
rect 3730 8726 3769 8760
rect 3803 8726 3842 8760
rect 3876 8726 3915 8760
rect 3949 8726 3988 8760
rect 4022 8726 4061 8760
rect 4095 8726 4134 8760
rect 4168 8726 4207 8760
rect 4241 8726 4280 8760
rect 4314 8726 4353 8760
rect 4387 8726 4426 8760
rect 4460 8726 4499 8760
rect 4533 8726 4572 8760
rect 4606 8726 4645 8760
rect 4679 8726 4718 8760
rect 4752 8726 4791 8760
rect 4825 8726 4864 8760
rect 4898 8726 4937 8760
rect 4971 8726 5010 8760
rect 5044 8726 5083 8760
rect 5117 8726 5156 8760
rect 5190 8726 5229 8760
rect 5263 8726 5302 8760
rect 5336 8726 5375 8760
rect 5409 8726 5448 8760
rect 5482 8726 5521 8760
rect 5555 8726 5594 8760
rect 5628 8726 5667 8760
rect 5701 8726 5740 8760
rect 5774 8726 5813 8760
rect 5847 8726 5886 8760
rect 5920 8726 5959 8760
rect 5993 8726 6032 8760
rect 6066 8726 6105 8760
rect 6139 8726 6178 8760
rect 6212 8726 6251 8760
rect 6285 8726 6324 8760
rect 6358 8726 6397 8760
rect 6431 8726 6470 8760
rect 6504 8726 6543 8760
rect 6577 8726 6616 8760
rect 6650 8726 6689 8760
rect 6723 8726 6762 8760
rect 6796 8726 6835 8760
rect 6869 8726 6908 8760
rect 6942 8726 6981 8760
rect 7015 8726 7054 8760
rect 7088 8726 7127 8760
rect 7161 8726 7200 8760
rect 7234 8726 7273 8760
rect 7307 8726 7346 8760
rect 7380 8726 7419 8760
rect 7453 8726 7492 8760
rect 7526 8726 7565 8760
rect 7599 8726 7638 8760
rect 7672 8726 7711 8760
rect 7745 8726 7784 8760
rect 7818 8726 7857 8760
rect 7891 8726 7930 8760
rect 7964 8726 8003 8760
rect 8037 8726 8075 8760
rect 8109 8726 8147 8760
rect 8181 8726 8219 8760
rect 8253 8726 8291 8760
rect 8325 8726 8363 8760
rect 8397 8726 8435 8760
rect 8469 8726 8507 8760
rect 8541 8726 8579 8760
rect 8613 8726 8651 8760
rect 8685 8726 8723 8760
rect 8757 8726 8795 8760
rect 8829 8726 8867 8760
rect 8901 8726 8939 8760
rect 8973 8726 9011 8760
rect 9045 8726 9083 8760
rect 9117 8726 9155 8760
rect 9189 8726 9227 8760
rect 9261 8726 9299 8760
rect 9333 8726 9371 8760
rect 9405 8726 9443 8760
rect 9477 8726 9515 8760
rect 9549 8726 9587 8760
rect 9621 8726 9659 8760
rect 9693 8726 9731 8760
rect 9765 8726 9803 8760
rect 9837 8726 9875 8760
rect 9909 8726 9947 8760
rect 9981 8726 10019 8760
rect 10053 8726 10091 8760
rect 10125 8726 10163 8760
rect 10197 8726 10235 8760
rect 10269 8726 10307 8760
rect 10341 8726 10379 8760
rect 10413 8726 10451 8760
rect 10485 8726 10523 8760
rect 10557 8726 10595 8760
rect 10629 8726 10667 8760
rect 10701 8726 10739 8760
rect 10773 8726 10811 8760
rect 10845 8726 10883 8760
rect 10917 8726 10955 8760
rect 10989 8726 11027 8760
rect 11061 8726 11099 8760
rect 11133 8726 11171 8760
rect 11205 8726 11243 8760
rect 11277 8726 11315 8760
rect 11349 8726 11387 8760
rect 11421 8726 11459 8760
rect 11493 8726 11531 8760
rect 11565 8726 11603 8760
rect 11637 8726 11675 8760
rect 11709 8726 11747 8760
rect 11781 8726 11819 8760
rect 11853 8726 11891 8760
rect 11925 8726 11963 8760
rect 11997 8726 12035 8760
rect 12069 8726 12107 8760
rect 12141 8726 12179 8760
rect 12213 8726 12251 8760
rect 12285 8726 12323 8760
rect 12357 8726 12395 8760
rect 12429 8726 12467 8760
rect 12501 8726 12539 8760
rect 12573 8726 12611 8760
rect 12645 8726 12683 8760
rect 12717 8726 12755 8760
rect 12789 8726 12827 8760
rect 12861 8726 12899 8760
rect 12933 8726 12971 8760
rect 13005 8726 13043 8760
rect 13077 8726 13115 8760
rect 13149 8726 13187 8760
rect 13221 8726 13259 8760
rect 13293 8726 13331 8760
rect 13365 8726 13403 8760
rect 13437 8726 13475 8760
rect 13509 8726 13547 8760
rect 13581 8726 13619 8760
rect 13653 8726 13691 8760
rect 13725 8726 13763 8760
rect 13797 8726 13835 8760
rect 13869 8726 13907 8760
rect 13941 8726 13979 8760
rect 14013 8726 14051 8760
rect 14085 8726 14123 8760
rect 14157 8726 14195 8760
rect 14229 8758 14240 8760
rect 14301 8758 14312 8760
rect 14373 8758 14384 8760
rect 14445 8758 14456 8760
rect 14517 8758 14528 8760
rect 14589 8758 14600 8760
rect 14229 8745 14267 8758
rect 14301 8745 14339 8758
rect 14373 8745 14411 8758
rect 14445 8745 14483 8758
rect 14517 8745 14555 8758
rect 14589 8745 14627 8758
rect 14229 8726 14240 8745
rect 14301 8726 14312 8745
rect 14373 8726 14384 8745
rect 14445 8726 14456 8745
rect 14517 8726 14528 8745
rect 14589 8726 14600 8745
rect 14661 8726 14699 8760
rect 14733 8726 14771 8760
rect 14805 8726 14843 8760
rect 14877 8726 15114 8760
rect 3045 8719 14240 8726
rect 964 8713 14240 8719
rect 964 8699 2306 8713
tri 2306 8699 2320 8713 nw
tri 3344 8699 3358 8713 ne
rect 3358 8699 14240 8713
tri 728 8693 734 8699 ne
rect 734 8693 2243 8699
tri 734 8636 791 8693 ne
rect 791 8670 2243 8693
rect 791 8636 842 8670
tri 791 8602 825 8636 ne
rect 825 8618 842 8636
rect 894 8618 912 8670
rect 964 8636 2243 8670
tri 2243 8636 2306 8699 nw
tri 3358 8636 3421 8699 ne
rect 3421 8693 14240 8699
rect 14292 8693 14312 8726
rect 14364 8693 14384 8726
rect 14436 8693 14456 8726
rect 14508 8693 14528 8726
rect 14580 8693 14600 8726
rect 14652 8693 15114 8726
rect 3421 8680 15114 8693
rect 3421 8636 14240 8680
rect 14292 8636 14312 8680
rect 14364 8636 14384 8680
rect 14436 8636 14456 8680
rect 14508 8636 14528 8680
rect 14580 8636 14600 8680
rect 14652 8636 15114 8680
rect 964 8618 984 8636
rect 825 8602 912 8618
rect 946 8602 984 8618
rect 1018 8602 1056 8636
rect 1090 8602 1128 8636
rect 1162 8602 1200 8636
rect 1234 8602 1272 8636
rect 1306 8602 1344 8636
rect 1378 8602 1416 8636
rect 1450 8602 1488 8636
rect 1522 8602 1560 8636
rect 1594 8602 1632 8636
rect 1666 8602 1704 8636
rect 1738 8602 1776 8636
rect 1810 8602 1849 8636
rect 1883 8602 1922 8636
rect 1956 8602 1995 8636
rect 2029 8602 2068 8636
rect 2102 8602 2141 8636
rect 2175 8602 2209 8636
tri 2209 8602 2243 8636 nw
tri 3421 8602 3455 8636 ne
rect 3455 8602 3477 8636
rect 3511 8602 3550 8636
rect 3584 8602 3623 8636
rect 3657 8602 3696 8636
rect 3730 8602 3769 8636
rect 3803 8602 3842 8636
rect 3876 8602 3915 8636
rect 3949 8602 3988 8636
rect 4022 8602 4061 8636
rect 4095 8602 4134 8636
rect 4168 8602 4207 8636
rect 4241 8602 4280 8636
rect 4314 8602 4353 8636
rect 4387 8602 4426 8636
rect 4460 8602 4499 8636
rect 4533 8602 4572 8636
rect 4606 8602 4645 8636
rect 4679 8602 4718 8636
rect 4752 8602 4791 8636
rect 4825 8602 4864 8636
rect 4898 8602 4937 8636
rect 4971 8602 5010 8636
rect 5044 8602 5083 8636
rect 5117 8602 5156 8636
rect 5190 8602 5229 8636
rect 5263 8602 5302 8636
rect 5336 8602 5375 8636
rect 5409 8602 5448 8636
rect 5482 8602 5521 8636
rect 5555 8602 5594 8636
rect 5628 8602 5667 8636
rect 5701 8602 5740 8636
rect 5774 8602 5813 8636
rect 5847 8602 5886 8636
rect 5920 8602 5959 8636
rect 5993 8602 6032 8636
rect 6066 8602 6105 8636
rect 6139 8602 6178 8636
rect 6212 8602 6251 8636
rect 6285 8602 6324 8636
rect 6358 8602 6397 8636
rect 6431 8602 6470 8636
rect 6504 8602 6543 8636
rect 6577 8602 6616 8636
rect 6650 8602 6689 8636
rect 6723 8602 6762 8636
rect 6796 8602 6835 8636
rect 6869 8602 6908 8636
rect 6942 8602 6981 8636
rect 7015 8602 7054 8636
rect 7088 8602 7127 8636
rect 7161 8602 7200 8636
rect 7234 8602 7273 8636
rect 7307 8602 7346 8636
rect 7380 8602 7419 8636
rect 7453 8602 7492 8636
rect 7526 8602 7565 8636
rect 7599 8602 7638 8636
rect 7672 8602 7711 8636
rect 7745 8602 7784 8636
rect 7818 8602 7857 8636
rect 7891 8602 7930 8636
rect 7964 8602 8003 8636
rect 8037 8602 8075 8636
rect 8109 8602 8147 8636
rect 8181 8602 8219 8636
rect 8253 8602 8291 8636
rect 8325 8602 8363 8636
rect 8397 8602 8435 8636
rect 8469 8602 8507 8636
rect 8541 8602 8579 8636
rect 8613 8602 8651 8636
rect 8685 8602 8723 8636
rect 8757 8602 8795 8636
rect 8829 8602 8867 8636
rect 8901 8602 8939 8636
rect 8973 8602 9011 8636
rect 9045 8602 9083 8636
rect 9117 8602 9155 8636
rect 9189 8602 9227 8636
rect 9261 8602 9299 8636
rect 9333 8602 9371 8636
rect 9405 8602 9443 8636
rect 9477 8602 9515 8636
rect 9549 8602 9587 8636
rect 9621 8602 9659 8636
rect 9693 8602 9731 8636
rect 9765 8602 9803 8636
rect 9837 8602 9875 8636
rect 9909 8602 9947 8636
rect 9981 8602 10019 8636
rect 10053 8602 10091 8636
rect 10125 8602 10163 8636
rect 10197 8602 10235 8636
rect 10269 8602 10307 8636
rect 10341 8602 10379 8636
rect 10413 8602 10451 8636
rect 10485 8602 10523 8636
rect 10557 8602 10595 8636
rect 10629 8602 10667 8636
rect 10701 8602 10739 8636
rect 10773 8602 10811 8636
rect 10845 8602 10883 8636
rect 10917 8602 10955 8636
rect 10989 8602 11027 8636
rect 11061 8602 11099 8636
rect 11133 8602 11171 8636
rect 11205 8602 11243 8636
rect 11277 8602 11315 8636
rect 11349 8602 11387 8636
rect 11421 8602 11459 8636
rect 11493 8602 11531 8636
rect 11565 8602 11603 8636
rect 11637 8602 11675 8636
rect 11709 8602 11747 8636
rect 11781 8602 11819 8636
rect 11853 8602 11891 8636
rect 11925 8602 11963 8636
rect 11997 8602 12035 8636
rect 12069 8602 12107 8636
rect 12141 8602 12179 8636
rect 12213 8602 12251 8636
rect 12285 8602 12323 8636
rect 12357 8602 12395 8636
rect 12429 8602 12467 8636
rect 12501 8602 12539 8636
rect 12573 8602 12611 8636
rect 12645 8602 12683 8636
rect 12717 8602 12755 8636
rect 12789 8602 12827 8636
rect 12861 8602 12899 8636
rect 12933 8602 12971 8636
rect 13005 8602 13043 8636
rect 13077 8602 13115 8636
rect 13149 8602 13187 8636
rect 13221 8602 13259 8636
rect 13293 8602 13331 8636
rect 13365 8602 13403 8636
rect 13437 8602 13475 8636
rect 13509 8602 13547 8636
rect 13581 8602 13619 8636
rect 13653 8602 13691 8636
rect 13725 8602 13763 8636
rect 13797 8602 13835 8636
rect 13869 8602 13907 8636
rect 13941 8602 13979 8636
rect 14013 8602 14051 8636
rect 14085 8602 14123 8636
rect 14157 8602 14195 8636
rect 14229 8628 14240 8636
rect 14301 8628 14312 8636
rect 14373 8628 14384 8636
rect 14445 8628 14456 8636
rect 14517 8628 14528 8636
rect 14589 8628 14600 8636
rect 14229 8615 14267 8628
rect 14301 8615 14339 8628
rect 14373 8615 14411 8628
rect 14445 8615 14483 8628
rect 14517 8615 14555 8628
rect 14589 8615 14627 8628
rect 14229 8602 14240 8615
rect 14301 8602 14312 8615
rect 14373 8602 14384 8615
rect 14445 8602 14456 8615
rect 14517 8602 14528 8615
rect 14589 8602 14600 8615
rect 14661 8602 14699 8636
rect 14733 8602 14771 8636
rect 14805 8602 14843 8636
rect 14877 8602 15114 8636
tri 825 8595 832 8602 ne
rect 832 8595 2194 8602
tri 832 8587 840 8595 ne
rect 840 8587 2194 8595
tri 2194 8587 2209 8602 nw
tri 3455 8596 3461 8602 ne
rect 3461 8596 14240 8602
tri 3461 8587 3470 8596 ne
rect 3470 8587 14240 8596
tri 13739 8558 13768 8587 ne
rect 13768 8563 14240 8587
rect 14292 8563 14312 8602
rect 14364 8563 14384 8602
rect 14436 8563 14456 8602
rect 14508 8563 14528 8602
rect 14580 8563 14600 8602
rect 14652 8563 15114 8602
rect 13768 8558 15114 8563
tri 13768 8546 13780 8558 ne
rect 13780 8550 15114 8558
rect 13780 8546 14240 8550
tri 13780 8512 13814 8546 ne
rect 13814 8512 13992 8546
rect 14026 8512 14076 8546
rect 14110 8512 14240 8546
tri 13814 8478 13848 8512 ne
rect 13848 8478 14185 8512
rect 14219 8498 14240 8512
rect 14292 8498 14312 8550
rect 14364 8498 14384 8550
rect 14436 8498 14456 8550
rect 14508 8498 14528 8550
rect 14580 8498 14600 8550
rect 14652 8498 15114 8550
rect 14219 8485 14257 8498
rect 14291 8485 14329 8498
rect 14363 8485 14401 8498
rect 14435 8485 14473 8498
rect 14507 8485 15114 8498
rect 14219 8478 14240 8485
tri 13848 8474 13852 8478 ne
rect 13852 8474 14240 8478
tri 13852 8440 13886 8474 ne
rect 13886 8440 13992 8474
rect 14026 8440 14076 8474
rect 14110 8440 14240 8474
tri 13886 8435 13891 8440 ne
rect 13891 8435 14240 8440
tri 13891 8401 13925 8435 ne
rect 13925 8401 14185 8435
rect 14219 8433 14240 8435
rect 14292 8433 14312 8485
rect 14364 8433 14384 8485
rect 14436 8433 14456 8485
rect 14508 8433 14528 8485
rect 14580 8433 14600 8485
rect 14652 8462 15114 8485
rect 14652 8433 14692 8462
rect 14219 8420 14257 8433
rect 14291 8420 14329 8433
rect 14363 8420 14401 8433
rect 14435 8420 14473 8433
rect 14507 8428 14614 8433
rect 14648 8428 14692 8433
rect 14726 8428 14770 8462
rect 14804 8428 14848 8462
rect 14882 8428 14926 8462
rect 14960 8428 15004 8462
rect 15038 8428 15114 8462
rect 14507 8420 15114 8428
rect 14219 8401 14240 8420
tri 13925 8367 13959 8401 ne
rect 13959 8367 13992 8401
rect 14026 8367 14076 8401
rect 14110 8368 14240 8401
rect 14292 8368 14312 8420
rect 14364 8368 14384 8420
rect 14436 8368 14456 8420
rect 14508 8368 14528 8420
rect 14580 8368 14600 8420
rect 14652 8388 15114 8420
rect 14652 8368 14692 8388
rect 14110 8367 14614 8368
tri 13959 8360 13966 8367 ne
rect 13966 8360 14614 8367
rect 2496 8314 2549 8360
tri 13966 8358 13968 8360 ne
rect 13968 8358 14614 8360
tri 13968 8355 13971 8358 ne
rect 13971 8355 14185 8358
tri 13971 8324 14002 8355 ne
rect 14002 8324 14185 8355
rect 14219 8354 14257 8358
rect 14291 8354 14329 8358
rect 14363 8354 14401 8358
rect 14435 8354 14473 8358
rect 14507 8354 14614 8358
rect 14648 8354 14692 8368
rect 14726 8354 14770 8388
rect 14804 8354 14848 8388
rect 14882 8354 14926 8388
rect 14960 8354 15004 8388
rect 15038 8354 15114 8388
rect 14219 8324 14240 8354
tri 14002 8314 14012 8324 ne
rect 14012 8314 14240 8324
tri 14012 8287 14039 8314 ne
rect 14039 8302 14240 8314
rect 14292 8302 14312 8354
rect 14364 8302 14384 8354
rect 14436 8302 14456 8354
rect 14508 8302 14528 8354
rect 14580 8302 14600 8354
rect 14652 8314 15114 8354
rect 14652 8302 14692 8314
rect 14039 8288 14614 8302
rect 14648 8288 14692 8302
rect 14039 8287 14240 8288
rect 10798 8281 11156 8287
tri 7008 8254 7014 8260 se
rect 7014 8254 8627 8260
tri 6686 7932 7008 8254 se
rect 7008 7932 8509 8254
rect 8615 7932 8627 8254
rect 9590 8247 9881 8259
rect 9883 8258 10183 8259
rect 9590 8213 9596 8247
rect 9630 8213 9678 8247
rect 9712 8213 9881 8247
rect 9590 8144 9881 8213
rect 9590 8110 9596 8144
rect 9630 8110 9678 8144
rect 9712 8110 9881 8144
rect 9590 8041 9881 8110
rect 9590 8007 9596 8041
rect 9630 8007 9678 8041
rect 9712 8007 9881 8041
rect 9590 7995 9881 8007
rect 9882 7996 10184 8258
rect 10185 8247 10436 8259
rect 10185 8213 10314 8247
rect 10348 8213 10396 8247
rect 10430 8213 10436 8247
rect 10185 8144 10436 8213
rect 10185 8110 10314 8144
rect 10348 8110 10396 8144
rect 10430 8110 10436 8144
rect 10185 8041 10436 8110
rect 10185 8007 10314 8041
rect 10348 8007 10396 8041
rect 10430 8007 10436 8041
rect 9883 7995 10183 7996
rect 10185 7995 10436 8007
rect 10798 8229 10800 8281
rect 10852 8229 10876 8281
rect 10928 8254 10952 8281
rect 10932 8229 10952 8254
rect 11004 8229 11028 8281
rect 11080 8229 11104 8281
rect 10798 8220 10804 8229
rect 10838 8220 10898 8229
rect 10932 8220 11156 8229
rect 10798 8214 11156 8220
rect 10798 8162 10800 8214
rect 10852 8162 10876 8214
rect 10928 8179 10952 8214
rect 10932 8162 10952 8179
rect 11004 8162 11028 8214
rect 11080 8162 11104 8214
rect 10798 8147 10804 8162
rect 10838 8147 10898 8162
rect 10932 8147 11156 8162
rect 10798 8095 10800 8147
rect 10852 8095 10876 8147
rect 10932 8145 10952 8147
rect 10928 8104 10952 8145
rect 10932 8095 10952 8104
rect 11004 8095 11028 8147
rect 11080 8095 11104 8147
rect 10798 8079 10804 8095
rect 10838 8079 10898 8095
rect 10932 8079 11156 8095
rect 10798 8027 10800 8079
rect 10852 8027 10876 8079
rect 10932 8070 10952 8079
rect 10928 8028 10952 8070
rect 10932 8027 10952 8028
rect 11004 8027 11028 8079
rect 11080 8027 11104 8079
rect 10798 8011 10804 8027
rect 10838 8011 10898 8027
rect 10932 8011 11156 8027
tri 6672 7918 6686 7932 se
rect 6686 7926 8627 7932
rect 10798 7959 10800 8011
rect 10852 7959 10876 8011
rect 10932 7994 10952 8011
rect 10928 7959 10952 7994
rect 11004 7959 11028 8011
rect 11080 7959 11104 8011
rect 10798 7952 11156 7959
rect 10798 7943 10804 7952
rect 10838 7943 10898 7952
rect 10932 7943 11156 7952
rect 6686 7918 7144 7926
tri 7144 7918 7152 7926 nw
tri 6670 7916 6672 7918 se
rect 6672 7916 7142 7918
tri 7142 7916 7144 7918 nw
tri 6664 7910 6670 7916 se
rect 6670 7910 7136 7916
tri 7136 7910 7142 7916 nw
tri 6660 7906 6664 7910 se
rect 6664 7906 7132 7910
tri 7132 7906 7136 7910 nw
tri 6624 7870 6660 7906 se
rect 6660 7870 7096 7906
tri 7096 7870 7132 7906 nw
rect 10798 7891 10800 7943
rect 10852 7891 10876 7943
rect 10932 7918 10952 7943
rect 10928 7891 10952 7918
rect 11004 7891 11028 7943
rect 11080 7891 11104 7943
rect 10798 7885 11156 7891
rect 12252 8281 12622 8287
rect 12252 8229 12255 8281
rect 12307 8229 12333 8281
rect 12385 8229 12411 8281
rect 12463 8229 12489 8281
rect 12541 8229 12567 8281
rect 12619 8229 12622 8281
tri 14039 8280 14046 8287 ne
rect 14046 8280 14240 8287
tri 14046 8257 14069 8280 ne
rect 14069 8257 14185 8280
rect 12252 8210 12622 8229
rect 12252 8158 12255 8210
rect 12307 8158 12333 8210
rect 12385 8158 12411 8210
rect 12463 8158 12489 8210
rect 12541 8158 12567 8210
rect 12619 8158 12622 8210
rect 12252 8139 12622 8158
rect 12252 8087 12255 8139
rect 12307 8087 12333 8139
rect 12385 8087 12411 8139
rect 12463 8087 12489 8139
rect 12541 8087 12567 8139
rect 12619 8087 12622 8139
rect 12252 8068 12622 8087
rect 12252 8016 12255 8068
rect 12307 8016 12333 8068
rect 12385 8016 12411 8068
rect 12463 8016 12489 8068
rect 12541 8016 12567 8068
rect 12619 8033 12622 8068
tri 12622 8033 12645 8056 sw
rect 12619 8016 12645 8033
rect 12252 7999 12645 8016
tri 12645 7999 12679 8033 sw
rect 12252 7997 12679 7999
rect 12252 7945 12255 7997
rect 12307 7945 12333 7997
rect 12385 7945 12411 7997
rect 12463 7945 12489 7997
rect 12541 7945 12567 7997
rect 12619 7984 12679 7997
tri 12679 7984 12694 7999 sw
rect 12619 7950 12694 7984
tri 12694 7950 12728 7984 sw
rect 12619 7945 12728 7950
rect 12252 7925 12728 7945
rect 12252 7873 12255 7925
rect 12307 7873 12333 7925
rect 12385 7873 12411 7925
rect 12463 7873 12489 7925
rect 12541 7873 12567 7925
rect 12619 7916 12728 7925
tri 12728 7916 12762 7950 sw
rect 13310 7924 13365 8257
tri 14069 8246 14080 8257 ne
rect 14080 8246 14185 8257
rect 14219 8246 14240 8280
tri 14080 8240 14086 8246 ne
rect 14086 8240 14240 8246
tri 14086 8206 14120 8240 ne
rect 14120 8236 14240 8240
rect 14292 8236 14312 8288
rect 14364 8236 14384 8288
rect 14436 8236 14456 8288
rect 14508 8236 14528 8288
rect 14580 8236 14600 8288
rect 14652 8280 14692 8288
rect 14726 8280 14770 8314
rect 14804 8280 14848 8314
rect 14882 8280 14926 8314
rect 14960 8280 15004 8314
rect 15038 8280 15114 8314
rect 14652 8240 15114 8280
rect 14652 8236 14692 8240
rect 14120 8222 14614 8236
rect 14648 8222 14692 8236
rect 14120 8206 14240 8222
tri 14120 8202 14124 8206 ne
rect 14124 8202 14240 8206
tri 14124 8168 14158 8202 ne
rect 14158 8168 14185 8202
rect 14219 8170 14240 8202
rect 14292 8170 14312 8222
rect 14364 8170 14384 8222
rect 14436 8170 14456 8222
rect 14508 8170 14528 8222
rect 14580 8170 14600 8222
rect 14652 8206 14692 8222
rect 14726 8206 14770 8240
rect 14804 8206 14848 8240
rect 14882 8206 14926 8240
rect 14960 8206 15004 8240
rect 15038 8206 15114 8240
rect 14652 8170 15114 8206
rect 14219 8168 14257 8170
rect 14291 8168 14329 8170
rect 14363 8168 14401 8170
rect 14435 8168 14473 8170
rect 14507 8168 15114 8170
tri 14158 8166 14160 8168 ne
rect 14160 8166 15114 8168
tri 14160 8156 14170 8166 ne
rect 14170 8156 14614 8166
rect 14648 8156 14692 8166
tri 14170 8132 14194 8156 ne
rect 14194 8132 14240 8156
tri 14194 8115 14211 8132 ne
rect 14211 8115 14240 8132
tri 14211 8098 14228 8115 ne
rect 14228 8104 14240 8115
rect 14292 8104 14312 8156
rect 14364 8104 14384 8156
rect 14436 8115 14456 8156
rect 14508 8115 14528 8156
rect 14508 8104 14511 8115
rect 14580 8104 14600 8156
rect 14652 8132 14692 8156
rect 14726 8132 14770 8166
rect 14804 8132 14848 8166
rect 14882 8132 14926 8166
rect 14960 8132 15004 8166
rect 15038 8132 15114 8166
rect 14652 8104 15114 8132
rect 14228 8098 14431 8104
tri 14228 8081 14245 8098 ne
rect 14245 8081 14431 8098
rect 14465 8081 14511 8104
rect 14545 8092 15114 8104
rect 14545 8081 14614 8092
tri 14245 8058 14268 8081 ne
rect 14268 8058 14614 8081
rect 14648 8058 14692 8092
rect 14726 8058 14770 8092
rect 14804 8058 14848 8092
rect 14882 8058 14926 8092
rect 14960 8058 15004 8092
rect 15038 8058 15114 8092
tri 14268 8056 14270 8058 ne
rect 14270 8056 15114 8058
tri 14270 8033 14293 8056 ne
rect 14293 8033 15114 8056
tri 14293 7999 14327 8033 ne
rect 14327 7999 14431 8033
rect 14465 7999 14511 8033
rect 14545 8018 15114 8033
rect 14545 7999 14614 8018
tri 14327 7984 14342 7999 ne
rect 14342 7984 14614 7999
rect 14648 7984 14692 8018
rect 14726 7984 14770 8018
rect 14804 7984 14848 8018
rect 14882 7984 14926 8018
rect 14960 7984 15004 8018
rect 15038 7984 15114 8018
tri 14342 7950 14376 7984 ne
rect 14376 7950 15114 7984
tri 14376 7924 14402 7950 ne
rect 14402 7924 14431 7950
tri 14402 7916 14410 7924 ne
rect 14410 7916 14431 7924
rect 14465 7916 14511 7950
rect 14545 7944 15114 7950
rect 14545 7916 14614 7944
rect 12619 7910 12762 7916
tri 12762 7910 12768 7916 sw
tri 14410 7910 14416 7916 ne
rect 14416 7910 14614 7916
rect 14648 7910 14692 7944
rect 14726 7910 14770 7944
rect 14804 7910 14848 7944
rect 14882 7910 14926 7944
rect 14960 7910 15004 7944
rect 15038 7910 15114 7944
rect 12619 7904 12768 7910
tri 12768 7904 12774 7910 sw
tri 14416 7904 14422 7910 ne
rect 14422 7904 15114 7910
rect 12619 7885 12774 7904
tri 12774 7885 12793 7904 sw
tri 14422 7885 14441 7904 ne
rect 14441 7885 15114 7904
rect 12619 7873 12793 7885
rect 12252 7870 12793 7873
tri 12793 7870 12808 7885 sw
tri 14441 7870 14456 7885 ne
rect 14456 7870 15114 7885
tri 6611 7857 6624 7870 se
rect 6624 7857 7083 7870
tri 7083 7857 7096 7870 nw
rect 12252 7867 12808 7870
tri 12808 7867 12811 7870 sw
tri 14456 7867 14459 7870 ne
rect 14459 7867 14614 7870
tri 12563 7857 12573 7867 ne
rect 12573 7857 12811 7867
tri 12811 7857 12821 7867 sw
tri 14459 7857 14469 7867 ne
rect 14469 7857 14614 7867
rect 278 7851 7062 7857
rect 330 7836 7062 7851
tri 7062 7836 7083 7857 nw
tri 12573 7836 12594 7857 ne
rect 12594 7836 12821 7857
tri 12821 7836 12842 7857 sw
tri 14469 7836 14490 7857 ne
rect 14490 7836 14614 7857
rect 14648 7836 14692 7870
rect 14726 7836 14770 7870
rect 14804 7836 14848 7870
rect 14882 7836 14926 7870
rect 14960 7836 15004 7870
rect 15038 7836 15114 7870
rect 330 7799 7022 7836
rect 278 7796 7022 7799
tri 7022 7796 7062 7836 nw
tri 12594 7796 12634 7836 ne
rect 12634 7796 12842 7836
tri 12842 7796 12882 7836 sw
tri 14490 7796 14530 7836 ne
rect 14530 7796 15114 7836
rect 278 7785 6988 7796
rect 330 7762 6988 7785
tri 6988 7762 7022 7796 nw
tri 12634 7785 12645 7796 ne
rect 12645 7785 12882 7796
tri 12882 7785 12893 7796 sw
tri 14530 7785 14541 7796 ne
rect 14541 7785 14614 7796
tri 12645 7762 12668 7785 ne
rect 12668 7762 12893 7785
tri 12893 7762 12916 7785 sw
tri 14541 7762 14564 7785 ne
rect 14564 7762 14614 7785
rect 14648 7762 14692 7796
rect 14726 7762 14770 7796
rect 14804 7762 14848 7796
rect 14882 7762 14926 7796
rect 14960 7762 15004 7796
rect 15038 7762 15114 7796
rect 330 7733 6948 7762
rect 278 7722 6948 7733
tri 6948 7722 6988 7762 nw
tri 12668 7722 12708 7762 ne
rect 12708 7722 12916 7762
tri 12916 7722 12956 7762 sw
tri 14564 7722 14604 7762 ne
rect 14604 7722 15114 7762
rect 278 7718 6914 7722
rect 330 7688 6914 7718
tri 6914 7688 6948 7722 nw
tri 12708 7688 12742 7722 ne
rect 12742 7718 12956 7722
tri 12956 7718 12960 7722 sw
tri 14604 7718 14608 7722 ne
rect 12742 7688 12960 7718
tri 12960 7688 12990 7718 sw
rect 14608 7688 14614 7722
rect 14648 7688 14692 7722
rect 14726 7688 14770 7722
rect 14804 7688 14848 7722
rect 14882 7688 14926 7722
rect 14960 7688 15004 7722
rect 15038 7688 15114 7722
rect 330 7666 6874 7688
rect 278 7651 6874 7666
tri 25 7614 27 7616 sw
rect 25 7574 27 7614
tri 27 7574 67 7614 sw
rect 330 7648 6874 7651
tri 6874 7648 6914 7688 nw
tri 12742 7648 12782 7688 ne
rect 12782 7648 12990 7688
tri 12990 7648 13030 7688 sw
rect 14608 7648 15114 7688
rect 330 7614 6840 7648
tri 6840 7614 6874 7648 nw
tri 12782 7614 12816 7648 ne
rect 12816 7614 13030 7648
tri 13030 7614 13064 7648 sw
rect 14608 7614 14614 7648
rect 14648 7614 14692 7648
rect 14726 7614 14770 7648
rect 14804 7614 14848 7648
rect 14882 7614 14926 7648
rect 14960 7614 15004 7648
rect 15038 7614 15114 7648
rect 330 7599 6800 7614
rect 278 7584 6800 7599
rect 25 7540 67 7574
tri 67 7540 101 7574 sw
rect 25 7526 101 7540
tri 101 7526 115 7540 sw
rect 330 7574 6800 7584
tri 6800 7574 6840 7614 nw
tri 12816 7574 12856 7614 ne
rect 12856 7574 13064 7614
tri 13064 7574 13104 7614 sw
rect 14608 7574 15114 7614
rect 330 7561 6787 7574
tri 6787 7561 6800 7574 nw
tri 12856 7561 12869 7574 ne
rect 12869 7561 13104 7574
tri 13104 7561 13117 7574 sw
rect 330 7540 6766 7561
tri 6766 7540 6787 7561 nw
rect 330 7532 6752 7540
rect 278 7526 6752 7532
tri 6752 7526 6766 7540 nw
rect 25 7499 115 7526
tri 115 7499 142 7526 sw
rect 11129 7509 11135 7561
rect 11187 7509 11208 7561
rect 11260 7509 11280 7561
rect 11332 7509 11338 7561
tri 12869 7540 12890 7561 ne
rect 12890 7540 13117 7561
tri 13117 7540 13138 7561 sw
rect 14608 7540 14614 7574
rect 14648 7540 14692 7574
rect 14726 7540 14770 7574
rect 14804 7540 14848 7574
rect 14882 7540 14926 7574
rect 14960 7540 15004 7574
rect 15038 7540 15114 7574
tri 12890 7537 12893 7540 ne
rect 25 7465 142 7499
tri 142 7465 176 7499 sw
rect 11129 7481 11338 7509
rect 25 7429 176 7465
tri 176 7429 212 7465 sw
rect 11129 7429 11135 7481
rect 11187 7429 11208 7481
rect 11260 7429 11280 7481
rect 11332 7429 11338 7481
rect 12893 7499 13138 7540
tri 13138 7499 13179 7540 sw
rect 14608 7499 15114 7540
rect 12893 7465 13179 7499
tri 13179 7465 13213 7499 sw
rect 14608 7465 14614 7499
rect 14648 7465 14692 7499
rect 14726 7465 14770 7499
rect 14804 7465 14848 7499
rect 14882 7465 14926 7499
rect 14960 7465 15004 7499
rect 15038 7465 15114 7499
rect 12893 7435 13213 7465
tri 13213 7435 13243 7465 sw
rect 25 7424 212 7429
tri 212 7424 217 7429 sw
rect 25 7390 217 7424
tri 217 7390 251 7424 sw
rect 25 7381 251 7390
tri 251 7381 260 7390 sw
rect 25 7374 1405 7381
rect 25 7340 57 7374
rect 91 7340 132 7374
rect 166 7340 207 7374
rect 241 7340 282 7374
rect 316 7340 357 7374
rect 391 7340 432 7374
rect 466 7340 507 7374
rect 541 7340 582 7374
rect 616 7340 657 7374
rect 691 7340 732 7374
rect 766 7340 807 7374
rect 841 7340 882 7374
rect 916 7340 957 7374
rect 991 7340 1032 7374
rect 1066 7340 1107 7374
rect 1141 7340 1182 7374
rect 1216 7340 1256 7374
rect 1290 7340 1330 7374
rect 1364 7349 1405 7374
tri 1405 7349 1437 7381 sw
rect 1364 7340 1437 7349
rect 25 7315 1437 7340
tri 1437 7315 1471 7349 sw
rect 25 7290 1471 7315
rect 25 7256 57 7290
rect 91 7256 132 7290
rect 166 7256 207 7290
rect 241 7256 282 7290
rect 316 7256 357 7290
rect 391 7256 432 7290
rect 466 7256 507 7290
rect 541 7256 582 7290
rect 616 7256 657 7290
rect 691 7256 732 7290
rect 766 7256 807 7290
rect 841 7256 882 7290
rect 916 7256 957 7290
rect 991 7256 1032 7290
rect 1066 7256 1107 7290
rect 1141 7256 1182 7290
rect 1216 7256 1256 7290
rect 1290 7256 1330 7290
rect 1364 7274 1471 7290
tri 1471 7274 1512 7315 sw
rect 1364 7256 1512 7274
rect 25 7240 1512 7256
tri 1512 7240 1546 7274 sw
rect 25 7226 1546 7240
tri 1546 7226 1560 7240 sw
rect 25 7220 7162 7226
rect 25 7206 1431 7220
rect 25 7172 57 7206
rect 91 7172 132 7206
rect 166 7172 207 7206
rect 241 7172 282 7206
rect 316 7172 357 7206
rect 391 7172 432 7206
rect 466 7172 507 7206
rect 541 7172 582 7206
rect 616 7172 657 7206
rect 691 7172 732 7206
rect 766 7172 807 7206
rect 841 7172 882 7206
rect 916 7172 957 7206
rect 991 7172 1032 7206
rect 1066 7172 1107 7206
rect 1141 7172 1182 7206
rect 1216 7172 1256 7206
rect 1290 7172 1330 7206
rect 1364 7186 1431 7206
rect 1465 7186 1504 7220
rect 1538 7186 1577 7220
rect 1611 7186 1650 7220
rect 1684 7186 1723 7220
rect 1757 7186 1796 7220
rect 1830 7186 1869 7220
rect 1903 7186 1942 7220
rect 1976 7186 2015 7220
rect 2049 7186 2088 7220
rect 2122 7186 2161 7220
rect 2195 7186 2234 7220
rect 2268 7186 2307 7220
rect 2341 7186 2380 7220
rect 2414 7186 2453 7220
rect 2487 7186 2526 7220
rect 2560 7186 2599 7220
rect 2633 7186 2672 7220
rect 2706 7186 2745 7220
rect 2779 7186 2818 7220
rect 2852 7186 2891 7220
rect 2925 7186 2964 7220
rect 2998 7186 3037 7220
rect 3071 7186 3110 7220
rect 3144 7186 3183 7220
rect 3217 7186 3256 7220
rect 3290 7186 3329 7220
rect 3363 7186 3402 7220
rect 3436 7186 3475 7220
rect 3509 7186 3548 7220
rect 3582 7186 3621 7220
rect 3655 7186 3694 7220
rect 3728 7186 3767 7220
rect 3801 7186 3840 7220
rect 3874 7186 3913 7220
rect 3947 7186 3986 7220
rect 4020 7186 4059 7220
rect 4093 7186 4132 7220
rect 4166 7186 4205 7220
rect 4239 7186 4278 7220
rect 4312 7186 4351 7220
rect 4385 7186 4424 7220
rect 4458 7186 4497 7220
rect 4531 7186 4570 7220
rect 4604 7186 4643 7220
rect 4677 7186 4716 7220
rect 4750 7186 4789 7220
rect 4823 7186 4862 7220
rect 4896 7186 4935 7220
rect 4969 7186 5008 7220
rect 5042 7186 5081 7220
rect 5115 7186 5154 7220
rect 5188 7186 5227 7220
rect 5261 7186 5300 7220
rect 5334 7186 5373 7220
rect 5407 7186 5446 7220
rect 5480 7186 5519 7220
rect 5553 7186 5592 7220
rect 5626 7186 5665 7220
rect 5699 7186 5738 7220
rect 5772 7186 5811 7220
rect 5845 7186 5884 7220
rect 5918 7186 5957 7220
rect 5991 7186 6030 7220
rect 6064 7186 6103 7220
rect 6137 7186 6176 7220
rect 6210 7186 6249 7220
rect 6283 7186 6322 7220
rect 6356 7186 6395 7220
rect 6429 7186 6468 7220
rect 6502 7186 6540 7220
rect 6574 7186 6612 7220
rect 6646 7186 6684 7220
rect 6718 7186 6756 7220
rect 6790 7186 6828 7220
rect 6862 7186 6900 7220
rect 6934 7186 6972 7220
rect 7006 7186 7044 7220
rect 7078 7186 7116 7220
rect 7150 7186 7162 7220
rect 1364 7180 7162 7186
rect 1364 7172 1564 7180
rect 25 7165 1564 7172
tri 1564 7165 1579 7180 nw
rect 25 7125 1524 7165
tri 1524 7125 1564 7165 nw
rect 25 7124 1523 7125
tri 1523 7124 1524 7125 nw
tri 7474 7124 7475 7125 se
rect 7475 7124 7873 7125
rect 25 7122 1489 7124
rect 25 7088 57 7122
rect 91 7088 132 7122
rect 166 7088 207 7122
rect 241 7088 282 7122
rect 316 7088 357 7122
rect 391 7088 432 7122
rect 466 7088 507 7122
rect 541 7088 582 7122
rect 616 7088 657 7122
rect 691 7088 732 7122
rect 766 7088 807 7122
rect 841 7088 882 7122
rect 916 7088 957 7122
rect 991 7088 1032 7122
rect 1066 7088 1107 7122
rect 1141 7088 1182 7122
rect 1216 7088 1256 7122
rect 1290 7088 1330 7122
rect 1364 7090 1489 7122
tri 1489 7090 1523 7124 nw
tri 7440 7090 7474 7124 se
rect 7474 7090 7873 7124
rect 1364 7088 1396 7090
rect 25 7038 1396 7088
rect 25 7004 57 7038
rect 91 7004 132 7038
rect 166 7004 207 7038
rect 241 7004 282 7038
rect 316 7004 357 7038
rect 391 7004 432 7038
rect 466 7004 507 7038
rect 541 7004 582 7038
rect 616 7004 657 7038
rect 691 7004 732 7038
rect 766 7004 807 7038
rect 841 7004 882 7038
rect 916 7004 957 7038
rect 991 7004 1032 7038
rect 1066 7004 1107 7038
rect 1141 7004 1182 7038
rect 1216 7004 1256 7038
rect 1290 7004 1330 7038
rect 1364 7004 1396 7038
rect 25 6997 1396 7004
tri 1396 6997 1489 7090 nw
tri 7347 6997 7440 7090 se
rect 7440 6997 7873 7090
tri 7291 6941 7347 6997 se
rect 7347 6995 7873 6997
rect 7347 6941 7475 6995
tri 7475 6941 7529 6995 nw
tri 7230 6880 7291 6941 se
rect 7291 6880 7414 6941
tri 7414 6880 7475 6941 nw
rect 338 6874 7359 6880
rect 390 6825 7359 6874
tri 7359 6825 7414 6880 nw
rect 390 6822 7325 6825
rect 338 6808 7325 6822
rect 390 6791 7325 6808
tri 7325 6791 7359 6825 nw
rect 390 6756 7287 6791
rect 338 6753 7287 6756
tri 7287 6753 7325 6791 nw
rect 338 6750 7284 6753
tri 7284 6750 7287 6753 nw
tri 12882 6647 12893 6658 se
rect 12893 6647 13243 7435
rect 14608 7424 15114 7465
rect 14608 7390 14614 7424
rect 14648 7390 14692 7424
rect 14726 7390 14770 7424
rect 14804 7390 14848 7424
rect 14882 7390 14926 7424
rect 14960 7390 15004 7424
rect 15038 7390 15114 7424
rect 14608 7349 15114 7390
rect 14608 7315 14614 7349
rect 14648 7315 14692 7349
rect 14726 7315 14770 7349
rect 14804 7315 14848 7349
rect 14882 7315 14926 7349
rect 14960 7315 15004 7349
rect 15038 7315 15114 7349
rect 14608 7274 15114 7315
rect 14608 7240 14614 7274
rect 14648 7240 14692 7274
rect 14726 7240 14770 7274
rect 14804 7240 14848 7274
rect 14882 7240 14926 7274
rect 14960 7240 15004 7274
rect 15038 7240 15114 7274
rect 14608 7199 15114 7240
rect 14608 7165 14614 7199
rect 14648 7165 14692 7199
rect 14726 7165 14770 7199
rect 14804 7165 14848 7199
rect 14882 7165 14926 7199
rect 14960 7165 15004 7199
rect 15038 7165 15114 7199
rect 14608 7124 15114 7165
rect 14608 7090 14614 7124
rect 14648 7090 14692 7124
rect 14726 7090 14770 7124
rect 14804 7090 14848 7124
rect 14882 7090 14926 7124
rect 14960 7090 15004 7124
rect 15038 7090 15114 7124
rect 14608 7053 15114 7090
rect 15062 6825 15108 6837
rect 15062 6791 15068 6825
rect 15102 6791 15108 6825
rect 15062 6753 15108 6791
rect 15062 6719 15068 6753
rect 15102 6719 15108 6753
rect 15062 6681 15108 6719
tri 13243 6647 13254 6658 sw
rect 15062 6647 15068 6681
rect 15102 6647 15108 6681
tri 12844 6609 12882 6647 se
rect 12882 6609 13254 6647
tri 13254 6609 13292 6647 sw
rect 15062 6609 15108 6647
tri 12810 6575 12844 6609 se
rect 12844 6575 13292 6609
tri 13292 6575 13326 6609 sw
rect 15062 6575 15068 6609
rect 15102 6575 15108 6609
tri 12772 6537 12810 6575 se
rect 12810 6537 13326 6575
tri 13326 6537 13364 6575 sw
rect 15062 6537 15108 6575
tri 12738 6503 12772 6537 se
rect 12772 6503 13364 6537
tri 13364 6503 13398 6537 sw
rect 15062 6503 15068 6537
rect 15102 6503 15108 6537
tri 12700 6465 12738 6503 se
rect 12738 6465 13398 6503
tri 13398 6465 13436 6503 sw
rect 15062 6465 15108 6503
tri 12685 6450 12700 6465 se
rect 12700 6450 13436 6465
tri 13436 6450 13451 6465 sw
rect 15062 6450 15068 6465
rect 56 6439 15068 6450
rect 56 6405 68 6439
rect 102 6405 141 6439
rect 175 6405 214 6439
rect 248 6405 287 6439
rect 321 6405 360 6439
rect 394 6405 433 6439
rect 467 6405 506 6439
rect 540 6405 579 6439
rect 613 6405 652 6439
rect 686 6405 725 6439
rect 759 6405 798 6439
rect 832 6405 871 6439
rect 905 6405 944 6439
rect 978 6405 1017 6439
rect 1051 6405 1090 6439
rect 56 6367 1090 6405
rect 56 6333 68 6367
rect 102 6333 141 6367
rect 175 6333 214 6367
rect 248 6333 287 6367
rect 321 6333 360 6367
rect 394 6333 433 6367
rect 467 6333 506 6367
rect 540 6333 579 6367
rect 613 6333 652 6367
rect 686 6333 725 6367
rect 759 6333 798 6367
rect 832 6333 871 6367
rect 905 6333 944 6367
rect 978 6333 1017 6367
rect 1051 6333 1090 6367
rect 56 6295 1090 6333
rect 56 6261 68 6295
rect 102 6261 141 6295
rect 175 6261 214 6295
rect 248 6261 287 6295
rect 321 6261 360 6295
rect 394 6261 433 6295
rect 467 6261 506 6295
rect 540 6261 579 6295
rect 613 6261 652 6295
rect 686 6261 725 6295
rect 759 6261 798 6295
rect 832 6261 871 6295
rect 905 6261 944 6295
rect 978 6261 1017 6295
rect 1051 6261 1090 6295
rect 56 6223 1090 6261
rect 56 6189 68 6223
rect 102 6189 141 6223
rect 175 6189 214 6223
rect 248 6189 287 6223
rect 321 6189 360 6223
rect 394 6189 433 6223
rect 467 6189 506 6223
rect 540 6189 579 6223
rect 613 6189 652 6223
rect 686 6189 725 6223
rect 759 6189 798 6223
rect 832 6189 871 6223
rect 905 6189 944 6223
rect 978 6189 1017 6223
rect 1051 6189 1090 6223
rect 56 6151 1090 6189
rect 56 6117 68 6151
rect 102 6117 141 6151
rect 175 6117 214 6151
rect 248 6117 287 6151
rect 321 6117 360 6151
rect 394 6117 433 6151
rect 467 6117 506 6151
rect 540 6117 579 6151
rect 613 6117 652 6151
rect 686 6117 725 6151
rect 759 6117 798 6151
rect 832 6117 871 6151
rect 905 6117 944 6151
rect 978 6117 1017 6151
rect 1051 6117 1090 6151
rect 15020 6431 15068 6439
rect 15102 6450 15108 6465
rect 15102 6431 15114 6450
rect 15020 6393 15114 6431
rect 15020 6359 15068 6393
rect 15102 6359 15114 6393
rect 15020 6321 15114 6359
rect 15020 6287 15068 6321
rect 15102 6287 15114 6321
rect 15020 6249 15114 6287
rect 15020 6215 15068 6249
rect 15102 6215 15114 6249
rect 15020 6177 15114 6215
rect 15020 6143 15068 6177
rect 15102 6143 15114 6177
rect 15020 6117 15114 6143
rect 56 6105 15114 6117
rect 56 6086 15068 6105
rect 14974 6071 15068 6086
rect 15102 6071 15114 6105
rect 14974 6033 15114 6071
rect 14974 5999 15068 6033
rect 15102 5999 15114 6033
rect 14974 5961 15114 5999
rect 14974 5927 15068 5961
rect 15102 5927 15114 5961
rect 14974 5889 15114 5927
rect 14974 5855 15068 5889
rect 15102 5855 15114 5889
rect 14974 5817 15114 5855
rect 14974 5783 15068 5817
rect 15102 5783 15114 5817
rect 14974 5745 15114 5783
rect 14974 5711 15068 5745
rect 15102 5711 15114 5745
rect 14974 5673 15114 5711
rect 14974 5639 15068 5673
rect 15102 5639 15114 5673
rect 14974 5601 15114 5639
rect 510 5568 809 5586
rect 510 5516 516 5568
rect 568 5516 634 5568
rect 686 5516 751 5568
rect 803 5516 809 5568
rect 510 5498 809 5516
rect 14249 5565 14371 5583
rect 14249 5513 14313 5565
rect 14365 5513 14371 5565
rect 14249 5495 14371 5513
rect 14974 5567 15068 5601
rect 15102 5567 15114 5601
rect 14974 5529 15114 5567
rect 14974 5495 15068 5529
rect 15102 5495 15114 5529
rect 435 5465 703 5471
rect 487 5413 507 5465
rect 559 5413 579 5465
rect 631 5413 651 5465
rect 742 5427 748 5479
rect 800 5427 811 5479
rect 14241 5465 14495 5471
rect 435 5400 703 5413
rect 487 5348 507 5400
rect 559 5348 579 5400
rect 631 5348 651 5400
rect 435 5335 703 5348
rect 487 5283 507 5335
rect 559 5283 579 5335
rect 631 5283 651 5335
rect 435 5270 703 5283
rect 487 5218 507 5270
rect 559 5218 579 5270
rect 631 5218 651 5270
rect 435 5205 703 5218
rect 487 5153 507 5205
rect 559 5153 579 5205
rect 631 5153 651 5205
rect 435 5140 703 5153
rect 487 5088 507 5140
rect 559 5088 579 5140
rect 631 5088 651 5140
rect 435 5075 703 5088
rect 487 5023 507 5075
rect 559 5023 579 5075
rect 631 5023 651 5075
rect 435 5010 703 5023
rect 487 4958 507 5010
rect 559 4958 579 5010
rect 631 4958 651 5010
rect 435 4945 703 4958
rect 487 4893 507 4945
rect 559 4893 579 4945
rect 631 4893 651 4945
rect 435 4880 703 4893
rect 487 4828 507 4880
rect 559 4828 579 4880
rect 631 4828 651 4880
rect 435 4815 703 4828
rect 487 4763 507 4815
rect 559 4763 579 4815
rect 631 4763 651 4815
rect 435 4750 703 4763
rect 487 4698 507 4750
rect 559 4698 579 4750
rect 631 4698 651 4750
rect 435 4685 703 4698
rect 487 4633 507 4685
rect 559 4633 579 4685
rect 631 4633 651 4685
rect 435 4620 703 4633
rect 487 4568 507 4620
rect 559 4568 579 4620
rect 631 4568 651 4620
rect 435 4555 703 4568
rect 487 4503 507 4555
rect 559 4503 579 4555
rect 631 4503 651 4555
rect 435 4490 703 4503
rect 487 4438 507 4490
rect 559 4438 579 4490
rect 631 4438 651 4490
rect 435 4425 703 4438
rect 487 4373 507 4425
rect 559 4373 579 4425
rect 631 4373 651 4425
rect 435 4360 703 4373
rect 487 4308 507 4360
rect 559 4308 579 4360
rect 631 4308 651 4360
rect 435 4295 703 4308
rect 487 4243 507 4295
rect 559 4243 579 4295
rect 631 4243 651 4295
rect 435 4230 703 4243
rect 487 4178 507 4230
rect 559 4178 579 4230
rect 631 4178 651 4230
rect 435 4165 703 4178
rect 487 4113 507 4165
rect 559 4113 579 4165
rect 631 4113 651 4165
rect 435 4099 703 4113
rect 487 4047 507 4099
rect 559 4047 579 4099
rect 631 4047 651 4099
rect 435 4033 703 4047
rect 487 3981 507 4033
rect 559 3981 579 4033
rect 631 3981 651 4033
rect 435 3967 703 3981
rect 487 3915 507 3967
rect 559 3915 579 3967
rect 631 3915 651 3967
rect 435 3901 703 3915
rect 487 3849 507 3901
rect 559 3849 579 3901
rect 631 3849 651 3901
rect 435 3835 703 3849
rect 487 3783 507 3835
rect 559 3783 579 3835
rect 631 3783 651 3835
rect 435 3769 703 3783
rect 487 3717 507 3769
rect 559 3717 579 3769
rect 631 3717 651 3769
rect 435 3703 703 3717
rect 487 3651 507 3703
rect 559 3651 579 3703
rect 631 3651 651 3703
rect 435 1923 703 3651
rect 14241 5413 14243 5465
rect 14295 5413 14309 5465
rect 14361 5413 14375 5465
rect 14427 5413 14441 5465
rect 14493 5413 14495 5465
rect 14241 5400 14495 5413
rect 14241 5348 14243 5400
rect 14295 5348 14309 5400
rect 14361 5348 14375 5400
rect 14427 5348 14441 5400
rect 14493 5348 14495 5400
rect 14241 5335 14495 5348
rect 14241 5283 14243 5335
rect 14295 5283 14309 5335
rect 14361 5283 14375 5335
rect 14427 5283 14441 5335
rect 14493 5283 14495 5335
rect 14241 5270 14495 5283
rect 14241 5218 14243 5270
rect 14295 5218 14309 5270
rect 14361 5218 14375 5270
rect 14427 5218 14441 5270
rect 14493 5218 14495 5270
rect 14241 5205 14495 5218
rect 14241 5153 14243 5205
rect 14295 5153 14309 5205
rect 14361 5153 14375 5205
rect 14427 5153 14441 5205
rect 14493 5153 14495 5205
rect 14241 5140 14495 5153
rect 14241 5088 14243 5140
rect 14295 5088 14309 5140
rect 14361 5088 14375 5140
rect 14427 5088 14441 5140
rect 14493 5088 14495 5140
rect 14241 5075 14495 5088
rect 14241 5023 14243 5075
rect 14295 5023 14309 5075
rect 14361 5023 14375 5075
rect 14427 5023 14441 5075
rect 14493 5023 14495 5075
rect 14241 5010 14495 5023
rect 14241 4958 14243 5010
rect 14295 4958 14309 5010
rect 14361 4958 14375 5010
rect 14427 4958 14441 5010
rect 14493 4958 14495 5010
rect 14241 4945 14495 4958
rect 14241 4893 14243 4945
rect 14295 4893 14309 4945
rect 14361 4893 14375 4945
rect 14427 4893 14441 4945
rect 14493 4893 14495 4945
rect 14241 4880 14495 4893
rect 14241 4828 14243 4880
rect 14295 4828 14309 4880
rect 14361 4828 14375 4880
rect 14427 4828 14441 4880
rect 14493 4828 14495 4880
rect 14241 4815 14495 4828
rect 14241 4763 14243 4815
rect 14295 4763 14309 4815
rect 14361 4763 14375 4815
rect 14427 4763 14441 4815
rect 14493 4763 14495 4815
rect 14241 4750 14495 4763
rect 14241 4698 14243 4750
rect 14295 4698 14309 4750
rect 14361 4698 14375 4750
rect 14427 4698 14441 4750
rect 14493 4698 14495 4750
rect 14241 4685 14495 4698
rect 14241 4633 14243 4685
rect 14295 4633 14309 4685
rect 14361 4633 14375 4685
rect 14427 4633 14441 4685
rect 14493 4633 14495 4685
rect 14241 4620 14495 4633
rect 14241 4568 14243 4620
rect 14295 4568 14309 4620
rect 14361 4568 14375 4620
rect 14427 4568 14441 4620
rect 14493 4568 14495 4620
rect 14241 4555 14495 4568
rect 14241 4503 14243 4555
rect 14295 4503 14309 4555
rect 14361 4503 14375 4555
rect 14427 4503 14441 4555
rect 14493 4503 14495 4555
rect 14241 4490 14495 4503
rect 14241 4438 14243 4490
rect 14295 4438 14309 4490
rect 14361 4438 14375 4490
rect 14427 4438 14441 4490
rect 14493 4438 14495 4490
rect 14241 4425 14495 4438
rect 14241 4373 14243 4425
rect 14295 4373 14309 4425
rect 14361 4373 14375 4425
rect 14427 4373 14441 4425
rect 14493 4373 14495 4425
rect 14241 4359 14495 4373
rect 14241 4307 14243 4359
rect 14295 4307 14309 4359
rect 14361 4307 14375 4359
rect 14427 4307 14441 4359
rect 14493 4307 14495 4359
rect 14241 4293 14495 4307
rect 14241 4241 14243 4293
rect 14295 4241 14309 4293
rect 14361 4241 14375 4293
rect 14427 4241 14441 4293
rect 14493 4241 14495 4293
rect 14241 4227 14495 4241
rect 14241 4175 14243 4227
rect 14295 4175 14309 4227
rect 14361 4175 14375 4227
rect 14427 4175 14441 4227
rect 14493 4175 14495 4227
rect 14241 4161 14495 4175
rect 14241 4109 14243 4161
rect 14295 4109 14309 4161
rect 14361 4109 14375 4161
rect 14427 4109 14441 4161
rect 14493 4109 14495 4161
rect 14241 4095 14495 4109
rect 14241 4043 14243 4095
rect 14295 4043 14309 4095
rect 14361 4043 14375 4095
rect 14427 4043 14441 4095
rect 14493 4043 14495 4095
rect 14241 4029 14495 4043
rect 14241 3977 14243 4029
rect 14295 3977 14309 4029
rect 14361 3977 14375 4029
rect 14427 3977 14441 4029
rect 14493 3977 14495 4029
rect 14241 3963 14495 3977
rect 14241 3911 14243 3963
rect 14295 3911 14309 3963
rect 14361 3911 14375 3963
rect 14427 3911 14441 3963
rect 14493 3911 14495 3963
rect 14241 3897 14495 3911
rect 14241 3845 14243 3897
rect 14295 3845 14309 3897
rect 14361 3845 14375 3897
rect 14427 3845 14441 3897
rect 14493 3845 14495 3897
rect 14241 3831 14495 3845
rect 14241 3779 14243 3831
rect 14295 3779 14309 3831
rect 14361 3779 14375 3831
rect 14427 3779 14441 3831
rect 14493 3779 14495 3831
rect 14241 3765 14495 3779
rect 14241 3713 14243 3765
rect 14295 3713 14309 3765
rect 14361 3713 14375 3765
rect 14427 3713 14441 3765
rect 14493 3713 14495 3765
rect 14241 3699 14495 3713
rect 14241 3647 14243 3699
rect 14295 3647 14309 3699
rect 14361 3647 14375 3699
rect 14427 3647 14441 3699
rect 14493 3647 14495 3699
rect 14241 3641 14495 3647
rect 14974 5457 15114 5495
rect 14974 5423 15068 5457
rect 15102 5423 15114 5457
rect 14974 5385 15114 5423
rect 14974 5351 15068 5385
rect 15102 5351 15114 5385
rect 14974 5313 15114 5351
rect 14974 5279 15068 5313
rect 15102 5279 15114 5313
rect 14974 5241 15114 5279
rect 14974 5207 15068 5241
rect 15102 5207 15114 5241
rect 14974 5169 15114 5207
rect 14974 5135 15068 5169
rect 15102 5135 15114 5169
rect 14974 5097 15114 5135
rect 14974 5063 15068 5097
rect 15102 5063 15114 5097
rect 14974 5025 15114 5063
rect 14974 4991 15068 5025
rect 15102 4991 15114 5025
rect 14974 4953 15114 4991
rect 14974 4919 15068 4953
rect 15102 4919 15114 4953
rect 14974 4881 15114 4919
rect 14974 4847 15068 4881
rect 15102 4847 15114 4881
rect 14974 4809 15114 4847
rect 14974 4775 15068 4809
rect 15102 4775 15114 4809
rect 14974 4737 15114 4775
rect 14974 4703 15068 4737
rect 15102 4703 15114 4737
rect 14974 4665 15114 4703
rect 14974 4631 15068 4665
rect 15102 4631 15114 4665
rect 14974 4593 15114 4631
rect 14974 4559 15068 4593
rect 15102 4559 15114 4593
rect 14974 4521 15114 4559
rect 14974 4487 15068 4521
rect 15102 4487 15114 4521
rect 14974 4449 15114 4487
rect 14974 4415 15068 4449
rect 15102 4415 15114 4449
rect 14974 4377 15114 4415
rect 14974 4343 15068 4377
rect 15102 4343 15114 4377
rect 14974 4305 15114 4343
rect 14974 4271 15068 4305
rect 15102 4271 15114 4305
rect 14974 4233 15114 4271
rect 14974 4199 15068 4233
rect 15102 4199 15114 4233
rect 14974 4161 15114 4199
rect 14974 4127 15068 4161
rect 15102 4127 15114 4161
rect 14974 4089 15114 4127
rect 14974 4055 15068 4089
rect 15102 4055 15114 4089
rect 14974 4017 15114 4055
rect 14974 3983 15068 4017
rect 15102 3983 15114 4017
rect 14974 3945 15114 3983
rect 14974 3911 15068 3945
rect 15102 3911 15114 3945
rect 14974 3873 15114 3911
rect 14974 3839 15068 3873
rect 15102 3839 15114 3873
rect 14974 3801 15114 3839
rect 14974 3767 15068 3801
rect 15102 3767 15114 3801
rect 14974 3729 15114 3767
rect 14974 3695 15068 3729
rect 15102 3695 15114 3729
rect 14974 3657 15114 3695
rect 14974 3623 15068 3657
rect 15102 3623 15114 3657
rect 14974 3585 15114 3623
rect 14974 3551 15068 3585
rect 15102 3551 15114 3585
rect 14974 3513 15114 3551
rect 14974 3479 15068 3513
rect 15102 3479 15114 3513
rect 14974 3441 15114 3479
rect 14974 3407 15068 3441
rect 15102 3407 15114 3441
rect 14974 3369 15114 3407
rect 14974 3335 15068 3369
rect 15102 3335 15114 3369
rect 14974 3297 15114 3335
rect 14974 3263 15068 3297
rect 15102 3263 15114 3297
rect 14974 3225 15114 3263
rect 14974 3191 15068 3225
rect 15102 3191 15114 3225
rect 14974 3153 15114 3191
rect 14974 3119 15068 3153
rect 15102 3119 15114 3153
rect 14974 3081 15114 3119
rect 14974 3047 15068 3081
rect 15102 3047 15114 3081
rect 14974 3009 15114 3047
rect 14974 2975 15068 3009
rect 15102 2975 15114 3009
rect 14974 2937 15114 2975
rect 14974 2903 15068 2937
rect 15102 2903 15114 2937
rect 14974 2865 15114 2903
rect 14974 2831 15068 2865
rect 15102 2831 15114 2865
rect 14974 2793 15114 2831
rect 14974 2759 15068 2793
rect 15102 2759 15114 2793
rect 14974 2721 15114 2759
rect 14974 2687 15068 2721
rect 15102 2687 15114 2721
rect 14974 2649 15114 2687
rect 14974 2615 15068 2649
rect 15102 2615 15114 2649
rect 14974 2577 15114 2615
rect 14974 2543 15068 2577
rect 15102 2543 15114 2577
rect 14974 2505 15114 2543
rect 14974 2471 15068 2505
rect 15102 2471 15114 2505
rect 14974 2433 15114 2471
rect 14974 2399 15068 2433
rect 15102 2399 15114 2433
rect 14974 2361 15114 2399
rect 14974 2327 15068 2361
rect 15102 2327 15114 2361
rect 14974 2289 15114 2327
rect 14974 2255 15068 2289
rect 15102 2255 15114 2289
rect 14974 2217 15114 2255
rect 14974 2183 15068 2217
rect 15102 2183 15114 2217
rect 14974 2145 15114 2183
rect 14974 2111 15068 2145
rect 15102 2111 15114 2145
rect 14974 2073 15114 2111
rect 14974 2039 15068 2073
rect 15102 2039 15114 2073
rect 14974 2001 15114 2039
rect 14974 1967 15068 2001
rect 15102 1967 15114 2001
rect 14974 1929 15114 1967
rect 14974 1895 15068 1929
rect 15102 1895 15114 1929
rect 14974 1857 15114 1895
rect 14974 1823 15068 1857
rect 15102 1823 15114 1857
rect 14974 1785 15114 1823
rect 14974 1751 15068 1785
rect 15102 1751 15114 1785
rect 14974 1713 15114 1751
rect 14974 1679 15068 1713
rect 15102 1679 15114 1713
rect 14974 1641 15114 1679
rect 14974 1607 15068 1641
rect 15102 1607 15114 1641
rect 14974 1569 15114 1607
rect 14974 1535 15068 1569
rect 15102 1535 15114 1569
rect 14974 1497 15114 1535
rect 14974 1463 15068 1497
rect 15102 1463 15114 1497
rect 14974 1425 15114 1463
rect 14974 1391 15068 1425
rect 15102 1391 15114 1425
rect 14974 1353 15114 1391
rect 14974 1319 15068 1353
rect 15102 1319 15114 1353
rect 14974 1300 15114 1319
rect 7031 1281 15114 1300
rect 7031 1247 15068 1281
rect 15102 1247 15114 1281
rect 7031 1217 15114 1247
rect 7031 1183 7069 1217
rect 7103 1183 7142 1217
rect 7176 1183 7215 1217
rect 7249 1183 7288 1217
rect 7322 1183 7361 1217
rect 7395 1183 7434 1217
rect 7468 1183 7507 1217
rect 7541 1183 7580 1217
rect 7614 1183 7653 1217
rect 7687 1183 7726 1217
rect 7760 1183 7799 1217
rect 7833 1183 7872 1217
rect 7906 1183 7945 1217
rect 7979 1183 8018 1217
rect 8052 1183 8091 1217
rect 8125 1183 8164 1217
rect 8198 1183 8237 1217
rect 8271 1183 8310 1217
rect 8344 1183 8383 1217
rect 8417 1183 8456 1217
rect 8490 1183 8528 1217
rect 8562 1183 8600 1217
rect 8634 1183 8672 1217
rect 8706 1183 8744 1217
rect 8778 1183 8816 1217
rect 8850 1183 8888 1217
rect 8922 1183 8960 1217
rect 8994 1183 9032 1217
rect 9066 1183 9104 1217
rect 9138 1183 9176 1217
rect 9210 1183 9248 1217
rect 9282 1183 9320 1217
rect 9354 1183 9392 1217
rect 9426 1183 9464 1217
rect 9498 1183 9536 1217
rect 9570 1183 9608 1217
rect 9642 1183 9680 1217
rect 9714 1183 9752 1217
rect 9786 1183 9824 1217
rect 9858 1183 9896 1217
rect 9930 1183 9968 1217
rect 10002 1183 10040 1217
rect 10074 1183 10112 1217
rect 10146 1183 10184 1217
rect 10218 1183 10256 1217
rect 10290 1183 10328 1217
rect 10362 1183 10400 1217
rect 10434 1183 10472 1217
rect 10506 1183 10544 1217
rect 10578 1183 10616 1217
rect 10650 1183 10688 1217
rect 10722 1183 10760 1217
rect 10794 1183 10832 1217
rect 10866 1183 10904 1217
rect 10938 1183 10976 1217
rect 11010 1183 11048 1217
rect 11082 1183 11120 1217
rect 11154 1183 11192 1217
rect 11226 1183 11264 1217
rect 11298 1183 11336 1217
rect 11370 1183 11408 1217
rect 11442 1183 11480 1217
rect 11514 1183 11552 1217
rect 11586 1183 11624 1217
rect 11658 1183 11696 1217
rect 11730 1183 11768 1217
rect 11802 1183 11840 1217
rect 11874 1183 11912 1217
rect 11946 1183 11984 1217
rect 12018 1183 12056 1217
rect 12090 1183 12139 1217
rect 12173 1183 12212 1217
rect 12246 1183 12285 1217
rect 12319 1183 12358 1217
rect 12392 1183 12431 1217
rect 12465 1183 12504 1217
rect 12538 1183 12577 1217
rect 12611 1183 12650 1217
rect 12684 1183 12723 1217
rect 12757 1183 12796 1217
rect 12830 1183 12869 1217
rect 12903 1183 12942 1217
rect 12976 1183 13015 1217
rect 13049 1183 13088 1217
rect 13122 1183 13161 1217
rect 13195 1183 13234 1217
rect 13268 1183 13307 1217
rect 13341 1183 13380 1217
rect 13414 1183 13452 1217
rect 13486 1183 13524 1217
rect 13558 1183 13596 1217
rect 13630 1183 13668 1217
rect 13702 1183 13740 1217
rect 13774 1183 13812 1217
rect 13846 1183 13884 1217
rect 13918 1183 13956 1217
rect 13990 1183 14028 1217
rect 14062 1183 14100 1217
rect 14134 1183 14172 1217
rect 14206 1183 14244 1217
rect 14278 1183 14316 1217
rect 14350 1183 14388 1217
rect 14422 1183 14460 1217
rect 14494 1183 14532 1217
rect 14566 1183 14604 1217
rect 14638 1183 14676 1217
rect 14710 1183 14748 1217
rect 14782 1183 14820 1217
rect 14854 1183 14892 1217
rect 14926 1183 14964 1217
rect 14998 1209 15114 1217
rect 14998 1183 15068 1209
rect 7031 1175 15068 1183
rect 15102 1175 15114 1209
rect 7031 1139 15114 1175
rect 7031 1105 7069 1139
rect 7103 1105 7142 1139
rect 7176 1105 7215 1139
rect 7249 1105 7288 1139
rect 7322 1105 7361 1139
rect 7395 1105 7434 1139
rect 7468 1105 7507 1139
rect 7541 1105 7580 1139
rect 7614 1105 7653 1139
rect 7687 1105 7726 1139
rect 7760 1105 7799 1139
rect 7833 1105 7872 1139
rect 7906 1105 7945 1139
rect 7979 1105 8018 1139
rect 8052 1105 8091 1139
rect 8125 1105 8164 1139
rect 8198 1105 8237 1139
rect 8271 1105 8310 1139
rect 8344 1105 8383 1139
rect 8417 1105 8456 1139
rect 8490 1105 8528 1139
rect 8562 1105 8600 1139
rect 8634 1105 8672 1139
rect 8706 1105 8744 1139
rect 8778 1105 8816 1139
rect 8850 1105 8888 1139
rect 8922 1105 8960 1139
rect 8994 1105 9032 1139
rect 9066 1105 9104 1139
rect 9138 1105 9176 1139
rect 9210 1105 9248 1139
rect 9282 1105 9320 1139
rect 9354 1105 9392 1139
rect 9426 1105 9464 1139
rect 9498 1105 9536 1139
rect 9570 1105 9608 1139
rect 9642 1105 9680 1139
rect 9714 1105 9752 1139
rect 9786 1105 9824 1139
rect 9858 1105 9896 1139
rect 9930 1105 9968 1139
rect 10002 1105 10040 1139
rect 10074 1105 10112 1139
rect 10146 1105 10184 1139
rect 10218 1105 10256 1139
rect 10290 1105 10328 1139
rect 10362 1105 10400 1139
rect 10434 1105 10472 1139
rect 10506 1105 10544 1139
rect 10578 1105 10616 1139
rect 10650 1105 10688 1139
rect 10722 1105 10760 1139
rect 10794 1105 10832 1139
rect 10866 1105 10904 1139
rect 10938 1105 10976 1139
rect 11010 1105 11048 1139
rect 11082 1105 11120 1139
rect 11154 1105 11192 1139
rect 11226 1105 11264 1139
rect 11298 1105 11336 1139
rect 11370 1105 11408 1139
rect 11442 1105 11480 1139
rect 11514 1105 11552 1139
rect 11586 1105 11624 1139
rect 11658 1105 11696 1139
rect 11730 1105 11768 1139
rect 11802 1105 11840 1139
rect 11874 1105 11912 1139
rect 11946 1105 11984 1139
rect 12018 1105 12056 1139
rect 12090 1105 12139 1139
rect 12173 1105 12212 1139
rect 12246 1105 12285 1139
rect 12319 1105 12358 1139
rect 12392 1105 12431 1139
rect 12465 1105 12504 1139
rect 12538 1105 12577 1139
rect 12611 1105 12650 1139
rect 12684 1105 12723 1139
rect 12757 1105 12796 1139
rect 12830 1105 12869 1139
rect 12903 1105 12942 1139
rect 12976 1105 13015 1139
rect 13049 1105 13088 1139
rect 13122 1105 13161 1139
rect 13195 1105 13234 1139
rect 13268 1105 13307 1139
rect 13341 1105 13380 1139
rect 13414 1105 13452 1139
rect 13486 1105 13524 1139
rect 13558 1105 13596 1139
rect 13630 1105 13668 1139
rect 13702 1105 13740 1139
rect 13774 1105 13812 1139
rect 13846 1105 13884 1139
rect 13918 1105 13956 1139
rect 13990 1105 14028 1139
rect 14062 1105 14100 1139
rect 14134 1105 14172 1139
rect 14206 1105 14244 1139
rect 14278 1105 14316 1139
rect 14350 1105 14388 1139
rect 14422 1105 14460 1139
rect 14494 1105 14532 1139
rect 14566 1105 14604 1139
rect 14638 1105 14676 1139
rect 14710 1105 14748 1139
rect 14782 1105 14820 1139
rect 14854 1105 14892 1139
rect 14926 1105 14964 1139
rect 14998 1137 15114 1139
rect 14998 1105 15068 1137
rect 7031 1103 15068 1105
rect 15102 1103 15114 1137
rect 451 932 1620 1077
rect 7031 1065 15114 1103
rect 7031 1061 15068 1065
rect 7031 1027 7069 1061
rect 7103 1027 7142 1061
rect 7176 1027 7215 1061
rect 7249 1027 7288 1061
rect 7322 1027 7361 1061
rect 7395 1027 7434 1061
rect 7468 1027 7507 1061
rect 7541 1027 7580 1061
rect 7614 1027 7653 1061
rect 7687 1027 7726 1061
rect 7760 1027 7799 1061
rect 7833 1027 7872 1061
rect 7906 1027 7945 1061
rect 7979 1027 8018 1061
rect 8052 1027 8091 1061
rect 8125 1027 8164 1061
rect 8198 1027 8237 1061
rect 8271 1027 8310 1061
rect 8344 1027 8383 1061
rect 8417 1027 8456 1061
rect 8490 1027 8528 1061
rect 8562 1027 8600 1061
rect 8634 1027 8672 1061
rect 8706 1027 8744 1061
rect 8778 1027 8816 1061
rect 8850 1027 8888 1061
rect 8922 1027 8960 1061
rect 8994 1027 9032 1061
rect 9066 1027 9104 1061
rect 9138 1027 9176 1061
rect 9210 1027 9248 1061
rect 9282 1027 9320 1061
rect 9354 1027 9392 1061
rect 9426 1027 9464 1061
rect 9498 1027 9536 1061
rect 9570 1027 9608 1061
rect 9642 1027 9680 1061
rect 9714 1027 9752 1061
rect 9786 1027 9824 1061
rect 9858 1027 9896 1061
rect 9930 1027 9968 1061
rect 10002 1027 10040 1061
rect 10074 1027 10112 1061
rect 10146 1027 10184 1061
rect 10218 1027 10256 1061
rect 10290 1027 10328 1061
rect 10362 1027 10400 1061
rect 10434 1027 10472 1061
rect 10506 1027 10544 1061
rect 10578 1027 10616 1061
rect 10650 1027 10688 1061
rect 10722 1027 10760 1061
rect 10794 1027 10832 1061
rect 10866 1027 10904 1061
rect 10938 1027 10976 1061
rect 11010 1027 11048 1061
rect 11082 1027 11120 1061
rect 11154 1027 11192 1061
rect 11226 1027 11264 1061
rect 11298 1027 11336 1061
rect 11370 1027 11408 1061
rect 11442 1027 11480 1061
rect 11514 1027 11552 1061
rect 11586 1027 11624 1061
rect 11658 1027 11696 1061
rect 11730 1027 11768 1061
rect 11802 1027 11840 1061
rect 11874 1027 11912 1061
rect 11946 1027 11984 1061
rect 12018 1027 12056 1061
rect 12090 1027 12139 1061
rect 12173 1027 12212 1061
rect 12246 1027 12285 1061
rect 12319 1027 12358 1061
rect 12392 1027 12431 1061
rect 12465 1027 12504 1061
rect 12538 1027 12577 1061
rect 12611 1027 12650 1061
rect 12684 1027 12723 1061
rect 12757 1027 12796 1061
rect 12830 1027 12869 1061
rect 12903 1027 12942 1061
rect 12976 1027 13015 1061
rect 13049 1027 13088 1061
rect 13122 1027 13161 1061
rect 13195 1027 13234 1061
rect 13268 1027 13307 1061
rect 13341 1027 13380 1061
rect 13414 1027 13452 1061
rect 13486 1027 13524 1061
rect 13558 1027 13596 1061
rect 13630 1027 13668 1061
rect 13702 1027 13740 1061
rect 13774 1027 13812 1061
rect 13846 1027 13884 1061
rect 13918 1027 13956 1061
rect 13990 1027 14028 1061
rect 14062 1027 14100 1061
rect 14134 1027 14172 1061
rect 14206 1027 14244 1061
rect 14278 1027 14316 1061
rect 14350 1027 14388 1061
rect 14422 1027 14460 1061
rect 14494 1027 14532 1061
rect 14566 1027 14604 1061
rect 14638 1027 14676 1061
rect 14710 1027 14748 1061
rect 14782 1027 14820 1061
rect 14854 1027 14892 1061
rect 14926 1027 14964 1061
rect 14998 1031 15068 1061
rect 15102 1031 15114 1065
rect 14998 1027 15114 1031
rect 7031 1020 15114 1027
rect 7034 993 7295 1020
tri 7295 993 7322 1020 nw
tri 14305 993 14332 1020 ne
rect 14332 993 15114 1020
rect 7034 989 7291 993
tri 7291 989 7295 993 nw
tri 14332 989 14336 993 ne
rect 14336 989 15068 993
rect 7034 966 7268 989
tri 7268 966 7291 989 nw
tri 14336 966 14359 989 ne
rect 14359 966 14576 989
rect 7034 955 7257 966
tri 7257 955 7268 966 nw
tri 14359 955 14370 966 ne
rect 14370 955 14576 966
rect 14610 955 14654 989
rect 14688 955 14732 989
rect 14766 955 14810 989
rect 14844 955 14888 989
rect 14922 955 14966 989
rect 15000 959 15068 989
rect 15102 959 15114 993
rect 15000 955 15114 959
rect 3948 909 5117 955
rect 7034 930 7232 955
tri 7232 930 7257 955 nw
tri 14370 930 14395 955 ne
rect 14395 930 15114 955
rect 7034 923 7225 930
tri 7225 923 7232 930 nw
rect 9784 923 11347 930
rect 7034 918 7191 923
rect 7034 884 7104 918
rect 7138 889 7191 918
tri 7191 889 7225 923 nw
rect 9784 889 9796 923
rect 9830 889 9872 923
rect 9906 889 9948 923
rect 9982 889 10024 923
rect 10058 889 10100 923
rect 10134 889 10176 923
rect 10210 889 10251 923
rect 10285 889 10326 923
rect 10360 889 10401 923
rect 10435 889 10476 923
rect 10510 889 10551 923
rect 10585 889 10626 923
rect 10660 889 10701 923
rect 10735 889 10776 923
rect 10810 889 10851 923
rect 10885 889 10926 923
rect 10960 889 11001 923
rect 11035 889 11076 923
rect 11110 889 11151 923
rect 11185 889 11226 923
rect 11260 889 11301 923
rect 11335 889 11347 923
tri 14395 921 14404 930 ne
rect 14404 921 15114 930
tri 14404 916 14409 921 ne
rect 14409 916 15068 921
rect 7138 884 7184 889
rect 7034 882 7184 884
tri 7184 882 7191 889 nw
rect 7034 872 7174 882
tri 7174 872 7184 882 nw
rect 574 820 580 872
rect 632 820 648 872
rect 700 820 706 872
rect 7034 871 7173 872
tri 7173 871 7174 872 nw
rect 574 806 706 820
rect 574 754 580 806
rect 632 754 648 806
rect 700 754 706 806
rect 3710 819 3716 871
rect 3768 819 3796 871
rect 3848 819 3876 871
rect 3928 819 3934 871
rect 3710 805 3934 819
rect 3710 753 3716 805
rect 3768 753 3796 805
rect 3848 753 3876 805
rect 3928 753 3934 805
rect 7034 849 7151 871
tri 7151 849 7173 871 nw
rect 7034 843 7145 849
tri 7145 843 7151 849 nw
rect 7034 839 7141 843
tri 7141 839 7145 843 nw
rect 9784 839 11347 889
tri 14409 882 14443 916 ne
rect 14443 882 14576 916
rect 14610 882 14654 916
rect 14688 882 14732 916
rect 14766 882 14810 916
rect 14844 882 14888 916
rect 14922 882 14966 916
rect 15000 887 15068 916
rect 15102 887 15114 921
rect 15000 882 15114 887
tri 14443 872 14453 882 ne
rect 14453 872 15114 882
tri 14453 871 14454 872 ne
rect 14454 871 15114 872
tri 14454 849 14476 871 ne
rect 14476 849 15114 871
tri 14476 843 14482 849 ne
rect 14482 843 15068 849
rect 7034 805 7107 839
tri 7107 805 7141 839 nw
rect 9784 805 9796 839
rect 9830 805 9872 839
rect 9906 805 9948 839
rect 9982 805 10024 839
rect 10058 805 10100 839
rect 10134 805 10176 839
rect 10210 805 10251 839
rect 10285 805 10326 839
rect 10360 805 10401 839
rect 10435 805 10476 839
rect 10510 805 10551 839
rect 10585 805 10626 839
rect 10660 805 10701 839
rect 10735 805 10776 839
rect 10810 805 10851 839
rect 10885 805 10926 839
rect 10960 805 11001 839
rect 11035 805 11076 839
rect 11110 805 11151 839
rect 11185 805 11226 839
rect 11260 805 11301 839
rect 11335 805 11347 839
tri 14482 809 14516 843 ne
rect 14516 809 14576 843
rect 14610 809 14654 843
rect 14688 809 14732 843
rect 14766 809 14810 843
rect 14844 809 14888 843
rect 14922 809 14966 843
rect 15000 815 15068 843
rect 15102 815 15114 849
rect 15000 809 15114 815
rect 7034 777 7079 805
tri 7079 777 7107 805 nw
rect 7034 770 7072 777
tri 7072 770 7079 777 nw
rect 7034 755 7057 770
tri 7057 755 7072 770 nw
rect 9784 755 11347 805
tri 14516 794 14531 809 ne
rect 14531 794 15114 809
rect 7034 753 7055 755
tri 7055 753 7057 755 nw
tri 7034 732 7055 753 nw
rect 9784 721 9796 755
rect 9830 721 9872 755
rect 9906 721 9948 755
rect 9982 721 10024 755
rect 10058 721 10100 755
rect 10134 721 10176 755
rect 10210 721 10251 755
rect 10285 721 10326 755
rect 10360 721 10401 755
rect 10435 721 10476 755
rect 10510 721 10551 755
rect 10585 721 10626 755
rect 10660 721 10701 755
rect 10735 721 10776 755
rect 10810 721 10851 755
rect 10885 721 10926 755
rect 10960 721 11001 755
rect 11035 721 11076 755
rect 11110 721 11151 755
rect 11185 721 11226 755
rect 11260 721 11301 755
rect 11335 721 11347 755
rect 11799 736 11831 794
tri 14531 777 14548 794 ne
rect 14548 777 15114 794
tri 14548 770 14555 777 ne
rect 14555 770 15068 777
tri 14555 759 14566 770 ne
rect 14566 736 14576 770
rect 14610 736 14654 770
rect 14688 736 14732 770
rect 14766 736 14810 770
rect 14844 736 14888 770
rect 14922 736 14966 770
rect 15000 743 15068 770
rect 15102 743 15114 777
rect 15000 736 15114 743
rect 761 683 794 715
rect 6527 686 6583 719
rect 9784 671 11347 721
rect 9784 637 9796 671
rect 9830 637 9872 671
rect 9906 637 9948 671
rect 9982 637 10024 671
rect 10058 637 10100 671
rect 10134 637 10176 671
rect 10210 637 10251 671
rect 10285 637 10326 671
rect 10360 637 10401 671
rect 10435 637 10476 671
rect 10510 637 10551 671
rect 10585 637 10626 671
rect 10660 637 10701 671
rect 10735 637 10776 671
rect 10810 637 10851 671
rect 10885 637 10926 671
rect 10960 637 11001 671
rect 11035 637 11076 671
rect 11110 637 11151 671
rect 11185 637 11226 671
rect 11260 637 11301 671
rect 11335 637 11347 671
rect 9784 587 11347 637
rect 9784 553 9796 587
rect 9830 553 9872 587
rect 9906 553 9948 587
rect 9982 553 10024 587
rect 10058 553 10100 587
rect 10134 553 10176 587
rect 10210 553 10251 587
rect 10285 553 10326 587
rect 10360 553 10401 587
rect 10435 553 10476 587
rect 10510 553 10551 587
rect 10585 553 10626 587
rect 10660 553 10701 587
rect 10735 553 10776 587
rect 10810 553 10851 587
rect 10885 553 10926 587
rect 10960 553 11001 587
rect 11035 553 11076 587
rect 11110 553 11151 587
rect 11185 553 11226 587
rect 11260 553 11301 587
rect 11335 553 11347 587
rect 9784 503 11347 553
rect 574 435 580 487
rect 632 435 648 487
rect 700 435 706 487
rect 574 421 706 435
rect 574 369 580 421
rect 632 369 648 421
rect 700 369 706 421
rect 3710 435 3716 487
rect 3768 435 3796 487
rect 3848 435 3876 487
rect 3928 435 3934 487
rect 9784 469 9796 503
rect 9830 469 9872 503
rect 9906 469 9948 503
rect 9982 469 10024 503
rect 10058 469 10100 503
rect 10134 469 10176 503
rect 10210 469 10251 503
rect 10285 469 10326 503
rect 10360 469 10401 503
rect 10435 469 10476 503
rect 10510 469 10551 503
rect 10585 469 10626 503
rect 10660 469 10701 503
rect 10735 469 10776 503
rect 10810 469 10851 503
rect 10885 469 10926 503
rect 10960 469 11001 503
rect 11035 469 11076 503
rect 11110 469 11151 503
rect 11185 469 11226 503
rect 11260 469 11301 503
rect 11335 469 11347 503
rect 9784 462 11347 469
rect 14566 705 15114 736
rect 14566 697 15068 705
rect 14566 663 14576 697
rect 14610 663 14654 697
rect 14688 663 14732 697
rect 14766 663 14810 697
rect 14844 663 14888 697
rect 14922 663 14966 697
rect 15000 671 15068 697
rect 15102 671 15114 705
rect 15000 663 15114 671
rect 14566 633 15114 663
rect 14566 623 15068 633
rect 14566 589 14576 623
rect 14610 589 14654 623
rect 14688 589 14732 623
rect 14766 589 14810 623
rect 14844 589 14888 623
rect 14922 589 14966 623
rect 15000 599 15068 623
rect 15102 599 15114 633
rect 15000 589 15114 599
rect 14566 561 15114 589
rect 14566 549 15068 561
rect 14566 515 14576 549
rect 14610 515 14654 549
rect 14688 515 14732 549
rect 14766 515 14810 549
rect 14844 515 14888 549
rect 14922 515 14966 549
rect 15000 527 15068 549
rect 15102 527 15114 561
rect 15000 515 15114 527
rect 14566 489 15114 515
rect 14566 475 15068 489
rect 3710 421 3934 435
rect 3710 369 3716 421
rect 3768 369 3796 421
rect 3848 369 3876 421
rect 3928 369 3934 421
rect 14566 441 14576 475
rect 14610 441 14654 475
rect 14688 441 14732 475
rect 14766 441 14810 475
rect 14844 441 14888 475
rect 14922 441 14966 475
rect 15000 455 15068 475
rect 15102 455 15114 489
rect 15000 441 15114 455
rect 14566 429 15114 441
tri 14566 417 14578 429 ne
rect 14578 417 15114 429
tri 14578 402 14593 417 ne
rect 14593 402 15068 417
tri 14593 390 14605 402 ne
rect 14605 390 15068 402
tri 14605 369 14626 390 ne
rect 14626 369 14657 390
tri 14626 356 14639 369 ne
rect 14639 356 14657 369
rect 14691 356 14735 390
rect 14769 356 14813 390
rect 14847 356 14891 390
rect 14925 356 14969 390
rect 15003 383 15068 390
rect 15102 383 15114 417
rect 15003 356 15114 383
tri 14639 355 14640 356 ne
rect 14640 345 15114 356
rect 14167 280 14252 332
rect 14640 312 15068 345
rect 14640 278 14657 312
rect 14691 278 14735 312
rect 14769 278 14813 312
rect 14847 278 14891 312
rect 14925 278 14969 312
rect 15003 311 15068 312
rect 15102 311 15114 345
rect 15003 278 15114 311
rect 14640 272 15114 278
rect 14640 238 15068 272
rect 15102 238 15114 272
rect 14640 234 15114 238
rect 13921 168 14073 220
rect 14640 200 14657 234
rect 14691 200 14735 234
rect 14769 200 14813 234
rect 14847 200 14891 234
rect 14925 200 14969 234
rect 15003 200 15114 234
rect 14640 199 15114 200
rect 14640 165 15068 199
rect 15102 165 15114 199
rect 14640 156 15114 165
rect 278 83 284 135
rect 336 83 348 135
rect 400 83 3716 135
rect 3768 83 3796 135
rect 3848 83 3876 135
rect 3928 83 3934 135
rect 14164 88 14240 140
rect 14640 122 14657 156
rect 14691 122 14735 156
rect 14769 122 14813 156
rect 14847 122 14891 156
rect 14925 122 14969 156
rect 15003 126 15114 156
rect 15003 122 15068 126
rect 14640 92 15068 122
rect 15102 92 15114 126
rect 14640 77 15114 92
rect 14640 43 14657 77
rect 14691 43 14735 77
rect 14769 43 14813 77
rect 14847 43 14891 77
rect 14925 43 14969 77
rect 15003 53 15114 77
rect 15003 43 15068 53
rect 14640 19 15068 43
rect 15102 19 15114 53
rect 14640 -23 15114 19
rect 49 -1067 83 -1013
rect 167 -1074 205 -1007
rect 258 -1075 313 -1023
rect 377 -1075 415 -1020
rect 5878 -9151 5930 -9145
rect 5878 -9223 5930 -9203
rect 5878 -9281 5930 -9275
rect 5247 -9994 5253 -9942
rect 5305 -9994 5328 -9942
rect 5380 -9994 5403 -9942
rect 5455 -9994 5478 -9942
rect 5530 -9994 5553 -9942
rect 5605 -9994 5627 -9942
rect 5679 -9994 5685 -9942
rect 5247 -10017 5685 -9994
rect 5247 -10069 5253 -10017
rect 5305 -10069 5328 -10017
rect 5380 -10069 5403 -10017
rect 5455 -10069 5478 -10017
rect 5530 -10069 5553 -10017
rect 5605 -10069 5627 -10017
rect 5679 -10069 5685 -10017
rect 5247 -10092 5685 -10069
rect 5247 -10144 5253 -10092
rect 5305 -10144 5328 -10092
rect 5380 -10144 5403 -10092
rect 5455 -10144 5478 -10092
rect 5530 -10144 5553 -10092
rect 5605 -10144 5627 -10092
rect 5679 -10144 5685 -10092
rect 5247 -10985 5253 -10933
rect 5305 -10985 5328 -10933
rect 5380 -10985 5403 -10933
rect 5455 -10985 5478 -10933
rect 5530 -10985 5553 -10933
rect 5605 -10985 5627 -10933
rect 5679 -10985 5685 -10933
rect 5247 -11011 5685 -10985
rect 5247 -11063 5253 -11011
rect 5305 -11063 5328 -11011
rect 5380 -11063 5403 -11011
rect 5455 -11063 5478 -11011
rect 5530 -11063 5553 -11011
rect 5605 -11063 5627 -11011
rect 5679 -11063 5685 -11011
<< rmetal1 >>
rect 9881 8258 9883 8259
rect 10183 8258 10185 8259
rect 9881 7996 9882 8258
rect 10184 7996 10185 8258
rect 9881 7995 9883 7996
rect 10183 7995 10185 7996
<< via1 >>
rect 359 16093 411 16145
rect 359 16029 411 16081
rect 278 15937 330 15989
rect 278 15873 330 15925
rect 541 9978 593 10030
rect 616 9978 668 10030
rect 690 9978 742 10030
rect 764 9978 816 10030
rect 838 9978 890 10030
rect 912 9978 964 10030
rect 541 9904 593 9956
rect 616 9904 668 9956
rect 690 9904 742 9956
rect 764 9904 816 9956
rect 838 9904 890 9956
rect 912 9904 964 9956
rect 541 9830 593 9882
rect 616 9830 668 9882
rect 690 9830 742 9882
rect 764 9830 816 9882
rect 838 9830 890 9882
rect 912 9830 964 9882
rect 12258 9342 12310 9359
rect 12335 9342 12387 9359
rect 12412 9342 12464 9359
rect 12488 9342 12540 9359
rect 12258 9308 12287 9342
rect 12287 9308 12310 9342
rect 12335 9308 12359 9342
rect 12359 9308 12387 9342
rect 12412 9308 12431 9342
rect 12431 9308 12464 9342
rect 12488 9308 12503 9342
rect 12503 9308 12537 9342
rect 12537 9308 12540 9342
rect 12258 9307 12310 9308
rect 12335 9307 12387 9308
rect 12412 9307 12464 9308
rect 12488 9307 12540 9308
rect 12564 9342 12616 9359
rect 12564 9308 12575 9342
rect 12575 9308 12609 9342
rect 12609 9308 12616 9342
rect 12564 9307 12616 9308
rect 12258 9256 12310 9271
rect 12335 9256 12387 9271
rect 12412 9256 12464 9271
rect 12488 9256 12540 9271
rect 12258 9222 12287 9256
rect 12287 9222 12310 9256
rect 12335 9222 12359 9256
rect 12359 9222 12387 9256
rect 12412 9222 12431 9256
rect 12431 9222 12464 9256
rect 12488 9222 12503 9256
rect 12503 9222 12537 9256
rect 12537 9222 12540 9256
rect 12258 9219 12310 9222
rect 12335 9219 12387 9222
rect 12412 9219 12464 9222
rect 12488 9219 12540 9222
rect 12564 9256 12616 9271
rect 12564 9222 12575 9256
rect 12575 9222 12609 9256
rect 12609 9222 12616 9256
rect 12564 9219 12616 9222
rect 12258 9170 12310 9183
rect 12335 9170 12387 9183
rect 12412 9170 12464 9183
rect 12488 9170 12540 9183
rect 12258 9136 12287 9170
rect 12287 9136 12310 9170
rect 12335 9136 12359 9170
rect 12359 9136 12387 9170
rect 12412 9136 12431 9170
rect 12431 9136 12464 9170
rect 12488 9136 12503 9170
rect 12503 9136 12537 9170
rect 12537 9136 12540 9170
rect 12258 9131 12310 9136
rect 12335 9131 12387 9136
rect 12412 9131 12464 9136
rect 12488 9131 12540 9136
rect 12564 9170 12616 9183
rect 12564 9136 12575 9170
rect 12575 9136 12609 9170
rect 12609 9136 12616 9170
rect 12564 9131 12616 9136
rect 14240 9408 14292 9460
rect 14312 9408 14364 9460
rect 14384 9408 14436 9460
rect 14456 9408 14508 9460
rect 14528 9408 14580 9460
rect 14600 9408 14652 9460
rect 14240 9343 14292 9395
rect 14312 9343 14364 9395
rect 14384 9343 14436 9395
rect 14456 9343 14508 9395
rect 14528 9343 14580 9395
rect 14600 9343 14652 9395
rect 14240 9278 14292 9330
rect 14312 9278 14364 9330
rect 14384 9278 14436 9330
rect 14456 9278 14508 9330
rect 14528 9278 14580 9330
rect 14600 9278 14652 9330
rect 14240 9213 14292 9265
rect 14312 9213 14364 9265
rect 14384 9213 14436 9265
rect 14456 9213 14508 9265
rect 14528 9213 14580 9265
rect 14600 9213 14652 9265
rect 14240 9148 14292 9200
rect 14312 9148 14364 9200
rect 14384 9148 14436 9200
rect 14456 9148 14508 9200
rect 14528 9148 14580 9200
rect 14600 9148 14652 9200
rect 14240 9083 14292 9135
rect 14312 9083 14364 9135
rect 14384 9083 14436 9135
rect 14456 9083 14508 9135
rect 14528 9083 14580 9135
rect 14600 9083 14652 9135
rect 14240 9018 14292 9070
rect 14312 9018 14364 9070
rect 14384 9018 14436 9070
rect 14456 9018 14508 9070
rect 14528 9018 14580 9070
rect 14600 9018 14652 9070
rect 14240 8953 14292 9005
rect 14312 8953 14364 9005
rect 14384 8953 14436 9005
rect 14456 8953 14508 9005
rect 14528 8953 14580 9005
rect 14600 8953 14652 9005
rect 14240 8888 14292 8940
rect 14312 8888 14364 8940
rect 14384 8888 14436 8940
rect 14456 8888 14508 8940
rect 14528 8888 14580 8940
rect 14600 8888 14652 8940
rect 541 8775 593 8827
rect 616 8775 668 8827
rect 690 8775 742 8827
rect 764 8775 816 8827
rect 838 8775 890 8827
rect 912 8775 964 8827
rect 14240 8823 14292 8875
rect 14312 8823 14364 8875
rect 14384 8823 14436 8875
rect 14456 8823 14508 8875
rect 14528 8823 14580 8875
rect 14600 8823 14652 8875
rect 14240 8760 14292 8810
rect 14312 8760 14364 8810
rect 14384 8760 14436 8810
rect 14456 8760 14508 8810
rect 14528 8760 14580 8810
rect 14600 8760 14652 8810
rect 541 8719 544 8751
rect 544 8719 578 8751
rect 578 8719 593 8751
rect 541 8699 593 8719
rect 616 8719 618 8751
rect 618 8719 652 8751
rect 652 8719 668 8751
rect 616 8699 668 8719
rect 690 8719 691 8751
rect 691 8719 725 8751
rect 725 8719 742 8751
rect 690 8699 742 8719
rect 764 8719 798 8751
rect 798 8719 816 8751
rect 838 8719 871 8751
rect 871 8719 890 8751
rect 764 8699 816 8719
rect 838 8699 890 8719
rect 912 8726 946 8751
rect 946 8726 964 8751
rect 912 8699 964 8726
rect 14240 8758 14267 8760
rect 14267 8758 14292 8760
rect 14312 8758 14339 8760
rect 14339 8758 14364 8760
rect 14384 8758 14411 8760
rect 14411 8758 14436 8760
rect 14456 8758 14483 8760
rect 14483 8758 14508 8760
rect 14528 8758 14555 8760
rect 14555 8758 14580 8760
rect 14600 8758 14627 8760
rect 14627 8758 14652 8760
rect 14240 8726 14267 8745
rect 14267 8726 14292 8745
rect 14312 8726 14339 8745
rect 14339 8726 14364 8745
rect 14384 8726 14411 8745
rect 14411 8726 14436 8745
rect 14456 8726 14483 8745
rect 14483 8726 14508 8745
rect 14528 8726 14555 8745
rect 14555 8726 14580 8745
rect 14600 8726 14627 8745
rect 14627 8726 14652 8745
rect 842 8618 894 8670
rect 912 8636 964 8670
rect 14240 8693 14292 8726
rect 14312 8693 14364 8726
rect 14384 8693 14436 8726
rect 14456 8693 14508 8726
rect 14528 8693 14580 8726
rect 14600 8693 14652 8726
rect 14240 8636 14292 8680
rect 14312 8636 14364 8680
rect 14384 8636 14436 8680
rect 14456 8636 14508 8680
rect 14528 8636 14580 8680
rect 14600 8636 14652 8680
rect 912 8618 946 8636
rect 946 8618 964 8636
rect 14240 8628 14267 8636
rect 14267 8628 14292 8636
rect 14312 8628 14339 8636
rect 14339 8628 14364 8636
rect 14384 8628 14411 8636
rect 14411 8628 14436 8636
rect 14456 8628 14483 8636
rect 14483 8628 14508 8636
rect 14528 8628 14555 8636
rect 14555 8628 14580 8636
rect 14600 8628 14627 8636
rect 14627 8628 14652 8636
rect 14240 8602 14267 8615
rect 14267 8602 14292 8615
rect 14312 8602 14339 8615
rect 14339 8602 14364 8615
rect 14384 8602 14411 8615
rect 14411 8602 14436 8615
rect 14456 8602 14483 8615
rect 14483 8602 14508 8615
rect 14528 8602 14555 8615
rect 14555 8602 14580 8615
rect 14600 8602 14627 8615
rect 14627 8602 14652 8615
rect 14240 8563 14292 8602
rect 14312 8563 14364 8602
rect 14384 8563 14436 8602
rect 14456 8563 14508 8602
rect 14528 8563 14580 8602
rect 14600 8563 14652 8602
rect 14240 8512 14292 8550
rect 14240 8498 14257 8512
rect 14257 8498 14291 8512
rect 14291 8498 14292 8512
rect 14312 8512 14364 8550
rect 14312 8498 14329 8512
rect 14329 8498 14363 8512
rect 14363 8498 14364 8512
rect 14384 8512 14436 8550
rect 14384 8498 14401 8512
rect 14401 8498 14435 8512
rect 14435 8498 14436 8512
rect 14456 8512 14508 8550
rect 14456 8498 14473 8512
rect 14473 8498 14507 8512
rect 14507 8498 14508 8512
rect 14528 8498 14580 8550
rect 14600 8498 14652 8550
rect 14240 8478 14257 8485
rect 14257 8478 14291 8485
rect 14291 8478 14292 8485
rect 14240 8435 14292 8478
rect 14240 8433 14257 8435
rect 14257 8433 14291 8435
rect 14291 8433 14292 8435
rect 14312 8478 14329 8485
rect 14329 8478 14363 8485
rect 14363 8478 14364 8485
rect 14312 8435 14364 8478
rect 14312 8433 14329 8435
rect 14329 8433 14363 8435
rect 14363 8433 14364 8435
rect 14384 8478 14401 8485
rect 14401 8478 14435 8485
rect 14435 8478 14436 8485
rect 14384 8435 14436 8478
rect 14384 8433 14401 8435
rect 14401 8433 14435 8435
rect 14435 8433 14436 8435
rect 14456 8478 14473 8485
rect 14473 8478 14507 8485
rect 14507 8478 14508 8485
rect 14456 8435 14508 8478
rect 14456 8433 14473 8435
rect 14473 8433 14507 8435
rect 14507 8433 14508 8435
rect 14528 8433 14580 8485
rect 14600 8462 14652 8485
rect 14600 8433 14614 8462
rect 14614 8433 14648 8462
rect 14648 8433 14652 8462
rect 14240 8401 14257 8420
rect 14257 8401 14291 8420
rect 14291 8401 14292 8420
rect 14240 8368 14292 8401
rect 14312 8401 14329 8420
rect 14329 8401 14363 8420
rect 14363 8401 14364 8420
rect 14312 8368 14364 8401
rect 14384 8401 14401 8420
rect 14401 8401 14435 8420
rect 14435 8401 14436 8420
rect 14384 8368 14436 8401
rect 14456 8401 14473 8420
rect 14473 8401 14507 8420
rect 14507 8401 14508 8420
rect 14456 8368 14508 8401
rect 14528 8368 14580 8420
rect 14600 8388 14652 8420
rect 14600 8368 14614 8388
rect 14614 8368 14648 8388
rect 14648 8368 14652 8388
rect 14240 8324 14257 8354
rect 14257 8324 14291 8354
rect 14291 8324 14292 8354
rect 14240 8302 14292 8324
rect 14312 8324 14329 8354
rect 14329 8324 14363 8354
rect 14363 8324 14364 8354
rect 14312 8302 14364 8324
rect 14384 8324 14401 8354
rect 14401 8324 14435 8354
rect 14435 8324 14436 8354
rect 14384 8302 14436 8324
rect 14456 8324 14473 8354
rect 14473 8324 14507 8354
rect 14507 8324 14508 8354
rect 14456 8302 14508 8324
rect 14528 8302 14580 8354
rect 14600 8314 14652 8354
rect 14600 8302 14614 8314
rect 14614 8302 14648 8314
rect 14648 8302 14652 8314
rect 10800 8254 10852 8281
rect 10800 8229 10804 8254
rect 10804 8229 10838 8254
rect 10838 8229 10852 8254
rect 10876 8254 10928 8281
rect 10876 8229 10898 8254
rect 10898 8229 10928 8254
rect 10952 8229 11004 8281
rect 11028 8229 11080 8281
rect 11104 8229 11156 8281
rect 10800 8179 10852 8214
rect 10800 8162 10804 8179
rect 10804 8162 10838 8179
rect 10838 8162 10852 8179
rect 10876 8179 10928 8214
rect 10876 8162 10898 8179
rect 10898 8162 10928 8179
rect 10952 8162 11004 8214
rect 11028 8162 11080 8214
rect 11104 8162 11156 8214
rect 10800 8145 10804 8147
rect 10804 8145 10838 8147
rect 10838 8145 10852 8147
rect 10800 8104 10852 8145
rect 10800 8095 10804 8104
rect 10804 8095 10838 8104
rect 10838 8095 10852 8104
rect 10876 8145 10898 8147
rect 10898 8145 10928 8147
rect 10876 8104 10928 8145
rect 10876 8095 10898 8104
rect 10898 8095 10928 8104
rect 10952 8095 11004 8147
rect 11028 8095 11080 8147
rect 11104 8095 11156 8147
rect 10800 8070 10804 8079
rect 10804 8070 10838 8079
rect 10838 8070 10852 8079
rect 10800 8028 10852 8070
rect 10800 8027 10804 8028
rect 10804 8027 10838 8028
rect 10838 8027 10852 8028
rect 10876 8070 10898 8079
rect 10898 8070 10928 8079
rect 10876 8028 10928 8070
rect 10876 8027 10898 8028
rect 10898 8027 10928 8028
rect 10952 8027 11004 8079
rect 11028 8027 11080 8079
rect 11104 8027 11156 8079
rect 10800 7994 10804 8011
rect 10804 7994 10838 8011
rect 10838 7994 10852 8011
rect 10800 7959 10852 7994
rect 10876 7994 10898 8011
rect 10898 7994 10928 8011
rect 10876 7959 10928 7994
rect 10952 7959 11004 8011
rect 11028 7959 11080 8011
rect 11104 7959 11156 8011
rect 10800 7918 10804 7943
rect 10804 7918 10838 7943
rect 10838 7918 10852 7943
rect 10800 7891 10852 7918
rect 10876 7918 10898 7943
rect 10898 7918 10928 7943
rect 10876 7891 10928 7918
rect 10952 7891 11004 7943
rect 11028 7891 11080 7943
rect 11104 7891 11156 7943
rect 12255 8229 12307 8281
rect 12333 8229 12385 8281
rect 12411 8229 12463 8281
rect 12489 8229 12541 8281
rect 12567 8229 12619 8281
rect 14240 8280 14292 8288
rect 12255 8158 12307 8210
rect 12333 8158 12385 8210
rect 12411 8158 12463 8210
rect 12489 8158 12541 8210
rect 12567 8158 12619 8210
rect 12255 8087 12307 8139
rect 12333 8087 12385 8139
rect 12411 8087 12463 8139
rect 12489 8087 12541 8139
rect 12567 8087 12619 8139
rect 12255 8016 12307 8068
rect 12333 8016 12385 8068
rect 12411 8016 12463 8068
rect 12489 8016 12541 8068
rect 12567 8016 12619 8068
rect 12255 7945 12307 7997
rect 12333 7945 12385 7997
rect 12411 7945 12463 7997
rect 12489 7945 12541 7997
rect 12567 7945 12619 7997
rect 12255 7873 12307 7925
rect 12333 7873 12385 7925
rect 12411 7873 12463 7925
rect 12489 7873 12541 7925
rect 12567 7873 12619 7925
rect 14240 8246 14257 8280
rect 14257 8246 14291 8280
rect 14291 8246 14292 8280
rect 14240 8236 14292 8246
rect 14312 8280 14364 8288
rect 14312 8246 14329 8280
rect 14329 8246 14363 8280
rect 14363 8246 14364 8280
rect 14312 8236 14364 8246
rect 14384 8280 14436 8288
rect 14384 8246 14401 8280
rect 14401 8246 14435 8280
rect 14435 8246 14436 8280
rect 14384 8236 14436 8246
rect 14456 8280 14508 8288
rect 14456 8246 14473 8280
rect 14473 8246 14507 8280
rect 14507 8246 14508 8280
rect 14456 8236 14508 8246
rect 14528 8236 14580 8288
rect 14600 8280 14614 8288
rect 14614 8280 14648 8288
rect 14648 8280 14652 8288
rect 14600 8240 14652 8280
rect 14600 8236 14614 8240
rect 14614 8236 14648 8240
rect 14648 8236 14652 8240
rect 14240 8202 14292 8222
rect 14240 8170 14257 8202
rect 14257 8170 14291 8202
rect 14291 8170 14292 8202
rect 14312 8202 14364 8222
rect 14312 8170 14329 8202
rect 14329 8170 14363 8202
rect 14363 8170 14364 8202
rect 14384 8202 14436 8222
rect 14384 8170 14401 8202
rect 14401 8170 14435 8202
rect 14435 8170 14436 8202
rect 14456 8202 14508 8222
rect 14456 8170 14473 8202
rect 14473 8170 14507 8202
rect 14507 8170 14508 8202
rect 14528 8170 14580 8222
rect 14600 8206 14614 8222
rect 14614 8206 14648 8222
rect 14648 8206 14652 8222
rect 14600 8170 14652 8206
rect 14240 8104 14292 8156
rect 14312 8104 14364 8156
rect 14384 8115 14436 8156
rect 14456 8115 14508 8156
rect 14528 8115 14580 8156
rect 14384 8104 14431 8115
rect 14431 8104 14436 8115
rect 14456 8104 14465 8115
rect 14465 8104 14508 8115
rect 14528 8104 14545 8115
rect 14545 8104 14580 8115
rect 14600 8132 14614 8156
rect 14614 8132 14648 8156
rect 14648 8132 14652 8156
rect 14600 8104 14652 8132
rect 278 7799 330 7851
rect 278 7733 330 7785
rect 278 7666 330 7718
rect 278 7599 330 7651
rect 278 7532 330 7584
rect 11135 7509 11187 7561
rect 11208 7509 11260 7561
rect 11280 7509 11332 7561
rect 11135 7429 11187 7481
rect 11208 7429 11260 7481
rect 11280 7429 11332 7481
rect 338 6822 390 6874
rect 338 6756 390 6808
rect 516 5516 568 5568
rect 634 5516 686 5568
rect 751 5516 803 5568
rect 14313 5513 14365 5565
rect 435 5413 487 5465
rect 507 5413 559 5465
rect 579 5413 631 5465
rect 651 5413 703 5465
rect 748 5427 800 5479
rect 435 5348 487 5400
rect 507 5348 559 5400
rect 579 5348 631 5400
rect 651 5348 703 5400
rect 435 5283 487 5335
rect 507 5283 559 5335
rect 579 5283 631 5335
rect 651 5283 703 5335
rect 435 5218 487 5270
rect 507 5218 559 5270
rect 579 5218 631 5270
rect 651 5218 703 5270
rect 435 5153 487 5205
rect 507 5153 559 5205
rect 579 5153 631 5205
rect 651 5153 703 5205
rect 435 5088 487 5140
rect 507 5088 559 5140
rect 579 5088 631 5140
rect 651 5088 703 5140
rect 435 5023 487 5075
rect 507 5023 559 5075
rect 579 5023 631 5075
rect 651 5023 703 5075
rect 435 4958 487 5010
rect 507 4958 559 5010
rect 579 4958 631 5010
rect 651 4958 703 5010
rect 435 4893 487 4945
rect 507 4893 559 4945
rect 579 4893 631 4945
rect 651 4893 703 4945
rect 435 4828 487 4880
rect 507 4828 559 4880
rect 579 4828 631 4880
rect 651 4828 703 4880
rect 435 4763 487 4815
rect 507 4763 559 4815
rect 579 4763 631 4815
rect 651 4763 703 4815
rect 435 4698 487 4750
rect 507 4698 559 4750
rect 579 4698 631 4750
rect 651 4698 703 4750
rect 435 4633 487 4685
rect 507 4633 559 4685
rect 579 4633 631 4685
rect 651 4633 703 4685
rect 435 4568 487 4620
rect 507 4568 559 4620
rect 579 4568 631 4620
rect 651 4568 703 4620
rect 435 4503 487 4555
rect 507 4503 559 4555
rect 579 4503 631 4555
rect 651 4503 703 4555
rect 435 4438 487 4490
rect 507 4438 559 4490
rect 579 4438 631 4490
rect 651 4438 703 4490
rect 435 4373 487 4425
rect 507 4373 559 4425
rect 579 4373 631 4425
rect 651 4373 703 4425
rect 435 4308 487 4360
rect 507 4308 559 4360
rect 579 4308 631 4360
rect 651 4308 703 4360
rect 435 4243 487 4295
rect 507 4243 559 4295
rect 579 4243 631 4295
rect 651 4243 703 4295
rect 435 4178 487 4230
rect 507 4178 559 4230
rect 579 4178 631 4230
rect 651 4178 703 4230
rect 435 4113 487 4165
rect 507 4113 559 4165
rect 579 4113 631 4165
rect 651 4113 703 4165
rect 435 4047 487 4099
rect 507 4047 559 4099
rect 579 4047 631 4099
rect 651 4047 703 4099
rect 435 3981 487 4033
rect 507 3981 559 4033
rect 579 3981 631 4033
rect 651 3981 703 4033
rect 435 3915 487 3967
rect 507 3915 559 3967
rect 579 3915 631 3967
rect 651 3915 703 3967
rect 435 3849 487 3901
rect 507 3849 559 3901
rect 579 3849 631 3901
rect 651 3849 703 3901
rect 435 3783 487 3835
rect 507 3783 559 3835
rect 579 3783 631 3835
rect 651 3783 703 3835
rect 435 3717 487 3769
rect 507 3717 559 3769
rect 579 3717 631 3769
rect 651 3717 703 3769
rect 435 3651 487 3703
rect 507 3651 559 3703
rect 579 3651 631 3703
rect 651 3651 703 3703
rect 14243 5413 14295 5465
rect 14309 5413 14361 5465
rect 14375 5413 14427 5465
rect 14441 5413 14493 5465
rect 14243 5348 14295 5400
rect 14309 5348 14361 5400
rect 14375 5348 14427 5400
rect 14441 5348 14493 5400
rect 14243 5283 14295 5335
rect 14309 5283 14361 5335
rect 14375 5283 14427 5335
rect 14441 5283 14493 5335
rect 14243 5218 14295 5270
rect 14309 5218 14361 5270
rect 14375 5218 14427 5270
rect 14441 5218 14493 5270
rect 14243 5153 14295 5205
rect 14309 5153 14361 5205
rect 14375 5153 14427 5205
rect 14441 5153 14493 5205
rect 14243 5088 14295 5140
rect 14309 5088 14361 5140
rect 14375 5088 14427 5140
rect 14441 5088 14493 5140
rect 14243 5023 14295 5075
rect 14309 5023 14361 5075
rect 14375 5023 14427 5075
rect 14441 5023 14493 5075
rect 14243 4958 14295 5010
rect 14309 4958 14361 5010
rect 14375 4958 14427 5010
rect 14441 4958 14493 5010
rect 14243 4893 14295 4945
rect 14309 4893 14361 4945
rect 14375 4893 14427 4945
rect 14441 4893 14493 4945
rect 14243 4828 14295 4880
rect 14309 4828 14361 4880
rect 14375 4828 14427 4880
rect 14441 4828 14493 4880
rect 14243 4763 14295 4815
rect 14309 4763 14361 4815
rect 14375 4763 14427 4815
rect 14441 4763 14493 4815
rect 14243 4698 14295 4750
rect 14309 4698 14361 4750
rect 14375 4698 14427 4750
rect 14441 4698 14493 4750
rect 14243 4633 14295 4685
rect 14309 4633 14361 4685
rect 14375 4633 14427 4685
rect 14441 4633 14493 4685
rect 14243 4568 14295 4620
rect 14309 4568 14361 4620
rect 14375 4568 14427 4620
rect 14441 4568 14493 4620
rect 14243 4503 14295 4555
rect 14309 4503 14361 4555
rect 14375 4503 14427 4555
rect 14441 4503 14493 4555
rect 14243 4438 14295 4490
rect 14309 4438 14361 4490
rect 14375 4438 14427 4490
rect 14441 4438 14493 4490
rect 14243 4373 14295 4425
rect 14309 4373 14361 4425
rect 14375 4373 14427 4425
rect 14441 4373 14493 4425
rect 14243 4307 14295 4359
rect 14309 4307 14361 4359
rect 14375 4307 14427 4359
rect 14441 4307 14493 4359
rect 14243 4241 14295 4293
rect 14309 4241 14361 4293
rect 14375 4241 14427 4293
rect 14441 4241 14493 4293
rect 14243 4175 14295 4227
rect 14309 4175 14361 4227
rect 14375 4175 14427 4227
rect 14441 4175 14493 4227
rect 14243 4109 14295 4161
rect 14309 4109 14361 4161
rect 14375 4109 14427 4161
rect 14441 4109 14493 4161
rect 14243 4043 14295 4095
rect 14309 4043 14361 4095
rect 14375 4043 14427 4095
rect 14441 4043 14493 4095
rect 14243 3977 14295 4029
rect 14309 3977 14361 4029
rect 14375 3977 14427 4029
rect 14441 3977 14493 4029
rect 14243 3911 14295 3963
rect 14309 3911 14361 3963
rect 14375 3911 14427 3963
rect 14441 3911 14493 3963
rect 14243 3845 14295 3897
rect 14309 3845 14361 3897
rect 14375 3845 14427 3897
rect 14441 3845 14493 3897
rect 14243 3779 14295 3831
rect 14309 3779 14361 3831
rect 14375 3779 14427 3831
rect 14441 3779 14493 3831
rect 14243 3713 14295 3765
rect 14309 3713 14361 3765
rect 14375 3713 14427 3765
rect 14441 3713 14493 3765
rect 14243 3647 14295 3699
rect 14309 3647 14361 3699
rect 14375 3647 14427 3699
rect 14441 3647 14493 3699
rect 580 820 632 872
rect 648 820 700 872
rect 580 754 632 806
rect 648 754 700 806
rect 3716 819 3768 871
rect 3796 819 3848 871
rect 3876 819 3928 871
rect 3716 753 3768 805
rect 3796 753 3848 805
rect 3876 753 3928 805
rect 580 435 632 487
rect 648 435 700 487
rect 580 369 632 421
rect 648 369 700 421
rect 3716 435 3768 487
rect 3796 435 3848 487
rect 3876 435 3928 487
rect 3716 369 3768 421
rect 3796 369 3848 421
rect 3876 369 3928 421
rect 284 83 336 135
rect 348 83 400 135
rect 3716 83 3768 135
rect 3796 83 3848 135
rect 3876 83 3928 135
rect 5878 -9157 5930 -9151
rect 5878 -9191 5884 -9157
rect 5884 -9191 5918 -9157
rect 5918 -9191 5930 -9157
rect 5878 -9203 5930 -9191
rect 5878 -9229 5930 -9223
rect 5878 -9263 5884 -9229
rect 5884 -9263 5918 -9229
rect 5918 -9263 5930 -9229
rect 5878 -9275 5930 -9263
rect 5253 -9994 5305 -9942
rect 5328 -9994 5380 -9942
rect 5403 -9994 5455 -9942
rect 5478 -9994 5530 -9942
rect 5553 -9994 5605 -9942
rect 5627 -9994 5679 -9942
rect 5253 -10069 5305 -10017
rect 5328 -10069 5380 -10017
rect 5403 -10069 5455 -10017
rect 5478 -10069 5530 -10017
rect 5553 -10069 5605 -10017
rect 5627 -10069 5679 -10017
rect 5253 -10144 5305 -10092
rect 5328 -10144 5380 -10092
rect 5403 -10144 5455 -10092
rect 5478 -10144 5530 -10092
rect 5553 -10144 5605 -10092
rect 5627 -10144 5679 -10092
rect 5253 -10985 5305 -10933
rect 5328 -10985 5380 -10933
rect 5403 -10985 5455 -10933
rect 5478 -10985 5530 -10933
rect 5553 -10985 5605 -10933
rect 5627 -10985 5679 -10933
rect 5253 -11063 5305 -11011
rect 5328 -11063 5380 -11011
rect 5403 -11063 5455 -11011
rect 5478 -11063 5530 -11011
rect 5553 -11063 5605 -11011
rect 5627 -11063 5679 -11011
<< metal2 >>
tri 385 16276 406 16297 ne
rect 406 16204 437 16242
tri 406 16183 427 16204 ne
rect 427 16183 437 16204
tri 437 16183 469 16215 sw
tri 427 16173 437 16183 ne
rect 437 16173 469 16183
tri 437 16171 439 16173 ne
rect 359 16145 411 16151
rect 359 16081 411 16093
rect 359 16023 411 16029
rect 278 15989 330 15995
rect 278 15925 330 15937
rect 278 15867 330 15873
rect 278 15850 313 15867
tri 313 15850 330 15867 nw
rect 278 7873 310 15850
tri 310 15847 313 15850 nw
tri 356 15847 359 15850 se
rect 359 15847 399 16023
tri 399 16011 411 16023 nw
tri 341 15832 356 15847 se
rect 356 15832 399 15847
tri 338 15829 341 15832 se
rect 341 15829 378 15832
rect 338 7959 378 15829
tri 378 15811 399 15832 nw
tri 406 15769 439 15802 se
rect 439 15790 469 16173
rect 439 15769 448 15790
tri 448 15769 469 15790 nw
rect 406 15684 437 15769
tri 437 15758 448 15769 nw
rect 4395 12316 7294 13416
rect 11116 10850 12657 11943
rect 535 10030 970 10031
rect 535 9978 541 10030
rect 593 9978 616 10030
rect 668 9978 690 10030
rect 742 9978 764 10030
rect 816 9978 838 10030
rect 890 9978 912 10030
rect 964 9978 970 10030
rect 535 9956 970 9978
rect 535 9904 541 9956
rect 593 9904 616 9956
rect 668 9904 690 9956
rect 742 9904 764 9956
rect 816 9904 838 9956
rect 890 9904 912 9956
rect 964 9904 970 9956
rect 535 9882 970 9904
rect 535 9830 541 9882
rect 593 9830 616 9882
rect 668 9830 690 9882
rect 742 9830 764 9882
rect 816 9830 838 9882
rect 890 9830 912 9882
rect 964 9830 970 9882
rect 535 8827 970 9830
rect 14240 9460 14652 9466
rect 14292 9408 14312 9460
rect 14364 9408 14384 9460
rect 14436 9408 14456 9460
rect 14508 9408 14528 9460
rect 14580 9408 14600 9460
rect 14240 9395 14652 9408
rect 535 8775 541 8827
rect 593 8775 616 8827
rect 668 8775 690 8827
rect 742 8775 764 8827
rect 816 8775 838 8827
rect 890 8775 912 8827
rect 964 8775 970 8827
rect 535 8751 970 8775
rect 535 8699 541 8751
rect 593 8699 616 8751
rect 668 8699 690 8751
rect 742 8699 764 8751
rect 816 8699 838 8751
rect 890 8699 912 8751
rect 964 8699 970 8751
rect 535 8670 970 8699
rect 535 8618 842 8670
rect 894 8618 912 8670
rect 964 8618 970 8670
tri 378 7959 383 7964 sw
rect 338 7945 383 7959
tri 383 7945 397 7959 sw
rect 338 7943 397 7945
tri 397 7943 399 7945 sw
rect 338 7942 399 7943
tri 399 7942 400 7943 sw
rect 338 7913 400 7942
tri 338 7891 360 7913 ne
tri 310 7873 314 7877 sw
rect 278 7857 314 7873
tri 314 7857 330 7873 sw
rect 278 7851 330 7857
rect 278 7785 330 7799
rect 278 7718 330 7733
rect 278 7651 330 7666
rect 278 7584 330 7599
rect 278 7526 330 7532
rect 278 135 310 7526
tri 310 7509 327 7526 nw
tri 338 7347 360 7369 se
rect 360 7347 400 7913
rect 338 7338 400 7347
rect 338 6880 378 7338
tri 378 7316 400 7338 nw
tri 435 7071 535 7171 se
rect 535 7071 970 8618
rect 12252 9359 12622 9360
rect 12252 9307 12258 9359
rect 12310 9307 12335 9359
rect 12387 9307 12412 9359
rect 12464 9307 12488 9359
rect 12540 9307 12564 9359
rect 12616 9307 12622 9359
rect 12252 9271 12622 9307
rect 12252 9219 12258 9271
rect 12310 9219 12335 9271
rect 12387 9219 12412 9271
rect 12464 9219 12488 9271
rect 12540 9219 12564 9271
rect 12616 9219 12622 9271
rect 12252 9183 12622 9219
rect 12252 9131 12258 9183
rect 12310 9131 12335 9183
rect 12387 9131 12412 9183
rect 12464 9131 12488 9183
rect 12540 9131 12564 9183
rect 12616 9131 12622 9183
rect 10800 8281 11156 8287
rect 10852 8229 10876 8281
rect 10928 8229 10952 8281
rect 11004 8229 11028 8281
rect 11080 8229 11104 8281
rect 10800 8214 11156 8229
rect 10852 8162 10876 8214
rect 10928 8162 10952 8214
rect 11004 8162 11028 8214
rect 11080 8162 11104 8214
rect 10800 8147 11156 8162
rect 10852 8095 10876 8147
rect 10928 8095 10952 8147
rect 11004 8095 11028 8147
rect 11080 8095 11104 8147
rect 10800 8079 11156 8095
rect 10852 8027 10876 8079
rect 10928 8027 10952 8079
rect 11004 8027 11028 8079
rect 11080 8027 11104 8079
rect 10800 8011 11156 8027
rect 10852 7959 10876 8011
rect 10928 7959 10952 8011
rect 11004 7959 11028 8011
rect 11080 7959 11104 8011
rect 10800 7943 11156 7959
rect 10852 7891 10876 7943
rect 10928 7891 10952 7943
rect 11004 7891 11028 7943
rect 11080 7891 11104 7943
rect 10800 7561 11156 7891
rect 12252 8281 12622 9131
rect 12252 8229 12255 8281
rect 12307 8229 12333 8281
rect 12385 8229 12411 8281
rect 12463 8229 12489 8281
rect 12541 8229 12567 8281
rect 12619 8229 12622 8281
rect 12252 8210 12622 8229
rect 12252 8158 12255 8210
rect 12307 8158 12333 8210
rect 12385 8158 12411 8210
rect 12463 8158 12489 8210
rect 12541 8158 12567 8210
rect 12619 8158 12622 8210
rect 12252 8139 12622 8158
rect 12252 8087 12255 8139
rect 12307 8087 12333 8139
rect 12385 8087 12411 8139
rect 12463 8087 12489 8139
rect 12541 8087 12567 8139
rect 12619 8087 12622 8139
rect 12252 8068 12622 8087
rect 12252 8016 12255 8068
rect 12307 8016 12333 8068
rect 12385 8016 12411 8068
rect 12463 8016 12489 8068
rect 12541 8016 12567 8068
rect 12619 8016 12622 8068
rect 12252 7997 12622 8016
rect 12252 7945 12255 7997
rect 12307 7945 12333 7997
rect 12385 7945 12411 7997
rect 12463 7945 12489 7997
rect 12541 7945 12567 7997
rect 12619 7945 12622 7997
rect 12252 7925 12622 7945
rect 12252 7873 12255 7925
rect 12307 7873 12333 7925
rect 12385 7873 12411 7925
rect 12463 7873 12489 7925
rect 12541 7873 12567 7925
rect 12619 7873 12622 7925
rect 12252 7867 12622 7873
rect 14292 9343 14312 9395
rect 14364 9343 14384 9395
rect 14436 9343 14456 9395
rect 14508 9343 14528 9395
rect 14580 9343 14600 9395
rect 14240 9330 14652 9343
rect 14292 9278 14312 9330
rect 14364 9278 14384 9330
rect 14436 9278 14456 9330
rect 14508 9278 14528 9330
rect 14580 9278 14600 9330
rect 14240 9265 14652 9278
rect 14292 9213 14312 9265
rect 14364 9213 14384 9265
rect 14436 9213 14456 9265
rect 14508 9213 14528 9265
rect 14580 9213 14600 9265
rect 14240 9200 14652 9213
rect 14292 9148 14312 9200
rect 14364 9148 14384 9200
rect 14436 9148 14456 9200
rect 14508 9148 14528 9200
rect 14580 9148 14600 9200
rect 14240 9135 14652 9148
rect 14292 9083 14312 9135
rect 14364 9083 14384 9135
rect 14436 9083 14456 9135
rect 14508 9083 14528 9135
rect 14580 9083 14600 9135
rect 14240 9070 14652 9083
rect 14292 9018 14312 9070
rect 14364 9018 14384 9070
rect 14436 9018 14456 9070
rect 14508 9018 14528 9070
rect 14580 9018 14600 9070
rect 14240 9005 14652 9018
rect 14292 8953 14312 9005
rect 14364 8953 14384 9005
rect 14436 8953 14456 9005
rect 14508 8953 14528 9005
rect 14580 8953 14600 9005
rect 14240 8940 14652 8953
rect 14292 8888 14312 8940
rect 14364 8888 14384 8940
rect 14436 8888 14456 8940
rect 14508 8888 14528 8940
rect 14580 8888 14600 8940
rect 14240 8875 14652 8888
rect 14292 8823 14312 8875
rect 14364 8823 14384 8875
rect 14436 8823 14456 8875
rect 14508 8823 14528 8875
rect 14580 8823 14600 8875
rect 14240 8810 14652 8823
rect 14292 8758 14312 8810
rect 14364 8758 14384 8810
rect 14436 8758 14456 8810
rect 14508 8758 14528 8810
rect 14580 8758 14600 8810
rect 14240 8745 14652 8758
rect 14292 8693 14312 8745
rect 14364 8693 14384 8745
rect 14436 8693 14456 8745
rect 14508 8693 14528 8745
rect 14580 8693 14600 8745
rect 14240 8680 14652 8693
rect 14292 8628 14312 8680
rect 14364 8628 14384 8680
rect 14436 8628 14456 8680
rect 14508 8628 14528 8680
rect 14580 8628 14600 8680
rect 14240 8615 14652 8628
rect 14292 8563 14312 8615
rect 14364 8563 14384 8615
rect 14436 8563 14456 8615
rect 14508 8563 14528 8615
rect 14580 8563 14600 8615
rect 14240 8550 14652 8563
rect 14292 8498 14312 8550
rect 14364 8498 14384 8550
rect 14436 8498 14456 8550
rect 14508 8498 14528 8550
rect 14580 8498 14600 8550
rect 14240 8485 14652 8498
rect 14292 8433 14312 8485
rect 14364 8433 14384 8485
rect 14436 8433 14456 8485
rect 14508 8433 14528 8485
rect 14580 8433 14600 8485
rect 14240 8420 14652 8433
rect 14292 8368 14312 8420
rect 14364 8368 14384 8420
rect 14436 8368 14456 8420
rect 14508 8368 14528 8420
rect 14580 8368 14600 8420
rect 14240 8354 14652 8368
rect 14292 8302 14312 8354
rect 14364 8302 14384 8354
rect 14436 8302 14456 8354
rect 14508 8302 14528 8354
rect 14580 8302 14600 8354
rect 14240 8288 14652 8302
rect 14292 8236 14312 8288
rect 14364 8236 14384 8288
rect 14436 8236 14456 8288
rect 14508 8236 14528 8288
rect 14580 8236 14600 8288
rect 14240 8222 14652 8236
rect 14292 8170 14312 8222
rect 14364 8170 14384 8222
rect 14436 8170 14456 8222
rect 14508 8170 14528 8222
rect 14580 8170 14600 8222
rect 14240 8156 14652 8170
rect 14292 8104 14312 8156
rect 14364 8104 14384 8156
rect 14436 8104 14456 8156
rect 14508 8104 14528 8156
rect 14580 8104 14600 8156
tri 11156 7561 11338 7743 sw
rect 10800 7509 11135 7561
rect 11187 7509 11208 7561
rect 11260 7509 11280 7561
rect 11332 7509 11338 7561
rect 10800 7481 11338 7509
rect 10800 7429 11135 7481
rect 11187 7429 11208 7481
rect 11260 7429 11280 7481
rect 11332 7429 11338 7481
rect 435 6992 970 7071
rect 435 6892 870 6992
tri 870 6892 970 6992 nw
tri 378 6880 390 6892 sw
rect 338 6874 390 6880
rect 338 6808 390 6822
rect 338 6750 390 6756
rect 338 872 378 6750
tri 378 6738 390 6750 nw
rect 435 5568 823 6892
tri 823 6845 870 6892 nw
rect 435 5516 516 5568
rect 568 5516 634 5568
rect 686 5516 751 5568
rect 803 5516 823 5568
rect 435 5479 823 5516
rect 435 5465 748 5479
rect 487 5413 507 5465
rect 559 5413 579 5465
rect 631 5413 651 5465
rect 703 5427 748 5465
rect 800 5427 823 5479
rect 703 5413 823 5427
rect 435 5400 823 5413
rect 487 5348 507 5400
rect 559 5348 579 5400
rect 631 5348 651 5400
rect 703 5348 823 5400
rect 435 5335 823 5348
rect 487 5283 507 5335
rect 559 5283 579 5335
rect 631 5283 651 5335
rect 703 5283 823 5335
rect 435 5270 823 5283
rect 487 5218 507 5270
rect 559 5218 579 5270
rect 631 5218 651 5270
rect 703 5218 823 5270
rect 435 5205 823 5218
rect 487 5153 507 5205
rect 559 5153 579 5205
rect 631 5153 651 5205
rect 703 5153 823 5205
rect 435 5140 823 5153
rect 487 5088 507 5140
rect 559 5088 579 5140
rect 631 5088 651 5140
rect 703 5088 823 5140
rect 14240 5565 14652 8104
rect 14240 5513 14313 5565
rect 14365 5513 14652 5565
rect 14240 5465 14652 5513
rect 14240 5413 14243 5465
rect 14295 5413 14309 5465
rect 14361 5413 14375 5465
rect 14427 5413 14441 5465
rect 14493 5413 14652 5465
rect 14240 5400 14652 5413
rect 14240 5348 14243 5400
rect 14295 5348 14309 5400
rect 14361 5348 14375 5400
rect 14427 5348 14441 5400
rect 14493 5348 14652 5400
rect 14240 5335 14652 5348
rect 14240 5283 14243 5335
rect 14295 5283 14309 5335
rect 14361 5283 14375 5335
rect 14427 5283 14441 5335
rect 14493 5283 14652 5335
rect 14240 5270 14652 5283
rect 14240 5218 14243 5270
rect 14295 5218 14309 5270
rect 14361 5218 14375 5270
rect 14427 5218 14441 5270
rect 14493 5218 14652 5270
rect 14240 5205 14652 5218
rect 14240 5153 14243 5205
rect 14295 5153 14309 5205
rect 14361 5153 14375 5205
rect 14427 5153 14441 5205
rect 14493 5153 14652 5205
rect 14240 5140 14652 5153
rect 14240 5088 14243 5140
rect 14295 5088 14309 5140
rect 14361 5088 14375 5140
rect 14427 5088 14441 5140
rect 14493 5088 14652 5140
rect 435 5075 823 5088
rect 487 5023 507 5075
rect 559 5023 579 5075
rect 631 5023 651 5075
rect 703 5023 823 5075
rect 435 5010 823 5023
rect 487 4958 507 5010
rect 559 4958 579 5010
rect 631 4958 651 5010
rect 703 4958 823 5010
rect 435 4945 823 4958
rect 487 4893 507 4945
rect 559 4893 579 4945
rect 631 4893 651 4945
rect 703 4893 823 4945
rect 435 4880 823 4893
rect 487 4828 507 4880
rect 559 4828 579 4880
rect 631 4828 651 4880
rect 703 4828 823 4880
rect 435 4815 823 4828
rect 487 4763 507 4815
rect 559 4763 579 4815
rect 631 4763 651 4815
rect 703 4763 823 4815
rect 435 4750 823 4763
rect 487 4698 507 4750
rect 559 4698 579 4750
rect 631 4698 651 4750
rect 703 4698 823 4750
rect 435 4685 823 4698
rect 487 4633 507 4685
rect 559 4633 579 4685
rect 631 4633 651 4685
rect 703 4633 823 4685
rect 435 4620 823 4633
rect 487 4568 507 4620
rect 559 4568 579 4620
rect 631 4568 651 4620
rect 703 4568 823 4620
rect 435 4555 823 4568
rect 487 4503 507 4555
rect 559 4503 579 4555
rect 631 4503 651 4555
rect 703 4503 823 4555
rect 435 4490 823 4503
rect 487 4438 507 4490
rect 559 4438 579 4490
rect 631 4438 651 4490
rect 703 4438 823 4490
rect 435 4425 823 4438
rect 487 4373 507 4425
rect 559 4373 579 4425
rect 631 4373 651 4425
rect 703 4373 823 4425
rect 435 4360 823 4373
rect 487 4308 507 4360
rect 559 4308 579 4360
rect 631 4308 651 4360
rect 703 4308 823 4360
rect 435 4295 823 4308
rect 487 4243 507 4295
rect 559 4243 579 4295
rect 631 4243 651 4295
rect 703 4243 823 4295
rect 435 4230 823 4243
rect 487 4178 507 4230
rect 559 4178 579 4230
rect 631 4178 651 4230
rect 703 4178 823 4230
rect 435 4165 823 4178
rect 487 4113 507 4165
rect 559 4113 579 4165
rect 631 4113 651 4165
rect 703 4113 823 4165
rect 435 4099 823 4113
rect 487 4047 507 4099
rect 559 4047 579 4099
rect 631 4047 651 4099
rect 703 4047 823 4099
rect 435 4033 823 4047
rect 487 3981 507 4033
rect 559 3981 579 4033
rect 631 3981 651 4033
rect 703 3981 823 4033
rect 11116 3995 12657 5088
rect 14240 5075 14652 5088
rect 14240 5023 14243 5075
rect 14295 5023 14309 5075
rect 14361 5023 14375 5075
rect 14427 5023 14441 5075
rect 14493 5023 14652 5075
rect 14240 5010 14652 5023
rect 14240 4958 14243 5010
rect 14295 4958 14309 5010
rect 14361 4958 14375 5010
rect 14427 4958 14441 5010
rect 14493 4958 14652 5010
rect 14240 4945 14652 4958
rect 14240 4893 14243 4945
rect 14295 4893 14309 4945
rect 14361 4893 14375 4945
rect 14427 4893 14441 4945
rect 14493 4893 14652 4945
rect 14240 4880 14652 4893
rect 14240 4828 14243 4880
rect 14295 4828 14309 4880
rect 14361 4828 14375 4880
rect 14427 4828 14441 4880
rect 14493 4828 14652 4880
rect 14240 4815 14652 4828
rect 14240 4763 14243 4815
rect 14295 4763 14309 4815
rect 14361 4763 14375 4815
rect 14427 4763 14441 4815
rect 14493 4763 14652 4815
rect 14240 4750 14652 4763
rect 14240 4698 14243 4750
rect 14295 4698 14309 4750
rect 14361 4698 14375 4750
rect 14427 4698 14441 4750
rect 14493 4698 14652 4750
rect 14240 4685 14652 4698
rect 14240 4633 14243 4685
rect 14295 4633 14309 4685
rect 14361 4633 14375 4685
rect 14427 4633 14441 4685
rect 14493 4633 14652 4685
rect 14240 4620 14652 4633
rect 14240 4568 14243 4620
rect 14295 4568 14309 4620
rect 14361 4568 14375 4620
rect 14427 4568 14441 4620
rect 14493 4568 14652 4620
rect 14240 4555 14652 4568
rect 14240 4503 14243 4555
rect 14295 4503 14309 4555
rect 14361 4503 14375 4555
rect 14427 4503 14441 4555
rect 14493 4503 14652 4555
rect 14240 4490 14652 4503
rect 14240 4438 14243 4490
rect 14295 4438 14309 4490
rect 14361 4438 14375 4490
rect 14427 4438 14441 4490
rect 14493 4438 14652 4490
rect 14240 4425 14652 4438
rect 14240 4373 14243 4425
rect 14295 4373 14309 4425
rect 14361 4373 14375 4425
rect 14427 4373 14441 4425
rect 14493 4373 14652 4425
rect 14240 4359 14652 4373
rect 14240 4307 14243 4359
rect 14295 4307 14309 4359
rect 14361 4307 14375 4359
rect 14427 4307 14441 4359
rect 14493 4307 14652 4359
rect 14240 4293 14652 4307
rect 14240 4241 14243 4293
rect 14295 4241 14309 4293
rect 14361 4241 14375 4293
rect 14427 4241 14441 4293
rect 14493 4241 14652 4293
rect 14240 4227 14652 4241
rect 14240 4175 14243 4227
rect 14295 4175 14309 4227
rect 14361 4175 14375 4227
rect 14427 4175 14441 4227
rect 14493 4175 14652 4227
rect 14240 4161 14652 4175
rect 14240 4109 14243 4161
rect 14295 4109 14309 4161
rect 14361 4109 14375 4161
rect 14427 4109 14441 4161
rect 14493 4109 14652 4161
rect 14240 4095 14652 4109
rect 14240 4043 14243 4095
rect 14295 4043 14309 4095
rect 14361 4043 14375 4095
rect 14427 4043 14441 4095
rect 14493 4043 14652 4095
rect 14240 4029 14652 4043
rect 435 3967 823 3981
rect 487 3915 507 3967
rect 559 3915 579 3967
rect 631 3915 651 3967
rect 703 3915 823 3967
rect 435 3901 823 3915
rect 487 3849 507 3901
rect 559 3849 579 3901
rect 631 3849 651 3901
rect 703 3849 823 3901
rect 14240 3977 14243 4029
rect 14295 3977 14309 4029
rect 14361 3977 14375 4029
rect 14427 3977 14441 4029
rect 14493 3977 14652 4029
rect 14240 3963 14652 3977
rect 14240 3911 14243 3963
rect 14295 3911 14309 3963
rect 14361 3911 14375 3963
rect 14427 3911 14441 3963
rect 14493 3911 14652 3963
rect 14240 3897 14652 3911
tri 14234 3883 14240 3889 se
rect 14240 3883 14243 3897
rect 435 3845 823 3849
tri 823 3845 861 3883 sw
tri 14196 3845 14234 3883 se
rect 14234 3845 14243 3883
rect 14295 3845 14309 3897
rect 14361 3845 14375 3897
rect 14427 3845 14441 3897
rect 14493 3845 14652 3897
rect 435 3835 861 3845
rect 487 3783 507 3835
rect 559 3783 579 3835
rect 631 3783 651 3835
rect 703 3831 861 3835
tri 861 3831 875 3845 sw
tri 14182 3831 14196 3845 se
rect 14196 3831 14652 3845
rect 703 3783 875 3831
rect 435 3779 875 3783
tri 875 3779 927 3831 sw
tri 14130 3779 14182 3831 se
rect 14182 3779 14243 3831
rect 14295 3779 14309 3831
rect 14361 3779 14375 3831
rect 14427 3779 14441 3831
rect 14493 3779 14652 3831
rect 435 3769 927 3779
rect 487 3717 507 3769
rect 559 3717 579 3769
rect 631 3717 651 3769
rect 703 3765 927 3769
tri 927 3765 941 3779 sw
tri 14116 3765 14130 3779 se
rect 14130 3765 14652 3779
rect 703 3717 941 3765
rect 435 3713 941 3717
tri 941 3713 993 3765 sw
tri 14064 3713 14116 3765 se
rect 14116 3713 14243 3765
rect 14295 3713 14309 3765
rect 14361 3713 14375 3765
rect 14427 3713 14441 3765
rect 14493 3713 14652 3765
rect 435 3703 993 3713
rect 487 3651 507 3703
rect 559 3651 579 3703
rect 631 3651 651 3703
rect 703 3699 993 3703
tri 993 3699 1007 3713 sw
tri 14050 3699 14064 3713 se
rect 14064 3699 14652 3713
rect 703 3651 1007 3699
rect 435 3647 1007 3651
tri 1007 3647 1059 3699 sw
tri 13998 3647 14050 3699 se
rect 14050 3647 14243 3699
rect 14295 3647 14309 3699
rect 14361 3647 14375 3699
rect 14427 3647 14441 3699
rect 14493 3647 14652 3699
rect 435 3645 1059 3647
tri 1059 3645 1061 3647 sw
tri 13996 3645 13998 3647 se
rect 13998 3645 14652 3647
rect 435 3631 1061 3645
tri 1061 3631 1075 3645 sw
tri 13992 3641 13996 3645 se
rect 13996 3641 14652 3645
tri 13982 3631 13992 3641 se
rect 13992 3631 14652 3641
rect 435 2530 1090 3631
rect 14439 3628 14652 3631
rect 13300 2554 14652 3628
rect 14439 2530 14652 2554
tri 378 872 412 906 sw
rect 338 820 580 872
rect 632 820 648 872
rect 700 820 707 872
rect 338 806 707 820
rect 338 754 580 806
rect 632 754 648 806
rect 700 754 707 806
rect 338 753 707 754
rect 3710 871 3934 872
rect 3710 819 3716 871
rect 3768 819 3796 871
rect 3848 819 3876 871
rect 3928 819 3934 871
rect 3710 805 3934 819
rect 3710 753 3716 805
rect 3768 753 3796 805
rect 3848 753 3876 805
rect 3928 753 3934 805
rect 338 487 486 753
tri 486 661 578 753 nw
tri 486 487 551 552 sw
rect 3710 487 3934 753
rect 338 435 580 487
rect 632 435 648 487
rect 700 435 708 487
rect 338 421 708 435
rect 338 369 580 421
rect 632 369 648 421
rect 700 369 708 421
rect 338 368 708 369
rect 3710 435 3716 487
rect 3768 435 3796 487
rect 3848 435 3876 487
rect 3928 435 3934 487
rect 3710 421 3934 435
rect 3710 369 3716 421
rect 3768 369 3796 421
rect 3848 369 3876 421
rect 3928 369 3934 421
tri 310 135 352 177 sw
rect 3710 135 3934 369
rect 278 83 284 135
rect 336 83 348 135
rect 400 83 406 135
rect 3710 83 3716 135
rect 3768 83 3796 135
rect 3848 83 3876 135
rect 3928 83 3934 135
rect 14708 -6 14748 16057
rect 14788 -6 14828 16137
rect 14868 -6 14908 16246
rect 14948 -6 14988 16326
rect 15028 -6 15068 16406
rect 5247 -9151 5930 -9145
rect 5247 -9203 5878 -9151
rect 5247 -9223 5930 -9203
rect 5247 -9275 5878 -9223
rect 5247 -9281 5930 -9275
rect 5247 -9942 5685 -9281
tri 5685 -9474 5878 -9281 nw
rect 5247 -9994 5253 -9942
rect 5305 -9994 5328 -9942
rect 5380 -9994 5403 -9942
rect 5455 -9994 5478 -9942
rect 5530 -9994 5553 -9942
rect 5605 -9994 5627 -9942
rect 5679 -9994 5685 -9942
rect 5247 -10017 5685 -9994
rect 5247 -10069 5253 -10017
rect 5305 -10069 5328 -10017
rect 5380 -10069 5403 -10017
rect 5455 -10069 5478 -10017
rect 5530 -10069 5553 -10017
rect 5605 -10069 5627 -10017
rect 5679 -10069 5685 -10017
rect 5247 -10092 5685 -10069
rect 5247 -10144 5253 -10092
rect 5305 -10144 5328 -10092
rect 5380 -10144 5403 -10092
rect 5455 -10144 5478 -10092
rect 5530 -10144 5553 -10092
rect 5605 -10144 5627 -10092
rect 5679 -10144 5685 -10092
rect 5247 -10933 5685 -10144
rect 8191 -10933 8667 -9701
tri 8667 -10933 8773 -10827 sw
rect 5247 -10985 5253 -10933
rect 5305 -10985 5328 -10933
rect 5380 -10985 5403 -10933
rect 5455 -10985 5478 -10933
rect 5530 -10985 5553 -10933
rect 5605 -10985 5627 -10933
rect 5679 -10985 5685 -10933
rect 5247 -11011 5685 -10985
rect 5247 -11063 5253 -11011
rect 5305 -11063 5328 -11011
rect 5380 -11063 5403 -11011
rect 5455 -11063 5478 -11011
rect 5530 -11063 5553 -11011
rect 5605 -11063 5627 -11011
rect 5679 -11063 5685 -11011
<< metal3 >>
rect 4600 13425 5084 15087
rect 6107 13425 6811 15087
rect 9047 13425 9347 15087
use sky130_fd_io__com_pudrvr_strong_slowv2  sky130_fd_io__com_pudrvr_strong_slowv2_0
timestamp 1666464484
transform -1 0 7012 0 1 139
box -36 -176 3550 1143
use sky130_fd_io__com_pudrvr_weakv2  sky130_fd_io__com_pudrvr_weakv2_0
timestamp 1666464484
transform 1 0 78 0 1 139
box -36 -176 3550 1143
use sky130_fd_io__com_res_weak  sky130_fd_io__com_res_weak_0
timestamp 1666464484
transform 0 1 1833 1 0 6897
box -160 1014 679 10611
use sky130_fd_io__gpio_pddrvr_strong_slowv2  sky130_fd_io__gpio_pddrvr_strong_slowv2_0
timestamp 1666464484
transform 0 1 420 -1 0 15675
box -918 -419 1152 14752
use sky130_fd_io__gpio_pddrvr_weakv2  sky130_fd_io__gpio_pddrvr_weakv2_0
timestamp 1666464484
transform 0 1 5329 -1 0 15675
box -202 0 1152 7520
use sky130_fd_io__gpio_pudrvr_strongv2  sky130_fd_io__gpio_pudrvr_strongv2_0
timestamp 1666464484
transform 1 0 -580 0 1 622
box 467 -902 15583 5464
use sky130_fd_io__gpiov2_pddrvr_strong  sky130_fd_io__gpiov2_pddrvr_strong_0
timestamp 1666464484
transform 1 0 85 0 -1 17755
box -1000 1136 15088 31368
use sky130_fd_io__res250only_small  sky130_fd_io__res250only_small_0
timestamp 1666464484
transform -1 0 13372 0 -1 8288
box 0 0 2270 404
use sky130_fd_io__tk_em1s_cdns_5595914180852  sky130_fd_io__tk_em1s_cdns_5595914180852_0
timestamp 1666464484
transform -1 0 10237 0 -1 8259
box 0 0 1 1
use sky130_fd_pr__res_generic_po__example_5595914180853  sky130_fd_pr__res_generic_po__example_5595914180853_0
timestamp 1666464484
transform -1 0 10314 0 1 7886
box 15 31 585 32
use sky130_fd_pr__res_generic_po__example_5595914180855  sky130_fd_pr__res_generic_po__example_5595914180855_0
timestamp 1666464484
transform -1 0 9612 0 1 7886
box 15 31 985 32
use sky130_fd_pr__res_generic_po__example_5595914180856  sky130_fd_pr__res_generic_po__example_5595914180856_0
timestamp 1666464484
transform -1 0 10816 0 1 7886
box 15 31 385 32
use sky130_fd_pr__via_l1m1__example_5595914180832  sky130_fd_pr__via_l1m1__example_5595914180832_0
timestamp 1666464484
transform 1 0 8509 0 1 7932
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418080  sky130_fd_pr__via_pol1_centered__example_559591418080_0
timestamp 1666464484
transform 0 1 8561 1 0 8086
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418080  sky130_fd_pr__via_pol1_centered__example_559591418080_1
timestamp 1666464484
transform 0 -1 10867 1 0 8086
box 0 0 1 1
<< labels >>
flabel locali s 310 1322 402 1368 3 FreeSans 520 0 0 0 VGND
port 1 nsew
flabel comment s 1426 15454 1426 15454 0 FreeSans 440 0 0 0 CONDIODE
flabel comment s 6755 15452 6755 15452 0 FreeSans 440 0 0 0 CONDIODE
flabel metal2 s 14708 -6 14748 186 3 FreeSans 520 90 0 0 PD_H[0]
port 2 nsew
flabel metal2 s 14868 -6 14908 186 3 FreeSans 520 90 0 0 PD_H[2]
port 3 nsew
flabel metal2 s 14788 -6 14828 186 3 FreeSans 520 90 0 0 PD_H[1]
port 4 nsew
flabel metal2 s 14948 -6 14988 186 3 FreeSans 520 90 0 0 PD_H[3]
port 5 nsew
flabel metal2 s 13300 2554 14496 3628 3 FreeSans 520 0 0 0 VCC_IO
port 6 nsew
flabel metal2 s 11116 3995 12657 5088 3 FreeSans 520 0 0 0 PAD
port 7 nsew
flabel metal2 s 11116 10850 12657 11943 3 FreeSans 520 0 0 0 PAD
port 7 nsew
flabel metal2 s 15028 -6 15068 186 3 FreeSans 520 90 0 0 TIE_LO_ESD
port 8 nsew
flabel metal1 s 49 -1067 83 -1013 3 FreeSans 520 270 0 0 FORCE_HI_H_N
port 9 nsew
flabel metal1 s 377 -1075 415 -1020 3 FreeSans 520 270 0 0 FORCE_LO_H
port 10 nsew
flabel metal1 s 258 -1075 313 -1023 3 FreeSans 520 270 0 0 FORCE_LOVOL_H
port 11 nsew
flabel metal1 s 761 683 794 715 3 FreeSans 520 0 0 0 PU_H_N[0]
port 12 nsew
flabel metal1 s 6527 686 6583 719 3 FreeSans 520 0 0 0 PU_H_N[1]
port 13 nsew
flabel metal1 s 14167 280 14252 332 3 FreeSans 520 0 0 0 PU_H_N[2]
port 14 nsew
flabel metal1 s 13921 168 14073 220 3 FreeSans 520 0 0 0 PU_H_N[3]
port 15 nsew
flabel metal1 s 167 -1074 205 -1007 3 FreeSans 520 270 0 0 VSSIO_AMX
port 16 nsew
flabel metal1 s 2496 8314 2549 8360 3 FreeSans 520 0 0 0 VGND_IO
port 17 nsew
flabel metal1 s 14164 88 14240 140 3 FreeSans 520 0 0 0 TIE_HI_ESD
port 18 nsew
flabel metal1 s 13310 7924 13365 8257 3 FreeSans 520 0 0 0 PAD
port 7 nsew
flabel metal1 s 11799 736 11831 794 3 FreeSans 520 0 0 0 VCC_IO
port 6 nsew
flabel metal1 s 451 932 1620 1077 3 FreeSans 520 0 0 0 VCC_IO
port 6 nsew
flabel metal1 s 3948 909 5117 955 3 FreeSans 520 0 0 0 VCC_IO
port 6 nsew
<< properties >>
string GDS_END 48364804
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 47456218
<< end >>
