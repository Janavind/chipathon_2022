magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -66 377 1506 897
<< pwell >>
rect 53 43 1433 317
rect -26 -43 1466 43
<< mvnmos >>
rect 132 141 232 291
rect 288 141 388 291
rect 444 141 544 291
rect 600 141 700 291
rect 756 141 856 291
rect 912 141 1012 291
rect 1096 141 1196 291
rect 1252 141 1352 291
<< mvpmos >>
rect 160 443 260 743
rect 316 443 416 743
rect 472 443 572 743
rect 628 443 728 743
rect 784 443 884 743
rect 940 443 1040 743
rect 1096 443 1196 743
rect 1252 443 1352 743
<< mvndiff >>
rect 79 273 132 291
rect 79 239 87 273
rect 121 239 132 273
rect 79 205 132 239
rect 79 171 87 205
rect 121 171 132 205
rect 79 141 132 171
rect 232 264 288 291
rect 232 230 243 264
rect 277 230 288 264
rect 232 196 288 230
rect 232 162 243 196
rect 277 162 288 196
rect 232 141 288 162
rect 388 205 444 291
rect 388 171 399 205
rect 433 171 444 205
rect 388 141 444 171
rect 544 264 600 291
rect 544 230 555 264
rect 589 230 600 264
rect 544 196 600 230
rect 544 162 555 196
rect 589 162 600 196
rect 544 141 600 162
rect 700 205 756 291
rect 700 171 711 205
rect 745 171 756 205
rect 700 141 756 171
rect 856 264 912 291
rect 856 230 867 264
rect 901 230 912 264
rect 856 196 912 230
rect 856 162 867 196
rect 901 162 912 196
rect 856 141 912 162
rect 1012 205 1096 291
rect 1012 171 1023 205
rect 1057 171 1096 205
rect 1012 141 1096 171
rect 1196 264 1252 291
rect 1196 230 1207 264
rect 1241 230 1252 264
rect 1196 196 1252 230
rect 1196 162 1207 196
rect 1241 162 1252 196
rect 1196 141 1252 162
rect 1352 205 1407 291
rect 1352 171 1365 205
rect 1399 171 1407 205
rect 1352 141 1407 171
<< mvpdiff >>
rect 107 731 160 743
rect 107 697 115 731
rect 149 697 160 731
rect 107 663 160 697
rect 107 629 115 663
rect 149 629 160 663
rect 107 595 160 629
rect 107 561 115 595
rect 149 561 160 595
rect 107 527 160 561
rect 107 493 115 527
rect 149 493 160 527
rect 107 443 160 493
rect 260 689 316 743
rect 260 655 271 689
rect 305 655 316 689
rect 260 621 316 655
rect 260 587 271 621
rect 305 587 316 621
rect 260 553 316 587
rect 260 519 271 553
rect 305 519 316 553
rect 260 485 316 519
rect 260 451 271 485
rect 305 451 316 485
rect 260 443 316 451
rect 416 731 472 743
rect 416 697 427 731
rect 461 697 472 731
rect 416 663 472 697
rect 416 629 427 663
rect 461 629 472 663
rect 416 595 472 629
rect 416 561 427 595
rect 461 561 472 595
rect 416 527 472 561
rect 416 493 427 527
rect 461 493 472 527
rect 416 443 472 493
rect 572 689 628 743
rect 572 655 583 689
rect 617 655 628 689
rect 572 621 628 655
rect 572 587 583 621
rect 617 587 628 621
rect 572 553 628 587
rect 572 519 583 553
rect 617 519 628 553
rect 572 485 628 519
rect 572 451 583 485
rect 617 451 628 485
rect 572 443 628 451
rect 728 731 784 743
rect 728 697 739 731
rect 773 697 784 731
rect 728 663 784 697
rect 728 629 739 663
rect 773 629 784 663
rect 728 595 784 629
rect 728 561 739 595
rect 773 561 784 595
rect 728 527 784 561
rect 728 493 739 527
rect 773 493 784 527
rect 728 443 784 493
rect 884 689 940 743
rect 884 655 895 689
rect 929 655 940 689
rect 884 621 940 655
rect 884 587 895 621
rect 929 587 940 621
rect 884 553 940 587
rect 884 519 895 553
rect 929 519 940 553
rect 884 485 940 519
rect 884 451 895 485
rect 929 451 940 485
rect 884 443 940 451
rect 1040 731 1096 743
rect 1040 697 1051 731
rect 1085 697 1096 731
rect 1040 663 1096 697
rect 1040 629 1051 663
rect 1085 629 1096 663
rect 1040 595 1096 629
rect 1040 561 1051 595
rect 1085 561 1096 595
rect 1040 527 1096 561
rect 1040 493 1051 527
rect 1085 493 1096 527
rect 1040 443 1096 493
rect 1196 689 1252 743
rect 1196 655 1207 689
rect 1241 655 1252 689
rect 1196 621 1252 655
rect 1196 587 1207 621
rect 1241 587 1252 621
rect 1196 553 1252 587
rect 1196 519 1207 553
rect 1241 519 1252 553
rect 1196 485 1252 519
rect 1196 451 1207 485
rect 1241 451 1252 485
rect 1196 443 1252 451
rect 1352 731 1405 743
rect 1352 697 1363 731
rect 1397 697 1405 731
rect 1352 663 1405 697
rect 1352 629 1363 663
rect 1397 629 1405 663
rect 1352 595 1405 629
rect 1352 561 1363 595
rect 1397 561 1405 595
rect 1352 527 1405 561
rect 1352 493 1363 527
rect 1397 493 1405 527
rect 1352 443 1405 493
<< mvndiffc >>
rect 87 239 121 273
rect 87 171 121 205
rect 243 230 277 264
rect 243 162 277 196
rect 399 171 433 205
rect 555 230 589 264
rect 555 162 589 196
rect 711 171 745 205
rect 867 230 901 264
rect 867 162 901 196
rect 1023 171 1057 205
rect 1207 230 1241 264
rect 1207 162 1241 196
rect 1365 171 1399 205
<< mvpdiffc >>
rect 115 697 149 731
rect 115 629 149 663
rect 115 561 149 595
rect 115 493 149 527
rect 271 655 305 689
rect 271 587 305 621
rect 271 519 305 553
rect 271 451 305 485
rect 427 697 461 731
rect 427 629 461 663
rect 427 561 461 595
rect 427 493 461 527
rect 583 655 617 689
rect 583 587 617 621
rect 583 519 617 553
rect 583 451 617 485
rect 739 697 773 731
rect 739 629 773 663
rect 739 561 773 595
rect 739 493 773 527
rect 895 655 929 689
rect 895 587 929 621
rect 895 519 929 553
rect 895 451 929 485
rect 1051 697 1085 731
rect 1051 629 1085 663
rect 1051 561 1085 595
rect 1051 493 1085 527
rect 1207 655 1241 689
rect 1207 587 1241 621
rect 1207 519 1241 553
rect 1207 451 1241 485
rect 1363 697 1397 731
rect 1363 629 1397 663
rect 1363 561 1397 595
rect 1363 493 1397 527
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1440 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
<< poly >>
rect 160 743 260 769
rect 316 743 416 769
rect 472 743 572 769
rect 628 743 728 769
rect 784 743 884 769
rect 940 743 1040 769
rect 1096 743 1196 769
rect 1252 743 1352 769
rect 160 413 260 443
rect 316 413 416 443
rect 472 413 572 443
rect 628 413 728 443
rect 784 413 884 443
rect 940 413 1040 443
rect 1096 413 1196 443
rect 1252 413 1352 443
rect 62 363 1352 413
rect 62 329 78 363
rect 112 329 146 363
rect 180 329 214 363
rect 248 329 282 363
rect 316 329 350 363
rect 384 329 418 363
rect 452 329 486 363
rect 520 329 554 363
rect 588 329 622 363
rect 656 329 690 363
rect 724 329 758 363
rect 792 329 826 363
rect 860 329 894 363
rect 928 329 962 363
rect 996 329 1030 363
rect 1064 329 1098 363
rect 1132 329 1166 363
rect 1200 329 1234 363
rect 1268 329 1302 363
rect 1336 329 1352 363
rect 62 313 1352 329
rect 132 291 232 313
rect 288 291 388 313
rect 444 291 544 313
rect 600 291 700 313
rect 756 291 856 313
rect 912 291 1012 313
rect 1096 291 1196 313
rect 1252 291 1352 313
rect 132 115 232 141
rect 288 115 388 141
rect 444 115 544 141
rect 600 115 700 141
rect 756 115 856 141
rect 912 115 1012 141
rect 1096 115 1196 141
rect 1252 115 1352 141
<< polycont >>
rect 78 329 112 363
rect 146 329 180 363
rect 214 329 248 363
rect 282 329 316 363
rect 350 329 384 363
rect 418 329 452 363
rect 486 329 520 363
rect 554 329 588 363
rect 622 329 656 363
rect 690 329 724 363
rect 758 329 792 363
rect 826 329 860 363
rect 894 329 928 363
rect 962 329 996 363
rect 1030 329 1064 363
rect 1098 329 1132 363
rect 1166 329 1200 363
rect 1234 329 1268 363
rect 1302 329 1336 363
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1440 831
rect 19 731 1405 759
rect 19 729 115 731
rect 149 729 427 731
rect 461 729 739 731
rect 773 729 1051 731
rect 1085 729 1363 731
rect 1397 729 1405 731
rect 53 695 91 729
rect 149 697 163 729
rect 125 695 163 697
rect 197 725 355 729
rect 19 663 197 695
rect 389 695 427 729
rect 461 695 499 729
rect 533 725 667 729
rect 19 629 115 663
rect 149 629 197 663
rect 19 595 197 629
rect 19 561 115 595
rect 149 561 197 595
rect 19 527 197 561
rect 19 493 115 527
rect 149 493 197 527
rect 19 489 197 493
rect 255 655 271 689
rect 305 655 321 689
rect 255 621 321 655
rect 255 587 271 621
rect 305 587 321 621
rect 255 553 321 587
rect 255 519 271 553
rect 305 519 321 553
rect 255 485 321 519
rect 255 451 271 485
rect 305 451 321 485
rect 355 663 533 695
rect 701 695 739 729
rect 773 695 811 729
rect 845 725 979 729
rect 355 629 427 663
rect 461 629 533 663
rect 355 595 533 629
rect 355 561 427 595
rect 461 561 533 595
rect 355 527 533 561
rect 355 493 427 527
rect 461 493 533 527
rect 355 477 533 493
rect 567 655 583 689
rect 617 655 633 689
rect 567 621 633 655
rect 567 587 583 621
rect 617 587 633 621
rect 567 553 633 587
rect 567 519 583 553
rect 617 519 633 553
rect 567 485 633 519
rect 255 441 321 451
rect 567 451 583 485
rect 617 451 633 485
rect 667 663 845 695
rect 1013 695 1051 729
rect 1085 695 1123 729
rect 1157 725 1291 729
rect 667 629 739 663
rect 773 629 845 663
rect 667 595 845 629
rect 667 561 739 595
rect 773 561 845 595
rect 667 527 845 561
rect 667 493 739 527
rect 773 493 845 527
rect 667 477 845 493
rect 879 655 895 689
rect 929 655 945 689
rect 879 621 945 655
rect 879 587 895 621
rect 929 587 945 621
rect 879 553 945 587
rect 879 519 895 553
rect 929 519 945 553
rect 879 485 945 519
rect 567 441 633 451
rect 879 451 895 485
rect 929 451 945 485
rect 979 663 1157 695
rect 1325 697 1363 729
rect 1325 695 1371 697
rect 979 629 1051 663
rect 1085 629 1157 663
rect 979 595 1157 629
rect 979 561 1051 595
rect 1085 561 1157 595
rect 979 527 1157 561
rect 979 493 1051 527
rect 1085 493 1157 527
rect 979 477 1157 493
rect 1191 655 1207 689
rect 1241 655 1257 689
rect 1191 621 1257 655
rect 1191 587 1207 621
rect 1241 587 1257 621
rect 1191 553 1257 587
rect 1191 519 1207 553
rect 1241 519 1257 553
rect 1191 485 1257 519
rect 879 441 945 451
rect 1191 451 1207 485
rect 1241 451 1257 485
rect 1291 663 1405 695
rect 1291 629 1363 663
rect 1397 629 1405 663
rect 1291 595 1405 629
rect 1291 561 1363 595
rect 1397 561 1405 595
rect 1291 527 1405 561
rect 1291 493 1363 527
rect 1397 493 1405 527
rect 1291 477 1405 493
rect 1191 441 1257 451
rect 255 407 1422 441
rect 62 329 78 363
rect 112 329 146 363
rect 180 329 214 363
rect 248 329 282 363
rect 316 329 350 363
rect 384 329 418 363
rect 452 329 486 363
rect 520 329 554 363
rect 588 329 622 363
rect 656 329 690 363
rect 724 329 758 363
rect 792 329 826 363
rect 860 329 894 363
rect 928 329 962 363
rect 996 329 1030 363
rect 1064 329 1098 363
rect 1132 329 1166 363
rect 1200 329 1234 363
rect 1268 329 1302 363
rect 1336 329 1352 363
rect 62 316 1352 329
rect 239 279 1245 280
rect 1388 279 1422 407
rect 19 273 197 277
rect 19 239 87 273
rect 121 239 197 273
rect 19 205 197 239
rect 19 171 87 205
rect 121 171 197 205
rect 19 110 197 171
rect 239 264 1422 279
rect 239 230 243 264
rect 277 246 555 264
rect 277 230 281 246
rect 239 196 281 230
rect 551 230 555 246
rect 589 246 867 264
rect 589 230 593 246
rect 239 162 243 196
rect 277 162 281 196
rect 239 146 281 162
rect 315 205 517 209
rect 315 171 399 205
rect 433 171 517 205
rect 315 110 517 171
rect 551 196 593 230
rect 863 230 867 246
rect 901 246 1207 264
rect 901 230 905 246
rect 551 162 555 196
rect 589 162 593 196
rect 551 146 593 162
rect 627 205 829 209
rect 627 171 711 205
rect 745 171 829 205
rect 627 110 829 171
rect 863 196 905 230
rect 1183 230 1207 246
rect 1241 245 1422 264
rect 1241 230 1313 245
rect 863 162 867 196
rect 901 162 905 196
rect 863 146 905 162
rect 939 205 1149 209
rect 939 171 1023 205
rect 1057 171 1149 205
rect 939 110 1149 171
rect 1183 196 1313 230
rect 1183 162 1207 196
rect 1241 162 1313 196
rect 1183 146 1313 162
rect 1347 205 1421 209
rect 1347 171 1365 205
rect 1399 171 1421 205
rect 1347 110 1421 171
rect 53 76 91 110
rect 125 76 163 110
rect 197 76 235 110
rect 269 76 307 110
rect 341 76 379 110
rect 413 76 451 110
rect 485 76 523 110
rect 557 76 595 110
rect 629 76 667 110
rect 701 76 739 110
rect 773 76 811 110
rect 845 76 883 110
rect 917 76 955 110
rect 989 76 1027 110
rect 1061 76 1099 110
rect 1133 76 1171 110
rect 1205 76 1243 110
rect 1277 76 1315 110
rect 1349 76 1387 110
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 19 695 53 729
rect 91 697 115 729
rect 115 697 125 729
rect 91 695 125 697
rect 163 695 197 729
rect 355 695 389 729
rect 427 697 461 729
rect 427 695 461 697
rect 499 695 533 729
rect 667 695 701 729
rect 739 697 773 729
rect 739 695 773 697
rect 811 695 845 729
rect 979 695 1013 729
rect 1051 697 1085 729
rect 1051 695 1085 697
rect 1123 695 1157 729
rect 1291 695 1325 729
rect 1371 697 1397 729
rect 1397 697 1405 729
rect 1371 695 1405 697
rect 19 76 53 110
rect 91 76 125 110
rect 163 76 197 110
rect 235 76 269 110
rect 307 76 341 110
rect 379 76 413 110
rect 451 76 485 110
rect 523 76 557 110
rect 595 76 629 110
rect 667 76 701 110
rect 739 76 773 110
rect 811 76 845 110
rect 883 76 917 110
rect 955 76 989 110
rect 1027 76 1061 110
rect 1099 76 1133 110
rect 1171 76 1205 110
rect 1243 76 1277 110
rect 1315 76 1349 110
rect 1387 76 1421 110
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 831 1440 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1440 831
rect 0 791 1440 797
rect 0 729 1440 763
rect 0 695 19 729
rect 53 695 91 729
rect 125 695 163 729
rect 197 695 355 729
rect 389 695 427 729
rect 461 695 499 729
rect 533 695 667 729
rect 701 695 739 729
rect 773 695 811 729
rect 845 695 979 729
rect 1013 695 1051 729
rect 1085 695 1123 729
rect 1157 695 1291 729
rect 1325 695 1371 729
rect 1405 695 1440 729
rect 0 689 1440 695
rect 0 110 1440 125
rect 0 76 19 110
rect 53 76 91 110
rect 125 76 163 110
rect 197 76 235 110
rect 269 76 307 110
rect 341 76 379 110
rect 413 76 451 110
rect 485 76 523 110
rect 557 76 595 110
rect 629 76 667 110
rect 701 76 739 110
rect 773 76 811 110
rect 845 76 883 110
rect 917 76 955 110
rect 989 76 1027 110
rect 1061 76 1099 110
rect 1133 76 1171 110
rect 1205 76 1243 110
rect 1277 76 1315 110
rect 1349 76 1387 110
rect 1421 76 1440 110
rect 0 51 1440 76
rect 0 17 1440 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -23 1440 -17
<< labels >>
rlabel comment s 0 0 0 0 4 inv_8
flabel metal1 s 0 0 1440 23 0 FreeSans 340 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 0 51 1440 125 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 720 11 720 11 0 FreeSans 340 0 0 0 VNB
port 3 nsew
flabel metal1 s 0 689 1440 763 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 791 1440 814 0 FreeSans 340 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 720 802 720 802 0 FreeSans 340 0 0 0 VPB
port 4 nsew
flabel locali s 1183 168 1217 202 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 1279 168 1313 202 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1440 814
string GDS_END 59604
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 42586
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
