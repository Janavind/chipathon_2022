magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 825 203
rect 29 -17 63 21
rect 397 -17 431 21
<< locali >>
rect 27 324 78 492
rect 27 51 93 324
rect 303 258 344 493
rect 258 210 344 258
rect 378 210 444 493
rect 480 199 536 493
rect 581 199 658 265
rect 702 205 802 258
rect 597 169 658 199
rect 597 57 708 169
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 113 363 179 527
rect 227 329 269 492
rect 139 293 269 329
rect 139 165 183 293
rect 572 333 629 492
rect 665 367 708 527
rect 744 333 798 492
rect 572 299 798 333
rect 139 131 561 165
rect 139 130 383 131
rect 127 17 262 94
rect 317 52 383 130
rect 417 17 486 97
rect 520 52 561 131
rect 743 17 791 152
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 597 57 708 169 6 A1
port 1 nsew signal input
rlabel locali s 597 169 658 199 6 A1
port 1 nsew signal input
rlabel locali s 581 199 658 265 6 A1
port 1 nsew signal input
rlabel locali s 702 205 802 258 6 A2
port 2 nsew signal input
rlabel locali s 480 199 536 493 6 B1
port 3 nsew signal input
rlabel locali s 378 210 444 493 6 C1
port 4 nsew signal input
rlabel locali s 258 210 344 258 6 D1
port 5 nsew signal input
rlabel locali s 303 258 344 493 6 D1
port 5 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 397 -17 431 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 29 -17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 825 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 27 51 93 324 6 X
port 10 nsew signal output
rlabel locali s 27 324 78 492 6 X
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3761534
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3752842
<< end >>
