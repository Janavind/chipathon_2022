magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 273 157 556 203
rect 1 21 556 157
rect 28 -17 62 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 93 381 177
rect 448 47 478 177
<< scpmoshvt >>
rect 79 413 109 497
rect 163 413 193 497
rect 353 341 383 425
rect 448 297 478 497
<< ndiff >>
rect 299 165 351 177
rect 299 131 307 165
rect 341 131 351 165
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 93 245 131
rect 299 93 351 131
rect 381 93 448 177
rect 193 59 203 93
rect 237 59 245 93
rect 193 47 245 59
rect 396 59 404 93
rect 438 59 448 93
rect 396 47 448 59
rect 478 119 530 177
rect 478 85 488 119
rect 522 85 530 119
rect 478 47 530 85
<< pdiff >>
rect 27 459 79 497
rect 27 425 35 459
rect 69 425 79 459
rect 27 413 79 425
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 413 163 451
rect 193 485 245 497
rect 193 451 203 485
rect 237 451 245 485
rect 193 413 245 451
rect 398 425 448 497
rect 301 387 353 425
rect 301 353 309 387
rect 343 353 353 387
rect 301 341 353 353
rect 383 417 448 425
rect 383 383 404 417
rect 438 383 448 417
rect 383 341 448 383
rect 398 297 448 341
rect 478 459 530 497
rect 478 425 488 459
rect 522 425 530 459
rect 478 391 530 425
rect 478 357 488 391
rect 522 357 530 391
rect 478 297 530 357
<< ndiffc >>
rect 307 131 341 165
rect 35 85 69 119
rect 119 59 153 93
rect 203 59 237 93
rect 404 59 438 93
rect 488 85 522 119
<< pdiffc >>
rect 35 425 69 459
rect 119 451 153 485
rect 203 451 237 485
rect 309 353 343 387
rect 404 383 438 417
rect 488 425 522 459
rect 488 357 522 391
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 353 425 383 523
rect 448 497 478 523
rect 79 265 109 413
rect 163 265 193 413
rect 353 265 383 341
rect 448 265 478 297
rect 35 249 109 265
rect 35 215 45 249
rect 79 215 109 249
rect 35 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 293 249 386 265
rect 293 215 309 249
rect 343 215 386 249
rect 293 199 386 215
rect 428 249 488 265
rect 428 215 438 249
rect 472 215 488 249
rect 428 199 488 215
rect 79 131 109 199
rect 163 131 193 199
rect 351 177 381 199
rect 448 177 478 199
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 93
rect 448 21 478 47
<< polycont >>
rect 45 215 79 249
rect 161 215 195 249
rect 309 215 343 249
rect 438 215 472 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 459 76 493
rect 17 425 35 459
rect 69 425 76 459
rect 110 485 153 527
rect 110 451 119 485
rect 110 435 153 451
rect 187 485 264 493
rect 187 451 203 485
rect 237 451 264 485
rect 187 435 264 451
rect 17 401 76 425
rect 17 357 179 401
rect 17 249 111 323
rect 17 215 45 249
rect 79 215 111 249
rect 17 211 111 215
rect 145 265 179 357
rect 145 249 196 265
rect 145 215 161 249
rect 195 215 196 249
rect 145 199 196 215
rect 230 255 264 435
rect 303 387 348 486
rect 303 353 309 387
rect 343 353 348 387
rect 382 417 454 527
rect 382 383 404 417
rect 438 383 454 417
rect 488 459 540 493
rect 522 425 540 459
rect 488 391 540 425
rect 303 349 348 353
rect 522 357 540 391
rect 303 315 448 349
rect 414 265 448 315
rect 488 299 540 357
rect 230 249 380 255
rect 230 215 309 249
rect 343 215 380 249
rect 414 249 472 265
rect 414 215 438 249
rect 145 177 179 199
rect 19 143 179 177
rect 19 119 76 143
rect 19 85 35 119
rect 69 85 76 119
rect 230 109 264 215
rect 414 199 472 215
rect 414 181 448 199
rect 19 51 76 85
rect 110 93 153 109
rect 110 59 119 93
rect 110 17 153 59
rect 187 93 264 109
rect 187 59 203 93
rect 237 59 264 93
rect 187 51 264 59
rect 303 165 448 181
rect 506 165 540 299
rect 303 131 307 165
rect 341 147 448 165
rect 341 131 348 147
rect 303 51 348 131
rect 482 119 540 165
rect 382 93 448 113
rect 382 59 404 93
rect 438 59 448 93
rect 382 17 448 59
rect 482 85 488 119
rect 522 85 540 119
rect 482 51 540 85
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 28 289 62 323 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 493 425 527 459 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 493 357 527 391 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 493 85 527 119 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 28 221 62 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel metal1 s 28 527 62 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 28 -17 62 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel nwell s 28 527 62 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 28 -17 62 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 dlygate4sd1_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 2897510
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2892108
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 16.100 13.600 
<< end >>
