magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< locali >>
rect 400 1369 962 1388
rect 400 1263 412 1369
rect 950 1263 962 1369
rect 400 1251 962 1263
rect 400 125 962 137
rect 400 19 412 125
rect 950 19 962 125
rect 400 0 962 19
<< viali >>
rect 412 1263 950 1369
rect 412 19 950 125
<< obsli1 >>
rect 190 1225 256 1291
rect 1106 1225 1172 1291
rect 190 1203 230 1225
rect 1132 1203 1172 1225
rect 41 1179 230 1203
rect 41 1145 60 1179
rect 94 1145 230 1179
rect 41 1107 230 1145
rect 41 1073 60 1107
rect 94 1073 230 1107
rect 41 1035 230 1073
rect 41 1001 60 1035
rect 94 1001 230 1035
rect 41 963 230 1001
rect 41 929 60 963
rect 94 929 230 963
rect 41 891 230 929
rect 41 857 60 891
rect 94 857 230 891
rect 41 819 230 857
rect 41 785 60 819
rect 94 785 230 819
rect 41 747 230 785
rect 41 713 60 747
rect 94 713 230 747
rect 41 675 230 713
rect 41 641 60 675
rect 94 641 230 675
rect 41 603 230 641
rect 41 569 60 603
rect 94 569 230 603
rect 41 531 230 569
rect 41 497 60 531
rect 94 497 230 531
rect 41 459 230 497
rect 41 425 60 459
rect 94 425 230 459
rect 41 387 230 425
rect 41 353 60 387
rect 94 353 230 387
rect 41 315 230 353
rect 41 281 60 315
rect 94 281 230 315
rect 41 243 230 281
rect 41 209 60 243
rect 94 209 230 243
rect 41 185 230 209
rect 352 185 386 1203
rect 508 185 542 1203
rect 664 185 698 1203
rect 820 185 854 1203
rect 976 185 1010 1203
rect 1132 1179 1321 1203
rect 1132 1145 1268 1179
rect 1302 1145 1321 1179
rect 1132 1107 1321 1145
rect 1132 1073 1268 1107
rect 1302 1073 1321 1107
rect 1132 1035 1321 1073
rect 1132 1001 1268 1035
rect 1302 1001 1321 1035
rect 1132 963 1321 1001
rect 1132 929 1268 963
rect 1302 929 1321 963
rect 1132 891 1321 929
rect 1132 857 1268 891
rect 1302 857 1321 891
rect 1132 819 1321 857
rect 1132 785 1268 819
rect 1302 785 1321 819
rect 1132 747 1321 785
rect 1132 713 1268 747
rect 1302 713 1321 747
rect 1132 675 1321 713
rect 1132 641 1268 675
rect 1302 641 1321 675
rect 1132 603 1321 641
rect 1132 569 1268 603
rect 1302 569 1321 603
rect 1132 531 1321 569
rect 1132 497 1268 531
rect 1302 497 1321 531
rect 1132 459 1321 497
rect 1132 425 1268 459
rect 1302 425 1321 459
rect 1132 387 1321 425
rect 1132 353 1268 387
rect 1302 353 1321 387
rect 1132 315 1321 353
rect 1132 281 1268 315
rect 1302 281 1321 315
rect 1132 243 1321 281
rect 1132 209 1268 243
rect 1302 209 1321 243
rect 1132 185 1321 209
rect 190 163 230 185
rect 1132 163 1172 185
rect 190 97 256 163
rect 1106 97 1172 163
<< obsli1c >>
rect 60 1145 94 1179
rect 60 1073 94 1107
rect 60 1001 94 1035
rect 60 929 94 963
rect 60 857 94 891
rect 60 785 94 819
rect 60 713 94 747
rect 60 641 94 675
rect 60 569 94 603
rect 60 497 94 531
rect 60 425 94 459
rect 60 353 94 387
rect 60 281 94 315
rect 60 209 94 243
rect 1268 1145 1302 1179
rect 1268 1073 1302 1107
rect 1268 1001 1302 1035
rect 1268 929 1302 963
rect 1268 857 1302 891
rect 1268 785 1302 819
rect 1268 713 1302 747
rect 1268 641 1302 675
rect 1268 569 1302 603
rect 1268 497 1302 531
rect 1268 425 1302 459
rect 1268 353 1302 387
rect 1268 281 1302 315
rect 1268 209 1302 243
<< metal1 >>
rect 400 1369 962 1388
rect 400 1263 412 1369
rect 950 1263 962 1369
rect 400 1251 962 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 1262 1179 1321 1191
rect 1262 1145 1268 1179
rect 1302 1145 1321 1179
rect 1262 1107 1321 1145
rect 1262 1073 1268 1107
rect 1302 1073 1321 1107
rect 1262 1035 1321 1073
rect 1262 1001 1268 1035
rect 1302 1001 1321 1035
rect 1262 963 1321 1001
rect 1262 929 1268 963
rect 1302 929 1321 963
rect 1262 891 1321 929
rect 1262 857 1268 891
rect 1302 857 1321 891
rect 1262 819 1321 857
rect 1262 785 1268 819
rect 1302 785 1321 819
rect 1262 747 1321 785
rect 1262 713 1268 747
rect 1302 713 1321 747
rect 1262 675 1321 713
rect 1262 641 1268 675
rect 1302 641 1321 675
rect 1262 603 1321 641
rect 1262 569 1268 603
rect 1302 569 1321 603
rect 1262 531 1321 569
rect 1262 497 1268 531
rect 1302 497 1321 531
rect 1262 459 1321 497
rect 1262 425 1268 459
rect 1302 425 1321 459
rect 1262 387 1321 425
rect 1262 353 1268 387
rect 1302 353 1321 387
rect 1262 315 1321 353
rect 1262 281 1268 315
rect 1302 281 1321 315
rect 1262 243 1321 281
rect 1262 209 1268 243
rect 1302 209 1321 243
rect 1262 197 1321 209
rect 400 125 962 137
rect 400 19 412 125
rect 950 19 962 125
rect 400 0 962 19
<< obsm1 >>
rect 343 197 395 1191
rect 499 197 551 1191
rect 655 197 707 1191
rect 811 197 863 1191
rect 967 197 1019 1191
<< metal2 >>
rect 14 719 1348 1191
rect 14 197 1348 669
<< labels >>
rlabel metal2 s 14 719 1348 1191 6 DRAIN
port 1 nsew
rlabel viali s 412 1263 950 1369 6 GATE
port 2 nsew
rlabel viali s 412 19 950 125 6 GATE
port 2 nsew
rlabel locali s 400 1251 962 1388 6 GATE
port 2 nsew
rlabel locali s 400 0 962 137 6 GATE
port 2 nsew
rlabel metal1 s 400 1251 962 1388 6 GATE
port 2 nsew
rlabel metal1 s 400 0 962 137 6 GATE
port 2 nsew
rlabel metal2 s 14 197 1348 669 6 SOURCE
port 3 nsew
rlabel metal1 s 41 197 100 1191 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 1262 197 1321 1191 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 1348 1388
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8516152
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8485750
string device primitive
<< end >>
