magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -66 1201 102 1251
rect -66 419 1204 1201
rect -66 377 102 419
rect 1778 409 2142 1219
<< pwell >>
rect -26 1585 2810 1671
rect 162 1267 888 1585
rect 1819 1303 2029 1585
rect 162 309 746 359
rect 162 43 914 309
rect 1264 239 1718 1291
rect 1891 43 2101 325
rect -26 -43 2810 43
<< scnmos >>
rect 1902 1329 1932 1477
rect 1988 151 2018 299
<< scpmoshvt >>
rect 1904 959 1934 1183
rect 1986 445 2016 669
<< mvnmos >>
rect 241 1293 341 1493
rect 397 1293 497 1493
rect 553 1293 653 1493
rect 709 1293 809 1493
rect 241 183 341 333
rect 507 133 667 333
rect 735 133 835 283
rect 1343 265 1463 1265
rect 1519 265 1639 1265
<< mvpmos >>
rect 229 993 629 1077
rect 685 993 1085 1077
rect 241 485 341 635
rect 735 485 835 785
<< ndiff >>
rect 1845 1465 1902 1477
rect 1845 1431 1857 1465
rect 1891 1431 1902 1465
rect 1845 1375 1902 1431
rect 1845 1341 1857 1375
rect 1891 1341 1902 1375
rect 1845 1329 1902 1341
rect 1932 1465 2003 1477
rect 1932 1431 1957 1465
rect 1991 1431 2003 1465
rect 1932 1375 2003 1431
rect 1932 1341 1957 1375
rect 1991 1341 2003 1375
rect 1932 1329 2003 1341
rect 1917 287 1988 299
rect 1917 253 1929 287
rect 1963 253 1988 287
rect 1917 197 1988 253
rect 1917 163 1929 197
rect 1963 163 1988 197
rect 1917 151 1988 163
rect 2018 287 2075 299
rect 2018 253 2029 287
rect 2063 253 2075 287
rect 2018 197 2075 253
rect 2018 163 2029 197
rect 2063 163 2075 197
rect 2018 151 2075 163
<< pdiff >>
rect 1845 1171 1904 1183
rect 1845 1137 1857 1171
rect 1891 1137 1904 1171
rect 1845 1088 1904 1137
rect 1845 1054 1857 1088
rect 1891 1054 1904 1088
rect 1845 1005 1904 1054
rect 1845 971 1857 1005
rect 1891 971 1904 1005
rect 1845 959 1904 971
rect 1934 1145 2003 1183
rect 1934 1111 1957 1145
rect 1991 1111 2003 1145
rect 1934 1075 2003 1111
rect 1934 1041 1957 1075
rect 1991 1041 2003 1075
rect 1934 1005 2003 1041
rect 1934 971 1957 1005
rect 1991 971 2003 1005
rect 1934 959 2003 971
rect 1917 657 1986 669
rect 1917 623 1929 657
rect 1963 623 1986 657
rect 1917 587 1986 623
rect 1917 553 1929 587
rect 1963 553 1986 587
rect 1917 517 1986 553
rect 1917 483 1929 517
rect 1963 483 1986 517
rect 1917 445 1986 483
rect 2016 657 2075 669
rect 2016 623 2029 657
rect 2063 623 2075 657
rect 2016 574 2075 623
rect 2016 540 2029 574
rect 2063 540 2075 574
rect 2016 491 2075 540
rect 2016 457 2029 491
rect 2063 457 2075 491
rect 2016 445 2075 457
<< mvndiff >>
rect 188 1475 241 1493
rect 188 1441 196 1475
rect 230 1441 241 1475
rect 188 1407 241 1441
rect 188 1373 196 1407
rect 230 1373 241 1407
rect 188 1339 241 1373
rect 188 1305 196 1339
rect 230 1305 241 1339
rect 188 1293 241 1305
rect 341 1475 397 1493
rect 341 1441 352 1475
rect 386 1441 397 1475
rect 341 1407 397 1441
rect 341 1373 352 1407
rect 386 1373 397 1407
rect 341 1339 397 1373
rect 341 1305 352 1339
rect 386 1305 397 1339
rect 341 1293 397 1305
rect 497 1475 553 1493
rect 497 1441 508 1475
rect 542 1441 553 1475
rect 497 1407 553 1441
rect 497 1373 508 1407
rect 542 1373 553 1407
rect 497 1339 553 1373
rect 497 1305 508 1339
rect 542 1305 553 1339
rect 497 1293 553 1305
rect 653 1475 709 1493
rect 653 1441 664 1475
rect 698 1441 709 1475
rect 653 1407 709 1441
rect 653 1373 664 1407
rect 698 1373 709 1407
rect 653 1339 709 1373
rect 653 1305 664 1339
rect 698 1305 709 1339
rect 653 1293 709 1305
rect 809 1475 862 1493
rect 809 1441 820 1475
rect 854 1441 862 1475
rect 809 1407 862 1441
rect 809 1373 820 1407
rect 854 1373 862 1407
rect 809 1339 862 1373
rect 809 1305 820 1339
rect 854 1305 862 1339
rect 809 1293 862 1305
rect 1290 1195 1343 1265
rect 1290 1161 1298 1195
rect 1332 1161 1343 1195
rect 1290 1127 1343 1161
rect 1290 1093 1298 1127
rect 1332 1093 1343 1127
rect 1290 1059 1343 1093
rect 1290 1025 1298 1059
rect 1332 1025 1343 1059
rect 1290 991 1343 1025
rect 1290 957 1298 991
rect 1332 957 1343 991
rect 1290 923 1343 957
rect 1290 889 1298 923
rect 1332 889 1343 923
rect 1290 855 1343 889
rect 1290 821 1298 855
rect 1332 821 1343 855
rect 1290 787 1343 821
rect 1290 753 1298 787
rect 1332 753 1343 787
rect 1290 719 1343 753
rect 1290 685 1298 719
rect 1332 685 1343 719
rect 1290 651 1343 685
rect 1290 617 1298 651
rect 1332 617 1343 651
rect 1290 583 1343 617
rect 1290 549 1298 583
rect 1332 549 1343 583
rect 1290 515 1343 549
rect 1290 481 1298 515
rect 1332 481 1343 515
rect 1290 447 1343 481
rect 188 297 241 333
rect 188 263 196 297
rect 230 263 241 297
rect 188 229 241 263
rect 188 195 196 229
rect 230 195 241 229
rect 188 183 241 195
rect 341 297 394 333
rect 341 263 352 297
rect 386 263 394 297
rect 341 229 394 263
rect 341 195 352 229
rect 386 195 394 229
rect 341 183 394 195
rect 454 315 507 333
rect 454 281 462 315
rect 496 281 507 315
rect 454 247 507 281
rect 454 213 462 247
rect 496 213 507 247
rect 454 179 507 213
rect 454 145 462 179
rect 496 145 507 179
rect 454 133 507 145
rect 667 315 720 333
rect 667 281 678 315
rect 712 283 720 315
rect 712 281 735 283
rect 667 247 735 281
rect 667 213 678 247
rect 712 213 735 247
rect 667 179 735 213
rect 667 145 678 179
rect 712 145 735 179
rect 667 133 735 145
rect 835 247 888 283
rect 835 213 846 247
rect 880 213 888 247
rect 835 179 888 213
rect 835 145 846 179
rect 880 145 888 179
rect 1290 413 1298 447
rect 1332 413 1343 447
rect 1290 379 1343 413
rect 1290 345 1298 379
rect 1332 345 1343 379
rect 1290 311 1343 345
rect 1290 277 1298 311
rect 1332 277 1343 311
rect 1290 265 1343 277
rect 1463 1195 1519 1265
rect 1463 1161 1474 1195
rect 1508 1161 1519 1195
rect 1463 1127 1519 1161
rect 1463 1093 1474 1127
rect 1508 1093 1519 1127
rect 1463 1059 1519 1093
rect 1463 1025 1474 1059
rect 1508 1025 1519 1059
rect 1463 991 1519 1025
rect 1463 957 1474 991
rect 1508 957 1519 991
rect 1463 923 1519 957
rect 1463 889 1474 923
rect 1508 889 1519 923
rect 1463 855 1519 889
rect 1463 821 1474 855
rect 1508 821 1519 855
rect 1463 787 1519 821
rect 1463 753 1474 787
rect 1508 753 1519 787
rect 1463 719 1519 753
rect 1463 685 1474 719
rect 1508 685 1519 719
rect 1463 651 1519 685
rect 1463 617 1474 651
rect 1508 617 1519 651
rect 1463 583 1519 617
rect 1463 549 1474 583
rect 1508 549 1519 583
rect 1463 515 1519 549
rect 1463 481 1474 515
rect 1508 481 1519 515
rect 1463 447 1519 481
rect 1463 413 1474 447
rect 1508 413 1519 447
rect 1463 379 1519 413
rect 1463 345 1474 379
rect 1508 345 1519 379
rect 1463 311 1519 345
rect 1463 277 1474 311
rect 1508 277 1519 311
rect 1463 265 1519 277
rect 1639 1195 1692 1265
rect 1639 1161 1650 1195
rect 1684 1161 1692 1195
rect 1639 1127 1692 1161
rect 1639 1093 1650 1127
rect 1684 1093 1692 1127
rect 1639 1059 1692 1093
rect 1639 1025 1650 1059
rect 1684 1025 1692 1059
rect 1639 991 1692 1025
rect 1639 957 1650 991
rect 1684 957 1692 991
rect 1639 923 1692 957
rect 1639 889 1650 923
rect 1684 889 1692 923
rect 1639 855 1692 889
rect 1639 821 1650 855
rect 1684 821 1692 855
rect 1639 787 1692 821
rect 1639 753 1650 787
rect 1684 753 1692 787
rect 1639 719 1692 753
rect 1639 685 1650 719
rect 1684 685 1692 719
rect 1639 651 1692 685
rect 1639 617 1650 651
rect 1684 617 1692 651
rect 1639 583 1692 617
rect 1639 549 1650 583
rect 1684 549 1692 583
rect 1639 515 1692 549
rect 1639 481 1650 515
rect 1684 481 1692 515
rect 1639 447 1692 481
rect 1639 413 1650 447
rect 1684 413 1692 447
rect 1639 379 1692 413
rect 1639 345 1650 379
rect 1684 345 1692 379
rect 1639 311 1692 345
rect 1639 277 1650 311
rect 1684 277 1692 311
rect 1639 265 1692 277
rect 835 133 888 145
<< mvpdiff >>
rect 176 1039 229 1077
rect 176 1005 184 1039
rect 218 1005 229 1039
rect 176 993 229 1005
rect 629 1039 685 1077
rect 629 1005 640 1039
rect 674 1005 685 1039
rect 629 993 685 1005
rect 1085 1039 1138 1077
rect 1085 1005 1096 1039
rect 1130 1005 1138 1039
rect 1085 993 1138 1005
rect 682 735 735 785
rect 682 701 690 735
rect 724 701 735 735
rect 682 667 735 701
rect 188 599 241 635
rect 188 565 196 599
rect 230 565 241 599
rect 188 531 241 565
rect 188 497 196 531
rect 230 497 241 531
rect 188 485 241 497
rect 341 599 394 635
rect 341 565 352 599
rect 386 565 394 599
rect 341 531 394 565
rect 341 497 352 531
rect 386 497 394 531
rect 341 485 394 497
rect 682 633 690 667
rect 724 633 735 667
rect 682 599 735 633
rect 682 565 690 599
rect 724 565 735 599
rect 682 531 735 565
rect 682 497 690 531
rect 724 497 735 531
rect 682 485 735 497
rect 835 735 888 785
rect 835 701 846 735
rect 880 701 888 735
rect 835 667 888 701
rect 835 633 846 667
rect 880 633 888 667
rect 835 599 888 633
rect 835 565 846 599
rect 880 565 888 599
rect 835 531 888 565
rect 835 497 846 531
rect 880 497 888 531
rect 835 485 888 497
<< ndiffc >>
rect 1857 1431 1891 1465
rect 1857 1341 1891 1375
rect 1957 1431 1991 1465
rect 1957 1341 1991 1375
rect 1929 253 1963 287
rect 1929 163 1963 197
rect 2029 253 2063 287
rect 2029 163 2063 197
<< pdiffc >>
rect 1857 1137 1891 1171
rect 1857 1054 1891 1088
rect 1857 971 1891 1005
rect 1957 1111 1991 1145
rect 1957 1041 1991 1075
rect 1957 971 1991 1005
rect 1929 623 1963 657
rect 1929 553 1963 587
rect 1929 483 1963 517
rect 2029 623 2063 657
rect 2029 540 2063 574
rect 2029 457 2063 491
<< mvndiffc >>
rect 196 1441 230 1475
rect 196 1373 230 1407
rect 196 1305 230 1339
rect 352 1441 386 1475
rect 352 1373 386 1407
rect 352 1305 386 1339
rect 508 1441 542 1475
rect 508 1373 542 1407
rect 508 1305 542 1339
rect 664 1441 698 1475
rect 664 1373 698 1407
rect 664 1305 698 1339
rect 820 1441 854 1475
rect 820 1373 854 1407
rect 820 1305 854 1339
rect 1298 1161 1332 1195
rect 1298 1093 1332 1127
rect 1298 1025 1332 1059
rect 1298 957 1332 991
rect 1298 889 1332 923
rect 1298 821 1332 855
rect 1298 753 1332 787
rect 1298 685 1332 719
rect 1298 617 1332 651
rect 1298 549 1332 583
rect 1298 481 1332 515
rect 196 263 230 297
rect 196 195 230 229
rect 352 263 386 297
rect 352 195 386 229
rect 462 281 496 315
rect 462 213 496 247
rect 462 145 496 179
rect 678 281 712 315
rect 678 213 712 247
rect 678 145 712 179
rect 846 213 880 247
rect 846 145 880 179
rect 1298 413 1332 447
rect 1298 345 1332 379
rect 1298 277 1332 311
rect 1474 1161 1508 1195
rect 1474 1093 1508 1127
rect 1474 1025 1508 1059
rect 1474 957 1508 991
rect 1474 889 1508 923
rect 1474 821 1508 855
rect 1474 753 1508 787
rect 1474 685 1508 719
rect 1474 617 1508 651
rect 1474 549 1508 583
rect 1474 481 1508 515
rect 1474 413 1508 447
rect 1474 345 1508 379
rect 1474 277 1508 311
rect 1650 1161 1684 1195
rect 1650 1093 1684 1127
rect 1650 1025 1684 1059
rect 1650 957 1684 991
rect 1650 889 1684 923
rect 1650 821 1684 855
rect 1650 753 1684 787
rect 1650 685 1684 719
rect 1650 617 1684 651
rect 1650 549 1684 583
rect 1650 481 1684 515
rect 1650 413 1684 447
rect 1650 345 1684 379
rect 1650 277 1684 311
<< mvpdiffc >>
rect 184 1005 218 1039
rect 640 1005 674 1039
rect 1096 1005 1130 1039
rect 690 701 724 735
rect 196 565 230 599
rect 196 497 230 531
rect 352 565 386 599
rect 352 497 386 531
rect 690 633 724 667
rect 690 565 724 599
rect 690 497 724 531
rect 846 701 880 735
rect 846 633 880 667
rect 846 565 880 599
rect 846 497 880 531
<< nsubdiff >>
rect 1820 797 1850 831
rect 1884 797 1922 831
rect 1956 797 1987 831
<< mvpsubdiff >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2143 1645
rect 2177 1611 2239 1645
rect 2273 1611 2335 1645
rect 2369 1611 2431 1645
rect 2465 1611 2527 1645
rect 2561 1611 2623 1645
rect 2657 1611 2719 1645
rect 2753 1611 2784 1645
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< mvnsubdiff >>
rect 72 1004 106 1056
rect 72 831 106 970
rect 0 797 31 831
rect 65 797 137 831
<< nsubdiffcont >>
rect 1850 797 1884 831
rect 1922 797 1956 831
<< mvpsubdiffcont >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 1663 1611 1697 1645
rect 1759 1611 1793 1645
rect 1855 1611 1889 1645
rect 1951 1611 1985 1645
rect 2047 1611 2081 1645
rect 2143 1611 2177 1645
rect 2239 1611 2273 1645
rect 2335 1611 2369 1645
rect 2431 1611 2465 1645
rect 2527 1611 2561 1645
rect 2623 1611 2657 1645
rect 2719 1611 2753 1645
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< mvnsubdiffcont >>
rect 72 970 106 1004
rect 31 797 65 831
<< poly >>
rect 241 1493 341 1519
rect 397 1493 497 1519
rect 553 1493 653 1519
rect 709 1493 809 1519
rect 1040 1465 1684 1481
rect 1902 1477 1932 1504
rect 1040 1445 1566 1465
rect 241 1261 341 1293
rect 397 1261 497 1293
rect 241 1225 497 1261
rect 553 1261 653 1293
rect 709 1261 809 1293
rect 1040 1261 1076 1445
rect 1550 1431 1566 1445
rect 1600 1431 1634 1465
rect 1668 1431 1684 1465
rect 1550 1415 1684 1431
rect 553 1225 1076 1261
rect 1118 1333 1786 1369
rect 461 1183 497 1225
rect 1118 1183 1154 1333
rect 1750 1291 1786 1333
rect 1902 1291 1932 1329
rect 1343 1265 1463 1291
rect 1519 1265 1639 1291
rect 1750 1275 2075 1291
rect 229 1161 407 1177
rect 229 1127 289 1161
rect 323 1127 357 1161
rect 391 1127 407 1161
rect 461 1147 1154 1183
rect 229 1103 407 1127
rect 229 1077 629 1103
rect 685 1077 1085 1103
rect 229 967 629 993
rect 241 635 341 967
rect 685 925 1085 993
rect 422 909 1085 925
rect 422 875 438 909
rect 472 875 506 909
rect 540 875 1085 909
rect 422 859 1085 875
rect 735 785 835 811
rect 241 333 341 485
rect 735 432 835 485
rect 507 416 667 432
rect 507 382 546 416
rect 580 382 614 416
rect 648 382 667 416
rect 507 333 667 382
rect 735 416 1080 432
rect 735 382 962 416
rect 996 382 1030 416
rect 1064 382 1080 416
rect 735 366 1080 382
rect 241 157 341 183
rect 735 283 835 366
rect 1014 239 1080 366
rect 1750 1255 1957 1275
rect 1901 1241 1957 1255
rect 1991 1241 2025 1275
rect 2059 1241 2075 1275
rect 1901 1225 2075 1241
rect 1901 1198 1937 1225
rect 1904 1183 1934 1198
rect 1904 933 1934 959
rect 1986 669 2016 695
rect 1986 430 2016 445
rect 1983 403 2019 430
rect 1845 387 2019 403
rect 1845 353 1861 387
rect 1895 353 1929 387
rect 1963 353 2019 387
rect 1845 337 2019 353
rect 1988 299 2018 337
rect 1343 239 1463 265
rect 1519 239 1639 265
rect 1014 173 1639 239
rect 507 107 667 133
rect 735 107 835 133
rect 1988 125 2018 151
<< polycont >>
rect 1566 1431 1600 1465
rect 1634 1431 1668 1465
rect 289 1127 323 1161
rect 357 1127 391 1161
rect 438 875 472 909
rect 506 875 540 909
rect 546 382 580 416
rect 614 382 648 416
rect 962 382 996 416
rect 1030 382 1064 416
rect 1957 1241 1991 1275
rect 2025 1241 2059 1275
rect 1861 353 1895 387
rect 1929 353 1963 387
<< locali >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2143 1645
rect 2177 1611 2239 1645
rect 2273 1611 2335 1645
rect 2369 1611 2431 1645
rect 2465 1611 2527 1645
rect 2561 1611 2623 1645
rect 2657 1611 2719 1645
rect 2753 1611 2784 1645
rect 191 1525 980 1569
rect 191 1475 235 1525
rect 191 1441 196 1475
rect 230 1441 235 1475
rect 191 1407 235 1441
rect 191 1373 196 1407
rect 230 1373 235 1407
rect 191 1339 235 1373
rect 191 1305 196 1339
rect 230 1305 235 1339
rect 191 1289 235 1305
rect 347 1475 391 1491
rect 347 1441 352 1475
rect 386 1441 391 1475
rect 347 1407 391 1441
rect 347 1373 352 1407
rect 386 1373 391 1407
rect 347 1339 391 1373
rect 347 1305 352 1339
rect 386 1305 391 1339
rect 347 1255 391 1305
rect 503 1475 547 1525
rect 503 1441 508 1475
rect 542 1441 547 1475
rect 503 1407 547 1441
rect 503 1373 508 1407
rect 542 1373 547 1407
rect 503 1339 547 1373
rect 503 1305 508 1339
rect 542 1305 547 1339
rect 503 1289 547 1305
rect 659 1475 703 1491
rect 659 1441 664 1475
rect 698 1441 703 1475
rect 659 1407 703 1441
rect 659 1373 664 1407
rect 698 1373 703 1407
rect 659 1339 703 1373
rect 659 1305 664 1339
rect 698 1305 703 1339
rect 179 1211 391 1255
rect 72 1004 106 1056
rect 72 831 106 970
rect 179 1039 223 1211
rect 659 1177 703 1305
rect 815 1475 859 1525
rect 815 1441 820 1475
rect 854 1441 859 1475
rect 815 1407 859 1441
rect 815 1373 820 1407
rect 854 1373 859 1407
rect 815 1339 859 1373
rect 815 1305 820 1339
rect 854 1305 859 1339
rect 815 1289 859 1305
rect 936 1303 980 1525
rect 1941 1544 2059 1550
rect 1941 1510 1947 1544
rect 1981 1510 2019 1544
rect 2053 1510 2059 1544
rect 1941 1504 2059 1510
rect 1550 1465 1907 1481
rect 1550 1431 1566 1465
rect 1600 1431 1634 1465
rect 1668 1431 1857 1465
rect 1891 1431 1907 1465
rect 1550 1415 1907 1431
rect 1841 1375 1907 1415
rect 1841 1341 1857 1375
rect 1891 1341 1907 1375
rect 936 1259 1689 1303
rect 1293 1195 1337 1259
rect 273 1161 1135 1177
rect 273 1127 289 1161
rect 323 1127 357 1161
rect 391 1133 1135 1161
rect 391 1127 407 1133
rect 273 1111 407 1127
rect 179 1005 184 1039
rect 218 1005 223 1039
rect 179 959 223 1005
rect 635 1039 679 1081
rect 635 1005 640 1039
rect 674 1005 679 1039
rect 179 915 556 959
rect 422 909 556 915
rect 422 875 438 909
rect 472 875 506 909
rect 540 875 556 909
rect 635 926 679 1005
rect 1091 1039 1135 1133
rect 1091 1005 1096 1039
rect 1130 1005 1135 1039
rect 1091 989 1135 1005
rect 1293 1161 1298 1195
rect 1332 1161 1337 1195
rect 1293 1127 1337 1161
rect 1293 1093 1298 1127
rect 1332 1093 1337 1127
rect 1293 1059 1337 1093
rect 1293 1025 1298 1059
rect 1332 1025 1337 1059
rect 1293 991 1337 1025
rect 1293 957 1298 991
rect 1332 957 1337 991
rect 635 882 729 926
rect 422 859 556 875
rect 0 797 31 831
rect 65 797 103 831
rect 352 735 470 747
rect 352 701 358 735
rect 392 701 430 735
rect 464 701 470 735
rect 352 689 470 701
rect 191 599 235 615
rect 191 565 196 599
rect 230 565 235 599
rect 191 539 235 565
rect 151 531 235 539
rect 151 497 196 531
rect 230 497 235 531
rect 151 481 235 497
rect 352 599 386 689
rect 512 617 556 859
rect 685 747 729 882
rect 1293 923 1337 957
rect 1293 889 1298 923
rect 1332 889 1337 923
rect 1293 855 1337 889
rect 1293 821 1298 855
rect 1332 821 1337 855
rect 1293 787 1337 821
rect 1293 753 1298 787
rect 1332 753 1337 787
rect 612 735 729 747
rect 612 701 618 735
rect 652 701 690 735
rect 724 701 729 735
rect 612 689 729 701
rect 352 531 386 565
rect 352 481 386 497
rect 452 572 556 617
rect 685 667 729 689
rect 685 633 690 667
rect 724 633 729 667
rect 685 599 729 633
rect 151 321 195 481
rect 151 297 235 321
rect 452 315 496 572
rect 685 565 690 599
rect 724 565 729 599
rect 685 531 729 565
rect 685 497 690 531
rect 724 497 729 531
rect 685 481 729 497
rect 841 735 885 751
rect 841 701 846 735
rect 880 701 885 735
rect 841 667 885 701
rect 841 633 846 667
rect 880 633 885 667
rect 841 599 885 633
rect 841 565 846 599
rect 880 565 885 599
rect 841 531 885 565
rect 841 497 846 531
rect 880 497 885 531
rect 841 432 885 497
rect 1293 719 1337 753
rect 1293 685 1298 719
rect 1332 685 1337 719
rect 1293 651 1337 685
rect 1293 617 1298 651
rect 1332 617 1337 651
rect 1293 583 1337 617
rect 1293 549 1298 583
rect 1332 549 1337 583
rect 1293 515 1337 549
rect 1293 481 1298 515
rect 1332 481 1337 515
rect 1293 447 1337 481
rect 530 416 885 432
rect 530 382 546 416
rect 580 382 614 416
rect 648 388 885 416
rect 648 382 664 388
rect 530 366 664 382
rect 151 263 196 297
rect 230 263 235 297
rect 191 229 235 263
rect 191 195 196 229
rect 230 195 235 229
rect 191 179 235 195
rect 352 297 398 313
rect 386 263 398 297
rect 352 229 398 263
rect 386 195 398 229
rect 352 125 398 195
rect 452 281 462 315
rect 452 247 496 281
rect 452 213 462 247
rect 452 179 496 213
rect 452 145 462 179
rect 452 129 496 145
rect 672 315 718 331
rect 672 281 678 315
rect 712 281 718 315
rect 672 247 718 281
rect 672 213 678 247
rect 712 213 718 247
rect 672 179 718 213
rect 672 145 678 179
rect 712 145 718 179
rect 672 125 718 145
rect 841 247 885 388
rect 946 416 1080 432
rect 946 382 962 416
rect 996 382 1030 416
rect 1064 382 1080 416
rect 946 366 1080 382
rect 1293 413 1298 447
rect 1332 413 1337 447
rect 1293 379 1337 413
rect 1293 345 1298 379
rect 1332 345 1337 379
rect 1293 311 1337 345
rect 1293 277 1298 311
rect 1332 277 1337 311
rect 1293 261 1337 277
rect 1468 1195 1514 1211
rect 1468 1161 1474 1195
rect 1508 1161 1514 1195
rect 1468 1127 1514 1161
rect 1468 1093 1474 1127
rect 1508 1093 1514 1127
rect 1468 1059 1514 1093
rect 1468 1025 1474 1059
rect 1508 1025 1514 1059
rect 1468 991 1514 1025
rect 1468 957 1474 991
rect 1508 957 1514 991
rect 1468 923 1514 957
rect 1468 889 1474 923
rect 1508 889 1514 923
rect 1468 855 1514 889
rect 1468 821 1474 855
rect 1508 821 1514 855
rect 1468 787 1514 821
rect 1468 753 1474 787
rect 1508 753 1514 787
rect 1468 719 1514 753
rect 1468 685 1474 719
rect 1508 685 1514 719
rect 1468 651 1514 685
rect 1468 617 1474 651
rect 1508 617 1514 651
rect 1468 583 1514 617
rect 1468 549 1474 583
rect 1508 549 1514 583
rect 1468 515 1514 549
rect 1468 481 1474 515
rect 1508 481 1514 515
rect 1468 447 1514 481
rect 1468 413 1474 447
rect 1508 413 1514 447
rect 1468 379 1514 413
rect 1468 345 1474 379
rect 1508 345 1514 379
rect 1468 311 1514 345
rect 1468 277 1474 311
rect 1508 277 1514 311
rect 841 213 846 247
rect 880 213 885 247
rect 841 179 885 213
rect 841 145 846 179
rect 880 145 885 179
rect 841 129 885 145
rect 1468 125 1514 277
rect 1645 1195 1689 1259
rect 1645 1161 1650 1195
rect 1684 1161 1689 1195
rect 1645 1127 1689 1161
rect 1645 1093 1650 1127
rect 1684 1093 1689 1127
rect 1645 1059 1689 1093
rect 1645 1025 1650 1059
rect 1684 1025 1689 1059
rect 1645 991 1689 1025
rect 1645 957 1650 991
rect 1684 957 1689 991
rect 1645 923 1689 957
rect 1841 1171 1907 1341
rect 1941 1465 2007 1504
rect 1941 1431 1957 1465
rect 1991 1431 2007 1465
rect 1941 1375 2007 1431
rect 1941 1341 1957 1375
rect 1991 1341 2007 1375
rect 1941 1325 2007 1341
rect 1941 1275 2107 1291
rect 1941 1241 1957 1275
rect 1991 1241 2025 1275
rect 2059 1241 2107 1275
rect 1941 1225 2107 1241
rect 1841 1137 1857 1171
rect 1891 1137 1907 1171
rect 1841 1088 1907 1137
rect 1841 1054 1857 1088
rect 1891 1054 1907 1088
rect 1841 1005 1907 1054
rect 1841 971 1857 1005
rect 1891 971 1907 1005
rect 1841 955 1907 971
rect 1941 1145 2007 1161
rect 1941 1111 1957 1145
rect 1991 1111 2007 1145
rect 1941 1075 2007 1111
rect 1941 1041 1957 1075
rect 1991 1041 2007 1075
rect 1941 1005 2007 1041
rect 1941 971 1957 1005
rect 1991 971 2007 1005
rect 1645 889 1650 923
rect 1684 889 1689 923
rect 1645 855 1689 889
rect 1645 821 1650 855
rect 1684 821 1689 855
rect 1941 847 2007 971
rect 1645 787 1689 821
rect 1645 753 1650 787
rect 1684 753 1689 787
rect 1820 831 2007 847
rect 1820 797 1850 831
rect 1884 797 1922 831
rect 1956 797 2007 831
rect 1820 781 2007 797
rect 1645 719 1689 753
rect 1645 685 1650 719
rect 1684 685 1689 719
rect 1645 651 1689 685
rect 1913 673 1979 781
rect 2041 673 2107 1225
rect 1645 617 1650 651
rect 1684 617 1689 651
rect 1645 583 1689 617
rect 1861 657 1979 673
rect 1861 650 1929 657
rect 1963 650 1979 657
rect 1861 616 1867 650
rect 1901 623 1929 650
rect 1901 616 1939 623
rect 1973 616 1979 650
rect 1861 604 1979 616
rect 1645 549 1650 583
rect 1684 549 1689 583
rect 1645 515 1689 549
rect 1645 481 1650 515
rect 1684 481 1689 515
rect 1645 447 1689 481
rect 1913 587 1979 604
rect 1913 553 1929 587
rect 1963 553 1979 587
rect 1913 517 1979 553
rect 1913 483 1929 517
rect 1963 483 1979 517
rect 1913 467 1979 483
rect 2013 657 2107 673
rect 2013 623 2029 657
rect 2063 623 2107 657
rect 2013 607 2107 623
rect 2013 574 2079 607
rect 2013 540 2029 574
rect 2063 540 2079 574
rect 2013 491 2079 540
rect 1645 413 1650 447
rect 1684 413 1689 447
rect 1645 379 1689 413
rect 2013 457 2029 491
rect 2063 457 2079 491
rect 1645 345 1650 379
rect 1684 345 1689 379
rect 1645 311 1689 345
rect 1841 387 1979 403
rect 1841 353 1861 387
rect 1895 353 1929 387
rect 1963 353 1979 387
rect 1841 337 1979 353
rect 1645 277 1650 311
rect 1684 277 1689 311
rect 1645 261 1689 277
rect 1913 287 1979 303
rect 1913 253 1929 287
rect 1963 253 1979 287
rect 1913 197 1979 253
rect 1913 163 1929 197
rect 1963 163 1979 197
rect 1913 125 1979 163
rect 2013 287 2079 457
rect 2013 253 2029 287
rect 2063 253 2079 287
rect 2013 197 2079 253
rect 2013 163 2029 197
rect 2063 163 2079 197
rect 2013 147 2079 163
rect 280 119 398 125
rect 280 85 286 119
rect 320 85 358 119
rect 392 85 398 119
rect 280 79 398 85
rect 635 119 753 125
rect 635 85 641 119
rect 675 85 713 119
rect 747 85 753 119
rect 635 79 753 85
rect 1431 119 1549 125
rect 1431 85 1437 119
rect 1471 85 1509 119
rect 1543 85 1549 119
rect 1431 79 1549 85
rect 1861 119 1979 125
rect 1861 85 1867 119
rect 1901 85 1939 119
rect 1973 85 1979 119
rect 1861 79 1979 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 1663 1611 1697 1645
rect 1759 1611 1793 1645
rect 1855 1611 1889 1645
rect 1951 1611 1985 1645
rect 2047 1611 2081 1645
rect 2143 1611 2177 1645
rect 2239 1611 2273 1645
rect 2335 1611 2369 1645
rect 2431 1611 2465 1645
rect 2527 1611 2561 1645
rect 2623 1611 2657 1645
rect 2719 1611 2753 1645
rect 1947 1510 1981 1544
rect 2019 1510 2053 1544
rect 31 797 65 831
rect 103 797 137 831
rect 358 701 392 735
rect 430 701 464 735
rect 618 701 652 735
rect 690 701 724 735
rect 1867 616 1901 650
rect 1939 623 1963 650
rect 1963 623 1973 650
rect 1939 616 1973 623
rect 286 85 320 119
rect 358 85 392 119
rect 641 85 675 119
rect 713 85 747 119
rect 1437 85 1471 119
rect 1509 85 1543 119
rect 1867 85 1901 119
rect 1939 85 1973 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 1645 2784 1651
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2143 1645
rect 2177 1611 2239 1645
rect 2273 1611 2335 1645
rect 2369 1611 2431 1645
rect 2465 1611 2527 1645
rect 2561 1611 2623 1645
rect 2657 1611 2719 1645
rect 2753 1611 2784 1645
rect 0 1605 2784 1611
rect 0 1544 2784 1577
rect 0 1510 1947 1544
rect 1981 1510 2019 1544
rect 2053 1510 2784 1544
rect 0 1503 2784 1510
rect 0 865 2784 939
rect 0 831 2784 837
rect 0 797 31 831
rect 65 797 103 831
rect 137 797 2784 831
rect 0 791 2784 797
rect 0 735 2784 763
rect 0 701 358 735
rect 392 701 430 735
rect 464 701 618 735
rect 652 701 690 735
rect 724 701 2784 735
rect 0 689 2784 701
rect 14 650 2770 661
rect 14 616 1867 650
rect 1901 616 1939 650
rect 1973 616 2770 650
rect 14 604 2770 616
rect 0 119 2784 125
rect 0 85 286 119
rect 320 85 358 119
rect 392 85 641 119
rect 675 85 713 119
rect 747 85 1437 119
rect 1471 85 1509 119
rect 1543 85 1867 119
rect 1901 85 1939 119
rect 1973 85 2784 119
rect 0 51 2784 85
rect 0 17 2784 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -23 2784 -17
<< labels >>
flabel locali s 996 382 1030 416 0 FreeSans 400 0 0 0 SLEEP_B
port 2 nsew signal input
flabel locali s 1895 353 1929 387 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 156 382 190 416 0 FreeSans 400 90 0 0 X
port 8 nsew signal output
flabel metal1 s 0 1605 2784 1628 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 0 2784 23 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 51 2784 125 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 1503 2784 1577 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 791 2784 837 0 FreeSans 520 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 0 865 2784 939 0 FreeSans 520 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 689 2784 763 0 FreeSans 520 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 14 604 2770 661 0 FreeSans 520 0 0 0 LVPWR
port 3 nsew power bidirectional
flabel comment s 885 1048 885 1048 0 FreeSans 200 0 0 0 M3
flabel comment s 291 246 291 246 0 FreeSans 200 0 0 0 M7
flabel comment s 291 548 291 548 0 FreeSans 200 0 0 0 M8
flabel comment s 447 1390 447 1390 0 FreeSans 200 0 0 0 I16
flabel comment s 785 208 785 208 0 FreeSans 200 0 0 0 I6
flabel comment s 603 1390 603 1390 0 FreeSans 200 0 0 0 I15
flabel comment s 1225 1463 1225 1463 0 FreeSans 200 0 0 0 t4
flabel comment s 1315 736 1315 736 0 FreeSans 300 0 0 0 D
flabel comment s 1491 736 1491 736 0 FreeSans 300 0 0 0 S
flabel comment s 1667 736 1667 736 0 FreeSans 300 0 0 0 D
flabel comment s 863 196 863 196 0 FreeSans 300 0 0 0 D
flabel comment s 479 230 479 230 0 FreeSans 300 0 0 0 D
flabel comment s 695 230 695 230 0 FreeSans 300 0 0 0 S
flabel comment s 369 246 369 246 0 FreeSans 300 180 0 0 S
flabel comment s 213 246 213 246 0 FreeSans 300 180 0 0 D
flabel comment s 1423 736 1423 736 0 FreeSans 200 0 0 0 I23
flabel comment s 707 616 707 616 0 FreeSans 300 0 0 0 S
flabel comment s 863 616 863 616 0 FreeSans 300 0 0 0 D
flabel comment s 369 548 369 548 0 FreeSans 300 180 0 0 S
flabel comment s 213 548 213 548 0 FreeSans 300 180 0 0 D
flabel comment s 429 1048 429 1048 0 FreeSans 200 0 0 0 M4
flabel comment s 291 1390 291 1390 0 FreeSans 200 0 0 0 I16
flabel comment s 657 1022 657 1022 0 FreeSans 300 180 0 0 S
flabel comment s 201 1022 201 1022 0 FreeSans 300 180 0 0 D
flabel comment s 657 1022 657 1022 0 FreeSans 300 0 0 0 S
flabel comment s 1113 1022 1113 1022 0 FreeSans 300 0 0 0 D
flabel comment s 759 1390 759 1390 0 FreeSans 200 0 0 0 I15
flabel comment s 785 616 785 616 0 FreeSans 200 0 0 0 I7
flabel comment s 587 230 587 230 0 FreeSans 200 0 0 0 M9
flabel comment s 525 1390 525 1390 0 FreeSans 300 0 0 0 S
flabel comment s 681 1390 681 1390 0 FreeSans 300 0 0 0 D
flabel comment s 837 1390 837 1390 0 FreeSans 300 0 0 0 S
flabel comment s 681 1233 681 1233 0 FreeSans 200 0 0 0 t1
flabel comment s 525 1390 525 1390 0 FreeSans 300 180 0 0 S
flabel comment s 369 1390 369 1390 0 FreeSans 300 180 0 0 D
flabel comment s 1579 736 1579 736 0 FreeSans 200 0 0 0 I23
flabel comment s 213 1390 213 1390 0 FreeSans 300 180 0 0 S
flabel comment s 369 1233 369 1233 0 FreeSans 200 0 0 0 t2
flabel comment s 1225 1351 1225 1351 0 FreeSans 200 0 0 0 t3
rlabel viali s 1939 616 1973 650 1 LVPWR
port 3 nsew power bidirectional
rlabel viali s 1867 616 1901 650 1 LVPWR
port 3 nsew power bidirectional
rlabel metal1 s 14 604 2770 661 1 LVPWR
port 3 nsew power bidirectional
rlabel locali s 672 125 718 331 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 635 79 753 125 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 1468 125 1514 1211 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 1431 79 1549 125 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 1913 125 1979 303 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 1861 79 1979 125 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 1941 1504 2059 1550 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 1941 1325 2007 1504 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 2019 1510 2053 1544 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1947 1510 1981 1544 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1939 85 1973 119 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1867 85 1901 119 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1509 85 1543 119 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1437 85 1471 119 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 713 85 747 119 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 641 85 675 119 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 358 85 392 119 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 286 85 320 119 1 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 51 2784 125 1 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 1503 2784 1577 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 0 1611 2784 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2719 1611 2753 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2719 -17 2753 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2623 1611 2657 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2623 -17 2657 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2527 1611 2561 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2527 -17 2561 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2431 1611 2465 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2431 -17 2465 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2335 1611 2369 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2335 -17 2369 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2239 1611 2273 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2239 -17 2273 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2143 1611 2177 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2143 -17 2177 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2047 1611 2081 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2047 -17 2081 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1951 1611 1985 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1951 -17 1985 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1855 1611 1889 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1855 -17 1889 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1759 1611 1793 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1759 -17 1793 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1663 1611 1697 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1663 -17 1697 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1567 1611 1601 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1567 -17 1601 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1471 1611 1505 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1471 -17 1505 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1375 1611 1409 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1375 -17 1409 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1279 1611 1313 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1279 -17 1313 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1183 1611 1217 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1183 -17 1217 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1087 1611 1121 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1087 -17 1121 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 991 1611 1025 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 991 -17 1025 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 895 1611 929 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 895 -17 929 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 799 1611 833 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 799 -17 833 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 703 1611 737 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 703 -17 737 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 607 1611 641 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 607 -17 641 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 511 1611 545 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 511 -17 545 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 415 1611 449 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 415 -17 449 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 319 1611 353 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 319 -17 353 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 223 1611 257 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 223 -17 257 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 127 1611 161 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 127 -17 161 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 31 1611 65 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 31 -17 65 17 1 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 -23 2784 23 1 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 1605 2784 1651 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 103 797 137 831 1 VPB
port 6 nsew power bidirectional
rlabel viali s 31 797 65 831 1 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 791 2784 837 1 VPB
port 6 nsew power bidirectional
rlabel locali s 685 747 729 882 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 685 481 729 689 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 635 926 679 1081 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 635 882 729 926 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 612 689 729 747 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 690 701 724 735 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 618 701 652 735 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 430 701 464 735 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 358 701 392 735 1 VPWR
port 7 nsew power bidirectional
rlabel metal1 s 0 689 2784 763 1 VPWR
port 7 nsew power bidirectional
rlabel metal1 s 0 865 2784 939 1 VPWR
port 7 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 2784 1628
string GDS_END 301864
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 272604
string LEFclass CORE
string LEFsite unithvdbl
string LEFsymmetry X Y
<< end >>
