magic
tech sky130B
magscale 1 2
timestamp 1666199351
use sky130_fd_io__gpio_ovtv2_amux_switch_pmos  sky130_fd_io__gpio_ovtv2_amux_switch_pmos_0
timestamp 1666199351
transform -1 0 8611 0 1 -353
box -80 769 4262 1263
use sky130_fd_io__gpio_ovtv2_amux_switch_pmos  sky130_fd_io__gpio_ovtv2_amux_switch_pmos_1
timestamp 1666199351
transform 1 0 47 0 1 -353
box -80 769 4262 1263
<< properties >>
string GDS_END 28873430
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 28873276
<< end >>
