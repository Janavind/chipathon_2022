magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 9 21 643 203
rect 29 -17 63 21
<< scnmos >>
rect 87 47 117 177
rect 171 47 201 177
rect 255 47 285 177
rect 339 47 369 177
rect 523 47 553 177
<< scpmoshvt >>
rect 87 297 117 497
rect 171 297 201 497
rect 255 297 285 497
rect 339 297 369 497
rect 527 297 557 497
<< ndiff >>
rect 35 95 87 177
rect 35 61 43 95
rect 77 61 87 95
rect 35 47 87 61
rect 117 117 171 177
rect 117 83 127 117
rect 161 83 171 117
rect 117 47 171 83
rect 201 95 255 177
rect 201 61 211 95
rect 245 61 255 95
rect 201 47 255 61
rect 285 47 339 177
rect 369 97 523 177
rect 369 63 379 97
rect 413 63 479 97
rect 513 63 523 97
rect 369 47 523 63
rect 553 168 617 177
rect 553 134 569 168
rect 603 134 617 168
rect 553 100 617 134
rect 553 66 569 100
rect 603 66 617 100
rect 553 47 617 66
<< pdiff >>
rect 35 485 87 497
rect 35 451 43 485
rect 77 451 87 485
rect 35 417 87 451
rect 35 383 43 417
rect 77 383 87 417
rect 35 297 87 383
rect 117 297 171 497
rect 201 475 255 497
rect 201 441 211 475
rect 245 441 255 475
rect 201 407 255 441
rect 201 373 211 407
rect 245 373 255 407
rect 201 297 255 373
rect 285 475 339 497
rect 285 441 295 475
rect 329 441 339 475
rect 285 407 339 441
rect 285 373 295 407
rect 329 373 339 407
rect 285 297 339 373
rect 369 475 421 497
rect 369 441 379 475
rect 413 441 421 475
rect 369 297 421 441
rect 475 475 527 497
rect 475 441 483 475
rect 517 441 527 475
rect 475 407 527 441
rect 475 373 483 407
rect 517 373 527 407
rect 475 297 527 373
rect 557 477 617 497
rect 557 443 567 477
rect 601 443 617 477
rect 557 409 617 443
rect 557 375 567 409
rect 601 375 617 409
rect 557 341 617 375
rect 557 307 567 341
rect 601 307 617 341
rect 557 297 617 307
<< ndiffc >>
rect 43 61 77 95
rect 127 83 161 117
rect 211 61 245 95
rect 379 63 413 97
rect 479 63 513 97
rect 569 134 603 168
rect 569 66 603 100
<< pdiffc >>
rect 43 451 77 485
rect 43 383 77 417
rect 211 441 245 475
rect 211 373 245 407
rect 295 441 329 475
rect 295 373 329 407
rect 379 441 413 475
rect 483 441 517 475
rect 483 373 517 407
rect 567 443 601 477
rect 567 375 601 409
rect 567 307 601 341
<< poly >>
rect 87 497 117 523
rect 171 497 201 523
rect 255 497 285 523
rect 339 497 369 523
rect 527 497 557 523
rect 87 265 117 297
rect 171 265 201 297
rect 255 265 285 297
rect 339 265 369 297
rect 527 265 557 297
rect 75 249 129 265
rect 75 215 85 249
rect 119 215 129 249
rect 75 199 129 215
rect 171 249 285 265
rect 171 215 202 249
rect 236 215 285 249
rect 171 199 285 215
rect 327 249 381 265
rect 327 215 337 249
rect 371 215 381 249
rect 327 199 381 215
rect 423 249 557 265
rect 423 215 433 249
rect 467 232 557 249
rect 467 215 553 232
rect 423 199 553 215
rect 87 177 117 199
rect 171 177 201 199
rect 255 177 285 199
rect 339 177 369 199
rect 523 177 553 199
rect 87 21 117 47
rect 171 21 201 47
rect 255 21 285 47
rect 339 21 369 47
rect 523 21 553 47
<< polycont >>
rect 85 215 119 249
rect 202 215 236 249
rect 337 215 371 249
rect 433 215 467 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 485 93 493
rect 17 451 43 485
rect 77 451 93 485
rect 17 417 93 451
rect 17 383 43 417
rect 77 383 93 417
rect 17 357 93 383
rect 211 475 245 527
rect 211 407 245 441
rect 211 357 245 373
rect 279 475 345 493
rect 279 441 295 475
rect 329 441 345 475
rect 279 407 345 441
rect 379 475 413 527
rect 379 425 413 441
rect 447 475 527 493
rect 447 441 483 475
rect 517 441 527 475
rect 279 373 295 407
rect 329 391 345 407
rect 447 407 527 441
rect 447 391 483 407
rect 329 373 483 391
rect 517 373 527 407
rect 279 357 527 373
rect 563 477 627 493
rect 563 443 567 477
rect 601 443 627 477
rect 563 409 627 443
rect 563 375 567 409
rect 601 375 627 409
rect 17 165 51 357
rect 563 341 627 375
rect 85 289 346 323
rect 563 307 567 341
rect 601 307 627 341
rect 85 249 134 289
rect 119 215 134 249
rect 168 249 278 255
rect 168 215 202 249
rect 236 215 278 249
rect 312 249 346 289
rect 501 273 627 307
rect 421 249 467 265
rect 312 215 337 249
rect 371 215 387 249
rect 421 215 433 249
rect 85 199 134 215
rect 421 165 467 215
rect 17 131 467 165
rect 127 117 161 131
rect 27 61 43 95
rect 77 61 93 95
rect 501 97 535 273
rect 127 67 161 83
rect 27 17 93 61
rect 195 61 211 95
rect 245 61 261 95
rect 344 63 379 97
rect 413 63 479 97
rect 513 63 535 97
rect 569 168 627 184
rect 603 134 627 168
rect 569 100 627 134
rect 603 66 627 100
rect 195 17 261 61
rect 569 17 627 66
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 121 289 155 323 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 581 289 615 323 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 xor2_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 637768
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 632386
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 2.720 3.220 2.720 
<< end >>
