magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< locali >>
rect 0 1397 2682 1431
rect 430 724 464 1167
rect 430 690 559 724
rect 1525 690 1559 724
rect 345 485 379 551
rect 212 361 246 427
rect 79 237 113 303
rect 0 -17 2682 17
use sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_4  sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_4_0
timestamp 1666199351
transform 1 0 478 0 1 0
box -36 -17 2240 1471
use sky130_sram_1kbyte_1rw1r_32x256_8_pnand3  sky130_sram_1kbyte_1rw1r_32x256_8_pnand3_0
timestamp 1666199351
transform 1 0 0 0 1 0
box -36 -17 514 1471
<< labels >>
rlabel locali s 1542 707 1542 707 4 Z
port 1 nsew
rlabel locali s 96 270 96 270 4 A
port 2 nsew
rlabel locali s 229 394 229 394 4 B
port 3 nsew
rlabel locali s 362 518 362 518 4 C
port 4 nsew
rlabel locali s 1341 0 1341 0 4 gnd
port 5 nsew
rlabel locali s 1341 1414 1341 1414 4 vdd
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 2682 1414
string GDS_END 6268862
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 6267614
<< end >>
