magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -66 377 3906 897
<< pwell >>
rect 1843 236 3125 291
rect 111 221 3125 236
rect 3399 221 3836 283
rect 111 43 3836 221
rect -26 -43 3866 43
<< mvnmos >>
rect 194 126 294 210
rect 336 126 436 210
rect 492 126 592 210
rect 634 126 734 210
rect 790 126 890 210
rect 946 126 1046 210
rect 1212 126 1312 210
rect 1368 126 1468 210
rect 1510 126 1610 210
rect 1652 126 1752 210
rect 1922 181 2022 265
rect 2104 115 2204 265
rect 2260 115 2360 265
rect 2439 181 2539 265
rect 2646 181 2746 265
rect 2804 181 2904 265
rect 2946 181 3046 265
rect 3212 111 3312 195
rect 3482 173 3582 257
rect 3657 107 3757 257
<< mvpmos >>
rect 122 649 222 733
rect 264 649 364 733
rect 424 649 524 733
rect 566 649 666 733
rect 722 649 822 733
rect 936 649 1036 733
rect 1212 641 1312 725
rect 1368 641 1468 725
rect 1510 641 1610 725
rect 1682 641 1782 725
rect 1952 543 2052 693
rect 2127 543 2227 743
rect 2283 543 2383 743
rect 2474 543 2574 627
rect 2616 543 2716 627
rect 2804 543 2904 627
rect 2960 543 3060 627
rect 3158 543 3258 693
rect 3474 443 3574 593
rect 3653 443 3753 743
<< mvndiff >>
rect 1869 240 1922 265
rect 137 185 194 210
rect 137 151 149 185
rect 183 151 194 185
rect 137 126 194 151
rect 294 126 336 210
rect 436 181 492 210
rect 436 147 447 181
rect 481 147 492 181
rect 436 126 492 147
rect 592 126 634 210
rect 734 185 790 210
rect 734 151 745 185
rect 779 151 790 185
rect 734 126 790 151
rect 890 185 946 210
rect 890 151 901 185
rect 935 151 946 185
rect 890 126 946 151
rect 1046 185 1099 210
rect 1046 151 1057 185
rect 1091 151 1099 185
rect 1046 126 1099 151
rect 1159 185 1212 210
rect 1159 151 1167 185
rect 1201 151 1212 185
rect 1159 126 1212 151
rect 1312 189 1368 210
rect 1312 155 1323 189
rect 1357 155 1368 189
rect 1312 126 1368 155
rect 1468 126 1510 210
rect 1610 126 1652 210
rect 1752 189 1809 210
rect 1752 155 1763 189
rect 1797 155 1809 189
rect 1869 206 1877 240
rect 1911 206 1922 240
rect 1869 181 1922 206
rect 2022 253 2104 265
rect 2022 219 2052 253
rect 2086 219 2104 253
rect 2022 181 2104 219
rect 2044 161 2104 181
rect 1752 126 1809 155
rect 2044 127 2052 161
rect 2086 127 2104 161
rect 2044 115 2104 127
rect 2204 257 2260 265
rect 2204 223 2215 257
rect 2249 223 2260 257
rect 2204 157 2260 223
rect 2204 123 2215 157
rect 2249 123 2260 157
rect 2204 115 2260 123
rect 2360 257 2439 265
rect 2360 223 2371 257
rect 2405 223 2439 257
rect 2360 181 2439 223
rect 2539 181 2646 265
rect 2746 240 2804 265
rect 2746 206 2757 240
rect 2791 206 2804 240
rect 2746 181 2804 206
rect 2904 181 2946 265
rect 3046 240 3099 265
rect 3046 206 3057 240
rect 3091 206 3099 240
rect 3046 181 3099 206
rect 3425 215 3482 257
rect 2360 157 2417 181
rect 2360 123 2371 157
rect 2405 123 2417 157
rect 3159 170 3212 195
rect 2360 115 2417 123
rect 3159 136 3167 170
rect 3201 136 3212 170
rect 3159 111 3212 136
rect 3312 170 3365 195
rect 3425 181 3437 215
rect 3471 181 3482 215
rect 3425 173 3482 181
rect 3582 245 3657 257
rect 3582 211 3612 245
rect 3646 211 3657 245
rect 3582 173 3657 211
rect 3312 136 3323 170
rect 3357 136 3365 170
rect 3604 153 3657 173
rect 3312 111 3365 136
rect 3604 119 3612 153
rect 3646 119 3657 153
rect 3604 107 3657 119
rect 3757 245 3810 257
rect 3757 211 3768 245
rect 3802 211 3810 245
rect 3757 153 3810 211
rect 3757 119 3768 153
rect 3802 119 3810 153
rect 3757 107 3810 119
<< mvpdiff >>
rect 65 708 122 733
rect 65 674 77 708
rect 111 674 122 708
rect 65 649 122 674
rect 222 649 264 733
rect 364 725 424 733
rect 364 691 375 725
rect 409 691 424 725
rect 364 649 424 691
rect 524 649 566 733
rect 666 708 722 733
rect 666 674 677 708
rect 711 674 722 708
rect 666 649 722 674
rect 822 720 936 733
rect 822 686 834 720
rect 868 686 936 720
rect 822 649 936 686
rect 1036 691 1093 733
rect 2074 731 2127 743
rect 1036 657 1047 691
rect 1081 657 1093 691
rect 1036 649 1093 657
rect 1155 700 1212 725
rect 1155 666 1167 700
rect 1201 666 1212 700
rect 1155 641 1212 666
rect 1312 687 1368 725
rect 1312 653 1323 687
rect 1357 653 1368 687
rect 1312 641 1368 653
rect 1468 641 1510 725
rect 1610 717 1682 725
rect 1610 683 1621 717
rect 1655 683 1682 717
rect 1610 641 1682 683
rect 1782 687 1839 725
rect 2074 697 2082 731
rect 2116 697 2127 731
rect 2074 693 2127 697
rect 1782 653 1793 687
rect 1827 653 1839 687
rect 1782 641 1839 653
rect 1899 681 1952 693
rect 1899 647 1907 681
rect 1941 647 1952 681
rect 1899 589 1952 647
rect 1899 555 1907 589
rect 1941 555 1952 589
rect 1899 543 1952 555
rect 2052 543 2127 693
rect 2227 588 2283 743
rect 2227 554 2238 588
rect 2272 554 2283 588
rect 2227 543 2283 554
rect 2383 627 2452 743
rect 3596 735 3653 743
rect 2731 708 2789 716
rect 2731 674 2743 708
rect 2777 674 2789 708
rect 3596 701 3608 735
rect 3642 701 3653 735
rect 2731 627 2789 674
rect 3101 685 3158 693
rect 3101 651 3113 685
rect 3147 651 3158 685
rect 3101 627 3158 651
rect 2383 590 2474 627
rect 2383 556 2410 590
rect 2444 556 2474 590
rect 2383 543 2474 556
rect 2574 543 2616 627
rect 2716 543 2804 627
rect 2904 602 2960 627
rect 2904 568 2915 602
rect 2949 568 2960 602
rect 2904 543 2960 568
rect 3060 585 3158 627
rect 3060 551 3113 585
rect 3147 551 3158 585
rect 3060 543 3158 551
rect 3258 685 3315 693
rect 3258 651 3269 685
rect 3303 651 3315 685
rect 3258 585 3315 651
rect 3596 652 3653 701
rect 3596 618 3608 652
rect 3642 618 3653 652
rect 3596 593 3653 618
rect 3258 551 3269 585
rect 3303 551 3315 585
rect 3258 543 3315 551
rect 3417 585 3474 593
rect 3417 551 3429 585
rect 3463 551 3474 585
rect 3417 495 3474 551
rect 3417 461 3429 495
rect 3463 461 3474 495
rect 3417 443 3474 461
rect 3574 568 3653 593
rect 3574 534 3608 568
rect 3642 534 3653 568
rect 3574 485 3653 534
rect 3574 451 3608 485
rect 3642 451 3653 485
rect 3574 443 3653 451
rect 3753 735 3810 743
rect 3753 701 3764 735
rect 3798 701 3810 735
rect 3753 652 3810 701
rect 3753 618 3764 652
rect 3798 618 3810 652
rect 3753 568 3810 618
rect 3753 534 3764 568
rect 3798 534 3810 568
rect 3753 485 3810 534
rect 3753 451 3764 485
rect 3798 451 3810 485
rect 3753 443 3810 451
<< mvndiffc >>
rect 149 151 183 185
rect 447 147 481 181
rect 745 151 779 185
rect 901 151 935 185
rect 1057 151 1091 185
rect 1167 151 1201 185
rect 1323 155 1357 189
rect 1763 155 1797 189
rect 1877 206 1911 240
rect 2052 219 2086 253
rect 2052 127 2086 161
rect 2215 223 2249 257
rect 2215 123 2249 157
rect 2371 223 2405 257
rect 2757 206 2791 240
rect 3057 206 3091 240
rect 2371 123 2405 157
rect 3167 136 3201 170
rect 3437 181 3471 215
rect 3612 211 3646 245
rect 3323 136 3357 170
rect 3612 119 3646 153
rect 3768 211 3802 245
rect 3768 119 3802 153
<< mvpdiffc >>
rect 77 674 111 708
rect 375 691 409 725
rect 677 674 711 708
rect 834 686 868 720
rect 1047 657 1081 691
rect 1167 666 1201 700
rect 1323 653 1357 687
rect 1621 683 1655 717
rect 2082 697 2116 731
rect 1793 653 1827 687
rect 1907 647 1941 681
rect 1907 555 1941 589
rect 2238 554 2272 588
rect 2743 674 2777 708
rect 3608 701 3642 735
rect 3113 651 3147 685
rect 2410 556 2444 590
rect 2915 568 2949 602
rect 3113 551 3147 585
rect 3269 651 3303 685
rect 3608 618 3642 652
rect 3269 551 3303 585
rect 3429 551 3463 585
rect 3429 461 3463 495
rect 3608 534 3642 568
rect 3608 451 3642 485
rect 3764 701 3798 735
rect 3764 618 3798 652
rect 3764 534 3798 568
rect 3764 451 3798 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3840 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3840 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
<< poly >>
rect 122 733 222 759
rect 264 733 364 759
rect 424 733 524 759
rect 566 733 666 759
rect 722 733 822 759
rect 936 733 1036 759
rect 1212 725 1312 751
rect 1368 725 1468 751
rect 1510 725 1610 751
rect 1682 725 1782 751
rect 2127 743 2227 769
rect 2283 743 2383 769
rect 3653 743 3753 769
rect 122 623 222 649
rect 116 569 222 623
rect 116 535 162 569
rect 196 535 222 569
rect 116 523 222 535
rect 116 501 212 523
rect 116 467 162 501
rect 196 467 212 501
rect 264 481 364 649
rect 424 535 524 649
rect 116 451 212 467
rect 254 409 364 481
rect 194 397 364 409
rect 406 515 524 535
rect 406 481 426 515
rect 460 481 524 515
rect 406 447 524 481
rect 406 413 426 447
rect 460 435 524 447
rect 566 582 666 649
rect 566 548 595 582
rect 629 548 666 582
rect 566 461 666 548
rect 722 623 822 649
rect 722 509 864 623
rect 790 505 864 509
rect 790 471 810 505
rect 844 471 864 505
rect 566 435 734 461
rect 460 413 480 435
rect 406 397 480 413
rect 194 313 294 397
rect 21 286 294 313
rect 21 252 37 286
rect 71 252 105 286
rect 139 252 173 286
rect 207 252 294 286
rect 21 232 294 252
rect 194 210 294 232
rect 336 339 450 355
rect 336 305 399 339
rect 433 305 450 339
rect 336 255 450 305
rect 492 331 566 351
rect 492 297 512 331
rect 546 313 566 331
rect 546 297 592 313
rect 336 210 436 255
rect 492 210 592 297
rect 634 210 734 435
rect 790 437 864 471
rect 790 403 810 437
rect 844 403 864 437
rect 936 509 1036 649
rect 1952 693 2052 719
rect 1212 593 1312 641
rect 1212 559 1237 593
rect 1271 559 1312 593
rect 1212 525 1312 559
rect 1368 527 1468 641
rect 936 489 1046 509
rect 936 455 992 489
rect 1026 455 1046 489
rect 1212 491 1237 525
rect 1271 491 1312 525
rect 1212 471 1312 491
rect 1360 507 1468 527
rect 1360 473 1406 507
rect 1440 473 1468 507
rect 936 421 1046 455
rect 1360 439 1468 473
rect 1360 423 1406 439
rect 936 409 992 421
rect 790 313 864 403
rect 946 387 992 409
rect 1026 387 1046 421
rect 790 210 890 313
rect 946 210 1046 387
rect 1212 405 1406 423
rect 1440 427 1468 439
rect 1510 512 1610 641
rect 1510 492 1627 512
rect 1510 458 1573 492
rect 1607 458 1627 492
rect 1440 405 1460 427
rect 1212 389 1460 405
rect 1510 424 1627 458
rect 1510 390 1573 424
rect 1607 390 1627 424
rect 1212 210 1312 389
rect 1510 370 1627 390
rect 1682 493 1782 641
rect 3158 693 3258 719
rect 2474 627 2574 653
rect 2616 627 2716 653
rect 2804 627 2904 653
rect 2960 627 3060 653
rect 3474 593 3574 619
rect 1952 517 2052 543
rect 2127 521 2227 543
rect 1682 459 1702 493
rect 1736 459 1782 493
rect 1368 331 1468 347
rect 1368 297 1413 331
rect 1447 297 1468 331
rect 1368 210 1468 297
rect 1510 210 1610 370
rect 1682 317 1782 459
rect 1652 225 1782 317
rect 1846 417 2052 517
rect 2094 495 2227 521
rect 2094 461 2114 495
rect 2148 470 2227 495
rect 2283 521 2383 543
rect 2283 470 2432 521
rect 2148 461 2194 470
rect 2094 421 2194 461
rect 2380 431 2432 470
rect 1846 339 2022 417
rect 1846 305 1866 339
rect 1900 305 1968 339
rect 2002 305 2022 339
rect 1846 287 2022 305
rect 1922 265 2022 287
rect 2104 391 2194 421
rect 2246 411 2316 428
rect 2104 265 2204 391
rect 2246 377 2262 411
rect 2296 389 2316 411
rect 2296 377 2360 389
rect 2246 343 2360 377
rect 2246 309 2262 343
rect 2296 309 2360 343
rect 2246 289 2360 309
rect 2402 367 2432 431
rect 2474 495 2574 543
rect 2474 461 2512 495
rect 2546 461 2574 495
rect 2474 421 2574 461
rect 2616 517 2716 543
rect 2616 495 2746 517
rect 2616 461 2692 495
rect 2726 461 2746 495
rect 2616 427 2746 461
rect 2616 417 2692 427
rect 2646 393 2692 417
rect 2726 393 2746 427
rect 2402 347 2604 367
rect 2402 313 2418 347
rect 2452 313 2486 347
rect 2520 313 2554 347
rect 2588 313 2604 347
rect 2402 291 2604 313
rect 2260 265 2360 289
rect 2439 265 2539 291
rect 2646 265 2746 393
rect 2804 490 2904 543
rect 2804 456 2824 490
rect 2858 456 2904 490
rect 2960 459 3060 543
rect 2804 422 2904 456
rect 2804 388 2824 422
rect 2858 388 2904 422
rect 2804 265 2904 388
rect 2946 439 3060 459
rect 2946 405 3001 439
rect 3035 405 3060 439
rect 2946 371 3060 405
rect 2946 337 3001 371
rect 3035 337 3060 371
rect 2946 291 3060 337
rect 3158 495 3258 543
rect 3158 461 3178 495
rect 3212 461 3258 495
rect 3158 427 3258 461
rect 3158 393 3178 427
rect 3212 393 3258 427
rect 3474 417 3574 443
rect 3653 417 3753 443
rect 2946 265 3046 291
rect 1652 210 1752 225
rect 1922 155 2022 181
rect 194 100 294 126
rect 336 100 436 126
rect 492 100 592 126
rect 634 100 734 126
rect 790 58 890 126
rect 946 100 1046 126
rect 1212 100 1312 126
rect 1368 100 1468 126
rect 1510 100 1610 126
rect 1652 58 1752 126
rect 3158 253 3258 393
rect 3300 355 3582 417
rect 3300 321 3320 355
rect 3354 321 3582 355
rect 3300 301 3582 321
rect 3482 257 3582 301
rect 3653 347 3757 417
rect 3653 313 3673 347
rect 3707 313 3757 347
rect 3653 283 3757 313
rect 3657 257 3757 283
rect 3158 219 3312 253
rect 3212 195 3312 219
rect 2439 155 2539 181
rect 2646 155 2746 181
rect 2804 155 2904 181
rect 2946 155 3046 181
rect 2104 89 2204 115
rect 2260 89 2360 115
rect 3482 147 3582 173
rect 3212 85 3312 111
rect 3657 81 3757 107
rect 790 28 1752 58
<< polycont >>
rect 162 535 196 569
rect 162 467 196 501
rect 426 481 460 515
rect 426 413 460 447
rect 595 548 629 582
rect 810 471 844 505
rect 37 252 71 286
rect 105 252 139 286
rect 173 252 207 286
rect 399 305 433 339
rect 512 297 546 331
rect 810 403 844 437
rect 1237 559 1271 593
rect 992 455 1026 489
rect 1237 491 1271 525
rect 1406 473 1440 507
rect 992 387 1026 421
rect 1406 405 1440 439
rect 1573 458 1607 492
rect 1573 390 1607 424
rect 1702 459 1736 493
rect 1413 297 1447 331
rect 2114 461 2148 495
rect 1866 305 1900 339
rect 1968 305 2002 339
rect 2262 377 2296 411
rect 2262 309 2296 343
rect 2512 461 2546 495
rect 2692 461 2726 495
rect 2692 393 2726 427
rect 2418 313 2452 347
rect 2486 313 2520 347
rect 2554 313 2588 347
rect 2824 456 2858 490
rect 2824 388 2858 422
rect 3001 405 3035 439
rect 3001 337 3035 371
rect 3178 461 3212 495
rect 3178 393 3212 427
rect 3320 321 3354 355
rect 3673 313 3707 347
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3840 831
rect 61 708 127 741
rect 61 674 77 708
rect 111 674 127 708
rect 284 735 474 741
rect 284 701 290 735
rect 324 701 362 735
rect 396 725 434 735
rect 409 701 434 725
rect 468 701 474 735
rect 284 691 375 701
rect 409 691 474 701
rect 512 708 711 741
rect 512 707 677 708
rect 61 655 127 674
rect 512 655 546 707
rect 61 621 546 655
rect 747 735 925 741
rect 781 701 819 735
rect 853 720 891 735
rect 868 701 891 720
rect 747 686 834 701
rect 868 686 925 701
rect 747 681 925 686
rect 961 727 1201 761
rect 61 372 95 621
rect 146 569 546 585
rect 146 535 162 569
rect 196 551 546 569
rect 196 535 212 551
rect 146 501 212 535
rect 146 467 162 501
rect 196 467 212 501
rect 146 451 212 467
rect 61 338 293 372
rect 21 286 223 302
rect 21 252 37 286
rect 71 252 105 286
rect 139 252 173 286
rect 207 252 223 286
rect 21 236 223 252
rect 133 185 199 199
rect 133 151 149 185
rect 183 151 199 185
rect 133 87 199 151
rect 259 183 293 338
rect 329 253 363 551
rect 399 481 426 515
rect 460 481 476 515
rect 399 447 476 481
rect 512 496 546 551
rect 582 582 641 652
rect 677 645 711 674
rect 961 645 995 727
rect 1151 700 1201 727
rect 677 611 995 645
rect 1031 657 1047 691
rect 1081 657 1097 691
rect 582 548 595 582
rect 629 548 641 582
rect 1031 575 1097 657
rect 1151 666 1167 700
rect 1151 633 1201 666
rect 582 532 641 548
rect 677 541 1097 575
rect 677 496 711 541
rect 512 462 711 496
rect 793 471 810 505
rect 844 498 935 505
rect 844 471 895 498
rect 793 464 895 471
rect 929 464 935 498
rect 399 413 426 447
rect 460 413 476 447
rect 399 401 476 413
rect 793 458 935 464
rect 976 489 1127 505
rect 793 437 860 458
rect 793 403 810 437
rect 844 403 860 437
rect 976 455 992 489
rect 1026 455 1127 489
rect 976 421 1127 455
rect 399 367 635 401
rect 976 387 992 421
rect 1026 387 1127 421
rect 976 367 1127 387
rect 399 339 449 367
rect 433 305 449 339
rect 399 289 449 305
rect 496 297 512 331
rect 546 297 562 331
rect 601 310 1127 367
rect 496 269 562 297
rect 496 253 1107 269
rect 329 235 1107 253
rect 329 219 562 235
rect 729 185 795 199
rect 259 181 497 183
rect 259 147 447 181
rect 481 147 497 181
rect 259 123 497 147
rect 729 151 745 185
rect 779 151 795 185
rect 729 87 795 151
rect 133 53 795 87
rect 831 185 1021 199
rect 831 151 901 185
rect 935 151 1021 185
rect 831 113 1021 151
rect 831 79 837 113
rect 871 79 909 113
rect 943 79 981 113
rect 1015 79 1021 113
rect 1057 185 1107 235
rect 1167 201 1201 633
rect 1091 151 1107 185
rect 1057 103 1107 151
rect 1151 185 1201 201
rect 1151 151 1167 185
rect 1151 103 1201 151
rect 1237 727 1443 761
rect 1237 593 1271 727
rect 1237 525 1271 559
rect 831 73 1021 79
rect 1237 87 1271 491
rect 1307 687 1373 691
rect 1307 653 1323 687
rect 1357 653 1373 687
rect 1307 577 1373 653
rect 1409 647 1443 727
rect 1481 735 1671 741
rect 1481 701 1487 735
rect 1521 701 1559 735
rect 1593 717 1631 735
rect 1593 701 1621 717
rect 1665 701 1671 735
rect 1481 683 1621 701
rect 1655 683 1671 701
rect 1707 727 1957 761
rect 1707 647 1741 727
rect 1409 613 1741 647
rect 1777 687 1843 691
rect 1777 653 1793 687
rect 1827 653 1843 687
rect 1777 577 1843 653
rect 1307 543 1843 577
rect 1307 199 1341 543
rect 1390 473 1406 507
rect 1440 473 1456 507
rect 1390 439 1456 473
rect 1390 405 1406 439
rect 1440 417 1456 439
rect 1557 492 1623 507
rect 1557 458 1573 492
rect 1607 458 1623 492
rect 1557 424 1623 458
rect 1659 498 1752 507
rect 1659 464 1663 498
rect 1697 493 1752 498
rect 1697 464 1702 493
rect 1659 459 1702 464
rect 1736 459 1752 493
rect 1659 445 1752 459
rect 1809 479 1843 543
rect 1891 681 1957 727
rect 1993 737 2183 747
rect 1993 703 1999 737
rect 2033 703 2071 737
rect 2105 731 2143 737
rect 2116 703 2143 731
rect 2177 703 2183 737
rect 1993 697 2082 703
rect 2116 697 2183 703
rect 2603 735 2793 741
rect 2603 701 2609 735
rect 2643 701 2681 735
rect 2715 708 2753 735
rect 2715 701 2743 708
rect 2787 701 2793 735
rect 3055 735 3233 741
rect 1891 647 1907 681
rect 1941 661 1957 681
rect 2603 674 2743 701
rect 2777 674 2793 701
rect 2829 671 3019 705
rect 1941 647 2562 661
rect 1891 627 2562 647
rect 2829 638 2863 671
rect 1891 589 1957 627
rect 1891 555 1907 589
rect 1941 555 1957 589
rect 1891 539 1957 555
rect 2192 588 2288 591
rect 2192 554 2238 588
rect 2272 554 2288 588
rect 2192 535 2288 554
rect 2098 495 2156 511
rect 2098 479 2114 495
rect 1809 461 2114 479
rect 2148 461 2156 495
rect 1809 445 2156 461
rect 1440 405 1521 417
rect 1390 383 1521 405
rect 1409 331 1451 347
rect 1409 297 1413 331
rect 1447 297 1451 331
rect 1487 339 1521 383
rect 1557 390 1573 424
rect 1607 409 1623 424
rect 2192 409 2226 535
rect 2324 491 2358 627
rect 1607 390 2226 409
rect 1557 375 2226 390
rect 1487 305 1866 339
rect 1900 305 1968 339
rect 2002 305 2156 339
rect 1409 269 1451 297
rect 1409 240 1927 269
rect 1409 235 1877 240
rect 1307 189 1373 199
rect 1307 155 1323 189
rect 1357 155 1373 189
rect 1307 123 1373 155
rect 1409 87 1451 235
rect 1861 206 1877 235
rect 1911 206 1927 240
rect 1237 53 1451 87
rect 1623 189 1813 199
rect 1623 155 1763 189
rect 1797 155 1813 189
rect 1861 177 1927 206
rect 1968 253 2086 269
rect 1968 219 2052 253
rect 1623 113 1813 155
rect 1623 79 1629 113
rect 1663 79 1701 113
rect 1735 79 1773 113
rect 1807 79 1813 113
rect 1623 73 1813 79
rect 1968 161 2086 219
rect 1968 127 2052 161
rect 1968 113 2086 127
rect 1968 79 1974 113
rect 2008 79 2046 113
rect 2080 79 2086 113
rect 1968 73 2086 79
rect 2122 87 2156 305
rect 2192 257 2226 375
rect 2262 457 2358 491
rect 2394 590 2460 591
rect 2394 556 2410 590
rect 2444 556 2460 590
rect 2262 411 2296 457
rect 2394 421 2460 556
rect 2496 495 2562 627
rect 2496 461 2512 495
rect 2546 461 2562 495
rect 2496 457 2562 461
rect 2606 604 2863 638
rect 2606 421 2640 604
rect 2899 602 2949 635
rect 2899 568 2915 602
rect 2262 343 2296 377
rect 2262 293 2296 309
rect 2332 387 2640 421
rect 2676 534 2949 568
rect 2676 495 2742 534
rect 2676 461 2692 495
rect 2726 461 2742 495
rect 2676 427 2742 461
rect 2676 393 2692 427
rect 2726 393 2742 427
rect 2332 273 2366 387
rect 2676 379 2742 393
rect 2808 464 2815 498
rect 2849 490 2874 498
rect 2808 456 2824 464
rect 2858 456 2874 490
rect 2808 422 2874 456
rect 2808 388 2824 422
rect 2858 388 2874 422
rect 2808 379 2874 388
rect 2402 347 2604 351
rect 2402 313 2418 347
rect 2452 313 2486 347
rect 2520 313 2554 347
rect 2588 343 2604 347
rect 2588 313 2879 343
rect 2402 309 2879 313
rect 2332 257 2421 273
rect 2192 223 2215 257
rect 2249 223 2265 257
rect 2192 157 2265 223
rect 2192 123 2215 157
rect 2249 123 2265 157
rect 2332 223 2371 257
rect 2405 223 2421 257
rect 2332 157 2421 223
rect 2332 123 2371 157
rect 2405 123 2421 157
rect 2457 87 2491 309
rect 2122 53 2491 87
rect 2617 240 2807 273
rect 2617 206 2757 240
rect 2791 206 2807 240
rect 2617 113 2807 206
rect 2617 79 2623 113
rect 2657 79 2695 113
rect 2729 79 2767 113
rect 2801 79 2807 113
rect 2845 141 2879 309
rect 2915 269 2949 534
rect 2985 455 3019 671
rect 3089 701 3127 735
rect 3161 701 3199 735
rect 3546 735 3728 751
rect 3546 701 3548 735
rect 3582 701 3608 735
rect 3654 701 3692 735
rect 3726 701 3728 735
rect 3055 685 3233 701
rect 3055 651 3113 685
rect 3147 651 3233 685
rect 3055 585 3233 651
rect 3055 551 3113 585
rect 3147 551 3233 585
rect 3055 535 3233 551
rect 3269 685 3319 701
rect 3303 651 3319 685
rect 3269 585 3319 651
rect 3546 652 3728 701
rect 3546 618 3608 652
rect 3642 618 3728 652
rect 3303 551 3319 585
rect 3097 495 3228 499
rect 3097 461 3178 495
rect 3212 461 3228 495
rect 2985 439 3051 455
rect 2985 405 3001 439
rect 3035 405 3051 439
rect 2985 371 3051 405
rect 3097 427 3228 461
rect 3097 393 3178 427
rect 3212 393 3228 427
rect 3097 391 3228 393
rect 3269 425 3319 551
rect 3413 585 3510 601
rect 3413 551 3429 585
rect 3463 551 3510 585
rect 3413 495 3510 551
rect 3413 461 3429 495
rect 3463 461 3510 495
rect 3269 391 3440 425
rect 2985 337 3001 371
rect 3035 355 3051 371
rect 3035 337 3320 355
rect 2985 321 3320 337
rect 3354 321 3370 355
rect 3406 285 3440 391
rect 2915 240 3107 269
rect 2915 235 3057 240
rect 3041 206 3057 235
rect 3091 206 3107 240
rect 3041 177 3107 206
rect 3151 251 3440 285
rect 3476 363 3510 461
rect 3546 568 3728 618
rect 3546 534 3608 568
rect 3642 534 3728 568
rect 3546 485 3728 534
rect 3546 451 3608 485
rect 3642 451 3728 485
rect 3546 435 3728 451
rect 3764 735 3815 751
rect 3798 701 3815 735
rect 3764 652 3815 701
rect 3798 618 3815 652
rect 3764 568 3815 618
rect 3798 534 3815 568
rect 3764 485 3815 534
rect 3798 451 3815 485
rect 3476 347 3723 363
rect 3476 313 3673 347
rect 3707 313 3723 347
rect 3476 297 3723 313
rect 3151 170 3217 251
rect 3476 215 3510 297
rect 3151 141 3167 170
rect 2845 136 3167 141
rect 3201 136 3217 170
rect 2845 107 3217 136
rect 3255 170 3373 199
rect 3255 136 3323 170
rect 3357 136 3373 170
rect 3421 181 3437 215
rect 3471 181 3510 215
rect 3421 165 3510 181
rect 3546 245 3728 261
rect 3546 211 3612 245
rect 3646 211 3728 245
rect 3255 113 3373 136
rect 2617 73 2807 79
rect 3255 79 3261 113
rect 3295 79 3333 113
rect 3367 79 3373 113
rect 3255 73 3373 79
rect 3546 153 3728 211
rect 3546 119 3612 153
rect 3646 119 3728 153
rect 3546 113 3728 119
rect 3546 79 3548 113
rect 3582 79 3620 113
rect 3654 79 3692 113
rect 3726 79 3728 113
rect 3764 245 3815 451
rect 3764 211 3768 245
rect 3802 211 3815 245
rect 3764 153 3815 211
rect 3764 119 3768 153
rect 3802 119 3815 153
rect 3764 103 3815 119
rect 3546 73 3728 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3840 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 290 701 324 735
rect 362 725 396 735
rect 362 701 375 725
rect 375 701 396 725
rect 434 701 468 735
rect 747 701 781 735
rect 819 720 853 735
rect 819 701 834 720
rect 834 701 853 720
rect 891 701 925 735
rect 895 464 929 498
rect 837 79 871 113
rect 909 79 943 113
rect 981 79 1015 113
rect 1487 701 1521 735
rect 1559 701 1593 735
rect 1631 717 1665 735
rect 1631 701 1655 717
rect 1655 701 1665 717
rect 1663 464 1697 498
rect 1999 703 2033 737
rect 2071 731 2105 737
rect 2071 703 2082 731
rect 2082 703 2105 731
rect 2143 703 2177 737
rect 2609 701 2643 735
rect 2681 701 2715 735
rect 2753 708 2787 735
rect 2753 701 2777 708
rect 2777 701 2787 708
rect 1629 79 1663 113
rect 1701 79 1735 113
rect 1773 79 1807 113
rect 1974 79 2008 113
rect 2046 79 2080 113
rect 2815 490 2849 498
rect 2815 464 2824 490
rect 2824 464 2849 490
rect 2623 79 2657 113
rect 2695 79 2729 113
rect 2767 79 2801 113
rect 3055 701 3089 735
rect 3127 701 3161 735
rect 3199 701 3233 735
rect 3548 701 3582 735
rect 3620 701 3642 735
rect 3642 701 3654 735
rect 3692 701 3726 735
rect 3261 79 3295 113
rect 3333 79 3367 113
rect 3548 79 3582 113
rect 3620 79 3654 113
rect 3692 79 3726 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
<< metal1 >>
rect 0 831 3840 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3840 831
rect 0 791 3840 797
rect 0 737 3840 763
rect 0 735 1999 737
rect 0 701 290 735
rect 324 701 362 735
rect 396 701 434 735
rect 468 701 747 735
rect 781 701 819 735
rect 853 701 891 735
rect 925 701 1487 735
rect 1521 701 1559 735
rect 1593 701 1631 735
rect 1665 703 1999 735
rect 2033 703 2071 737
rect 2105 703 2143 737
rect 2177 735 3840 737
rect 2177 703 2609 735
rect 1665 701 2609 703
rect 2643 701 2681 735
rect 2715 701 2753 735
rect 2787 701 3055 735
rect 3089 701 3127 735
rect 3161 701 3199 735
rect 3233 701 3548 735
rect 3582 701 3620 735
rect 3654 701 3692 735
rect 3726 701 3840 735
rect 0 689 3840 701
rect 883 498 941 504
rect 883 464 895 498
rect 929 495 941 498
rect 1651 498 1709 504
rect 1651 495 1663 498
rect 929 467 1663 495
rect 929 464 941 467
rect 883 458 941 464
rect 1651 464 1663 467
rect 1697 495 1709 498
rect 2803 498 2861 504
rect 2803 495 2815 498
rect 1697 467 2815 495
rect 1697 464 1709 467
rect 1651 458 1709 464
rect 2803 464 2815 467
rect 2849 464 2861 498
rect 2803 458 2861 464
rect 0 113 3840 125
rect 0 79 837 113
rect 871 79 909 113
rect 943 79 981 113
rect 1015 79 1629 113
rect 1663 79 1701 113
rect 1735 79 1773 113
rect 1807 79 1974 113
rect 2008 79 2046 113
rect 2080 79 2623 113
rect 2657 79 2695 113
rect 2729 79 2767 113
rect 2801 79 3261 113
rect 3295 79 3333 113
rect 3367 79 3548 113
rect 3582 79 3620 113
rect 3654 79 3692 113
rect 3726 79 3840 113
rect 0 51 3840 79
rect 0 17 3840 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3840 17
rect 0 -23 3840 -17
<< labels >>
flabel comment s 1256 43 1256 43 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfrtp_1
flabel metal1 s 0 51 3840 125 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 0 0 3840 23 0 FreeSans 340 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 0 689 3840 763 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 791 3840 814 0 FreeSans 340 0 0 0 VPB
port 8 nsew power bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 607 612 641 646 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 3103 464 3137 498 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 3775 168 3809 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3775 242 3809 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3775 316 3809 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3775 390 3809 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3775 464 3809 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3775 538 3809 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3775 612 3809 646 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 3840 814
string GDS_END 444346
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 407998
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
