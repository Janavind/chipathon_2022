magic
tech sky130B
magscale 1 2
timestamp 1669700202
<< viali >>
rect 5457 47209 5491 47243
rect 7297 47209 7331 47243
rect 7941 47209 7975 47243
rect 8401 47209 8435 47243
rect 9689 47209 9723 47243
rect 10793 47209 10827 47243
rect 11897 47209 11931 47243
rect 13001 47209 13035 47243
rect 14381 47209 14415 47243
rect 15209 47209 15243 47243
rect 16129 47209 16163 47243
rect 17233 47209 17267 47243
rect 17969 47209 18003 47243
rect 21373 47209 21407 47243
rect 23397 47209 23431 47243
rect 24777 47209 24811 47243
rect 26433 47209 26467 47243
rect 42717 47209 42751 47243
rect 43453 47209 43487 47243
rect 44281 47209 44315 47243
rect 46673 47209 46707 47243
rect 18705 47141 18739 47175
rect 20729 47141 20763 47175
rect 41337 47141 41371 47175
rect 4077 47073 4111 47107
rect 4353 47073 4387 47107
rect 19533 47073 19567 47107
rect 23673 47073 23707 47107
rect 23857 47073 23891 47107
rect 31401 47073 31435 47107
rect 32597 47073 32631 47107
rect 33977 47073 34011 47107
rect 34069 47073 34103 47107
rect 37841 47073 37875 47107
rect 38669 47073 38703 47107
rect 40049 47073 40083 47107
rect 45293 47073 45327 47107
rect 5641 47005 5675 47039
rect 9873 47005 9907 47039
rect 10977 47005 11011 47039
rect 12081 47005 12115 47039
rect 13185 47005 13219 47039
rect 14565 47005 14599 47039
rect 15393 47005 15427 47039
rect 16313 47005 16347 47039
rect 17417 47005 17451 47039
rect 18153 47005 18187 47039
rect 18889 47005 18923 47039
rect 19441 47005 19475 47039
rect 19960 47005 19994 47039
rect 21189 47005 21223 47039
rect 22017 47005 22051 47039
rect 22201 47005 22235 47039
rect 22385 47005 22419 47039
rect 22937 47005 22971 47039
rect 23581 47005 23615 47039
rect 23765 47005 23799 47039
rect 24041 47005 24075 47039
rect 24593 47005 24627 47039
rect 25697 47005 25731 47039
rect 25881 47005 25915 47039
rect 25973 47005 26007 47039
rect 27169 47005 27203 47039
rect 27445 47005 27479 47039
rect 29009 47005 29043 47039
rect 29837 47005 29871 47039
rect 30113 47005 30147 47039
rect 32321 47005 32355 47039
rect 33793 47005 33827 47039
rect 35909 47005 35943 47039
rect 36185 47005 36219 47039
rect 37657 47005 37691 47039
rect 37933 47005 37967 47039
rect 38945 47005 38979 47039
rect 40325 47005 40359 47039
rect 42901 47005 42935 47039
rect 43637 47005 43671 47039
rect 44465 47005 44499 47039
rect 45477 47005 45511 47039
rect 46029 47005 46063 47039
rect 29193 46937 29227 46971
rect 31585 46937 31619 46971
rect 31769 46937 31803 46971
rect 36829 46937 36863 46971
rect 41981 46937 42015 46971
rect 19901 46869 19935 46903
rect 20085 46869 20119 46903
rect 25513 46869 25547 46903
rect 28825 46869 28859 46903
rect 33609 46869 33643 46903
rect 36737 46869 36771 46903
rect 37473 46869 37507 46903
rect 3985 46665 4019 46699
rect 18429 46665 18463 46699
rect 19165 46665 19199 46699
rect 21281 46665 21315 46699
rect 23857 46665 23891 46699
rect 25881 46665 25915 46699
rect 26065 46665 26099 46699
rect 33977 46665 34011 46699
rect 34161 46665 34195 46699
rect 22201 46597 22235 46631
rect 25237 46597 25271 46631
rect 30205 46597 30239 46631
rect 38577 46597 38611 46631
rect 4813 46529 4847 46563
rect 6009 46529 6043 46563
rect 7021 46529 7055 46563
rect 9229 46529 9263 46563
rect 10333 46529 10367 46563
rect 11713 46529 11747 46563
rect 12541 46529 12575 46563
rect 13645 46529 13679 46563
rect 14749 46529 14783 46563
rect 15853 46529 15887 46563
rect 17233 46529 17267 46563
rect 18613 46529 18647 46563
rect 19349 46529 19383 46563
rect 19993 46529 20027 46563
rect 21340 46529 21374 46563
rect 22385 46529 22419 46563
rect 22477 46529 22511 46563
rect 22753 46529 22787 46563
rect 23397 46529 23431 46563
rect 24041 46529 24075 46563
rect 24225 46529 24259 46563
rect 24409 46527 24443 46561
rect 24593 46529 24627 46563
rect 25421 46529 25455 46563
rect 26006 46529 26040 46563
rect 27353 46529 27387 46563
rect 28273 46529 28307 46563
rect 28457 46529 28491 46563
rect 28549 46529 28583 46563
rect 29377 46529 29411 46563
rect 29561 46529 29595 46563
rect 30665 46529 30699 46563
rect 30849 46529 30883 46563
rect 31585 46529 31619 46563
rect 34158 46529 34192 46563
rect 35081 46529 35115 46563
rect 36185 46529 36219 46563
rect 36645 46529 36679 46563
rect 37657 46529 37691 46563
rect 38393 46529 38427 46563
rect 38669 46529 38703 46563
rect 39129 46529 39163 46563
rect 39773 46529 39807 46563
rect 40877 46529 40911 46563
rect 43269 46529 43303 46563
rect 43913 46529 43947 46563
rect 45201 46529 45235 46563
rect 45845 46529 45879 46563
rect 19809 46461 19843 46495
rect 20821 46461 20855 46495
rect 22661 46461 22695 46495
rect 24317 46461 24351 46495
rect 26433 46461 26467 46495
rect 26525 46461 26559 46495
rect 27629 46461 27663 46495
rect 29009 46461 29043 46495
rect 29193 46461 29227 46495
rect 30113 46461 30147 46495
rect 30297 46461 30331 46495
rect 31769 46461 31803 46495
rect 32321 46461 32355 46495
rect 32597 46461 32631 46495
rect 34621 46461 34655 46495
rect 35817 46461 35851 46495
rect 36461 46461 36495 46495
rect 37933 46461 37967 46495
rect 41153 46461 41187 46495
rect 44557 46461 44591 46495
rect 27169 46393 27203 46427
rect 36553 46393 36587 46427
rect 42625 46393 42659 46427
rect 17877 46325 17911 46359
rect 20177 46325 20211 46359
rect 20913 46325 20947 46359
rect 21465 46325 21499 46359
rect 25053 46325 25087 46359
rect 27537 46325 27571 46359
rect 28089 46325 28123 46359
rect 31401 46325 31435 46359
rect 34529 46325 34563 46359
rect 37473 46325 37507 46359
rect 37841 46325 37875 46359
rect 38393 46325 38427 46359
rect 5917 46121 5951 46155
rect 16957 46121 16991 46155
rect 18061 46121 18095 46155
rect 18705 46121 18739 46155
rect 22753 46121 22787 46155
rect 24961 46121 24995 46155
rect 28641 46121 28675 46155
rect 31585 46121 31619 46155
rect 38117 46121 38151 46155
rect 40693 46121 40727 46155
rect 41981 46121 42015 46155
rect 42625 46121 42659 46155
rect 43269 46121 43303 46155
rect 43821 46121 43855 46155
rect 44373 46121 44407 46155
rect 45201 46121 45235 46155
rect 20913 46053 20947 46087
rect 30297 46053 30331 46087
rect 32965 46053 32999 46087
rect 37105 46053 37139 46087
rect 38485 46053 38519 46087
rect 41337 46053 41371 46087
rect 19625 45985 19659 46019
rect 23673 45985 23707 46019
rect 25329 45985 25363 46019
rect 25421 45985 25455 46019
rect 28733 45985 28767 46019
rect 31861 45985 31895 46019
rect 31953 45985 31987 46019
rect 33141 45985 33175 46019
rect 33425 45985 33459 46019
rect 34989 45985 35023 46019
rect 36553 45985 36587 46019
rect 37565 45985 37599 46019
rect 38393 45985 38427 46019
rect 40049 45985 40083 46019
rect 18245 45917 18279 45951
rect 18889 45917 18923 45951
rect 19809 45917 19843 45951
rect 19993 45917 20027 45951
rect 20821 45917 20855 45951
rect 20913 45917 20947 45951
rect 21373 45917 21407 45951
rect 21557 45917 21591 45951
rect 23857 45917 23891 45951
rect 24041 45917 24075 45951
rect 25145 45917 25179 45951
rect 25237 45917 25271 45951
rect 26525 45917 26559 45951
rect 26709 45917 26743 45951
rect 26801 45917 26835 45951
rect 27445 45895 27479 45929
rect 27537 45917 27571 45951
rect 27733 45917 27767 45951
rect 27823 45927 27857 45961
rect 28273 45917 28307 45951
rect 28457 45917 28491 45951
rect 29837 45917 29871 45951
rect 30481 45917 30515 45951
rect 30757 45917 30791 45951
rect 31769 45917 31803 45951
rect 32045 45917 32079 45951
rect 33241 45917 33275 45951
rect 33334 45917 33368 45951
rect 35633 45917 35667 45951
rect 35725 45917 35759 45951
rect 35909 45917 35943 45951
rect 36001 45917 36035 45951
rect 36645 45917 36679 45951
rect 37473 45917 37507 45951
rect 38313 45917 38347 45951
rect 38589 45917 38623 45951
rect 39129 45917 39163 45951
rect 20637 45849 20671 45883
rect 22937 45849 22971 45883
rect 23121 45849 23155 45883
rect 26341 45849 26375 45883
rect 27261 45849 27295 45883
rect 30665 45849 30699 45883
rect 34161 45849 34195 45883
rect 34345 45849 34379 45883
rect 10057 45781 10091 45815
rect 21741 45781 21775 45815
rect 22293 45781 22327 45815
rect 33977 45781 34011 45815
rect 35449 45781 35483 45815
rect 20729 45577 20763 45611
rect 23121 45577 23155 45611
rect 26249 45577 26283 45611
rect 27537 45577 27571 45611
rect 28089 45577 28123 45611
rect 30757 45577 30791 45611
rect 17785 45509 17819 45543
rect 19717 45509 19751 45543
rect 25881 45509 25915 45543
rect 25973 45509 26007 45543
rect 27169 45509 27203 45543
rect 31677 45509 31711 45543
rect 33425 45509 33459 45543
rect 33793 45509 33827 45543
rect 33931 45509 33965 45543
rect 34529 45509 34563 45543
rect 38393 45509 38427 45543
rect 18521 45441 18555 45475
rect 20726 45441 20760 45475
rect 22201 45441 22235 45475
rect 23397 45441 23431 45475
rect 24133 45441 24167 45475
rect 24777 45441 24811 45475
rect 24961 45441 24995 45475
rect 25763 45441 25797 45475
rect 26065 45441 26099 45475
rect 27353 45441 27387 45475
rect 27629 45441 27663 45475
rect 28457 45441 28491 45475
rect 29285 45441 29319 45475
rect 29561 45441 29595 45475
rect 30389 45441 30423 45475
rect 31309 45441 31343 45475
rect 31493 45441 31527 45475
rect 31769 45441 31803 45475
rect 32321 45441 32355 45475
rect 32413 45441 32447 45475
rect 32597 45441 32631 45475
rect 32689 45441 32723 45475
rect 33609 45441 33643 45475
rect 33701 45441 33735 45475
rect 35265 45441 35299 45475
rect 35449 45441 35483 45475
rect 35541 45441 35575 45475
rect 36001 45441 36035 45475
rect 36093 45441 36127 45475
rect 36277 45441 36311 45475
rect 37657 45441 37691 45475
rect 38668 45441 38702 45475
rect 38761 45441 38795 45475
rect 39865 45441 39899 45475
rect 41153 45441 41187 45475
rect 19165 45373 19199 45407
rect 21189 45373 21223 45407
rect 22017 45373 22051 45407
rect 23305 45373 23339 45407
rect 23489 45373 23523 45407
rect 23581 45373 23615 45407
rect 25605 45373 25639 45407
rect 28549 45373 28583 45407
rect 29101 45373 29135 45407
rect 29469 45373 29503 45407
rect 30481 45373 30515 45407
rect 34069 45373 34103 45407
rect 37473 45373 37507 45407
rect 37933 45373 37967 45407
rect 39221 45373 39255 45407
rect 40509 45373 40543 45407
rect 25145 45305 25179 45339
rect 29377 45305 29411 45339
rect 36461 45305 36495 45339
rect 19993 45237 20027 45271
rect 20545 45237 20579 45271
rect 21097 45237 21131 45271
rect 22385 45237 22419 45271
rect 24317 45237 24351 45271
rect 32873 45237 32907 45271
rect 35081 45237 35115 45271
rect 37841 45237 37875 45271
rect 19901 45033 19935 45067
rect 22569 45033 22603 45067
rect 25973 45033 26007 45067
rect 31309 45033 31343 45067
rect 33149 45033 33183 45067
rect 33977 45033 34011 45067
rect 37105 45033 37139 45067
rect 38025 45033 38059 45067
rect 39313 45033 39347 45067
rect 40049 45033 40083 45067
rect 40785 45033 40819 45067
rect 23489 44965 23523 44999
rect 28733 44965 28767 44999
rect 30573 44965 30607 44999
rect 31401 44965 31435 44999
rect 34897 44965 34931 44999
rect 20545 44897 20579 44931
rect 21649 44897 21683 44931
rect 23765 44897 23799 44931
rect 31769 44897 31803 44931
rect 32873 44897 32907 44931
rect 36093 44897 36127 44931
rect 37473 44897 37507 44931
rect 38669 44897 38703 44931
rect 20085 44829 20119 44863
rect 20729 44829 20763 44863
rect 21373 44829 21407 44863
rect 22569 44829 22603 44863
rect 22753 44829 22787 44863
rect 22845 44829 22879 44863
rect 24593 44829 24627 44863
rect 24685 44829 24719 44863
rect 24869 44829 24903 44863
rect 24961 44829 24995 44863
rect 25881 44829 25915 44863
rect 27077 44829 27111 44863
rect 27353 44829 27387 44863
rect 27997 44829 28031 44863
rect 28089 44829 28123 44863
rect 28181 44829 28215 44863
rect 28733 44829 28767 44863
rect 29009 44829 29043 44863
rect 29959 44829 29993 44863
rect 30113 44829 30147 44863
rect 30757 44829 30791 44863
rect 30849 44829 30883 44863
rect 32781 44829 32815 44863
rect 33885 44829 33919 44863
rect 35081 44829 35115 44863
rect 35265 44829 35299 44863
rect 35357 44829 35391 44863
rect 36185 44829 36219 44863
rect 37381 44829 37415 44863
rect 38209 44829 38243 44863
rect 25145 44761 25179 44795
rect 28917 44761 28951 44795
rect 30573 44761 30607 44795
rect 18889 44693 18923 44727
rect 20913 44693 20947 44727
rect 23305 44693 23339 44727
rect 26341 44693 26375 44727
rect 26893 44693 26927 44727
rect 27261 44693 27295 44727
rect 27813 44693 27847 44727
rect 29745 44693 29779 44727
rect 34345 44693 34379 44727
rect 35909 44693 35943 44727
rect 36553 44693 36587 44727
rect 20269 44489 20303 44523
rect 21005 44489 21039 44523
rect 22753 44489 22787 44523
rect 23765 44489 23799 44523
rect 25697 44489 25731 44523
rect 28273 44489 28307 44523
rect 32321 44489 32355 44523
rect 33701 44489 33735 44523
rect 35081 44489 35115 44523
rect 36461 44489 36495 44523
rect 37473 44489 37507 44523
rect 38393 44489 38427 44523
rect 26525 44421 26559 44455
rect 33149 44421 33183 44455
rect 33885 44421 33919 44455
rect 20821 44353 20855 44387
rect 22569 44353 22603 44387
rect 23397 44353 23431 44387
rect 24685 44353 24719 44387
rect 24777 44353 24811 44387
rect 25329 44353 25363 44387
rect 25513 44353 25547 44387
rect 26341 44353 26375 44387
rect 26617 44353 26651 44387
rect 27813 44353 27847 44387
rect 27905 44353 27939 44387
rect 29101 44353 29135 44387
rect 32505 44353 32539 44387
rect 34069 44353 34103 44387
rect 34713 44353 34747 44387
rect 35541 44353 35575 44387
rect 36645 44353 36679 44387
rect 36737 44375 36771 44409
rect 36829 44353 36863 44387
rect 37657 44353 37691 44387
rect 23305 44285 23339 44319
rect 26157 44285 26191 44319
rect 29193 44285 29227 44319
rect 30205 44285 30239 44319
rect 31401 44285 31435 44319
rect 31585 44285 31619 44319
rect 32689 44285 32723 44319
rect 34621 44285 34655 44319
rect 36001 44285 36035 44319
rect 37933 44285 37967 44319
rect 22109 44217 22143 44251
rect 28733 44217 28767 44251
rect 37841 44217 37875 44251
rect 19809 44149 19843 44183
rect 24501 44149 24535 44183
rect 27629 44149 27663 44183
rect 35633 44149 35667 44183
rect 20453 43945 20487 43979
rect 22201 43945 22235 43979
rect 23305 43945 23339 43979
rect 23765 43945 23799 43979
rect 25789 43945 25823 43979
rect 26525 43945 26559 43979
rect 27537 43945 27571 43979
rect 30205 43945 30239 43979
rect 30849 43945 30883 43979
rect 32229 43945 32263 43979
rect 33609 43945 33643 43979
rect 35541 43945 35575 43979
rect 35725 43945 35759 43979
rect 36185 43945 36219 43979
rect 36829 43945 36863 43979
rect 21557 43877 21591 43911
rect 29837 43877 29871 43911
rect 31309 43877 31343 43911
rect 25053 43809 25087 43843
rect 25329 43809 25363 43843
rect 26709 43809 26743 43843
rect 27905 43809 27939 43843
rect 29009 43809 29043 43843
rect 29745 43809 29779 43843
rect 34069 43809 34103 43843
rect 21741 43741 21775 43775
rect 22385 43741 22419 43775
rect 23121 43741 23155 43775
rect 23305 43741 23339 43775
rect 23765 43741 23799 43775
rect 24041 43741 24075 43775
rect 24961 43741 24995 43775
rect 26801 43741 26835 43775
rect 27445 43741 27479 43775
rect 28825 43741 28859 43775
rect 30021 43741 30055 43775
rect 32597 43741 32631 43775
rect 33333 43741 33367 43775
rect 33425 43741 33459 43775
rect 33609 43741 33643 43775
rect 19901 43673 19935 43707
rect 32413 43673 32447 43707
rect 35357 43673 35391 43707
rect 35573 43673 35607 43707
rect 21097 43605 21131 43639
rect 23949 43605 23983 43639
rect 21189 43401 21223 43435
rect 23857 43401 23891 43435
rect 24501 43401 24535 43435
rect 25605 43401 25639 43435
rect 27429 43401 27463 43435
rect 28181 43401 28215 43435
rect 33793 43401 33827 43435
rect 35081 43401 35115 43435
rect 24685 43333 24719 43367
rect 27629 43333 27663 43367
rect 22477 43265 22511 43299
rect 23305 43265 23339 43299
rect 23765 43265 23799 43299
rect 23949 43265 23983 43299
rect 24869 43265 24903 43299
rect 25513 43265 25547 43299
rect 25789 43265 25823 43299
rect 26341 43265 26375 43299
rect 28273 43265 28307 43299
rect 29377 43265 29411 43299
rect 30021 43265 30055 43299
rect 31309 43265 31343 43299
rect 32965 43265 32999 43299
rect 33609 43265 33643 43299
rect 34897 43265 34931 43299
rect 35541 43265 35575 43299
rect 28733 43197 28767 43231
rect 32321 43197 32355 43231
rect 34253 43197 34287 43231
rect 25789 43129 25823 43163
rect 27261 43129 27295 43163
rect 27445 43061 27479 43095
rect 30665 43061 30699 43095
rect 25329 42857 25363 42891
rect 26157 42857 26191 42891
rect 26801 42857 26835 42891
rect 27905 42857 27939 42891
rect 33425 42857 33459 42891
rect 22845 42721 22879 42755
rect 24685 42721 24719 42755
rect 27261 42721 27295 42755
rect 28549 42721 28583 42755
rect 32229 42721 32263 42755
rect 28089 42653 28123 42687
rect 30389 42653 30423 42687
rect 29745 42585 29779 42619
rect 21925 42517 21959 42551
rect 23489 42517 23523 42551
rect 24041 42517 24075 42551
rect 24777 42313 24811 42347
rect 27169 42313 27203 42347
rect 27721 42313 27755 42347
rect 29009 42313 29043 42347
rect 29469 42313 29503 42347
rect 28457 42245 28491 42279
rect 23765 42041 23799 42075
rect 27813 41769 27847 41803
rect 25145 7497 25179 7531
rect 24501 7361 24535 7395
rect 26525 7361 26559 7395
rect 23121 7157 23155 7191
rect 23765 7157 23799 7191
rect 24593 7157 24627 7191
rect 25697 7157 25731 7191
rect 26433 7157 26467 7191
rect 25329 6817 25363 6851
rect 21189 6749 21223 6783
rect 22293 6749 22327 6783
rect 22937 6749 22971 6783
rect 23857 6749 23891 6783
rect 25145 6749 25179 6783
rect 26249 6749 26283 6783
rect 26709 6749 26743 6783
rect 27629 6749 27663 6783
rect 28457 6749 28491 6783
rect 22385 6613 22419 6647
rect 23029 6613 23063 6647
rect 23949 6613 23983 6647
rect 24685 6613 24719 6647
rect 28365 6613 28399 6647
rect 24501 6341 24535 6375
rect 27721 6341 27755 6375
rect 21281 6273 21315 6307
rect 27537 6273 27571 6307
rect 21373 6205 21407 6239
rect 23857 6205 23891 6239
rect 24317 6205 24351 6239
rect 24961 6205 24995 6239
rect 29193 6205 29227 6239
rect 22937 6137 22971 6171
rect 18981 6069 19015 6103
rect 19533 6069 19567 6103
rect 20269 6069 20303 6103
rect 22293 6069 22327 6103
rect 21465 5729 21499 5763
rect 22201 5729 22235 5763
rect 22385 5729 22419 5763
rect 22937 5729 22971 5763
rect 27629 5729 27663 5763
rect 18705 5661 18739 5695
rect 19993 5661 20027 5695
rect 20821 5661 20855 5695
rect 21281 5661 21315 5695
rect 24869 5661 24903 5695
rect 28089 5661 28123 5695
rect 28917 5661 28951 5695
rect 29929 5661 29963 5695
rect 25145 5593 25179 5627
rect 25789 5593 25823 5627
rect 27445 5593 27479 5627
rect 28181 5593 28215 5627
rect 19441 5525 19475 5559
rect 20085 5525 20119 5559
rect 29837 5525 29871 5559
rect 22293 5253 22327 5287
rect 24593 5253 24627 5287
rect 29653 5253 29687 5287
rect 18981 5185 19015 5219
rect 19625 5185 19659 5219
rect 22109 5185 22143 5219
rect 29009 5185 29043 5219
rect 19809 5117 19843 5151
rect 21373 5117 21407 5151
rect 23489 5117 23523 5151
rect 24409 5117 24443 5151
rect 25237 5117 25271 5151
rect 27813 5117 27847 5151
rect 28825 5117 28859 5151
rect 29469 5117 29503 5151
rect 30021 5117 30055 5151
rect 18521 5049 18555 5083
rect 17049 4981 17083 5015
rect 17877 4981 17911 5015
rect 19073 4981 19107 5015
rect 27997 4777 28031 4811
rect 29745 4777 29779 4811
rect 17601 4641 17635 4675
rect 19901 4641 19935 4675
rect 20085 4641 20119 4675
rect 21097 4641 21131 4675
rect 22201 4641 22235 4675
rect 22385 4641 22419 4675
rect 23581 4641 23615 4675
rect 25605 4641 25639 4675
rect 26341 4641 26375 4675
rect 30573 4641 30607 4675
rect 15117 4573 15151 4607
rect 15945 4573 15979 4607
rect 16957 4573 16991 4607
rect 18061 4573 18095 4607
rect 18889 4573 18923 4607
rect 24961 4573 24995 4607
rect 27905 4573 27939 4607
rect 28733 4573 28767 4607
rect 31217 4573 31251 4607
rect 31861 4573 31895 4607
rect 32321 4573 32355 4607
rect 25053 4505 25087 4539
rect 25789 4505 25823 4539
rect 31769 4437 31803 4471
rect 17049 4097 17083 4131
rect 17693 4097 17727 4131
rect 18337 4097 18371 4131
rect 19625 4097 19659 4131
rect 23673 4097 23707 4131
rect 29009 4097 29043 4131
rect 31309 4097 31343 4131
rect 32505 4097 32539 4131
rect 15669 4029 15703 4063
rect 18429 4029 18463 4063
rect 19809 4029 19843 4063
rect 21465 4029 21499 4063
rect 22385 4029 22419 4063
rect 24133 4029 24167 4063
rect 24317 4029 24351 4063
rect 24685 4029 24719 4063
rect 27445 4029 27479 4063
rect 28825 4029 28859 4063
rect 29469 4029 29503 4063
rect 31125 4029 31159 4063
rect 32965 4029 32999 4063
rect 16313 3961 16347 3995
rect 34897 3961 34931 3995
rect 12357 3893 12391 3927
rect 13185 3893 13219 3927
rect 14013 3893 14047 3927
rect 15025 3893 15059 3927
rect 17141 3893 17175 3927
rect 17785 3893 17819 3927
rect 19165 3893 19199 3927
rect 23029 3893 23063 3927
rect 26433 3893 26467 3927
rect 32413 3893 32447 3927
rect 33609 3893 33643 3927
rect 34253 3893 34287 3927
rect 35541 3893 35575 3927
rect 47777 3893 47811 3927
rect 16865 3689 16899 3723
rect 18797 3689 18831 3723
rect 20361 3689 20395 3723
rect 27905 3689 27939 3723
rect 33333 3689 33367 3723
rect 15025 3621 15059 3655
rect 34897 3621 34931 3655
rect 36185 3621 36219 3655
rect 38117 3621 38151 3655
rect 41337 3621 41371 3655
rect 47133 3621 47167 3655
rect 15669 3553 15703 3587
rect 17601 3553 17635 3587
rect 21557 3553 21591 3587
rect 21741 3553 21775 3587
rect 22201 3553 22235 3587
rect 25513 3553 25547 3587
rect 26065 3553 26099 3587
rect 31585 3553 31619 3587
rect 35541 3553 35575 3587
rect 36829 3553 36863 3587
rect 41981 3553 42015 3587
rect 47777 3553 47811 3587
rect 4353 3485 4387 3519
rect 4997 3485 5031 3519
rect 5825 3485 5859 3519
rect 6653 3485 6687 3519
rect 7481 3485 7515 3519
rect 8309 3485 8343 3519
rect 9137 3485 9171 3519
rect 9965 3485 9999 3519
rect 10793 3485 10827 3519
rect 11621 3485 11655 3519
rect 12449 3485 12483 3519
rect 13093 3485 13127 3519
rect 13737 3485 13771 3519
rect 16129 3485 16163 3519
rect 16773 3485 16807 3519
rect 18245 3485 18279 3519
rect 18705 3485 18739 3519
rect 19809 3485 19843 3519
rect 20269 3485 20303 3519
rect 20913 3485 20947 3519
rect 24041 3485 24075 3519
rect 24869 3485 24903 3519
rect 27813 3485 27847 3519
rect 28641 3485 28675 3519
rect 32229 3485 32263 3519
rect 32689 3485 32723 3519
rect 33977 3485 34011 3519
rect 37473 3485 37507 3519
rect 38761 3485 38795 3519
rect 40049 3485 40083 3519
rect 40693 3485 40727 3519
rect 42717 3485 42751 3519
rect 43361 3485 43395 3519
rect 45201 3485 45235 3519
rect 45845 3485 45879 3519
rect 46489 3485 46523 3519
rect 18153 3417 18187 3451
rect 24961 3417 24995 3451
rect 25697 3417 25731 3451
rect 29745 3417 29779 3451
rect 31401 3417 31435 3451
rect 16221 3349 16255 3383
rect 21005 3349 21039 3383
rect 23949 3349 23983 3383
rect 32137 3349 32171 3383
rect 17509 3077 17543 3111
rect 22661 3077 22695 3111
rect 24961 3077 24995 3111
rect 28825 3077 28859 3111
rect 31125 3077 31159 3111
rect 13093 3009 13127 3043
rect 15025 3009 15059 3043
rect 16129 3009 16163 3043
rect 19625 3009 19659 3043
rect 22477 3009 22511 3043
rect 24777 3009 24811 3043
rect 29009 3009 29043 3043
rect 33609 3009 33643 3043
rect 35541 3009 35575 3043
rect 37473 3009 37507 3043
rect 4077 2941 4111 2975
rect 5365 2941 5399 2975
rect 14381 2941 14415 2975
rect 17325 2941 17359 2975
rect 18981 2941 19015 2975
rect 19809 2941 19843 2975
rect 21465 2941 21499 2975
rect 24317 2941 24351 2975
rect 25513 2941 25547 2975
rect 27169 2941 27203 2975
rect 29469 2941 29503 2975
rect 31309 2941 31343 2975
rect 32965 2941 32999 2975
rect 38761 2941 38795 2975
rect 40693 2941 40727 2975
rect 43269 2941 43303 2975
rect 45201 2941 45235 2975
rect 12449 2873 12483 2907
rect 15669 2873 15703 2907
rect 34253 2873 34287 2907
rect 36185 2873 36219 2907
rect 38117 2873 38151 2907
rect 39405 2873 39439 2907
rect 41337 2873 41371 2907
rect 43913 2873 43947 2907
rect 45845 2873 45879 2907
rect 3433 2805 3467 2839
rect 4721 2805 4755 2839
rect 6009 2805 6043 2839
rect 7297 2805 7331 2839
rect 7941 2805 7975 2839
rect 8585 2805 8619 2839
rect 9229 2805 9263 2839
rect 9873 2805 9907 2839
rect 10517 2805 10551 2839
rect 11161 2805 11195 2839
rect 13737 2805 13771 2839
rect 16221 2805 16255 2839
rect 32321 2805 32355 2839
rect 34897 2805 34931 2839
rect 40049 2805 40083 2839
rect 42625 2805 42659 2839
rect 44557 2805 44591 2839
rect 46489 2805 46523 2839
rect 47777 2805 47811 2839
rect 13737 2601 13771 2635
rect 32413 2601 32447 2635
rect 33057 2601 33091 2635
rect 33609 2601 33643 2635
rect 34897 2601 34931 2635
rect 36185 2601 36219 2635
rect 37473 2601 37507 2635
rect 5365 2533 5399 2567
rect 7297 2533 7331 2567
rect 9873 2533 9907 2567
rect 12449 2533 12483 2567
rect 40049 2533 40083 2567
rect 43913 2533 43947 2567
rect 46489 2533 46523 2567
rect 4721 2465 4755 2499
rect 8585 2465 8619 2499
rect 11161 2465 11195 2499
rect 13093 2465 13127 2499
rect 17233 2465 17267 2499
rect 19809 2465 19843 2499
rect 21465 2465 21499 2499
rect 25789 2465 25823 2499
rect 26433 2465 26467 2499
rect 26617 2465 26651 2499
rect 28825 2465 28859 2499
rect 29009 2465 29043 2499
rect 31585 2465 31619 2499
rect 38761 2465 38795 2499
rect 40693 2465 40727 2499
rect 42625 2465 42659 2499
rect 45201 2465 45235 2499
rect 2145 2397 2179 2431
rect 2789 2397 2823 2431
rect 3433 2397 3467 2431
rect 6009 2397 6043 2431
rect 7941 2397 7975 2431
rect 10517 2397 10551 2431
rect 15025 2397 15059 2431
rect 15669 2397 15703 2431
rect 16313 2397 16347 2431
rect 17049 2397 17083 2431
rect 19625 2397 19659 2431
rect 22201 2397 22235 2431
rect 32505 2397 32539 2431
rect 32965 2397 32999 2431
rect 35541 2397 35575 2431
rect 38117 2397 38151 2431
rect 41337 2397 41371 2431
rect 43269 2397 43303 2431
rect 45845 2397 45879 2431
rect 47777 2397 47811 2431
rect 18889 2329 18923 2363
rect 22385 2329 22419 2363
rect 24041 2329 24075 2363
rect 27169 2329 27203 2363
rect 29745 2329 29779 2363
rect 31401 2329 31435 2363
<< metal1 >>
rect 10962 47812 10968 47864
rect 11020 47852 11026 47864
rect 20714 47852 20720 47864
rect 11020 47824 20720 47852
rect 11020 47812 11026 47824
rect 20714 47812 20720 47824
rect 20772 47812 20778 47864
rect 15378 47744 15384 47796
rect 15436 47784 15442 47796
rect 23382 47784 23388 47796
rect 15436 47756 23388 47784
rect 15436 47744 15442 47756
rect 23382 47744 23388 47756
rect 23440 47744 23446 47796
rect 18874 47608 18880 47660
rect 18932 47648 18938 47660
rect 20898 47648 20904 47660
rect 18932 47620 20904 47648
rect 18932 47608 18938 47620
rect 20898 47608 20904 47620
rect 20956 47608 20962 47660
rect 23658 47608 23664 47660
rect 23716 47648 23722 47660
rect 25682 47648 25688 47660
rect 23716 47620 25688 47648
rect 23716 47608 23722 47620
rect 25682 47608 25688 47620
rect 25740 47608 25746 47660
rect 14550 47540 14556 47592
rect 14608 47580 14614 47592
rect 20346 47580 20352 47592
rect 14608 47552 20352 47580
rect 14608 47540 14614 47552
rect 20346 47540 20352 47552
rect 20404 47540 20410 47592
rect 13170 47472 13176 47524
rect 13228 47512 13234 47524
rect 21450 47512 21456 47524
rect 13228 47484 21456 47512
rect 13228 47472 13234 47484
rect 21450 47472 21456 47484
rect 21508 47472 21514 47524
rect 23750 47472 23756 47524
rect 23808 47512 23814 47524
rect 30282 47512 30288 47524
rect 23808 47484 30288 47512
rect 23808 47472 23814 47484
rect 30282 47472 30288 47484
rect 30340 47472 30346 47524
rect 37826 47472 37832 47524
rect 37884 47512 37890 47524
rect 38378 47512 38384 47524
rect 37884 47484 38384 47512
rect 37884 47472 37890 47484
rect 38378 47472 38384 47484
rect 38436 47472 38442 47524
rect 11698 47404 11704 47456
rect 11756 47444 11762 47456
rect 17770 47444 17776 47456
rect 11756 47416 17776 47444
rect 11756 47404 11762 47416
rect 17770 47404 17776 47416
rect 17828 47404 17834 47456
rect 18138 47404 18144 47456
rect 18196 47444 18202 47456
rect 24026 47444 24032 47456
rect 18196 47416 24032 47444
rect 18196 47404 18202 47416
rect 24026 47404 24032 47416
rect 24084 47444 24090 47456
rect 29822 47444 29828 47456
rect 24084 47416 29828 47444
rect 24084 47404 24090 47416
rect 29822 47404 29828 47416
rect 29880 47404 29886 47456
rect 30006 47404 30012 47456
rect 30064 47444 30070 47456
rect 43438 47444 43444 47456
rect 30064 47416 43444 47444
rect 30064 47404 30070 47416
rect 43438 47404 43444 47416
rect 43496 47404 43502 47456
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 5074 47200 5080 47252
rect 5132 47240 5138 47252
rect 5445 47243 5503 47249
rect 5445 47240 5457 47243
rect 5132 47212 5457 47240
rect 5132 47200 5138 47212
rect 5445 47209 5457 47212
rect 5491 47209 5503 47243
rect 7282 47240 7288 47252
rect 7243 47212 7288 47240
rect 5445 47203 5503 47209
rect 7282 47200 7288 47212
rect 7340 47200 7346 47252
rect 7926 47240 7932 47252
rect 7887 47212 7932 47240
rect 7926 47200 7932 47212
rect 7984 47200 7990 47252
rect 8386 47240 8392 47252
rect 8347 47212 8392 47240
rect 8386 47200 8392 47212
rect 8444 47200 8450 47252
rect 9674 47240 9680 47252
rect 9635 47212 9680 47240
rect 9674 47200 9680 47212
rect 9732 47200 9738 47252
rect 10778 47240 10784 47252
rect 10739 47212 10784 47240
rect 10778 47200 10784 47212
rect 10836 47200 10842 47252
rect 11882 47240 11888 47252
rect 11843 47212 11888 47240
rect 11882 47200 11888 47212
rect 11940 47200 11946 47252
rect 12986 47240 12992 47252
rect 12947 47212 12992 47240
rect 12986 47200 12992 47212
rect 13044 47200 13050 47252
rect 13906 47200 13912 47252
rect 13964 47240 13970 47252
rect 14369 47243 14427 47249
rect 14369 47240 14381 47243
rect 13964 47212 14381 47240
rect 13964 47200 13970 47212
rect 14369 47209 14381 47212
rect 14415 47209 14427 47243
rect 15194 47240 15200 47252
rect 15155 47212 15200 47240
rect 14369 47203 14427 47209
rect 15194 47200 15200 47212
rect 15252 47200 15258 47252
rect 16114 47240 16120 47252
rect 16075 47212 16120 47240
rect 16114 47200 16120 47212
rect 16172 47200 16178 47252
rect 17218 47240 17224 47252
rect 17179 47212 17224 47240
rect 17218 47200 17224 47212
rect 17276 47200 17282 47252
rect 17957 47243 18015 47249
rect 17957 47209 17969 47243
rect 18003 47240 18015 47243
rect 19426 47240 19432 47252
rect 18003 47212 19432 47240
rect 18003 47209 18015 47212
rect 17957 47203 18015 47209
rect 19426 47200 19432 47212
rect 19484 47200 19490 47252
rect 21361 47243 21419 47249
rect 21361 47209 21373 47243
rect 21407 47240 21419 47243
rect 22738 47240 22744 47252
rect 21407 47212 22744 47240
rect 21407 47209 21419 47212
rect 21361 47203 21419 47209
rect 22738 47200 22744 47212
rect 22796 47200 22802 47252
rect 23382 47240 23388 47252
rect 23343 47212 23388 47240
rect 23382 47200 23388 47212
rect 23440 47200 23446 47252
rect 23842 47200 23848 47252
rect 23900 47240 23906 47252
rect 24765 47243 24823 47249
rect 24765 47240 24777 47243
rect 23900 47212 24777 47240
rect 23900 47200 23906 47212
rect 24765 47209 24777 47212
rect 24811 47209 24823 47243
rect 24765 47203 24823 47209
rect 26050 47200 26056 47252
rect 26108 47240 26114 47252
rect 26421 47243 26479 47249
rect 26421 47240 26433 47243
rect 26108 47212 26433 47240
rect 26108 47200 26114 47212
rect 26421 47209 26433 47212
rect 26467 47209 26479 47243
rect 26421 47203 26479 47209
rect 35434 47200 35440 47252
rect 35492 47240 35498 47252
rect 42705 47243 42763 47249
rect 42705 47240 42717 47243
rect 35492 47212 42717 47240
rect 35492 47200 35498 47212
rect 42705 47209 42717 47212
rect 42751 47209 42763 47243
rect 43438 47240 43444 47252
rect 43399 47212 43444 47240
rect 42705 47203 42763 47209
rect 43438 47200 43444 47212
rect 43496 47200 43502 47252
rect 44266 47240 44272 47252
rect 44227 47212 44272 47240
rect 44266 47200 44272 47212
rect 44324 47200 44330 47252
rect 45922 47200 45928 47252
rect 45980 47240 45986 47252
rect 46661 47243 46719 47249
rect 46661 47240 46673 47243
rect 45980 47212 46673 47240
rect 45980 47200 45986 47212
rect 46661 47209 46673 47212
rect 46707 47209 46719 47243
rect 46661 47203 46719 47209
rect 18693 47175 18751 47181
rect 12406 47144 18276 47172
rect 4062 47104 4068 47116
rect 4023 47076 4068 47104
rect 4062 47064 4068 47076
rect 4120 47064 4126 47116
rect 4341 47107 4399 47113
rect 4341 47073 4353 47107
rect 4387 47104 4399 47107
rect 11698 47104 11704 47116
rect 4387 47076 11704 47104
rect 4387 47073 4399 47076
rect 4341 47067 4399 47073
rect 11698 47064 11704 47076
rect 11756 47064 11762 47116
rect 5626 47036 5632 47048
rect 5587 47008 5632 47036
rect 5626 46996 5632 47008
rect 5684 46996 5690 47048
rect 9858 47036 9864 47048
rect 9819 47008 9864 47036
rect 9858 46996 9864 47008
rect 9916 46996 9922 47048
rect 10962 47036 10968 47048
rect 10923 47008 10968 47036
rect 10962 46996 10968 47008
rect 11020 46996 11026 47048
rect 12069 47039 12127 47045
rect 12069 47005 12081 47039
rect 12115 47005 12127 47039
rect 12069 46999 12127 47005
rect 12084 46968 12112 46999
rect 12406 46968 12434 47144
rect 18046 47104 18052 47116
rect 16316 47076 18052 47104
rect 13170 47036 13176 47048
rect 13131 47008 13176 47036
rect 13170 46996 13176 47008
rect 13228 46996 13234 47048
rect 14550 47036 14556 47048
rect 14511 47008 14556 47036
rect 14550 46996 14556 47008
rect 14608 46996 14614 47048
rect 15378 47036 15384 47048
rect 15339 47008 15384 47036
rect 15378 46996 15384 47008
rect 15436 46996 15442 47048
rect 16316 47045 16344 47076
rect 18046 47064 18052 47076
rect 18104 47064 18110 47116
rect 16301 47039 16359 47045
rect 16301 47005 16313 47039
rect 16347 47005 16359 47039
rect 16301 46999 16359 47005
rect 17405 47039 17463 47045
rect 17405 47005 17417 47039
rect 17451 47036 17463 47039
rect 18138 47036 18144 47048
rect 17451 47008 17816 47036
rect 18099 47008 18144 47036
rect 17451 47005 17463 47008
rect 17405 46999 17463 47005
rect 12084 46940 12434 46968
rect 17788 46900 17816 47008
rect 18138 46996 18144 47008
rect 18196 46996 18202 47048
rect 18248 46968 18276 47144
rect 18693 47141 18705 47175
rect 18739 47172 18751 47175
rect 20717 47175 20775 47181
rect 18739 47144 20208 47172
rect 18739 47141 18751 47144
rect 18693 47135 18751 47141
rect 18322 47064 18328 47116
rect 18380 47104 18386 47116
rect 18380 47076 19012 47104
rect 18380 47064 18386 47076
rect 18874 47036 18880 47048
rect 18835 47008 18880 47036
rect 18874 46996 18880 47008
rect 18932 46996 18938 47048
rect 18984 47036 19012 47076
rect 19334 47064 19340 47116
rect 19392 47104 19398 47116
rect 19521 47107 19579 47113
rect 19521 47104 19533 47107
rect 19392 47076 19533 47104
rect 19392 47064 19398 47076
rect 19521 47073 19533 47076
rect 19567 47073 19579 47107
rect 20180 47104 20208 47144
rect 20717 47141 20729 47175
rect 20763 47172 20775 47175
rect 26786 47172 26792 47184
rect 20763 47144 26792 47172
rect 20763 47141 20775 47144
rect 20717 47135 20775 47141
rect 26786 47132 26792 47144
rect 26844 47132 26850 47184
rect 35986 47132 35992 47184
rect 36044 47172 36050 47184
rect 41325 47175 41383 47181
rect 41325 47172 41337 47175
rect 36044 47144 41337 47172
rect 36044 47132 36050 47144
rect 41325 47141 41337 47144
rect 41371 47141 41383 47175
rect 41325 47135 41383 47141
rect 21634 47104 21640 47116
rect 20180 47076 21640 47104
rect 19521 47067 19579 47073
rect 21634 47064 21640 47076
rect 21692 47064 21698 47116
rect 23198 47064 23204 47116
rect 23256 47104 23262 47116
rect 23661 47107 23719 47113
rect 23661 47104 23673 47107
rect 23256 47076 23673 47104
rect 23256 47064 23262 47076
rect 23661 47073 23673 47076
rect 23707 47073 23719 47107
rect 23661 47067 23719 47073
rect 23842 47064 23848 47116
rect 23900 47104 23906 47116
rect 31389 47107 31447 47113
rect 23900 47076 24440 47104
rect 23900 47064 23906 47076
rect 19429 47039 19487 47045
rect 19429 47036 19441 47039
rect 18984 47008 19441 47036
rect 19429 47005 19441 47008
rect 19475 47005 19487 47039
rect 19429 46999 19487 47005
rect 19948 47039 20006 47045
rect 19948 47005 19960 47039
rect 19994 47036 20006 47039
rect 20254 47036 20260 47048
rect 19994 47008 20260 47036
rect 19994 47005 20006 47008
rect 19948 46999 20006 47005
rect 20254 46996 20260 47008
rect 20312 46996 20318 47048
rect 21082 46996 21088 47048
rect 21140 47036 21146 47048
rect 21177 47039 21235 47045
rect 21177 47036 21189 47039
rect 21140 47008 21189 47036
rect 21140 46996 21146 47008
rect 21177 47005 21189 47008
rect 21223 47005 21235 47039
rect 22005 47039 22063 47045
rect 22005 47036 22017 47039
rect 21177 46999 21235 47005
rect 21284 47008 22017 47036
rect 18248 46940 20116 46968
rect 18690 46900 18696 46912
rect 17788 46872 18696 46900
rect 18690 46860 18696 46872
rect 18748 46860 18754 46912
rect 19426 46860 19432 46912
rect 19484 46900 19490 46912
rect 20088 46909 20116 46940
rect 20438 46928 20444 46980
rect 20496 46968 20502 46980
rect 21284 46968 21312 47008
rect 22005 47005 22017 47008
rect 22051 47005 22063 47039
rect 22005 46999 22063 47005
rect 22094 46996 22100 47048
rect 22152 47036 22158 47048
rect 22189 47039 22247 47045
rect 22189 47036 22201 47039
rect 22152 47008 22201 47036
rect 22152 46996 22158 47008
rect 22189 47005 22201 47008
rect 22235 47005 22247 47039
rect 22189 46999 22247 47005
rect 22373 47039 22431 47045
rect 22373 47005 22385 47039
rect 22419 47005 22431 47039
rect 22373 46999 22431 47005
rect 22925 47039 22983 47045
rect 22925 47005 22937 47039
rect 22971 47036 22983 47039
rect 23290 47036 23296 47048
rect 22971 47008 23296 47036
rect 22971 47005 22983 47008
rect 22925 46999 22983 47005
rect 22388 46968 22416 46999
rect 23290 46996 23296 47008
rect 23348 46996 23354 47048
rect 23566 47036 23572 47048
rect 23527 47008 23572 47036
rect 23566 46996 23572 47008
rect 23624 46996 23630 47048
rect 23750 47036 23756 47048
rect 23711 47008 23756 47036
rect 23750 46996 23756 47008
rect 23808 46996 23814 47048
rect 24026 47036 24032 47048
rect 23987 47008 24032 47036
rect 24026 46996 24032 47008
rect 24084 46996 24090 47048
rect 24412 47036 24440 47076
rect 31389 47073 31401 47107
rect 31435 47104 31447 47107
rect 31754 47104 31760 47116
rect 31435 47076 31760 47104
rect 31435 47073 31447 47076
rect 31389 47067 31447 47073
rect 31754 47064 31760 47076
rect 31812 47064 31818 47116
rect 31938 47064 31944 47116
rect 31996 47104 32002 47116
rect 32585 47107 32643 47113
rect 32585 47104 32597 47107
rect 31996 47076 32597 47104
rect 31996 47064 32002 47076
rect 32585 47073 32597 47076
rect 32631 47073 32643 47107
rect 32585 47067 32643 47073
rect 33226 47064 33232 47116
rect 33284 47104 33290 47116
rect 33962 47104 33968 47116
rect 33284 47076 33968 47104
rect 33284 47064 33290 47076
rect 33962 47064 33968 47076
rect 34020 47064 34026 47116
rect 34057 47107 34115 47113
rect 34057 47073 34069 47107
rect 34103 47104 34115 47107
rect 34146 47104 34152 47116
rect 34103 47076 34152 47104
rect 34103 47073 34115 47076
rect 34057 47067 34115 47073
rect 34146 47064 34152 47076
rect 34204 47064 34210 47116
rect 37550 47064 37556 47116
rect 37608 47104 37614 47116
rect 37826 47104 37832 47116
rect 37608 47076 37832 47104
rect 37608 47064 37614 47076
rect 37826 47064 37832 47076
rect 37884 47064 37890 47116
rect 38657 47107 38715 47113
rect 38657 47104 38669 47107
rect 38580 47076 38669 47104
rect 24581 47039 24639 47045
rect 24412 47030 24532 47036
rect 24581 47030 24593 47039
rect 24412 47008 24593 47030
rect 24504 47005 24593 47008
rect 24627 47005 24639 47039
rect 25682 47036 25688 47048
rect 25643 47008 25688 47036
rect 24504 47002 24639 47005
rect 24581 46999 24639 47002
rect 25682 46996 25688 47008
rect 25740 46996 25746 47048
rect 25866 47036 25872 47048
rect 25827 47008 25872 47036
rect 25866 46996 25872 47008
rect 25924 46996 25930 47048
rect 25961 47039 26019 47045
rect 25961 47005 25973 47039
rect 26007 47036 26019 47039
rect 26142 47036 26148 47048
rect 26007 47008 26148 47036
rect 26007 47005 26019 47008
rect 25961 46999 26019 47005
rect 26142 46996 26148 47008
rect 26200 46996 26206 47048
rect 26418 46996 26424 47048
rect 26476 47036 26482 47048
rect 27154 47036 27160 47048
rect 26476 47008 27160 47036
rect 26476 46996 26482 47008
rect 27154 46996 27160 47008
rect 27212 46996 27218 47048
rect 27433 47039 27491 47045
rect 27433 47005 27445 47039
rect 27479 47036 27491 47039
rect 27614 47036 27620 47048
rect 27479 47008 27620 47036
rect 27479 47005 27491 47008
rect 27433 46999 27491 47005
rect 27614 46996 27620 47008
rect 27672 46996 27678 47048
rect 28997 47039 29055 47045
rect 28997 47005 29009 47039
rect 29043 47036 29055 47039
rect 29362 47036 29368 47048
rect 29043 47008 29368 47036
rect 29043 47005 29055 47008
rect 28997 46999 29055 47005
rect 29362 46996 29368 47008
rect 29420 46996 29426 47048
rect 29730 46996 29736 47048
rect 29788 47036 29794 47048
rect 29825 47039 29883 47045
rect 29825 47036 29837 47039
rect 29788 47008 29837 47036
rect 29788 46996 29794 47008
rect 29825 47005 29837 47008
rect 29871 47005 29883 47039
rect 29825 46999 29883 47005
rect 29914 46996 29920 47048
rect 29972 47036 29978 47048
rect 30101 47039 30159 47045
rect 30101 47036 30113 47039
rect 29972 47008 30113 47036
rect 29972 46996 29978 47008
rect 30101 47005 30113 47008
rect 30147 47005 30159 47039
rect 30101 46999 30159 47005
rect 32214 46996 32220 47048
rect 32272 47036 32278 47048
rect 32309 47039 32367 47045
rect 32309 47036 32321 47039
rect 32272 47008 32321 47036
rect 32272 46996 32278 47008
rect 32309 47005 32321 47008
rect 32355 47005 32367 47039
rect 33778 47036 33784 47048
rect 33739 47008 33784 47036
rect 32309 46999 32367 47005
rect 33778 46996 33784 47008
rect 33836 46996 33842 47048
rect 35897 47039 35955 47045
rect 35897 47005 35909 47039
rect 35943 47036 35955 47039
rect 36078 47036 36084 47048
rect 35943 47008 36084 47036
rect 35943 47005 35955 47008
rect 35897 46999 35955 47005
rect 36078 46996 36084 47008
rect 36136 46996 36142 47048
rect 36173 47039 36231 47045
rect 36173 47005 36185 47039
rect 36219 47005 36231 47039
rect 37642 47036 37648 47048
rect 37603 47008 37648 47036
rect 36173 46999 36231 47005
rect 24670 46968 24676 46980
rect 20496 46940 21312 46968
rect 22066 46940 24676 46968
rect 20496 46928 20502 46940
rect 19889 46903 19947 46909
rect 19889 46900 19901 46903
rect 19484 46872 19901 46900
rect 19484 46860 19490 46872
rect 19889 46869 19901 46872
rect 19935 46869 19947 46903
rect 19889 46863 19947 46869
rect 20073 46903 20131 46909
rect 20073 46869 20085 46903
rect 20119 46869 20131 46903
rect 20073 46863 20131 46869
rect 21910 46860 21916 46912
rect 21968 46900 21974 46912
rect 22066 46900 22094 46940
rect 24670 46928 24676 46940
rect 24728 46928 24734 46980
rect 29178 46968 29184 46980
rect 25332 46940 25636 46968
rect 29139 46940 29184 46968
rect 21968 46872 22094 46900
rect 21968 46860 21974 46872
rect 22922 46860 22928 46912
rect 22980 46900 22986 46912
rect 25332 46900 25360 46940
rect 25498 46900 25504 46912
rect 22980 46872 25360 46900
rect 25459 46872 25504 46900
rect 22980 46860 22986 46872
rect 25498 46860 25504 46872
rect 25556 46860 25562 46912
rect 25608 46900 25636 46940
rect 29178 46928 29184 46940
rect 29236 46928 29242 46980
rect 31573 46971 31631 46977
rect 31573 46937 31585 46971
rect 31619 46968 31631 46971
rect 31662 46968 31668 46980
rect 31619 46940 31668 46968
rect 31619 46937 31631 46940
rect 31573 46931 31631 46937
rect 31662 46928 31668 46940
rect 31720 46928 31726 46980
rect 31757 46971 31815 46977
rect 31757 46937 31769 46971
rect 31803 46968 31815 46971
rect 31846 46968 31852 46980
rect 31803 46940 31852 46968
rect 31803 46937 31815 46940
rect 31757 46931 31815 46937
rect 31846 46928 31852 46940
rect 31904 46928 31910 46980
rect 28813 46903 28871 46909
rect 28813 46900 28825 46903
rect 25608 46872 28825 46900
rect 28813 46869 28825 46872
rect 28859 46869 28871 46903
rect 28813 46863 28871 46869
rect 30834 46860 30840 46912
rect 30892 46900 30898 46912
rect 32214 46900 32220 46912
rect 30892 46872 32220 46900
rect 30892 46860 30898 46872
rect 32214 46860 32220 46872
rect 32272 46860 32278 46912
rect 33318 46860 33324 46912
rect 33376 46900 33382 46912
rect 33597 46903 33655 46909
rect 33597 46900 33609 46903
rect 33376 46872 33609 46900
rect 33376 46860 33382 46872
rect 33597 46869 33609 46872
rect 33643 46869 33655 46903
rect 33597 46863 33655 46869
rect 35342 46860 35348 46912
rect 35400 46900 35406 46912
rect 36188 46900 36216 46999
rect 37642 46996 37648 47008
rect 37700 46996 37706 47048
rect 37921 47039 37979 47045
rect 37921 47005 37933 47039
rect 37967 47005 37979 47039
rect 37921 46999 37979 47005
rect 36817 46971 36875 46977
rect 36817 46937 36829 46971
rect 36863 46968 36875 46971
rect 37274 46968 37280 46980
rect 36863 46940 37280 46968
rect 36863 46937 36875 46940
rect 36817 46931 36875 46937
rect 37274 46928 37280 46940
rect 37332 46928 37338 46980
rect 37366 46928 37372 46980
rect 37424 46968 37430 46980
rect 37936 46968 37964 46999
rect 37424 46940 37964 46968
rect 37424 46928 37430 46940
rect 38580 46934 38608 47076
rect 38657 47073 38669 47076
rect 38703 47073 38715 47107
rect 40034 47104 40040 47116
rect 39995 47076 40040 47104
rect 38657 47067 38715 47073
rect 40034 47064 40040 47076
rect 40092 47064 40098 47116
rect 41598 47064 41604 47116
rect 41656 47104 41662 47116
rect 45281 47107 45339 47113
rect 45281 47104 45293 47107
rect 41656 47076 45293 47104
rect 41656 47064 41662 47076
rect 45281 47073 45293 47076
rect 45327 47073 45339 47107
rect 45281 47067 45339 47073
rect 38838 46996 38844 47048
rect 38896 47036 38902 47048
rect 38933 47039 38991 47045
rect 38933 47036 38945 47039
rect 38896 47008 38945 47036
rect 38896 46996 38902 47008
rect 38933 47005 38945 47008
rect 38979 47005 38991 47039
rect 38933 46999 38991 47005
rect 40218 46996 40224 47048
rect 40276 47036 40282 47048
rect 40313 47039 40371 47045
rect 40313 47036 40325 47039
rect 40276 47008 40325 47036
rect 40276 46996 40282 47008
rect 40313 47005 40325 47008
rect 40359 47005 40371 47039
rect 40313 46999 40371 47005
rect 42889 47039 42947 47045
rect 42889 47005 42901 47039
rect 42935 47005 42947 47039
rect 42889 46999 42947 47005
rect 41966 46968 41972 46980
rect 41927 46940 41972 46968
rect 38580 46912 38700 46934
rect 41966 46928 41972 46940
rect 42024 46928 42030 46980
rect 42904 46968 42932 46999
rect 42978 46996 42984 47048
rect 43036 47036 43042 47048
rect 43625 47039 43683 47045
rect 43625 47036 43637 47039
rect 43036 47008 43637 47036
rect 43036 46996 43042 47008
rect 43625 47005 43637 47008
rect 43671 47036 43683 47039
rect 43806 47036 43812 47048
rect 43671 47008 43812 47036
rect 43671 47005 43683 47008
rect 43625 46999 43683 47005
rect 43806 46996 43812 47008
rect 43864 46996 43870 47048
rect 44174 46996 44180 47048
rect 44232 47036 44238 47048
rect 44453 47039 44511 47045
rect 44453 47036 44465 47039
rect 44232 47008 44465 47036
rect 44232 46996 44238 47008
rect 44453 47005 44465 47008
rect 44499 47005 44511 47039
rect 44453 46999 44511 47005
rect 45186 46996 45192 47048
rect 45244 47036 45250 47048
rect 45465 47039 45523 47045
rect 45465 47036 45477 47039
rect 45244 47008 45477 47036
rect 45244 46996 45250 47008
rect 45465 47005 45477 47008
rect 45511 47005 45523 47039
rect 45465 46999 45523 47005
rect 46017 47039 46075 47045
rect 46017 47005 46029 47039
rect 46063 47005 46075 47039
rect 46017 46999 46075 47005
rect 43254 46968 43260 46980
rect 42628 46940 43260 46968
rect 36630 46900 36636 46912
rect 35400 46872 36636 46900
rect 35400 46860 35406 46872
rect 36630 46860 36636 46872
rect 36688 46860 36694 46912
rect 36725 46903 36783 46909
rect 36725 46869 36737 46903
rect 36771 46900 36783 46903
rect 36906 46900 36912 46912
rect 36771 46872 36912 46900
rect 36771 46869 36783 46872
rect 36725 46863 36783 46869
rect 36906 46860 36912 46872
rect 36964 46860 36970 46912
rect 37458 46900 37464 46912
rect 37419 46872 37464 46900
rect 37458 46860 37464 46872
rect 37516 46860 37522 46912
rect 38580 46906 38660 46912
rect 38654 46860 38660 46906
rect 38712 46860 38718 46912
rect 42150 46860 42156 46912
rect 42208 46900 42214 46912
rect 42628 46900 42656 46940
rect 43254 46928 43260 46940
rect 43312 46928 43318 46980
rect 46032 46968 46060 46999
rect 45480 46940 46060 46968
rect 42208 46872 42656 46900
rect 42208 46860 42214 46872
rect 44818 46860 44824 46912
rect 44876 46900 44882 46912
rect 45480 46900 45508 46940
rect 44876 46872 45508 46900
rect 44876 46860 44882 46872
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 3973 46699 4031 46705
rect 3973 46665 3985 46699
rect 4019 46696 4031 46699
rect 4062 46696 4068 46708
rect 4019 46668 4068 46696
rect 4019 46665 4031 46668
rect 3973 46659 4031 46665
rect 4062 46656 4068 46668
rect 4120 46656 4126 46708
rect 18414 46696 18420 46708
rect 18375 46668 18420 46696
rect 18414 46656 18420 46668
rect 18472 46656 18478 46708
rect 19153 46699 19211 46705
rect 19153 46665 19165 46699
rect 19199 46696 19211 46699
rect 20530 46696 20536 46708
rect 19199 46668 20536 46696
rect 19199 46665 19211 46668
rect 19153 46659 19211 46665
rect 20530 46656 20536 46668
rect 20588 46656 20594 46708
rect 21269 46699 21327 46705
rect 21269 46665 21281 46699
rect 21315 46696 21327 46699
rect 22094 46696 22100 46708
rect 21315 46668 22100 46696
rect 21315 46665 21327 46668
rect 21269 46659 21327 46665
rect 22094 46656 22100 46668
rect 22152 46656 22158 46708
rect 23842 46696 23848 46708
rect 23803 46668 23848 46696
rect 23842 46656 23848 46668
rect 23900 46656 23906 46708
rect 25682 46656 25688 46708
rect 25740 46696 25746 46708
rect 25869 46699 25927 46705
rect 25869 46696 25881 46699
rect 25740 46668 25881 46696
rect 25740 46656 25746 46668
rect 25869 46665 25881 46668
rect 25915 46665 25927 46699
rect 25869 46659 25927 46665
rect 25958 46656 25964 46708
rect 26016 46696 26022 46708
rect 26053 46699 26111 46705
rect 26053 46696 26065 46699
rect 26016 46668 26065 46696
rect 26016 46656 26022 46668
rect 26053 46665 26065 46668
rect 26099 46665 26111 46699
rect 26053 46659 26111 46665
rect 30098 46656 30104 46708
rect 30156 46696 30162 46708
rect 30156 46668 33732 46696
rect 30156 46656 30162 46668
rect 22189 46631 22247 46637
rect 22189 46628 22201 46631
rect 6886 46600 22201 46628
rect 4798 46560 4804 46572
rect 4759 46532 4804 46560
rect 4798 46520 4804 46532
rect 4856 46520 4862 46572
rect 5994 46560 6000 46572
rect 5955 46532 6000 46560
rect 5994 46520 6000 46532
rect 6052 46520 6058 46572
rect 5626 46452 5632 46504
rect 5684 46492 5690 46504
rect 6886 46492 6914 46600
rect 22189 46597 22201 46600
rect 22235 46597 22247 46631
rect 22830 46628 22836 46640
rect 22189 46591 22247 46597
rect 22388 46600 22836 46628
rect 7006 46560 7012 46572
rect 6967 46532 7012 46560
rect 7006 46520 7012 46532
rect 7064 46520 7070 46572
rect 9214 46560 9220 46572
rect 9175 46532 9220 46560
rect 9214 46520 9220 46532
rect 9272 46520 9278 46572
rect 10318 46560 10324 46572
rect 10279 46532 10324 46560
rect 10318 46520 10324 46532
rect 10376 46520 10382 46572
rect 11330 46520 11336 46572
rect 11388 46560 11394 46572
rect 11701 46563 11759 46569
rect 11701 46560 11713 46563
rect 11388 46532 11713 46560
rect 11388 46520 11394 46532
rect 11701 46529 11713 46532
rect 11747 46529 11759 46563
rect 12526 46560 12532 46572
rect 12487 46532 12532 46560
rect 11701 46523 11759 46529
rect 12526 46520 12532 46532
rect 12584 46520 12590 46572
rect 13630 46560 13636 46572
rect 13591 46532 13636 46560
rect 13630 46520 13636 46532
rect 13688 46520 13694 46572
rect 14734 46560 14740 46572
rect 14695 46532 14740 46560
rect 14734 46520 14740 46532
rect 14792 46520 14798 46572
rect 15838 46560 15844 46572
rect 15799 46532 15844 46560
rect 15838 46520 15844 46532
rect 15896 46520 15902 46572
rect 17221 46563 17279 46569
rect 17221 46529 17233 46563
rect 17267 46560 17279 46563
rect 17954 46560 17960 46572
rect 17267 46532 17960 46560
rect 17267 46529 17279 46532
rect 17221 46523 17279 46529
rect 17954 46520 17960 46532
rect 18012 46520 18018 46572
rect 18601 46563 18659 46569
rect 18601 46529 18613 46563
rect 18647 46529 18659 46563
rect 19334 46560 19340 46572
rect 19295 46532 19340 46560
rect 18601 46523 18659 46529
rect 5684 46464 6914 46492
rect 18616 46492 18644 46523
rect 19334 46520 19340 46532
rect 19392 46520 19398 46572
rect 19981 46563 20039 46569
rect 19981 46529 19993 46563
rect 20027 46560 20039 46563
rect 20254 46560 20260 46572
rect 20027 46532 20260 46560
rect 20027 46529 20039 46532
rect 19981 46523 20039 46529
rect 20254 46520 20260 46532
rect 20312 46520 20318 46572
rect 20714 46520 20720 46572
rect 20772 46560 20778 46572
rect 21328 46563 21386 46569
rect 20772 46532 20944 46560
rect 20772 46520 20778 46532
rect 19518 46492 19524 46504
rect 18616 46464 19524 46492
rect 5684 46452 5690 46464
rect 19518 46452 19524 46464
rect 19576 46452 19582 46504
rect 19794 46492 19800 46504
rect 19755 46464 19800 46492
rect 19794 46452 19800 46464
rect 19852 46452 19858 46504
rect 20809 46495 20867 46501
rect 20809 46492 20821 46495
rect 19904 46464 20821 46492
rect 18690 46384 18696 46436
rect 18748 46424 18754 46436
rect 19904 46424 19932 46464
rect 20809 46461 20821 46464
rect 20855 46461 20867 46495
rect 20916 46492 20944 46532
rect 21328 46529 21340 46563
rect 21374 46560 21386 46563
rect 21542 46560 21548 46572
rect 21374 46532 21548 46560
rect 21374 46529 21386 46532
rect 21328 46523 21386 46529
rect 21542 46520 21548 46532
rect 21600 46520 21606 46572
rect 22278 46520 22284 46572
rect 22336 46560 22342 46572
rect 22388 46569 22416 46600
rect 22830 46588 22836 46600
rect 22888 46588 22894 46640
rect 23290 46588 23296 46640
rect 23348 46628 23354 46640
rect 24854 46628 24860 46640
rect 23348 46600 24860 46628
rect 23348 46588 23354 46600
rect 24854 46588 24860 46600
rect 24912 46588 24918 46640
rect 25222 46628 25228 46640
rect 25183 46600 25228 46628
rect 25222 46588 25228 46600
rect 25280 46588 25286 46640
rect 28074 46628 28080 46640
rect 25792 46600 28080 46628
rect 22373 46563 22431 46569
rect 22373 46560 22385 46563
rect 22336 46532 22385 46560
rect 22336 46520 22342 46532
rect 22373 46529 22385 46532
rect 22419 46529 22431 46563
rect 22373 46523 22431 46529
rect 22465 46563 22523 46569
rect 22465 46529 22477 46563
rect 22511 46529 22523 46563
rect 22738 46560 22744 46572
rect 22699 46532 22744 46560
rect 22465 46523 22523 46529
rect 22480 46492 22508 46523
rect 22738 46520 22744 46532
rect 22796 46520 22802 46572
rect 23385 46563 23443 46569
rect 23385 46529 23397 46563
rect 23431 46560 23443 46563
rect 23658 46560 23664 46572
rect 23431 46532 23664 46560
rect 23431 46529 23443 46532
rect 23385 46523 23443 46529
rect 23658 46520 23664 46532
rect 23716 46520 23722 46572
rect 24026 46560 24032 46572
rect 23987 46532 24032 46560
rect 24026 46520 24032 46532
rect 24084 46520 24090 46572
rect 24210 46520 24216 46572
rect 24268 46560 24274 46572
rect 24397 46561 24455 46567
rect 24268 46532 24313 46560
rect 24268 46520 24274 46532
rect 24397 46527 24409 46561
rect 24443 46560 24455 46561
rect 24486 46560 24492 46572
rect 24443 46532 24492 46560
rect 24443 46527 24455 46532
rect 24397 46521 24455 46527
rect 24486 46520 24492 46532
rect 24544 46520 24550 46572
rect 24581 46563 24639 46569
rect 24581 46529 24593 46563
rect 24627 46560 24639 46563
rect 24670 46560 24676 46572
rect 24627 46532 24676 46560
rect 24627 46529 24639 46532
rect 24581 46523 24639 46529
rect 24670 46520 24676 46532
rect 24728 46520 24734 46572
rect 24762 46520 24768 46572
rect 24820 46560 24826 46572
rect 25409 46563 25467 46569
rect 25409 46560 25421 46563
rect 24820 46532 25421 46560
rect 24820 46520 24826 46532
rect 25409 46529 25421 46532
rect 25455 46560 25467 46563
rect 25792 46560 25820 46600
rect 28074 46588 28080 46600
rect 28132 46588 28138 46640
rect 29086 46588 29092 46640
rect 29144 46628 29150 46640
rect 29144 46600 29592 46628
rect 29144 46588 29150 46600
rect 25455 46532 25820 46560
rect 25455 46529 25467 46532
rect 25409 46523 25467 46529
rect 25866 46520 25872 46572
rect 25924 46560 25930 46572
rect 25994 46563 26052 46569
rect 25994 46560 26006 46563
rect 25924 46532 26006 46560
rect 25924 46520 25930 46532
rect 25994 46529 26006 46532
rect 26040 46560 26052 46563
rect 26142 46560 26148 46572
rect 26040 46532 26148 46560
rect 26040 46529 26052 46532
rect 25994 46523 26052 46529
rect 26142 46520 26148 46532
rect 26200 46520 26206 46572
rect 27062 46560 27068 46572
rect 26252 46532 27068 46560
rect 20916 46464 22508 46492
rect 22649 46495 22707 46501
rect 20809 46455 20867 46461
rect 22649 46461 22661 46495
rect 22695 46492 22707 46495
rect 22922 46492 22928 46504
rect 22695 46464 22928 46492
rect 22695 46461 22707 46464
rect 22649 46455 22707 46461
rect 22922 46452 22928 46464
rect 22980 46452 22986 46504
rect 23014 46452 23020 46504
rect 23072 46492 23078 46504
rect 24302 46492 24308 46504
rect 23072 46464 24308 46492
rect 23072 46452 23078 46464
rect 24302 46452 24308 46464
rect 24360 46452 24366 46504
rect 24504 46492 24532 46520
rect 24504 46464 25084 46492
rect 18748 46396 19932 46424
rect 18748 46384 18754 46396
rect 20254 46384 20260 46436
rect 20312 46424 20318 46436
rect 24946 46424 24952 46436
rect 20312 46396 24952 46424
rect 20312 46384 20318 46396
rect 24946 46384 24952 46396
rect 25004 46384 25010 46436
rect 25056 46424 25084 46464
rect 25222 46452 25228 46504
rect 25280 46492 25286 46504
rect 26252 46492 26280 46532
rect 27062 46520 27068 46532
rect 27120 46560 27126 46572
rect 27341 46563 27399 46569
rect 27341 46560 27353 46563
rect 27120 46532 27353 46560
rect 27120 46520 27126 46532
rect 27341 46529 27353 46532
rect 27387 46529 27399 46563
rect 28166 46560 28172 46572
rect 27341 46523 27399 46529
rect 27432 46532 28172 46560
rect 26418 46492 26424 46504
rect 25280 46464 26280 46492
rect 26379 46464 26424 46492
rect 25280 46452 25286 46464
rect 26418 46452 26424 46464
rect 26476 46452 26482 46504
rect 26513 46495 26571 46501
rect 26513 46461 26525 46495
rect 26559 46492 26571 46495
rect 27432 46492 27460 46532
rect 28166 46520 28172 46532
rect 28224 46560 28230 46572
rect 28261 46563 28319 46569
rect 28261 46560 28273 46563
rect 28224 46532 28273 46560
rect 28224 46520 28230 46532
rect 28261 46529 28273 46532
rect 28307 46529 28319 46563
rect 28442 46560 28448 46572
rect 28403 46532 28448 46560
rect 28261 46523 28319 46529
rect 28442 46520 28448 46532
rect 28500 46520 28506 46572
rect 28534 46520 28540 46572
rect 28592 46560 28598 46572
rect 29362 46560 29368 46572
rect 28592 46532 28637 46560
rect 29323 46532 29368 46560
rect 28592 46520 28598 46532
rect 29362 46520 29368 46532
rect 29420 46520 29426 46572
rect 29564 46569 29592 46600
rect 29822 46588 29828 46640
rect 29880 46628 29886 46640
rect 30193 46631 30251 46637
rect 30193 46628 30205 46631
rect 29880 46600 30205 46628
rect 29880 46588 29886 46600
rect 30193 46597 30205 46600
rect 30239 46597 30251 46631
rect 31846 46628 31852 46640
rect 30193 46591 30251 46597
rect 31588 46600 31852 46628
rect 29549 46563 29607 46569
rect 29549 46529 29561 46563
rect 29595 46529 29607 46563
rect 30650 46560 30656 46572
rect 30611 46532 30656 46560
rect 29549 46523 29607 46529
rect 26559 46464 27460 46492
rect 27617 46495 27675 46501
rect 26559 46461 26571 46464
rect 26513 46455 26571 46461
rect 27617 46461 27629 46495
rect 27663 46492 27675 46495
rect 28460 46492 28488 46520
rect 27663 46464 28488 46492
rect 28997 46495 29055 46501
rect 27663 46461 27675 46464
rect 27617 46455 27675 46461
rect 28997 46461 29009 46495
rect 29043 46461 29055 46495
rect 29178 46492 29184 46504
rect 29139 46464 29184 46492
rect 28997 46455 29055 46461
rect 27157 46427 27215 46433
rect 27157 46424 27169 46427
rect 25056 46396 27169 46424
rect 27157 46393 27169 46396
rect 27203 46393 27215 46427
rect 29012 46424 29040 46455
rect 29178 46452 29184 46464
rect 29236 46452 29242 46504
rect 29564 46492 29592 46523
rect 30650 46520 30656 46532
rect 30708 46520 30714 46572
rect 30742 46520 30748 46572
rect 30800 46560 30806 46572
rect 31588 46569 31616 46600
rect 31846 46588 31852 46600
rect 31904 46628 31910 46640
rect 33704 46628 33732 46668
rect 33778 46656 33784 46708
rect 33836 46696 33842 46708
rect 33965 46699 34023 46705
rect 33965 46696 33977 46699
rect 33836 46668 33977 46696
rect 33836 46656 33842 46668
rect 33965 46665 33977 46668
rect 34011 46665 34023 46699
rect 33965 46659 34023 46665
rect 34054 46656 34060 46708
rect 34112 46696 34118 46708
rect 34149 46699 34207 46705
rect 34149 46696 34161 46699
rect 34112 46668 34161 46696
rect 34112 46656 34118 46668
rect 34149 46665 34161 46668
rect 34195 46665 34207 46699
rect 34149 46659 34207 46665
rect 34790 46656 34796 46708
rect 34848 46696 34854 46708
rect 34848 46668 39804 46696
rect 34848 46656 34854 46668
rect 37366 46628 37372 46640
rect 31904 46600 31984 46628
rect 33704 46600 35112 46628
rect 31904 46588 31910 46600
rect 30837 46563 30895 46569
rect 30837 46560 30849 46563
rect 30800 46532 30849 46560
rect 30800 46520 30806 46532
rect 30837 46529 30849 46532
rect 30883 46529 30895 46563
rect 30837 46523 30895 46529
rect 31573 46563 31631 46569
rect 31573 46529 31585 46563
rect 31619 46529 31631 46563
rect 31956 46560 31984 46600
rect 33778 46560 33784 46572
rect 31956 46532 33784 46560
rect 31573 46523 31631 46529
rect 33778 46520 33784 46532
rect 33836 46520 33842 46572
rect 34146 46560 34152 46572
rect 34107 46532 34152 46560
rect 34146 46520 34152 46532
rect 34204 46520 34210 46572
rect 35084 46569 35112 46600
rect 36188 46600 37372 46628
rect 36188 46569 36216 46600
rect 37366 46588 37372 46600
rect 37424 46628 37430 46640
rect 38565 46631 38623 46637
rect 38565 46628 38577 46631
rect 37424 46600 38577 46628
rect 37424 46588 37430 46600
rect 38565 46597 38577 46600
rect 38611 46597 38623 46631
rect 38565 46591 38623 46597
rect 35069 46563 35127 46569
rect 35069 46529 35081 46563
rect 35115 46529 35127 46563
rect 36173 46563 36231 46569
rect 35069 46523 35127 46529
rect 35452 46532 36032 46560
rect 30101 46495 30159 46501
rect 30101 46492 30113 46495
rect 29564 46464 30113 46492
rect 30101 46461 30113 46464
rect 30147 46461 30159 46495
rect 30101 46455 30159 46461
rect 30285 46495 30343 46501
rect 30285 46461 30297 46495
rect 30331 46461 30343 46495
rect 30285 46455 30343 46461
rect 27157 46387 27215 46393
rect 27264 46396 29040 46424
rect 30300 46424 30328 46455
rect 31662 46452 31668 46504
rect 31720 46492 31726 46504
rect 31757 46495 31815 46501
rect 31757 46492 31769 46495
rect 31720 46464 31769 46492
rect 31720 46452 31726 46464
rect 31757 46461 31769 46464
rect 31803 46492 31815 46495
rect 31846 46492 31852 46504
rect 31803 46464 31852 46492
rect 31803 46461 31815 46464
rect 31757 46455 31815 46461
rect 31846 46452 31852 46464
rect 31904 46452 31910 46504
rect 32030 46452 32036 46504
rect 32088 46492 32094 46504
rect 32309 46495 32367 46501
rect 32309 46492 32321 46495
rect 32088 46464 32321 46492
rect 32088 46452 32094 46464
rect 32309 46461 32321 46464
rect 32355 46461 32367 46495
rect 32582 46492 32588 46504
rect 32543 46464 32588 46492
rect 32309 46455 32367 46461
rect 32582 46452 32588 46464
rect 32640 46452 32646 46504
rect 33502 46452 33508 46504
rect 33560 46492 33566 46504
rect 34609 46495 34667 46501
rect 34609 46492 34621 46495
rect 33560 46464 34621 46492
rect 33560 46452 33566 46464
rect 34609 46461 34621 46464
rect 34655 46492 34667 46495
rect 35452 46492 35480 46532
rect 34655 46464 35480 46492
rect 34655 46461 34667 46464
rect 34609 46455 34667 46461
rect 35526 46452 35532 46504
rect 35584 46492 35590 46504
rect 35805 46495 35863 46501
rect 35805 46492 35817 46495
rect 35584 46464 35817 46492
rect 35584 46452 35590 46464
rect 35805 46461 35817 46464
rect 35851 46461 35863 46495
rect 36004 46492 36032 46532
rect 36173 46529 36185 46563
rect 36219 46529 36231 46563
rect 36173 46523 36231 46529
rect 36262 46520 36268 46572
rect 36320 46560 36326 46572
rect 36633 46563 36691 46569
rect 36320 46532 36584 46560
rect 36320 46520 36326 46532
rect 36446 46492 36452 46504
rect 36004 46464 36452 46492
rect 35805 46455 35863 46461
rect 36446 46452 36452 46464
rect 36504 46452 36510 46504
rect 36556 46492 36584 46532
rect 36633 46529 36645 46563
rect 36679 46560 36691 46563
rect 37458 46560 37464 46572
rect 36679 46532 37464 46560
rect 36679 46529 36691 46532
rect 36633 46523 36691 46529
rect 37458 46520 37464 46532
rect 37516 46520 37522 46572
rect 37645 46563 37703 46569
rect 37645 46529 37657 46563
rect 37691 46529 37703 46563
rect 37645 46523 37703 46529
rect 37660 46492 37688 46523
rect 38102 46520 38108 46572
rect 38160 46560 38166 46572
rect 38381 46563 38439 46569
rect 38381 46560 38393 46563
rect 38160 46532 38393 46560
rect 38160 46520 38166 46532
rect 38381 46529 38393 46532
rect 38427 46529 38439 46563
rect 38381 46523 38439 46529
rect 36556 46464 37688 46492
rect 37921 46495 37979 46501
rect 37921 46461 37933 46495
rect 37967 46492 37979 46495
rect 38470 46492 38476 46504
rect 37967 46464 38476 46492
rect 37967 46461 37979 46464
rect 37921 46455 37979 46461
rect 38470 46452 38476 46464
rect 38528 46452 38534 46504
rect 38580 46492 38608 46591
rect 38657 46563 38715 46569
rect 38657 46529 38669 46563
rect 38703 46560 38715 46563
rect 38838 46560 38844 46572
rect 38703 46532 38844 46560
rect 38703 46529 38715 46532
rect 38657 46523 38715 46529
rect 38838 46520 38844 46532
rect 38896 46520 38902 46572
rect 39114 46560 39120 46572
rect 39075 46532 39120 46560
rect 39114 46520 39120 46532
rect 39172 46520 39178 46572
rect 39776 46569 39804 46668
rect 39761 46563 39819 46569
rect 39761 46529 39773 46563
rect 39807 46529 39819 46563
rect 40862 46560 40868 46572
rect 40823 46532 40868 46560
rect 39761 46523 39819 46529
rect 40862 46520 40868 46532
rect 40920 46520 40926 46572
rect 42610 46520 42616 46572
rect 42668 46560 42674 46572
rect 43257 46563 43315 46569
rect 43257 46560 43269 46563
rect 42668 46532 43269 46560
rect 42668 46520 42674 46532
rect 43257 46529 43269 46532
rect 43303 46529 43315 46563
rect 43257 46523 43315 46529
rect 43346 46520 43352 46572
rect 43404 46560 43410 46572
rect 43901 46563 43959 46569
rect 43901 46560 43913 46563
rect 43404 46532 43913 46560
rect 43404 46520 43410 46532
rect 43901 46529 43913 46532
rect 43947 46529 43959 46563
rect 43901 46523 43959 46529
rect 44450 46520 44456 46572
rect 44508 46560 44514 46572
rect 45189 46563 45247 46569
rect 45189 46560 45201 46563
rect 44508 46532 45201 46560
rect 44508 46520 44514 46532
rect 45189 46529 45201 46532
rect 45235 46529 45247 46563
rect 45830 46560 45836 46572
rect 45791 46532 45836 46560
rect 45189 46523 45247 46529
rect 45830 46520 45836 46532
rect 45888 46520 45894 46572
rect 41141 46495 41199 46501
rect 41141 46492 41153 46495
rect 38580 46464 41153 46492
rect 41141 46461 41153 46464
rect 41187 46461 41199 46495
rect 41141 46455 41199 46461
rect 43714 46452 43720 46504
rect 43772 46492 43778 46504
rect 44545 46495 44603 46501
rect 44545 46492 44557 46495
rect 43772 46464 44557 46492
rect 43772 46452 43778 46464
rect 44545 46461 44557 46464
rect 44591 46461 44603 46495
rect 44545 46455 44603 46461
rect 30466 46424 30472 46436
rect 30300 46396 30472 46424
rect 17865 46359 17923 46365
rect 17865 46325 17877 46359
rect 17911 46356 17923 46359
rect 18782 46356 18788 46368
rect 17911 46328 18788 46356
rect 17911 46325 17923 46328
rect 17865 46319 17923 46325
rect 18782 46316 18788 46328
rect 18840 46316 18846 46368
rect 20070 46316 20076 46368
rect 20128 46356 20134 46368
rect 20165 46359 20223 46365
rect 20165 46356 20177 46359
rect 20128 46328 20177 46356
rect 20128 46316 20134 46328
rect 20165 46325 20177 46328
rect 20211 46325 20223 46359
rect 20898 46356 20904 46368
rect 20859 46328 20904 46356
rect 20165 46319 20223 46325
rect 20898 46316 20904 46328
rect 20956 46316 20962 46368
rect 21450 46356 21456 46368
rect 21411 46328 21456 46356
rect 21450 46316 21456 46328
rect 21508 46316 21514 46368
rect 23750 46316 23756 46368
rect 23808 46356 23814 46368
rect 25041 46359 25099 46365
rect 25041 46356 25053 46359
rect 23808 46328 25053 46356
rect 23808 46316 23814 46328
rect 25041 46325 25053 46328
rect 25087 46325 25099 46359
rect 25041 46319 25099 46325
rect 25130 46316 25136 46368
rect 25188 46356 25194 46368
rect 27264 46356 27292 46396
rect 30466 46384 30472 46396
rect 30524 46424 30530 46436
rect 36541 46427 36599 46433
rect 36541 46424 36553 46427
rect 30524 46396 36553 46424
rect 30524 46384 30530 46396
rect 36541 46393 36553 46396
rect 36587 46393 36599 46427
rect 36541 46387 36599 46393
rect 37090 46384 37096 46436
rect 37148 46424 37154 46436
rect 38746 46424 38752 46436
rect 37148 46396 38752 46424
rect 37148 46384 37154 46396
rect 38746 46384 38752 46396
rect 38804 46384 38810 46436
rect 41506 46384 41512 46436
rect 41564 46424 41570 46436
rect 42613 46427 42671 46433
rect 42613 46424 42625 46427
rect 41564 46396 42625 46424
rect 41564 46384 41570 46396
rect 42613 46393 42625 46396
rect 42659 46393 42671 46427
rect 42613 46387 42671 46393
rect 25188 46328 27292 46356
rect 25188 46316 25194 46328
rect 27338 46316 27344 46368
rect 27396 46356 27402 46368
rect 27525 46359 27583 46365
rect 27525 46356 27537 46359
rect 27396 46328 27537 46356
rect 27396 46316 27402 46328
rect 27525 46325 27537 46328
rect 27571 46325 27583 46359
rect 27525 46319 27583 46325
rect 27798 46316 27804 46368
rect 27856 46356 27862 46368
rect 28077 46359 28135 46365
rect 28077 46356 28089 46359
rect 27856 46328 28089 46356
rect 27856 46316 27862 46328
rect 28077 46325 28089 46328
rect 28123 46325 28135 46359
rect 28077 46319 28135 46325
rect 31389 46359 31447 46365
rect 31389 46325 31401 46359
rect 31435 46356 31447 46359
rect 31846 46356 31852 46368
rect 31435 46328 31852 46356
rect 31435 46325 31447 46328
rect 31389 46319 31447 46325
rect 31846 46316 31852 46328
rect 31904 46316 31910 46368
rect 32030 46316 32036 46368
rect 32088 46356 32094 46368
rect 34330 46356 34336 46368
rect 32088 46328 34336 46356
rect 32088 46316 32094 46328
rect 34330 46316 34336 46328
rect 34388 46316 34394 46368
rect 34517 46359 34575 46365
rect 34517 46325 34529 46359
rect 34563 46356 34575 46359
rect 34790 46356 34796 46368
rect 34563 46328 34796 46356
rect 34563 46325 34575 46328
rect 34517 46319 34575 46325
rect 34790 46316 34796 46328
rect 34848 46356 34854 46368
rect 35526 46356 35532 46368
rect 34848 46328 35532 46356
rect 34848 46316 34854 46328
rect 35526 46316 35532 46328
rect 35584 46316 35590 46368
rect 35986 46316 35992 46368
rect 36044 46356 36050 46368
rect 37461 46359 37519 46365
rect 37461 46356 37473 46359
rect 36044 46328 37473 46356
rect 36044 46316 36050 46328
rect 37461 46325 37473 46328
rect 37507 46325 37519 46359
rect 37461 46319 37519 46325
rect 37550 46316 37556 46368
rect 37608 46356 37614 46368
rect 37829 46359 37887 46365
rect 37829 46356 37841 46359
rect 37608 46328 37841 46356
rect 37608 46316 37614 46328
rect 37829 46325 37841 46328
rect 37875 46325 37887 46359
rect 37829 46319 37887 46325
rect 37918 46316 37924 46368
rect 37976 46356 37982 46368
rect 38381 46359 38439 46365
rect 38381 46356 38393 46359
rect 37976 46328 38393 46356
rect 37976 46316 37982 46328
rect 38381 46325 38393 46328
rect 38427 46325 38439 46359
rect 38381 46319 38439 46325
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 5902 46152 5908 46164
rect 5863 46124 5908 46152
rect 5902 46112 5908 46124
rect 5960 46112 5966 46164
rect 16942 46152 16948 46164
rect 16903 46124 16948 46152
rect 16942 46112 16948 46124
rect 17000 46112 17006 46164
rect 18046 46152 18052 46164
rect 18007 46124 18052 46152
rect 18046 46112 18052 46124
rect 18104 46112 18110 46164
rect 18690 46152 18696 46164
rect 18651 46124 18696 46152
rect 18690 46112 18696 46124
rect 18748 46112 18754 46164
rect 18782 46112 18788 46164
rect 18840 46152 18846 46164
rect 21266 46152 21272 46164
rect 18840 46124 21272 46152
rect 18840 46112 18846 46124
rect 21266 46112 21272 46124
rect 21324 46112 21330 46164
rect 22738 46152 22744 46164
rect 22699 46124 22744 46152
rect 22738 46112 22744 46124
rect 22796 46112 22802 46164
rect 22830 46112 22836 46164
rect 22888 46152 22894 46164
rect 24946 46152 24952 46164
rect 22888 46124 24072 46152
rect 24907 46124 24952 46152
rect 22888 46112 22894 46124
rect 20714 46044 20720 46096
rect 20772 46084 20778 46096
rect 20901 46087 20959 46093
rect 20901 46084 20913 46087
rect 20772 46056 20913 46084
rect 20772 46044 20778 46056
rect 20901 46053 20913 46056
rect 20947 46053 20959 46087
rect 20901 46047 20959 46053
rect 22646 46044 22652 46096
rect 22704 46084 22710 46096
rect 23934 46084 23940 46096
rect 22704 46056 23940 46084
rect 22704 46044 22710 46056
rect 23934 46044 23940 46056
rect 23992 46044 23998 46096
rect 24044 46084 24072 46124
rect 24946 46112 24952 46124
rect 25004 46112 25010 46164
rect 27338 46112 27344 46164
rect 27396 46152 27402 46164
rect 28534 46152 28540 46164
rect 27396 46124 28540 46152
rect 27396 46112 27402 46124
rect 28534 46112 28540 46124
rect 28592 46152 28598 46164
rect 28629 46155 28687 46161
rect 28629 46152 28641 46155
rect 28592 46124 28641 46152
rect 28592 46112 28598 46124
rect 28629 46121 28641 46124
rect 28675 46152 28687 46155
rect 28675 46124 29132 46152
rect 28675 46121 28687 46124
rect 28629 46115 28687 46121
rect 25130 46084 25136 46096
rect 24044 46056 25136 46084
rect 25130 46044 25136 46056
rect 25188 46044 25194 46096
rect 25222 46044 25228 46096
rect 25280 46044 25286 46096
rect 25866 46084 25872 46096
rect 25332 46056 25872 46084
rect 19613 46019 19671 46025
rect 19613 46016 19625 46019
rect 18248 45988 19625 46016
rect 18248 45957 18276 45988
rect 19613 45985 19625 45988
rect 19659 45985 19671 46019
rect 20438 46016 20444 46028
rect 19613 45979 19671 45985
rect 19720 45988 20444 46016
rect 18233 45951 18291 45957
rect 18233 45917 18245 45951
rect 18279 45917 18291 45951
rect 18233 45911 18291 45917
rect 18877 45951 18935 45957
rect 18877 45917 18889 45951
rect 18923 45948 18935 45951
rect 19720 45948 19748 45988
rect 20438 45976 20444 45988
rect 20496 45976 20502 46028
rect 23106 46016 23112 46028
rect 20916 45988 23112 46016
rect 18923 45920 19748 45948
rect 18923 45917 18935 45920
rect 18877 45911 18935 45917
rect 19794 45908 19800 45960
rect 19852 45948 19858 45960
rect 19852 45920 19897 45948
rect 19852 45908 19858 45920
rect 19978 45908 19984 45960
rect 20036 45948 20042 45960
rect 20916 45957 20944 45988
rect 23106 45976 23112 45988
rect 23164 45976 23170 46028
rect 23658 46016 23664 46028
rect 23619 45988 23664 46016
rect 23658 45976 23664 45988
rect 23716 45976 23722 46028
rect 24762 46016 24768 46028
rect 23860 45988 24768 46016
rect 20809 45951 20867 45957
rect 20036 45920 20081 45948
rect 20036 45908 20042 45920
rect 20809 45917 20821 45951
rect 20855 45917 20867 45951
rect 20809 45911 20867 45917
rect 20901 45951 20959 45957
rect 20901 45917 20913 45951
rect 20947 45917 20959 45951
rect 21358 45948 21364 45960
rect 21319 45920 21364 45948
rect 20901 45911 20959 45917
rect 20625 45883 20683 45889
rect 20625 45849 20637 45883
rect 20671 45849 20683 45883
rect 20824 45880 20852 45911
rect 21358 45908 21364 45920
rect 21416 45908 21422 45960
rect 21542 45948 21548 45960
rect 21503 45920 21548 45948
rect 21542 45908 21548 45920
rect 21600 45948 21606 45960
rect 23860 45957 23888 45988
rect 24762 45976 24768 45988
rect 24820 45976 24826 46028
rect 25240 46016 25268 46044
rect 25332 46025 25360 46056
rect 25866 46044 25872 46056
rect 25924 46044 25930 46096
rect 28166 46084 28172 46096
rect 27724 46056 28172 46084
rect 24964 45988 25268 46016
rect 25317 46019 25375 46025
rect 23845 45951 23903 45957
rect 21600 45920 23796 45948
rect 21600 45908 21606 45920
rect 22554 45880 22560 45892
rect 20824 45852 22560 45880
rect 20625 45843 20683 45849
rect 9858 45772 9864 45824
rect 9916 45812 9922 45824
rect 10045 45815 10103 45821
rect 10045 45812 10057 45815
rect 9916 45784 10057 45812
rect 9916 45772 9922 45784
rect 10045 45781 10057 45784
rect 10091 45812 10103 45815
rect 20254 45812 20260 45824
rect 10091 45784 20260 45812
rect 10091 45781 10103 45784
rect 10045 45775 10103 45781
rect 20254 45772 20260 45784
rect 20312 45772 20318 45824
rect 20640 45812 20668 45843
rect 22554 45840 22560 45852
rect 22612 45880 22618 45892
rect 22925 45883 22983 45889
rect 22925 45880 22937 45883
rect 22612 45852 22937 45880
rect 22612 45840 22618 45852
rect 22925 45849 22937 45852
rect 22971 45849 22983 45883
rect 23106 45880 23112 45892
rect 23067 45852 23112 45880
rect 22925 45843 22983 45849
rect 23106 45840 23112 45852
rect 23164 45840 23170 45892
rect 23768 45880 23796 45920
rect 23845 45917 23857 45951
rect 23891 45917 23903 45951
rect 23845 45911 23903 45917
rect 24029 45951 24087 45957
rect 24029 45917 24041 45951
rect 24075 45948 24087 45951
rect 24964 45948 24992 45988
rect 25317 45985 25329 46019
rect 25363 45985 25375 46019
rect 25317 45979 25375 45985
rect 25409 46019 25467 46025
rect 25409 45985 25421 46019
rect 25455 46016 25467 46019
rect 25498 46016 25504 46028
rect 25455 45988 25504 46016
rect 25455 45985 25467 45988
rect 25409 45979 25467 45985
rect 25498 45976 25504 45988
rect 25556 45976 25562 46028
rect 25130 45948 25136 45960
rect 24075 45920 24992 45948
rect 25091 45920 25136 45948
rect 24075 45917 24087 45920
rect 24029 45911 24087 45917
rect 25130 45908 25136 45920
rect 25188 45908 25194 45960
rect 25225 45951 25283 45957
rect 25225 45917 25237 45951
rect 25271 45948 25283 45951
rect 26050 45948 26056 45960
rect 25271 45920 26056 45948
rect 25271 45917 25283 45920
rect 25225 45911 25283 45917
rect 26050 45908 26056 45920
rect 26108 45908 26114 45960
rect 26513 45951 26571 45957
rect 26513 45917 26525 45951
rect 26559 45917 26571 45951
rect 26694 45948 26700 45960
rect 26655 45920 26700 45948
rect 26513 45911 26571 45917
rect 26329 45883 26387 45889
rect 26329 45880 26341 45883
rect 23768 45852 26341 45880
rect 26329 45849 26341 45852
rect 26375 45849 26387 45883
rect 26528 45880 26556 45911
rect 26694 45908 26700 45920
rect 26752 45908 26758 45960
rect 26786 45908 26792 45960
rect 26844 45948 26850 45960
rect 27724 45957 27752 46056
rect 28166 46044 28172 46056
rect 28224 46044 28230 46096
rect 28442 46044 28448 46096
rect 28500 46084 28506 46096
rect 29104 46084 29132 46124
rect 29178 46112 29184 46164
rect 29236 46152 29242 46164
rect 31573 46155 31631 46161
rect 31573 46152 31585 46155
rect 29236 46124 31585 46152
rect 29236 46112 29242 46124
rect 31573 46121 31585 46124
rect 31619 46121 31631 46155
rect 32582 46152 32588 46164
rect 31573 46115 31631 46121
rect 31680 46124 32588 46152
rect 29822 46084 29828 46096
rect 28500 46056 28856 46084
rect 29104 46056 29828 46084
rect 28500 46044 28506 46056
rect 28718 46016 28724 46028
rect 28679 45988 28724 46016
rect 28718 45976 28724 45988
rect 28776 45976 28782 46028
rect 28828 46016 28856 46056
rect 29822 46044 29828 46056
rect 29880 46044 29886 46096
rect 30282 46084 30288 46096
rect 30243 46056 30288 46084
rect 30282 46044 30288 46056
rect 30340 46044 30346 46096
rect 31680 46016 31708 46124
rect 32582 46112 32588 46124
rect 32640 46112 32646 46164
rect 37918 46152 37924 46164
rect 33060 46124 37924 46152
rect 31754 46044 31760 46096
rect 31812 46084 31818 46096
rect 32030 46084 32036 46096
rect 31812 46056 32036 46084
rect 31812 46044 31818 46056
rect 32030 46044 32036 46056
rect 32088 46044 32094 46096
rect 32950 46084 32956 46096
rect 32911 46056 32956 46084
rect 32950 46044 32956 46056
rect 33008 46044 33014 46096
rect 28828 45988 31708 46016
rect 31772 46016 31800 46044
rect 31849 46019 31907 46025
rect 31849 46016 31861 46019
rect 31772 45988 31861 46016
rect 31849 45985 31861 45988
rect 31895 45985 31907 46019
rect 31849 45979 31907 45985
rect 31941 46019 31999 46025
rect 31941 45985 31953 46019
rect 31987 46016 31999 46019
rect 32122 46016 32128 46028
rect 31987 45988 32128 46016
rect 31987 45985 31999 45988
rect 31941 45979 31999 45985
rect 32122 45976 32128 45988
rect 32180 46016 32186 46028
rect 33060 46016 33088 46124
rect 37918 46112 37924 46124
rect 37976 46112 37982 46164
rect 38102 46152 38108 46164
rect 38063 46124 38108 46152
rect 38102 46112 38108 46124
rect 38160 46112 38166 46164
rect 38378 46112 38384 46164
rect 38436 46152 38442 46164
rect 38436 46124 38884 46152
rect 38436 46112 38442 46124
rect 33226 46044 33232 46096
rect 33284 46044 33290 46096
rect 33318 46044 33324 46096
rect 33376 46044 33382 46096
rect 33778 46044 33784 46096
rect 33836 46084 33842 46096
rect 37093 46087 37151 46093
rect 37093 46084 37105 46087
rect 33836 46056 37105 46084
rect 33836 46044 33842 46056
rect 37093 46053 37105 46056
rect 37139 46053 37151 46087
rect 37093 46047 37151 46053
rect 32180 45988 33088 46016
rect 33129 46019 33187 46025
rect 32180 45976 32186 45988
rect 33129 45985 33141 46019
rect 33175 46016 33187 46019
rect 33244 46016 33272 46044
rect 33175 45988 33272 46016
rect 33336 46016 33364 46044
rect 33413 46019 33471 46025
rect 33413 46016 33425 46019
rect 33336 45988 33425 46016
rect 33175 45985 33187 45988
rect 33129 45979 33187 45985
rect 33413 45985 33425 45988
rect 33459 45985 33471 46019
rect 33413 45979 33471 45985
rect 34974 45976 34980 46028
rect 35032 46016 35038 46028
rect 35434 46016 35440 46028
rect 35032 45988 35440 46016
rect 35032 45976 35038 45988
rect 35434 45976 35440 45988
rect 35492 45976 35498 46028
rect 35526 45976 35532 46028
rect 35584 46016 35590 46028
rect 35802 46016 35808 46028
rect 35584 45988 35808 46016
rect 35584 45976 35590 45988
rect 27811 45961 27869 45967
rect 27525 45951 27583 45957
rect 26844 45920 26889 45948
rect 27433 45929 27491 45935
rect 26844 45908 26850 45920
rect 27433 45895 27445 45929
rect 27479 45895 27491 45929
rect 27525 45917 27537 45951
rect 27571 45917 27583 45951
rect 27525 45911 27583 45917
rect 27721 45951 27779 45957
rect 27721 45917 27733 45951
rect 27767 45917 27779 45951
rect 27811 45927 27823 45961
rect 27857 45958 27869 45961
rect 27857 45948 27936 45958
rect 28261 45951 28319 45957
rect 28261 45948 28273 45951
rect 27857 45930 28273 45948
rect 27857 45927 27869 45930
rect 27811 45921 27869 45927
rect 27908 45920 28273 45930
rect 27721 45911 27779 45917
rect 28261 45917 28273 45920
rect 28307 45917 28319 45951
rect 28261 45911 28319 45917
rect 27433 45889 27491 45895
rect 27249 45883 27307 45889
rect 27249 45880 27261 45883
rect 26528 45852 27261 45880
rect 26329 45843 26387 45849
rect 27249 45849 27261 45852
rect 27295 45849 27307 45883
rect 27249 45843 27307 45849
rect 21542 45812 21548 45824
rect 20640 45784 21548 45812
rect 21542 45772 21548 45784
rect 21600 45772 21606 45824
rect 21726 45812 21732 45824
rect 21687 45784 21732 45812
rect 21726 45772 21732 45784
rect 21784 45772 21790 45824
rect 22281 45815 22339 45821
rect 22281 45781 22293 45815
rect 22327 45812 22339 45815
rect 24026 45812 24032 45824
rect 22327 45784 24032 45812
rect 22327 45781 22339 45784
rect 22281 45775 22339 45781
rect 24026 45772 24032 45784
rect 24084 45772 24090 45824
rect 27338 45772 27344 45824
rect 27396 45812 27402 45824
rect 27448 45812 27476 45889
rect 27396 45784 27476 45812
rect 27540 45812 27568 45911
rect 28350 45908 28356 45960
rect 28408 45948 28414 45960
rect 28445 45951 28503 45957
rect 28445 45948 28457 45951
rect 28408 45920 28457 45948
rect 28408 45908 28414 45920
rect 28445 45917 28457 45920
rect 28491 45917 28503 45951
rect 28445 45911 28503 45917
rect 29825 45951 29883 45957
rect 29825 45917 29837 45951
rect 29871 45948 29883 45951
rect 30006 45948 30012 45960
rect 29871 45920 30012 45948
rect 29871 45917 29883 45920
rect 29825 45911 29883 45917
rect 27982 45840 27988 45892
rect 28040 45880 28046 45892
rect 29840 45880 29868 45911
rect 30006 45908 30012 45920
rect 30064 45908 30070 45960
rect 30466 45948 30472 45960
rect 30427 45920 30472 45948
rect 30466 45908 30472 45920
rect 30524 45908 30530 45960
rect 30742 45948 30748 45960
rect 30703 45920 30748 45948
rect 30742 45908 30748 45920
rect 30800 45908 30806 45960
rect 31754 45908 31760 45960
rect 31812 45948 31818 45960
rect 32033 45951 32091 45957
rect 31812 45920 31857 45948
rect 31812 45908 31818 45920
rect 32033 45917 32045 45951
rect 32079 45948 32091 45951
rect 32950 45948 32956 45960
rect 32079 45920 32956 45948
rect 32079 45917 32091 45920
rect 32033 45911 32091 45917
rect 32950 45908 32956 45920
rect 33008 45948 33014 45960
rect 33229 45951 33287 45957
rect 33229 45948 33241 45951
rect 33008 45920 33241 45948
rect 33008 45908 33014 45920
rect 33229 45917 33241 45920
rect 33275 45917 33287 45951
rect 33229 45911 33287 45917
rect 33322 45951 33380 45957
rect 33322 45917 33334 45951
rect 33368 45950 33380 45951
rect 33368 45948 33548 45950
rect 34054 45948 34060 45960
rect 33368 45922 34060 45948
rect 33368 45917 33380 45922
rect 33520 45920 34060 45922
rect 33322 45911 33380 45917
rect 34054 45908 34060 45920
rect 34112 45908 34118 45960
rect 34514 45908 34520 45960
rect 34572 45948 34578 45960
rect 35636 45957 35664 45988
rect 35802 45976 35808 45988
rect 35860 45976 35866 46028
rect 36538 46016 36544 46028
rect 35912 45988 36544 46016
rect 35621 45951 35679 45957
rect 34572 45920 35572 45948
rect 34572 45908 34578 45920
rect 30650 45880 30656 45892
rect 28040 45852 29868 45880
rect 30611 45852 30656 45880
rect 28040 45840 28046 45852
rect 30650 45840 30656 45852
rect 30708 45840 30714 45892
rect 33502 45840 33508 45892
rect 33560 45880 33566 45892
rect 34149 45883 34207 45889
rect 34149 45880 34161 45883
rect 33560 45852 34161 45880
rect 33560 45840 33566 45852
rect 34149 45849 34161 45852
rect 34195 45849 34207 45883
rect 34149 45843 34207 45849
rect 34333 45883 34391 45889
rect 34333 45849 34345 45883
rect 34379 45880 34391 45883
rect 34606 45880 34612 45892
rect 34379 45852 34612 45880
rect 34379 45849 34391 45852
rect 34333 45843 34391 45849
rect 34606 45840 34612 45852
rect 34664 45840 34670 45892
rect 35544 45880 35572 45920
rect 35621 45917 35633 45951
rect 35667 45917 35679 45951
rect 35621 45911 35679 45917
rect 35710 45908 35716 45960
rect 35768 45948 35774 45960
rect 35912 45957 35940 45988
rect 36538 45976 36544 45988
rect 36596 45976 36602 46028
rect 37553 46019 37611 46025
rect 37553 45985 37565 46019
rect 37599 46016 37611 46019
rect 38120 46016 38148 46112
rect 38286 46044 38292 46096
rect 38344 46044 38350 46096
rect 38470 46084 38476 46096
rect 38431 46056 38476 46084
rect 38470 46044 38476 46056
rect 38528 46044 38534 46096
rect 38562 46044 38568 46096
rect 38620 46044 38626 46096
rect 37599 45988 38148 46016
rect 38304 46016 38332 46044
rect 38381 46019 38439 46025
rect 38381 46016 38393 46019
rect 38304 45988 38393 46016
rect 37599 45985 37611 45988
rect 37553 45979 37611 45985
rect 38381 45985 38393 45988
rect 38427 45985 38439 46019
rect 38381 45979 38439 45985
rect 35897 45951 35955 45957
rect 35768 45920 35813 45948
rect 35768 45908 35774 45920
rect 35897 45917 35909 45951
rect 35943 45917 35955 45951
rect 35897 45911 35955 45917
rect 35986 45908 35992 45960
rect 36044 45948 36050 45960
rect 36044 45920 36089 45948
rect 36044 45908 36050 45920
rect 36446 45908 36452 45960
rect 36504 45948 36510 45960
rect 36633 45951 36691 45957
rect 36633 45948 36645 45951
rect 36504 45920 36645 45948
rect 36504 45908 36510 45920
rect 36633 45917 36645 45920
rect 36679 45917 36691 45951
rect 36633 45911 36691 45917
rect 37366 45908 37372 45960
rect 37424 45948 37430 45960
rect 37461 45951 37519 45957
rect 37461 45948 37473 45951
rect 37424 45920 37473 45948
rect 37424 45908 37430 45920
rect 37461 45917 37473 45920
rect 37507 45917 37519 45951
rect 37461 45911 37519 45917
rect 38010 45908 38016 45960
rect 38068 45948 38074 45960
rect 38580 45957 38608 46044
rect 38856 46016 38884 46124
rect 38930 46112 38936 46164
rect 38988 46152 38994 46164
rect 40681 46155 40739 46161
rect 40681 46152 40693 46155
rect 38988 46124 40693 46152
rect 38988 46112 38994 46124
rect 40681 46121 40693 46124
rect 40727 46121 40739 46155
rect 40681 46115 40739 46121
rect 41138 46112 41144 46164
rect 41196 46152 41202 46164
rect 41969 46155 42027 46161
rect 41969 46152 41981 46155
rect 41196 46124 41981 46152
rect 41196 46112 41202 46124
rect 41969 46121 41981 46124
rect 42015 46121 42027 46155
rect 41969 46115 42027 46121
rect 42242 46112 42248 46164
rect 42300 46152 42306 46164
rect 42613 46155 42671 46161
rect 42613 46152 42625 46155
rect 42300 46124 42625 46152
rect 42300 46112 42306 46124
rect 42613 46121 42625 46124
rect 42659 46121 42671 46155
rect 43254 46152 43260 46164
rect 43215 46124 43260 46152
rect 42613 46115 42671 46121
rect 43254 46112 43260 46124
rect 43312 46112 43318 46164
rect 43806 46152 43812 46164
rect 43767 46124 43812 46152
rect 43806 46112 43812 46124
rect 43864 46112 43870 46164
rect 44174 46112 44180 46164
rect 44232 46152 44238 46164
rect 44361 46155 44419 46161
rect 44361 46152 44373 46155
rect 44232 46124 44373 46152
rect 44232 46112 44238 46124
rect 44361 46121 44373 46124
rect 44407 46121 44419 46155
rect 45186 46152 45192 46164
rect 45147 46124 45192 46152
rect 44361 46115 44419 46121
rect 45186 46112 45192 46124
rect 45244 46112 45250 46164
rect 40310 46044 40316 46096
rect 40368 46084 40374 46096
rect 41325 46087 41383 46093
rect 41325 46084 41337 46087
rect 40368 46056 41337 46084
rect 40368 46044 40374 46056
rect 41325 46053 41337 46056
rect 41371 46053 41383 46087
rect 41325 46047 41383 46053
rect 40037 46019 40095 46025
rect 40037 46016 40049 46019
rect 38856 45988 40049 46016
rect 40037 45985 40049 45988
rect 40083 45985 40095 46019
rect 40037 45979 40095 45985
rect 38301 45951 38359 45957
rect 38301 45948 38313 45951
rect 38068 45920 38313 45948
rect 38068 45908 38074 45920
rect 38301 45917 38313 45920
rect 38347 45917 38359 45951
rect 38577 45951 38635 45957
rect 38577 45948 38589 45951
rect 38487 45920 38589 45948
rect 38301 45911 38359 45917
rect 38577 45917 38589 45920
rect 38623 45948 38635 45951
rect 38838 45948 38844 45960
rect 38623 45920 38844 45948
rect 38623 45917 38635 45920
rect 38577 45911 38635 45917
rect 38838 45908 38844 45920
rect 38896 45908 38902 45960
rect 39117 45951 39175 45957
rect 39117 45917 39129 45951
rect 39163 45948 39175 45951
rect 39163 45920 39344 45948
rect 39163 45917 39175 45920
rect 39117 45911 39175 45917
rect 35544 45852 36676 45880
rect 28718 45812 28724 45824
rect 27540 45784 28724 45812
rect 27396 45772 27402 45784
rect 28718 45772 28724 45784
rect 28776 45772 28782 45824
rect 31386 45772 31392 45824
rect 31444 45812 31450 45824
rect 31938 45812 31944 45824
rect 31444 45784 31944 45812
rect 31444 45772 31450 45784
rect 31938 45772 31944 45784
rect 31996 45772 32002 45824
rect 33962 45812 33968 45824
rect 33923 45784 33968 45812
rect 33962 45772 33968 45784
rect 34020 45772 34026 45824
rect 35437 45815 35495 45821
rect 35437 45781 35449 45815
rect 35483 45812 35495 45815
rect 35710 45812 35716 45824
rect 35483 45784 35716 45812
rect 35483 45781 35495 45784
rect 35437 45775 35495 45781
rect 35710 45772 35716 45784
rect 35768 45772 35774 45824
rect 36648 45812 36676 45852
rect 36722 45840 36728 45892
rect 36780 45880 36786 45892
rect 39206 45880 39212 45892
rect 36780 45852 39212 45880
rect 36780 45840 36786 45852
rect 39206 45840 39212 45852
rect 39264 45840 39270 45892
rect 39316 45812 39344 45920
rect 36648 45784 39344 45812
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 20717 45611 20775 45617
rect 20717 45577 20729 45611
rect 20763 45577 20775 45611
rect 23106 45608 23112 45620
rect 23067 45580 23112 45608
rect 20717 45571 20775 45577
rect 17770 45540 17776 45552
rect 17731 45512 17776 45540
rect 17770 45500 17776 45512
rect 17828 45540 17834 45552
rect 19705 45543 19763 45549
rect 19705 45540 19717 45543
rect 17828 45512 19717 45540
rect 17828 45500 17834 45512
rect 19705 45509 19717 45512
rect 19751 45540 19763 45543
rect 20530 45540 20536 45552
rect 19751 45512 20536 45540
rect 19751 45509 19763 45512
rect 19705 45503 19763 45509
rect 20530 45500 20536 45512
rect 20588 45500 20594 45552
rect 20732 45540 20760 45571
rect 23106 45568 23112 45580
rect 23164 45568 23170 45620
rect 24026 45608 24032 45620
rect 23939 45580 24032 45608
rect 24026 45568 24032 45580
rect 24084 45608 24090 45620
rect 26050 45608 26056 45620
rect 24084 45580 26056 45608
rect 24084 45568 24090 45580
rect 20806 45540 20812 45552
rect 20732 45512 20812 45540
rect 20806 45500 20812 45512
rect 20864 45500 20870 45552
rect 18509 45475 18567 45481
rect 18509 45441 18521 45475
rect 18555 45472 18567 45475
rect 19058 45472 19064 45484
rect 18555 45444 19064 45472
rect 18555 45441 18567 45444
rect 18509 45435 18567 45441
rect 19058 45432 19064 45444
rect 19116 45432 19122 45484
rect 20714 45475 20772 45481
rect 20714 45441 20726 45475
rect 20760 45472 20772 45475
rect 22189 45475 22247 45481
rect 22189 45472 22201 45475
rect 20760 45444 22201 45472
rect 20760 45441 20772 45444
rect 20714 45435 20772 45441
rect 22189 45441 22201 45444
rect 22235 45472 22247 45475
rect 22370 45472 22376 45484
rect 22235 45444 22376 45472
rect 22235 45441 22247 45444
rect 22189 45435 22247 45441
rect 22370 45432 22376 45444
rect 22428 45432 22434 45484
rect 23385 45475 23443 45481
rect 23385 45441 23397 45475
rect 23431 45472 23443 45475
rect 23750 45472 23756 45484
rect 23431 45444 23756 45472
rect 23431 45441 23443 45444
rect 23385 45435 23443 45441
rect 23750 45432 23756 45444
rect 23808 45432 23814 45484
rect 19153 45407 19211 45413
rect 19153 45373 19165 45407
rect 19199 45404 19211 45407
rect 20162 45404 20168 45416
rect 19199 45376 20168 45404
rect 19199 45373 19211 45376
rect 19153 45367 19211 45373
rect 20162 45364 20168 45376
rect 20220 45364 20226 45416
rect 21177 45407 21235 45413
rect 21177 45373 21189 45407
rect 21223 45373 21235 45407
rect 21177 45367 21235 45373
rect 19426 45296 19432 45348
rect 19484 45336 19490 45348
rect 21192 45336 21220 45367
rect 21358 45364 21364 45416
rect 21416 45404 21422 45416
rect 21910 45404 21916 45416
rect 21416 45376 21916 45404
rect 21416 45364 21422 45376
rect 21910 45364 21916 45376
rect 21968 45404 21974 45416
rect 22005 45407 22063 45413
rect 22005 45404 22017 45407
rect 21968 45376 22017 45404
rect 21968 45364 21974 45376
rect 22005 45373 22017 45376
rect 22051 45373 22063 45407
rect 23290 45404 23296 45416
rect 23251 45376 23296 45404
rect 22005 45367 22063 45373
rect 23290 45364 23296 45376
rect 23348 45364 23354 45416
rect 23474 45404 23480 45416
rect 23435 45376 23480 45404
rect 23474 45364 23480 45376
rect 23532 45364 23538 45416
rect 23569 45407 23627 45413
rect 23569 45373 23581 45407
rect 23615 45404 23627 45407
rect 24044 45404 24072 45568
rect 25314 45540 25320 45552
rect 24136 45512 25320 45540
rect 24136 45481 24164 45512
rect 25314 45500 25320 45512
rect 25372 45500 25378 45552
rect 25884 45549 25912 45580
rect 26050 45568 26056 45580
rect 26108 45568 26114 45620
rect 26234 45608 26240 45620
rect 26195 45580 26240 45608
rect 26234 45568 26240 45580
rect 26292 45568 26298 45620
rect 27338 45568 27344 45620
rect 27396 45608 27402 45620
rect 27525 45611 27583 45617
rect 27525 45608 27537 45611
rect 27396 45580 27537 45608
rect 27396 45568 27402 45580
rect 27525 45577 27537 45580
rect 27571 45577 27583 45611
rect 28074 45608 28080 45620
rect 28035 45580 28080 45608
rect 27525 45571 27583 45577
rect 28074 45568 28080 45580
rect 28132 45568 28138 45620
rect 30742 45608 30748 45620
rect 30703 45580 30748 45608
rect 30742 45568 30748 45580
rect 30800 45568 30806 45620
rect 34606 45608 34612 45620
rect 33244 45580 34612 45608
rect 25869 45543 25927 45549
rect 25869 45509 25881 45543
rect 25915 45509 25927 45543
rect 25869 45503 25927 45509
rect 25961 45543 26019 45549
rect 25961 45509 25973 45543
rect 26007 45540 26019 45543
rect 27157 45543 27215 45549
rect 27157 45540 27169 45543
rect 26007 45512 27169 45540
rect 26007 45509 26019 45512
rect 25961 45503 26019 45509
rect 27157 45509 27169 45512
rect 27203 45509 27215 45543
rect 31386 45540 31392 45552
rect 27157 45503 27215 45509
rect 27356 45512 31392 45540
rect 24121 45475 24179 45481
rect 24121 45441 24133 45475
rect 24167 45441 24179 45475
rect 24121 45435 24179 45441
rect 24765 45475 24823 45481
rect 24765 45441 24777 45475
rect 24811 45441 24823 45475
rect 24765 45435 24823 45441
rect 23615 45376 24072 45404
rect 23615 45373 23627 45376
rect 23569 45367 23627 45373
rect 19484 45308 21220 45336
rect 19484 45296 19490 45308
rect 21266 45296 21272 45348
rect 21324 45336 21330 45348
rect 22094 45336 22100 45348
rect 21324 45308 22100 45336
rect 21324 45296 21330 45308
rect 22094 45296 22100 45308
rect 22152 45296 22158 45348
rect 24780 45280 24808 45435
rect 24854 45432 24860 45484
rect 24912 45472 24918 45484
rect 25774 45481 25780 45484
rect 24949 45475 25007 45481
rect 24949 45472 24961 45475
rect 24912 45444 24961 45472
rect 24912 45432 24918 45444
rect 24949 45441 24961 45444
rect 24995 45441 25007 45475
rect 24949 45435 25007 45441
rect 25751 45475 25780 45481
rect 25751 45441 25763 45475
rect 25751 45435 25780 45441
rect 25774 45432 25780 45435
rect 25832 45432 25838 45484
rect 27356 45481 27384 45512
rect 29288 45484 29316 45512
rect 31386 45500 31392 45512
rect 31444 45500 31450 45552
rect 31665 45543 31723 45549
rect 31665 45509 31677 45543
rect 31711 45540 31723 45543
rect 31938 45540 31944 45552
rect 31711 45512 31944 45540
rect 31711 45509 31723 45512
rect 31665 45503 31723 45509
rect 31938 45500 31944 45512
rect 31996 45500 32002 45552
rect 33244 45540 33272 45580
rect 34606 45568 34612 45580
rect 34664 45568 34670 45620
rect 35526 45608 35532 45620
rect 35268 45580 35532 45608
rect 33410 45540 33416 45552
rect 32140 45512 33272 45540
rect 33371 45512 33416 45540
rect 26053 45475 26111 45481
rect 26053 45441 26065 45475
rect 26099 45441 26111 45475
rect 26053 45435 26111 45441
rect 27341 45475 27399 45481
rect 27341 45441 27353 45475
rect 27387 45441 27399 45475
rect 27614 45472 27620 45484
rect 27575 45444 27620 45472
rect 27341 45435 27399 45441
rect 25498 45364 25504 45416
rect 25556 45404 25562 45416
rect 25593 45407 25651 45413
rect 25593 45404 25605 45407
rect 25556 45376 25605 45404
rect 25556 45364 25562 45376
rect 25593 45373 25605 45376
rect 25639 45373 25651 45407
rect 25593 45367 25651 45373
rect 25133 45339 25191 45345
rect 25133 45305 25145 45339
rect 25179 45336 25191 45339
rect 26068 45336 26096 45435
rect 27614 45432 27620 45444
rect 27672 45432 27678 45484
rect 28442 45472 28448 45484
rect 28403 45444 28448 45472
rect 28442 45432 28448 45444
rect 28500 45432 28506 45484
rect 29270 45472 29276 45484
rect 29183 45444 29276 45472
rect 29270 45432 29276 45444
rect 29328 45432 29334 45484
rect 29546 45472 29552 45484
rect 29507 45444 29552 45472
rect 29546 45432 29552 45444
rect 29604 45432 29610 45484
rect 30377 45475 30435 45481
rect 30377 45441 30389 45475
rect 30423 45472 30435 45475
rect 31297 45475 31355 45481
rect 31297 45472 31309 45475
rect 30423 45444 31309 45472
rect 30423 45441 30435 45444
rect 30377 45435 30435 45441
rect 31297 45441 31309 45444
rect 31343 45441 31355 45475
rect 31297 45435 31355 45441
rect 31481 45475 31539 45481
rect 31481 45441 31493 45475
rect 31527 45441 31539 45475
rect 31481 45435 31539 45441
rect 31757 45475 31815 45481
rect 31757 45441 31769 45475
rect 31803 45472 31815 45475
rect 32140 45472 32168 45512
rect 32306 45472 32312 45484
rect 31803 45444 32168 45472
rect 32267 45444 32312 45472
rect 31803 45441 31815 45444
rect 31757 45435 31815 45441
rect 27632 45404 27660 45432
rect 25179 45308 26096 45336
rect 26160 45376 27660 45404
rect 28537 45407 28595 45413
rect 25179 45305 25191 45308
rect 25133 45299 25191 45305
rect 19978 45268 19984 45280
rect 19939 45240 19984 45268
rect 19978 45228 19984 45240
rect 20036 45228 20042 45280
rect 20346 45228 20352 45280
rect 20404 45268 20410 45280
rect 20533 45271 20591 45277
rect 20533 45268 20545 45271
rect 20404 45240 20545 45268
rect 20404 45228 20410 45240
rect 20533 45237 20545 45240
rect 20579 45237 20591 45271
rect 21082 45268 21088 45280
rect 21043 45240 21088 45268
rect 20533 45231 20591 45237
rect 21082 45228 21088 45240
rect 21140 45228 21146 45280
rect 22370 45268 22376 45280
rect 22331 45240 22376 45268
rect 22370 45228 22376 45240
rect 22428 45228 22434 45280
rect 24302 45268 24308 45280
rect 24263 45240 24308 45268
rect 24302 45228 24308 45240
rect 24360 45228 24366 45280
rect 24762 45268 24768 45280
rect 24675 45240 24768 45268
rect 24762 45228 24768 45240
rect 24820 45268 24826 45280
rect 26160 45268 26188 45376
rect 28537 45373 28549 45407
rect 28583 45404 28595 45407
rect 28718 45404 28724 45416
rect 28583 45376 28724 45404
rect 28583 45373 28595 45376
rect 28537 45367 28595 45373
rect 28718 45364 28724 45376
rect 28776 45404 28782 45416
rect 29089 45407 29147 45413
rect 29089 45404 29101 45407
rect 28776 45376 29101 45404
rect 28776 45364 28782 45376
rect 29089 45373 29101 45376
rect 29135 45373 29147 45407
rect 29457 45407 29515 45413
rect 29457 45404 29469 45407
rect 29089 45367 29147 45373
rect 29196 45376 29469 45404
rect 27614 45296 27620 45348
rect 27672 45336 27678 45348
rect 28350 45336 28356 45348
rect 27672 45308 28356 45336
rect 27672 45296 27678 45308
rect 28350 45296 28356 45308
rect 28408 45296 28414 45348
rect 28626 45296 28632 45348
rect 28684 45336 28690 45348
rect 29196 45336 29224 45376
rect 29457 45373 29469 45376
rect 29503 45404 29515 45407
rect 29914 45404 29920 45416
rect 29503 45376 29920 45404
rect 29503 45373 29515 45376
rect 29457 45367 29515 45373
rect 29914 45364 29920 45376
rect 29972 45364 29978 45416
rect 30466 45404 30472 45416
rect 30427 45376 30472 45404
rect 30466 45364 30472 45376
rect 30524 45364 30530 45416
rect 31496 45404 31524 45435
rect 32306 45432 32312 45444
rect 32364 45432 32370 45484
rect 32401 45475 32459 45481
rect 32401 45441 32413 45475
rect 32447 45441 32459 45475
rect 32582 45472 32588 45484
rect 32543 45444 32588 45472
rect 32401 45435 32459 45441
rect 32324 45404 32352 45432
rect 31496 45376 32352 45404
rect 28684 45308 29224 45336
rect 29365 45339 29423 45345
rect 28684 45296 28690 45308
rect 29365 45305 29377 45339
rect 29411 45305 29423 45339
rect 29365 45299 29423 45305
rect 24820 45240 26188 45268
rect 29380 45268 29408 45299
rect 31846 45296 31852 45348
rect 31904 45336 31910 45348
rect 32416 45336 32444 45435
rect 32582 45432 32588 45444
rect 32640 45432 32646 45484
rect 32692 45481 32720 45512
rect 33410 45500 33416 45512
rect 33468 45500 33474 45552
rect 33778 45540 33784 45552
rect 33520 45512 33784 45540
rect 32677 45475 32735 45481
rect 32677 45441 32689 45475
rect 32723 45441 32735 45475
rect 32677 45435 32735 45441
rect 32950 45432 32956 45484
rect 33008 45472 33014 45484
rect 33520 45472 33548 45512
rect 33778 45500 33784 45512
rect 33836 45500 33842 45552
rect 33962 45549 33968 45552
rect 33919 45543 33968 45549
rect 33919 45509 33931 45543
rect 33965 45509 33968 45543
rect 33919 45503 33968 45509
rect 33962 45500 33968 45503
rect 34020 45500 34026 45552
rect 34330 45500 34336 45552
rect 34388 45540 34394 45552
rect 34517 45543 34575 45549
rect 34517 45540 34529 45543
rect 34388 45512 34529 45540
rect 34388 45500 34394 45512
rect 34517 45509 34529 45512
rect 34563 45509 34575 45543
rect 34517 45503 34575 45509
rect 35268 45481 35296 45580
rect 35526 45568 35532 45580
rect 35584 45608 35590 45620
rect 36262 45608 36268 45620
rect 35584 45580 36268 45608
rect 35584 45568 35590 45580
rect 36262 45568 36268 45580
rect 36320 45568 36326 45620
rect 36354 45568 36360 45620
rect 36412 45608 36418 45620
rect 38102 45608 38108 45620
rect 36412 45580 38108 45608
rect 36412 45568 36418 45580
rect 38102 45568 38108 45580
rect 38160 45568 38166 45620
rect 38194 45568 38200 45620
rect 38252 45608 38258 45620
rect 38252 45580 39068 45608
rect 38252 45568 38258 45580
rect 35710 45500 35716 45552
rect 35768 45540 35774 45552
rect 38381 45543 38439 45549
rect 35768 45512 37688 45540
rect 35768 45500 35774 45512
rect 33008 45444 33548 45472
rect 33597 45475 33655 45481
rect 33008 45432 33014 45444
rect 33597 45441 33609 45475
rect 33643 45441 33655 45475
rect 33597 45435 33655 45441
rect 33689 45475 33747 45481
rect 33689 45441 33701 45475
rect 33735 45441 33747 45475
rect 33689 45435 33747 45441
rect 35253 45475 35311 45481
rect 35253 45441 35265 45475
rect 35299 45441 35311 45475
rect 35434 45472 35440 45484
rect 35395 45444 35440 45472
rect 35253 45435 35311 45441
rect 33612 45348 33640 45435
rect 31904 45308 32444 45336
rect 31904 45296 31910 45308
rect 33594 45296 33600 45348
rect 33652 45296 33658 45348
rect 33704 45336 33732 45435
rect 35434 45432 35440 45444
rect 35492 45432 35498 45484
rect 35529 45475 35587 45481
rect 35529 45441 35541 45475
rect 35575 45472 35587 45475
rect 35802 45472 35808 45484
rect 35575 45444 35808 45472
rect 35575 45441 35587 45444
rect 35529 45435 35587 45441
rect 35802 45432 35808 45444
rect 35860 45432 35866 45484
rect 35986 45472 35992 45484
rect 35947 45444 35992 45472
rect 35986 45432 35992 45444
rect 36044 45432 36050 45484
rect 36081 45475 36139 45481
rect 36081 45441 36093 45475
rect 36127 45472 36139 45475
rect 36170 45472 36176 45484
rect 36127 45444 36176 45472
rect 36127 45441 36139 45444
rect 36081 45435 36139 45441
rect 36170 45432 36176 45444
rect 36228 45432 36234 45484
rect 36265 45475 36323 45481
rect 36265 45441 36277 45475
rect 36311 45472 36323 45475
rect 37366 45472 37372 45484
rect 36311 45444 37372 45472
rect 36311 45441 36323 45444
rect 36265 45435 36323 45441
rect 37366 45432 37372 45444
rect 37424 45432 37430 45484
rect 37660 45481 37688 45512
rect 38381 45509 38393 45543
rect 38427 45540 38439 45543
rect 38562 45540 38568 45552
rect 38427 45512 38568 45540
rect 38427 45509 38439 45512
rect 38381 45503 38439 45509
rect 38562 45500 38568 45512
rect 38620 45500 38626 45552
rect 37645 45475 37703 45481
rect 37645 45441 37657 45475
rect 37691 45441 37703 45475
rect 38656 45475 38714 45481
rect 38656 45472 38668 45475
rect 37645 45435 37703 45441
rect 37752 45444 38668 45472
rect 34054 45404 34060 45416
rect 34015 45376 34060 45404
rect 34054 45364 34060 45376
rect 34112 45364 34118 45416
rect 37458 45404 37464 45416
rect 37419 45376 37464 45404
rect 37458 45364 37464 45376
rect 37516 45364 37522 45416
rect 37550 45364 37556 45416
rect 37608 45404 37614 45416
rect 37752 45404 37780 45444
rect 38656 45441 38668 45444
rect 38702 45441 38714 45475
rect 38656 45435 38714 45441
rect 38749 45475 38807 45481
rect 38749 45441 38761 45475
rect 38795 45441 38807 45475
rect 39040 45472 39068 45580
rect 39298 45568 39304 45620
rect 39356 45608 39362 45620
rect 39356 45580 40080 45608
rect 39356 45568 39362 45580
rect 39853 45475 39911 45481
rect 39853 45472 39865 45475
rect 39040 45444 39865 45472
rect 38749 45435 38807 45441
rect 39853 45441 39865 45444
rect 39899 45441 39911 45475
rect 39853 45435 39911 45441
rect 37608 45376 37780 45404
rect 37921 45407 37979 45413
rect 37608 45364 37614 45376
rect 37921 45373 37933 45407
rect 37967 45404 37979 45407
rect 38764 45404 38792 45435
rect 39206 45404 39212 45416
rect 37967 45376 38792 45404
rect 39167 45376 39212 45404
rect 37967 45373 37979 45376
rect 37921 45367 37979 45373
rect 36449 45339 36507 45345
rect 36449 45336 36461 45339
rect 33704 45308 36461 45336
rect 36449 45305 36461 45308
rect 36495 45305 36507 45339
rect 36449 45299 36507 45305
rect 36538 45296 36544 45348
rect 36596 45336 36602 45348
rect 37936 45336 37964 45367
rect 36596 45308 37964 45336
rect 38764 45336 38792 45376
rect 39206 45364 39212 45376
rect 39264 45364 39270 45416
rect 40052 45404 40080 45580
rect 40402 45432 40408 45484
rect 40460 45472 40466 45484
rect 41141 45475 41199 45481
rect 41141 45472 41153 45475
rect 40460 45444 41153 45472
rect 40460 45432 40466 45444
rect 41141 45441 41153 45444
rect 41187 45441 41199 45475
rect 41141 45435 41199 45441
rect 40497 45407 40555 45413
rect 40497 45404 40509 45407
rect 40052 45376 40509 45404
rect 40497 45373 40509 45376
rect 40543 45373 40555 45407
rect 41598 45404 41604 45416
rect 40497 45367 40555 45373
rect 41386 45376 41604 45404
rect 41386 45336 41414 45376
rect 41598 45364 41604 45376
rect 41656 45364 41662 45416
rect 38764 45308 41414 45336
rect 36596 45296 36602 45308
rect 29454 45268 29460 45280
rect 29380 45240 29460 45268
rect 24820 45228 24826 45240
rect 29454 45228 29460 45240
rect 29512 45228 29518 45280
rect 31754 45228 31760 45280
rect 31812 45268 31818 45280
rect 32861 45271 32919 45277
rect 32861 45268 32873 45271
rect 31812 45240 32873 45268
rect 31812 45228 31818 45240
rect 32861 45237 32873 45240
rect 32907 45237 32919 45271
rect 32861 45231 32919 45237
rect 35069 45271 35127 45277
rect 35069 45237 35081 45271
rect 35115 45268 35127 45271
rect 35342 45268 35348 45280
rect 35115 45240 35348 45268
rect 35115 45237 35127 45240
rect 35069 45231 35127 45237
rect 35342 45228 35348 45240
rect 35400 45228 35406 45280
rect 35710 45228 35716 45280
rect 35768 45268 35774 45280
rect 37829 45271 37887 45277
rect 37829 45268 37841 45271
rect 35768 45240 37841 45268
rect 35768 45228 35774 45240
rect 37829 45237 37841 45240
rect 37875 45237 37887 45271
rect 37829 45231 37887 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 19334 45024 19340 45076
rect 19392 45064 19398 45076
rect 19889 45067 19947 45073
rect 19889 45064 19901 45067
rect 19392 45036 19901 45064
rect 19392 45024 19398 45036
rect 19889 45033 19901 45036
rect 19935 45033 19947 45067
rect 22554 45064 22560 45076
rect 22515 45036 22560 45064
rect 19889 45027 19947 45033
rect 22554 45024 22560 45036
rect 22612 45024 22618 45076
rect 22738 45024 22744 45076
rect 22796 45064 22802 45076
rect 23750 45064 23756 45076
rect 22796 45036 23756 45064
rect 22796 45024 22802 45036
rect 20254 44956 20260 45008
rect 20312 44996 20318 45008
rect 21266 44996 21272 45008
rect 20312 44968 21272 44996
rect 20312 44956 20318 44968
rect 21266 44956 21272 44968
rect 21324 44956 21330 45008
rect 23492 45005 23520 45036
rect 23750 45024 23756 45036
rect 23808 45024 23814 45076
rect 25958 45064 25964 45076
rect 25919 45036 25964 45064
rect 25958 45024 25964 45036
rect 26016 45024 26022 45076
rect 26418 45024 26424 45076
rect 26476 45064 26482 45076
rect 29086 45064 29092 45076
rect 26476 45036 29092 45064
rect 26476 45024 26482 45036
rect 29086 45024 29092 45036
rect 29144 45024 29150 45076
rect 30466 45024 30472 45076
rect 30524 45064 30530 45076
rect 31297 45067 31355 45073
rect 31297 45064 31309 45067
rect 30524 45036 31309 45064
rect 30524 45024 30530 45036
rect 31297 45033 31309 45036
rect 31343 45033 31355 45067
rect 31297 45027 31355 45033
rect 31938 45024 31944 45076
rect 31996 45064 32002 45076
rect 32582 45064 32588 45076
rect 31996 45036 32588 45064
rect 31996 45024 32002 45036
rect 32582 45024 32588 45036
rect 32640 45024 32646 45076
rect 33137 45067 33195 45073
rect 33137 45033 33149 45067
rect 33183 45064 33195 45067
rect 33502 45064 33508 45076
rect 33183 45036 33508 45064
rect 33183 45033 33195 45036
rect 33137 45027 33195 45033
rect 33502 45024 33508 45036
rect 33560 45024 33566 45076
rect 33778 45024 33784 45076
rect 33836 45064 33842 45076
rect 33965 45067 34023 45073
rect 33965 45064 33977 45067
rect 33836 45036 33977 45064
rect 33836 45024 33842 45036
rect 33965 45033 33977 45036
rect 34011 45033 34023 45067
rect 37093 45067 37151 45073
rect 37093 45064 37105 45067
rect 33965 45027 34023 45033
rect 34072 45036 37105 45064
rect 23477 44999 23535 45005
rect 23477 44965 23489 44999
rect 23523 44965 23535 44999
rect 23477 44959 23535 44965
rect 26234 44956 26240 45008
rect 26292 44996 26298 45008
rect 28721 44999 28779 45005
rect 28721 44996 28733 44999
rect 26292 44968 28733 44996
rect 26292 44956 26298 44968
rect 28721 44965 28733 44968
rect 28767 44965 28779 44999
rect 28721 44959 28779 44965
rect 29362 44956 29368 45008
rect 29420 44996 29426 45008
rect 30561 44999 30619 45005
rect 30561 44996 30573 44999
rect 29420 44968 30573 44996
rect 29420 44956 29426 44968
rect 30561 44965 30573 44968
rect 30607 44965 30619 44999
rect 31389 44999 31447 45005
rect 31389 44996 31401 44999
rect 30561 44959 30619 44965
rect 30760 44968 31401 44996
rect 20530 44928 20536 44940
rect 20491 44900 20536 44928
rect 20530 44888 20536 44900
rect 20588 44928 20594 44940
rect 21634 44928 21640 44940
rect 20588 44900 21404 44928
rect 21595 44900 21640 44928
rect 20588 44888 20594 44900
rect 20070 44860 20076 44872
rect 20031 44832 20076 44860
rect 20070 44820 20076 44832
rect 20128 44820 20134 44872
rect 20717 44863 20775 44869
rect 20717 44829 20729 44863
rect 20763 44860 20775 44863
rect 20806 44860 20812 44872
rect 20763 44832 20812 44860
rect 20763 44829 20775 44832
rect 20717 44823 20775 44829
rect 20806 44820 20812 44832
rect 20864 44820 20870 44872
rect 21376 44869 21404 44900
rect 21634 44888 21640 44900
rect 21692 44888 21698 44940
rect 22572 44900 23520 44928
rect 22572 44869 22600 44900
rect 23492 44872 23520 44900
rect 23658 44888 23664 44940
rect 23716 44928 23722 44940
rect 23753 44931 23811 44937
rect 23753 44928 23765 44931
rect 23716 44900 23765 44928
rect 23716 44888 23722 44900
rect 23753 44897 23765 44900
rect 23799 44928 23811 44931
rect 27614 44928 27620 44940
rect 23799 44900 24716 44928
rect 23799 44897 23811 44900
rect 23753 44891 23811 44897
rect 21361 44863 21419 44869
rect 21361 44829 21373 44863
rect 21407 44829 21419 44863
rect 21361 44823 21419 44829
rect 22557 44863 22615 44869
rect 22557 44829 22569 44863
rect 22603 44829 22615 44863
rect 22738 44860 22744 44872
rect 22699 44832 22744 44860
rect 22557 44823 22615 44829
rect 22738 44820 22744 44832
rect 22796 44820 22802 44872
rect 22833 44863 22891 44869
rect 22833 44829 22845 44863
rect 22879 44829 22891 44863
rect 22833 44823 22891 44829
rect 22848 44792 22876 44823
rect 23290 44820 23296 44872
rect 23348 44820 23354 44872
rect 23474 44820 23480 44872
rect 23532 44820 23538 44872
rect 24578 44860 24584 44872
rect 24539 44832 24584 44860
rect 24578 44820 24584 44832
rect 24636 44820 24642 44872
rect 24688 44869 24716 44900
rect 27080 44900 27620 44928
rect 24673 44863 24731 44869
rect 24673 44829 24685 44863
rect 24719 44829 24731 44863
rect 24854 44860 24860 44872
rect 24815 44832 24860 44860
rect 24673 44823 24731 44829
rect 24854 44820 24860 44832
rect 24912 44820 24918 44872
rect 24949 44863 25007 44869
rect 24949 44829 24961 44863
rect 24995 44860 25007 44863
rect 25314 44860 25320 44872
rect 24995 44832 25320 44860
rect 24995 44829 25007 44832
rect 24949 44823 25007 44829
rect 25314 44820 25320 44832
rect 25372 44820 25378 44872
rect 25866 44860 25872 44872
rect 25827 44832 25872 44860
rect 25866 44820 25872 44832
rect 25924 44820 25930 44872
rect 27080 44869 27108 44900
rect 27614 44888 27620 44900
rect 27672 44888 27678 44940
rect 28000 44900 29040 44928
rect 27065 44863 27123 44869
rect 27065 44860 27077 44863
rect 26252 44832 27077 44860
rect 23308 44792 23336 44820
rect 25133 44795 25191 44801
rect 25133 44792 25145 44795
rect 22848 44764 25145 44792
rect 25133 44761 25145 44764
rect 25179 44761 25191 44795
rect 25133 44755 25191 44761
rect 18877 44727 18935 44733
rect 18877 44693 18889 44727
rect 18923 44724 18935 44727
rect 19978 44724 19984 44736
rect 18923 44696 19984 44724
rect 18923 44693 18935 44696
rect 18877 44687 18935 44693
rect 19978 44684 19984 44696
rect 20036 44684 20042 44736
rect 20806 44684 20812 44736
rect 20864 44724 20870 44736
rect 20901 44727 20959 44733
rect 20901 44724 20913 44727
rect 20864 44696 20913 44724
rect 20864 44684 20870 44696
rect 20901 44693 20913 44696
rect 20947 44693 20959 44727
rect 23290 44724 23296 44736
rect 23251 44696 23296 44724
rect 20901 44687 20959 44693
rect 23290 44684 23296 44696
rect 23348 44684 23354 44736
rect 24302 44684 24308 44736
rect 24360 44724 24366 44736
rect 26252 44724 26280 44832
rect 27065 44829 27077 44832
rect 27111 44829 27123 44863
rect 27065 44823 27123 44829
rect 27341 44863 27399 44869
rect 27341 44829 27353 44863
rect 27387 44860 27399 44863
rect 27522 44860 27528 44872
rect 27387 44832 27528 44860
rect 27387 44829 27399 44832
rect 27341 44823 27399 44829
rect 27522 44820 27528 44832
rect 27580 44820 27586 44872
rect 27798 44820 27804 44872
rect 27856 44860 27862 44872
rect 28000 44869 28028 44900
rect 27985 44863 28043 44869
rect 27985 44860 27997 44863
rect 27856 44832 27997 44860
rect 27856 44820 27862 44832
rect 27985 44829 27997 44832
rect 28031 44829 28043 44863
rect 27985 44823 28043 44829
rect 28077 44863 28135 44869
rect 28077 44829 28089 44863
rect 28123 44829 28135 44863
rect 28077 44823 28135 44829
rect 28169 44863 28227 44869
rect 28169 44829 28181 44863
rect 28215 44860 28227 44863
rect 28534 44860 28540 44872
rect 28215 44832 28540 44860
rect 28215 44829 28227 44832
rect 28169 44823 28227 44829
rect 28092 44736 28120 44823
rect 28534 44820 28540 44832
rect 28592 44820 28598 44872
rect 28718 44860 28724 44872
rect 28679 44832 28724 44860
rect 28718 44820 28724 44832
rect 28776 44820 28782 44872
rect 29012 44869 29040 44900
rect 28997 44863 29055 44869
rect 28997 44829 29009 44863
rect 29043 44860 29055 44863
rect 29546 44860 29552 44872
rect 29043 44832 29552 44860
rect 29043 44829 29055 44832
rect 28997 44823 29055 44829
rect 29546 44820 29552 44832
rect 29604 44860 29610 44872
rect 29604 44832 29776 44860
rect 29604 44820 29610 44832
rect 28442 44752 28448 44804
rect 28500 44792 28506 44804
rect 28905 44795 28963 44801
rect 28905 44792 28917 44795
rect 28500 44764 28917 44792
rect 28500 44752 28506 44764
rect 28905 44761 28917 44764
rect 28951 44761 28963 44795
rect 28905 44755 28963 44761
rect 24360 44696 26280 44724
rect 26329 44727 26387 44733
rect 24360 44684 24366 44696
rect 26329 44693 26341 44727
rect 26375 44724 26387 44727
rect 26602 44724 26608 44736
rect 26375 44696 26608 44724
rect 26375 44693 26387 44696
rect 26329 44687 26387 44693
rect 26602 44684 26608 44696
rect 26660 44684 26666 44736
rect 26878 44724 26884 44736
rect 26839 44696 26884 44724
rect 26878 44684 26884 44696
rect 26936 44684 26942 44736
rect 27249 44727 27307 44733
rect 27249 44693 27261 44727
rect 27295 44724 27307 44727
rect 27430 44724 27436 44736
rect 27295 44696 27436 44724
rect 27295 44693 27307 44696
rect 27249 44687 27307 44693
rect 27430 44684 27436 44696
rect 27488 44724 27494 44736
rect 27801 44727 27859 44733
rect 27801 44724 27813 44727
rect 27488 44696 27813 44724
rect 27488 44684 27494 44696
rect 27801 44693 27813 44696
rect 27847 44693 27859 44727
rect 27801 44687 27859 44693
rect 28074 44684 28080 44736
rect 28132 44684 28138 44736
rect 29748 44733 29776 44832
rect 29822 44820 29828 44872
rect 29880 44860 29886 44872
rect 29947 44863 30005 44869
rect 29947 44860 29959 44863
rect 29880 44832 29959 44860
rect 29880 44820 29886 44832
rect 29947 44829 29959 44832
rect 29993 44829 30005 44863
rect 29947 44823 30005 44829
rect 30098 44820 30104 44872
rect 30156 44860 30162 44872
rect 30760 44869 30788 44968
rect 31389 44965 31401 44968
rect 31435 44996 31447 44999
rect 32030 44996 32036 45008
rect 31435 44968 32036 44996
rect 31435 44965 31447 44968
rect 31389 44959 31447 44965
rect 32030 44956 32036 44968
rect 32088 44956 32094 45008
rect 33226 44956 33232 45008
rect 33284 44996 33290 45008
rect 33796 44996 33824 45024
rect 33284 44968 33824 44996
rect 33284 44956 33290 44968
rect 31757 44931 31815 44937
rect 31757 44897 31769 44931
rect 31803 44928 31815 44931
rect 31846 44928 31852 44940
rect 31803 44900 31852 44928
rect 31803 44897 31815 44900
rect 31757 44891 31815 44897
rect 31846 44888 31852 44900
rect 31904 44888 31910 44940
rect 32490 44888 32496 44940
rect 32548 44928 32554 44940
rect 32861 44931 32919 44937
rect 32861 44928 32873 44931
rect 32548 44900 32873 44928
rect 32548 44888 32554 44900
rect 32861 44897 32873 44900
rect 32907 44928 32919 44931
rect 34072 44928 34100 45036
rect 37093 45033 37105 45036
rect 37139 45033 37151 45067
rect 37093 45027 37151 45033
rect 37642 45024 37648 45076
rect 37700 45064 37706 45076
rect 38013 45067 38071 45073
rect 38013 45064 38025 45067
rect 37700 45036 38025 45064
rect 37700 45024 37706 45036
rect 38013 45033 38025 45036
rect 38059 45033 38071 45067
rect 38013 45027 38071 45033
rect 38654 45024 38660 45076
rect 38712 45064 38718 45076
rect 39301 45067 39359 45073
rect 39301 45064 39313 45067
rect 38712 45036 39313 45064
rect 38712 45024 38718 45036
rect 39301 45033 39313 45036
rect 39347 45033 39359 45067
rect 40034 45064 40040 45076
rect 39995 45036 40040 45064
rect 39301 45027 39359 45033
rect 40034 45024 40040 45036
rect 40092 45024 40098 45076
rect 40773 45067 40831 45073
rect 40773 45033 40785 45067
rect 40819 45064 40831 45067
rect 40862 45064 40868 45076
rect 40819 45036 40868 45064
rect 40819 45033 40831 45036
rect 40773 45027 40831 45033
rect 40862 45024 40868 45036
rect 40920 45024 40926 45076
rect 34606 44956 34612 45008
rect 34664 44996 34670 45008
rect 34885 44999 34943 45005
rect 34885 44996 34897 44999
rect 34664 44968 34897 44996
rect 34664 44956 34670 44968
rect 34885 44965 34897 44968
rect 34931 44965 34943 44999
rect 34885 44959 34943 44965
rect 35342 44956 35348 45008
rect 35400 44956 35406 45008
rect 35360 44928 35388 44956
rect 32907 44900 34100 44928
rect 35268 44900 35388 44928
rect 36081 44931 36139 44937
rect 32907 44897 32919 44900
rect 32861 44891 32919 44897
rect 30745 44863 30803 44869
rect 30156 44832 30201 44860
rect 30156 44820 30162 44832
rect 30745 44829 30757 44863
rect 30791 44829 30803 44863
rect 30745 44823 30803 44829
rect 30837 44863 30895 44869
rect 30837 44829 30849 44863
rect 30883 44860 30895 44863
rect 31662 44860 31668 44872
rect 30883 44832 31668 44860
rect 30883 44829 30895 44832
rect 30837 44823 30895 44829
rect 31662 44820 31668 44832
rect 31720 44820 31726 44872
rect 32766 44860 32772 44872
rect 32727 44832 32772 44860
rect 32766 44820 32772 44832
rect 32824 44820 32830 44872
rect 33873 44863 33931 44869
rect 33873 44829 33885 44863
rect 33919 44829 33931 44863
rect 35066 44860 35072 44872
rect 35027 44832 35072 44860
rect 33873 44823 33931 44829
rect 30561 44795 30619 44801
rect 30561 44761 30573 44795
rect 30607 44792 30619 44795
rect 32122 44792 32128 44804
rect 30607 44764 32128 44792
rect 30607 44761 30619 44764
rect 30561 44755 30619 44761
rect 32122 44752 32128 44764
rect 32180 44752 32186 44804
rect 33888 44792 33916 44823
rect 35066 44820 35072 44832
rect 35124 44820 35130 44872
rect 35268 44869 35296 44900
rect 36081 44897 36093 44931
rect 36127 44928 36139 44931
rect 36262 44928 36268 44940
rect 36127 44900 36268 44928
rect 36127 44897 36139 44900
rect 36081 44891 36139 44897
rect 36262 44888 36268 44900
rect 36320 44888 36326 44940
rect 37458 44928 37464 44940
rect 37419 44900 37464 44928
rect 37458 44888 37464 44900
rect 37516 44888 37522 44940
rect 38657 44931 38715 44937
rect 38657 44897 38669 44931
rect 38703 44928 38715 44931
rect 38746 44928 38752 44940
rect 38703 44900 38752 44928
rect 38703 44897 38715 44900
rect 38657 44891 38715 44897
rect 38746 44888 38752 44900
rect 38804 44888 38810 44940
rect 35253 44863 35311 44869
rect 35253 44829 35265 44863
rect 35299 44829 35311 44863
rect 35253 44823 35311 44829
rect 35345 44863 35403 44869
rect 35345 44829 35357 44863
rect 35391 44829 35403 44863
rect 36173 44863 36231 44869
rect 36173 44860 36185 44863
rect 35345 44823 35403 44829
rect 35452 44832 36185 44860
rect 34146 44792 34152 44804
rect 33888 44764 34152 44792
rect 34146 44752 34152 44764
rect 34204 44792 34210 44804
rect 34204 44764 34744 44792
rect 34204 44752 34210 44764
rect 29733 44727 29791 44733
rect 29733 44693 29745 44727
rect 29779 44724 29791 44727
rect 30006 44724 30012 44736
rect 29779 44696 30012 44724
rect 29779 44693 29791 44696
rect 29733 44687 29791 44693
rect 30006 44684 30012 44696
rect 30064 44684 30070 44736
rect 34333 44727 34391 44733
rect 34333 44693 34345 44727
rect 34379 44724 34391 44727
rect 34606 44724 34612 44736
rect 34379 44696 34612 44724
rect 34379 44693 34391 44696
rect 34333 44687 34391 44693
rect 34606 44684 34612 44696
rect 34664 44684 34670 44736
rect 34716 44724 34744 44764
rect 34974 44752 34980 44804
rect 35032 44792 35038 44804
rect 35360 44792 35388 44823
rect 35032 44764 35388 44792
rect 35032 44752 35038 44764
rect 35452 44724 35480 44832
rect 36173 44829 36185 44832
rect 36219 44860 36231 44863
rect 37366 44860 37372 44872
rect 36219 44832 36676 44860
rect 37279 44832 37372 44860
rect 36219 44829 36231 44832
rect 36173 44823 36231 44829
rect 35618 44752 35624 44804
rect 35676 44792 35682 44804
rect 36648 44792 36676 44832
rect 37366 44820 37372 44832
rect 37424 44860 37430 44872
rect 38010 44860 38016 44872
rect 37424 44832 38016 44860
rect 37424 44820 37430 44832
rect 38010 44820 38016 44832
rect 38068 44820 38074 44872
rect 38102 44820 38108 44872
rect 38160 44860 38166 44872
rect 38197 44863 38255 44869
rect 38197 44860 38209 44863
rect 38160 44832 38209 44860
rect 38160 44820 38166 44832
rect 38197 44829 38209 44832
rect 38243 44829 38255 44863
rect 38197 44823 38255 44829
rect 36906 44792 36912 44804
rect 35676 44764 36584 44792
rect 36648 44764 36912 44792
rect 35676 44752 35682 44764
rect 34716 44696 35480 44724
rect 35802 44684 35808 44736
rect 35860 44724 35866 44736
rect 36556 44733 36584 44764
rect 36906 44752 36912 44764
rect 36964 44792 36970 44804
rect 37918 44792 37924 44804
rect 36964 44764 37924 44792
rect 36964 44752 36970 44764
rect 37918 44752 37924 44764
rect 37976 44792 37982 44804
rect 38286 44792 38292 44804
rect 37976 44764 38292 44792
rect 37976 44752 37982 44764
rect 38286 44752 38292 44764
rect 38344 44752 38350 44804
rect 35897 44727 35955 44733
rect 35897 44724 35909 44727
rect 35860 44696 35909 44724
rect 35860 44684 35866 44696
rect 35897 44693 35909 44696
rect 35943 44693 35955 44727
rect 35897 44687 35955 44693
rect 36541 44727 36599 44733
rect 36541 44693 36553 44727
rect 36587 44724 36599 44727
rect 36814 44724 36820 44736
rect 36587 44696 36820 44724
rect 36587 44693 36599 44696
rect 36541 44687 36599 44693
rect 36814 44684 36820 44696
rect 36872 44724 36878 44736
rect 38470 44724 38476 44736
rect 36872 44696 38476 44724
rect 36872 44684 36878 44696
rect 38470 44684 38476 44696
rect 38528 44684 38534 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 20254 44520 20260 44532
rect 20215 44492 20260 44520
rect 20254 44480 20260 44492
rect 20312 44480 20318 44532
rect 20993 44523 21051 44529
rect 20993 44489 21005 44523
rect 21039 44489 21051 44523
rect 20993 44483 21051 44489
rect 22741 44523 22799 44529
rect 22741 44489 22753 44523
rect 22787 44489 22799 44523
rect 22741 44483 22799 44489
rect 23753 44523 23811 44529
rect 23753 44489 23765 44523
rect 23799 44520 23811 44523
rect 23842 44520 23848 44532
rect 23799 44492 23848 44520
rect 23799 44489 23811 44492
rect 23753 44483 23811 44489
rect 19426 44412 19432 44464
rect 19484 44452 19490 44464
rect 21008 44452 21036 44483
rect 19484 44424 21036 44452
rect 22756 44452 22784 44483
rect 23842 44480 23848 44492
rect 23900 44520 23906 44532
rect 24210 44520 24216 44532
rect 23900 44492 24216 44520
rect 23900 44480 23906 44492
rect 24210 44480 24216 44492
rect 24268 44480 24274 44532
rect 25685 44523 25743 44529
rect 25685 44489 25697 44523
rect 25731 44520 25743 44523
rect 25774 44520 25780 44532
rect 25731 44492 25780 44520
rect 25731 44489 25743 44492
rect 25685 44483 25743 44489
rect 25774 44480 25780 44492
rect 25832 44480 25838 44532
rect 25866 44480 25872 44532
rect 25924 44520 25930 44532
rect 28261 44523 28319 44529
rect 25924 44492 27936 44520
rect 25924 44480 25930 44492
rect 25130 44452 25136 44464
rect 22756 44424 25136 44452
rect 19484 44412 19490 44424
rect 25130 44412 25136 44424
rect 25188 44452 25194 44464
rect 25958 44452 25964 44464
rect 25188 44424 25964 44452
rect 25188 44412 25194 44424
rect 25958 44412 25964 44424
rect 26016 44412 26022 44464
rect 26513 44455 26571 44461
rect 26513 44421 26525 44455
rect 26559 44452 26571 44455
rect 26878 44452 26884 44464
rect 26559 44424 26884 44452
rect 26559 44421 26571 44424
rect 26513 44415 26571 44421
rect 26878 44412 26884 44424
rect 26936 44412 26942 44464
rect 27908 44452 27936 44492
rect 28261 44489 28273 44523
rect 28307 44520 28319 44523
rect 28534 44520 28540 44532
rect 28307 44492 28540 44520
rect 28307 44489 28319 44492
rect 28261 44483 28319 44489
rect 28534 44480 28540 44492
rect 28592 44480 28598 44532
rect 32306 44520 32312 44532
rect 32267 44492 32312 44520
rect 32306 44480 32312 44492
rect 32364 44480 32370 44532
rect 33594 44480 33600 44532
rect 33652 44520 33658 44532
rect 33689 44523 33747 44529
rect 33689 44520 33701 44523
rect 33652 44492 33701 44520
rect 33652 44480 33658 44492
rect 33689 44489 33701 44492
rect 33735 44489 33747 44523
rect 33689 44483 33747 44489
rect 34606 44480 34612 44532
rect 34664 44520 34670 44532
rect 34974 44520 34980 44532
rect 34664 44492 34980 44520
rect 34664 44480 34670 44492
rect 34974 44480 34980 44492
rect 35032 44480 35038 44532
rect 35069 44523 35127 44529
rect 35069 44489 35081 44523
rect 35115 44489 35127 44523
rect 35069 44483 35127 44489
rect 28074 44452 28080 44464
rect 27908 44424 28080 44452
rect 20806 44384 20812 44396
rect 20767 44356 20812 44384
rect 20806 44344 20812 44356
rect 20864 44344 20870 44396
rect 22557 44387 22615 44393
rect 22557 44353 22569 44387
rect 22603 44384 22615 44387
rect 22646 44384 22652 44396
rect 22603 44356 22652 44384
rect 22603 44353 22615 44356
rect 22557 44347 22615 44353
rect 22646 44344 22652 44356
rect 22704 44344 22710 44396
rect 23385 44387 23443 44393
rect 23385 44353 23397 44387
rect 23431 44384 23443 44387
rect 23750 44384 23756 44396
rect 23431 44356 23756 44384
rect 23431 44353 23443 44356
rect 23385 44347 23443 44353
rect 23750 44344 23756 44356
rect 23808 44344 23814 44396
rect 24673 44387 24731 44393
rect 24673 44353 24685 44387
rect 24719 44353 24731 44387
rect 24673 44347 24731 44353
rect 23290 44316 23296 44328
rect 23251 44288 23296 44316
rect 23290 44276 23296 44288
rect 23348 44276 23354 44328
rect 24688 44316 24716 44347
rect 24762 44344 24768 44396
rect 24820 44384 24826 44396
rect 25314 44384 25320 44396
rect 24820 44356 24865 44384
rect 25275 44356 25320 44384
rect 24820 44344 24826 44356
rect 25314 44344 25320 44356
rect 25372 44344 25378 44396
rect 25501 44387 25559 44393
rect 25501 44353 25513 44387
rect 25547 44384 25559 44387
rect 25590 44384 25596 44396
rect 25547 44356 25596 44384
rect 25547 44353 25559 44356
rect 25501 44347 25559 44353
rect 25590 44344 25596 44356
rect 25648 44344 25654 44396
rect 26329 44387 26387 44393
rect 26329 44353 26341 44387
rect 26375 44353 26387 44387
rect 26329 44347 26387 44353
rect 25332 44316 25360 44344
rect 26145 44319 26203 44325
rect 26145 44316 26157 44319
rect 24688 44288 25176 44316
rect 25332 44288 26157 44316
rect 25148 44260 25176 44288
rect 26145 44285 26157 44288
rect 26191 44285 26203 44319
rect 26344 44316 26372 44347
rect 26602 44344 26608 44396
rect 26660 44384 26666 44396
rect 27798 44384 27804 44396
rect 26660 44356 26705 44384
rect 27759 44356 27804 44384
rect 26660 44344 26666 44356
rect 27798 44344 27804 44356
rect 27856 44344 27862 44396
rect 27908 44393 27936 44424
rect 28074 44412 28080 44424
rect 28132 44452 28138 44464
rect 29454 44452 29460 44464
rect 28132 44424 29460 44452
rect 28132 44412 28138 44424
rect 29454 44412 29460 44424
rect 29512 44412 29518 44464
rect 29730 44412 29736 44464
rect 29788 44452 29794 44464
rect 33137 44455 33195 44461
rect 33137 44452 33149 44455
rect 29788 44424 33149 44452
rect 29788 44412 29794 44424
rect 33137 44421 33149 44424
rect 33183 44421 33195 44455
rect 33137 44415 33195 44421
rect 33873 44455 33931 44461
rect 33873 44421 33885 44455
rect 33919 44452 33931 44455
rect 34790 44452 34796 44464
rect 33919 44424 34796 44452
rect 33919 44421 33931 44424
rect 33873 44415 33931 44421
rect 34790 44412 34796 44424
rect 34848 44412 34854 44464
rect 35084 44452 35112 44483
rect 35434 44480 35440 44532
rect 35492 44520 35498 44532
rect 36449 44523 36507 44529
rect 36449 44520 36461 44523
rect 35492 44492 36461 44520
rect 35492 44480 35498 44492
rect 36449 44489 36461 44492
rect 36495 44489 36507 44523
rect 36906 44520 36912 44532
rect 36449 44483 36507 44489
rect 36740 44492 36912 44520
rect 35710 44452 35716 44464
rect 35084 44424 35716 44452
rect 35710 44412 35716 44424
rect 35768 44412 35774 44464
rect 36740 44415 36768 44492
rect 36906 44480 36912 44492
rect 36964 44480 36970 44532
rect 37458 44520 37464 44532
rect 37419 44492 37464 44520
rect 37458 44480 37464 44492
rect 37516 44480 37522 44532
rect 38102 44480 38108 44532
rect 38160 44520 38166 44532
rect 38381 44523 38439 44529
rect 38381 44520 38393 44523
rect 38160 44492 38393 44520
rect 38160 44480 38166 44492
rect 38381 44489 38393 44492
rect 38427 44489 38439 44523
rect 38381 44483 38439 44489
rect 36725 44409 36783 44415
rect 27893 44387 27951 44393
rect 27893 44353 27905 44387
rect 27939 44353 27951 44387
rect 27893 44347 27951 44353
rect 29089 44387 29147 44393
rect 29089 44353 29101 44387
rect 29135 44384 29147 44387
rect 29270 44384 29276 44396
rect 29135 44356 29276 44384
rect 29135 44353 29147 44356
rect 29089 44347 29147 44353
rect 29270 44344 29276 44356
rect 29328 44344 29334 44396
rect 32490 44384 32496 44396
rect 32451 44356 32496 44384
rect 32490 44344 32496 44356
rect 32548 44344 32554 44396
rect 34057 44387 34115 44393
rect 34057 44353 34069 44387
rect 34103 44353 34115 44387
rect 34057 44347 34115 44353
rect 34701 44387 34759 44393
rect 34701 44353 34713 44387
rect 34747 44353 34759 44387
rect 34701 44347 34759 44353
rect 27338 44316 27344 44328
rect 26344 44288 27344 44316
rect 26145 44279 26203 44285
rect 27338 44276 27344 44288
rect 27396 44276 27402 44328
rect 29178 44316 29184 44328
rect 29139 44288 29184 44316
rect 29178 44276 29184 44288
rect 29236 44276 29242 44328
rect 30190 44316 30196 44328
rect 30151 44288 30196 44316
rect 30190 44276 30196 44288
rect 30248 44276 30254 44328
rect 31389 44319 31447 44325
rect 31389 44285 31401 44319
rect 31435 44285 31447 44319
rect 31570 44316 31576 44328
rect 31531 44288 31576 44316
rect 31389 44279 31447 44285
rect 22097 44251 22155 44257
rect 22097 44217 22109 44251
rect 22143 44248 22155 44251
rect 22143 44220 24716 44248
rect 22143 44217 22155 44220
rect 22097 44211 22155 44217
rect 19797 44183 19855 44189
rect 19797 44149 19809 44183
rect 19843 44180 19855 44183
rect 19978 44180 19984 44192
rect 19843 44152 19984 44180
rect 19843 44149 19855 44152
rect 19797 44143 19855 44149
rect 19978 44140 19984 44152
rect 20036 44180 20042 44192
rect 20714 44180 20720 44192
rect 20036 44152 20720 44180
rect 20036 44140 20042 44152
rect 20714 44140 20720 44152
rect 20772 44140 20778 44192
rect 23934 44140 23940 44192
rect 23992 44180 23998 44192
rect 24489 44183 24547 44189
rect 24489 44180 24501 44183
rect 23992 44152 24501 44180
rect 23992 44140 23998 44152
rect 24489 44149 24501 44152
rect 24535 44180 24547 44183
rect 24578 44180 24584 44192
rect 24535 44152 24584 44180
rect 24535 44149 24547 44152
rect 24489 44143 24547 44149
rect 24578 44140 24584 44152
rect 24636 44140 24642 44192
rect 24688 44180 24716 44220
rect 25130 44208 25136 44260
rect 25188 44248 25194 44260
rect 28721 44251 28779 44257
rect 28721 44248 28733 44251
rect 25188 44220 28733 44248
rect 25188 44208 25194 44220
rect 28721 44217 28733 44220
rect 28767 44217 28779 44251
rect 28721 44211 28779 44217
rect 29086 44208 29092 44260
rect 29144 44248 29150 44260
rect 31404 44248 31432 44279
rect 31570 44276 31576 44288
rect 31628 44276 31634 44328
rect 32677 44319 32735 44325
rect 32677 44285 32689 44319
rect 32723 44316 32735 44319
rect 32766 44316 32772 44328
rect 32723 44288 32772 44316
rect 32723 44285 32735 44288
rect 32677 44279 32735 44285
rect 32766 44276 32772 44288
rect 32824 44316 32830 44328
rect 34072 44316 34100 44347
rect 34606 44316 34612 44328
rect 32824 44288 34100 44316
rect 34567 44288 34612 44316
rect 32824 44276 32830 44288
rect 29144 44220 31432 44248
rect 34072 44248 34100 44288
rect 34606 44276 34612 44288
rect 34664 44276 34670 44328
rect 34716 44316 34744 44347
rect 35342 44344 35348 44396
rect 35400 44384 35406 44396
rect 35529 44387 35587 44393
rect 35529 44384 35541 44387
rect 35400 44356 35541 44384
rect 35400 44344 35406 44356
rect 35529 44353 35541 44356
rect 35575 44353 35587 44387
rect 35529 44347 35587 44353
rect 36262 44344 36268 44396
rect 36320 44384 36326 44396
rect 36633 44387 36691 44393
rect 36633 44384 36645 44387
rect 36320 44356 36645 44384
rect 36320 44344 36326 44356
rect 36633 44353 36645 44356
rect 36679 44353 36691 44387
rect 36725 44375 36737 44409
rect 36771 44375 36783 44409
rect 36725 44369 36783 44375
rect 36817 44387 36875 44393
rect 36633 44347 36691 44353
rect 36817 44353 36829 44387
rect 36863 44382 36875 44387
rect 36906 44382 36912 44396
rect 36863 44354 36912 44382
rect 36863 44353 36875 44354
rect 36817 44347 36875 44353
rect 35989 44319 36047 44325
rect 35989 44316 36001 44319
rect 34716 44288 36001 44316
rect 35989 44285 36001 44288
rect 36035 44285 36047 44319
rect 36648 44316 36676 44347
rect 36906 44344 36912 44354
rect 36964 44344 36970 44396
rect 37645 44387 37703 44393
rect 37645 44353 37657 44387
rect 37691 44384 37703 44387
rect 38562 44384 38568 44396
rect 37691 44356 38568 44384
rect 37691 44353 37703 44356
rect 37645 44347 37703 44353
rect 36648 44288 36768 44316
rect 35989 44279 36047 44285
rect 36078 44248 36084 44260
rect 34072 44220 36084 44248
rect 29144 44208 29150 44220
rect 36078 44208 36084 44220
rect 36136 44208 36142 44260
rect 36740 44248 36768 44288
rect 37660 44248 37688 44347
rect 38562 44344 38568 44356
rect 38620 44344 38626 44396
rect 37918 44316 37924 44328
rect 37879 44288 37924 44316
rect 37918 44276 37924 44288
rect 37976 44276 37982 44328
rect 36740 44220 37688 44248
rect 37829 44251 37887 44257
rect 37829 44217 37841 44251
rect 37875 44248 37887 44251
rect 38470 44248 38476 44260
rect 37875 44220 38476 44248
rect 37875 44217 37887 44220
rect 37829 44211 37887 44217
rect 38470 44208 38476 44220
rect 38528 44208 38534 44260
rect 25406 44180 25412 44192
rect 24688 44152 25412 44180
rect 25406 44140 25412 44152
rect 25464 44140 25470 44192
rect 27522 44140 27528 44192
rect 27580 44180 27586 44192
rect 27617 44183 27675 44189
rect 27617 44180 27629 44183
rect 27580 44152 27629 44180
rect 27580 44140 27586 44152
rect 27617 44149 27629 44152
rect 27663 44149 27675 44183
rect 27617 44143 27675 44149
rect 35066 44140 35072 44192
rect 35124 44180 35130 44192
rect 35621 44183 35679 44189
rect 35621 44180 35633 44183
rect 35124 44152 35633 44180
rect 35124 44140 35130 44152
rect 35621 44149 35633 44152
rect 35667 44180 35679 44183
rect 35710 44180 35716 44192
rect 35667 44152 35716 44180
rect 35667 44149 35679 44152
rect 35621 44143 35679 44149
rect 35710 44140 35716 44152
rect 35768 44140 35774 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 20441 43979 20499 43985
rect 20441 43945 20453 43979
rect 20487 43976 20499 43979
rect 20530 43976 20536 43988
rect 20487 43948 20536 43976
rect 20487 43945 20499 43948
rect 20441 43939 20499 43945
rect 20530 43936 20536 43948
rect 20588 43936 20594 43988
rect 21082 43936 21088 43988
rect 21140 43976 21146 43988
rect 22189 43979 22247 43985
rect 22189 43976 22201 43979
rect 21140 43948 22201 43976
rect 21140 43936 21146 43948
rect 22189 43945 22201 43948
rect 22235 43945 22247 43979
rect 22189 43939 22247 43945
rect 23198 43936 23204 43988
rect 23256 43976 23262 43988
rect 23293 43979 23351 43985
rect 23293 43976 23305 43979
rect 23256 43948 23305 43976
rect 23256 43936 23262 43948
rect 23293 43945 23305 43948
rect 23339 43945 23351 43979
rect 23750 43976 23756 43988
rect 23711 43948 23756 43976
rect 23293 43939 23351 43945
rect 23750 43936 23756 43948
rect 23808 43936 23814 43988
rect 25038 43936 25044 43988
rect 25096 43976 25102 43988
rect 25777 43979 25835 43985
rect 25777 43976 25789 43979
rect 25096 43948 25789 43976
rect 25096 43936 25102 43948
rect 25777 43945 25789 43948
rect 25823 43945 25835 43979
rect 25777 43939 25835 43945
rect 26513 43979 26571 43985
rect 26513 43945 26525 43979
rect 26559 43976 26571 43979
rect 26694 43976 26700 43988
rect 26559 43948 26700 43976
rect 26559 43945 26571 43948
rect 26513 43939 26571 43945
rect 26694 43936 26700 43948
rect 26752 43936 26758 43988
rect 27338 43936 27344 43988
rect 27396 43976 27402 43988
rect 27525 43979 27583 43985
rect 27525 43976 27537 43979
rect 27396 43948 27537 43976
rect 27396 43936 27402 43948
rect 27525 43945 27537 43948
rect 27571 43945 27583 43979
rect 27525 43939 27583 43945
rect 29178 43936 29184 43988
rect 29236 43976 29242 43988
rect 30193 43979 30251 43985
rect 30193 43976 30205 43979
rect 29236 43948 30205 43976
rect 29236 43936 29242 43948
rect 30193 43945 30205 43948
rect 30239 43945 30251 43979
rect 30193 43939 30251 43945
rect 30837 43979 30895 43985
rect 30837 43945 30849 43979
rect 30883 43976 30895 43979
rect 31570 43976 31576 43988
rect 30883 43948 31576 43976
rect 30883 43945 30895 43948
rect 30837 43939 30895 43945
rect 31570 43936 31576 43948
rect 31628 43936 31634 43988
rect 32217 43979 32275 43985
rect 32217 43945 32229 43979
rect 32263 43976 32275 43979
rect 32582 43976 32588 43988
rect 32263 43948 32588 43976
rect 32263 43945 32275 43948
rect 32217 43939 32275 43945
rect 32582 43936 32588 43948
rect 32640 43936 32646 43988
rect 33597 43979 33655 43985
rect 33597 43945 33609 43979
rect 33643 43976 33655 43979
rect 34054 43976 34060 43988
rect 33643 43948 34060 43976
rect 33643 43945 33655 43948
rect 33597 43939 33655 43945
rect 34054 43936 34060 43948
rect 34112 43936 34118 43988
rect 35434 43936 35440 43988
rect 35492 43976 35498 43988
rect 35529 43979 35587 43985
rect 35529 43976 35541 43979
rect 35492 43948 35541 43976
rect 35492 43936 35498 43948
rect 35529 43945 35541 43948
rect 35575 43945 35587 43979
rect 35710 43976 35716 43988
rect 35671 43948 35716 43976
rect 35529 43939 35587 43945
rect 35710 43936 35716 43948
rect 35768 43936 35774 43988
rect 35894 43936 35900 43988
rect 35952 43976 35958 43988
rect 36173 43979 36231 43985
rect 36173 43976 36185 43979
rect 35952 43948 36185 43976
rect 35952 43936 35958 43948
rect 36173 43945 36185 43948
rect 36219 43945 36231 43979
rect 36173 43939 36231 43945
rect 36630 43936 36636 43988
rect 36688 43976 36694 43988
rect 36817 43979 36875 43985
rect 36817 43976 36829 43979
rect 36688 43948 36829 43976
rect 36688 43936 36694 43948
rect 36817 43945 36829 43948
rect 36863 43945 36875 43979
rect 36817 43939 36875 43945
rect 20898 43868 20904 43920
rect 20956 43908 20962 43920
rect 21545 43911 21603 43917
rect 21545 43908 21557 43911
rect 20956 43880 21557 43908
rect 20956 43868 20962 43880
rect 21545 43877 21557 43880
rect 21591 43877 21603 43911
rect 21545 43871 21603 43877
rect 29825 43911 29883 43917
rect 29825 43877 29837 43911
rect 29871 43908 29883 43911
rect 29914 43908 29920 43920
rect 29871 43880 29920 43908
rect 29871 43877 29883 43880
rect 29825 43871 29883 43877
rect 29914 43868 29920 43880
rect 29972 43868 29978 43920
rect 30558 43868 30564 43920
rect 30616 43908 30622 43920
rect 31297 43911 31355 43917
rect 31297 43908 31309 43911
rect 30616 43880 31309 43908
rect 30616 43868 30622 43880
rect 31297 43877 31309 43880
rect 31343 43877 31355 43911
rect 31297 43871 31355 43877
rect 24486 43840 24492 43852
rect 23124 43812 24492 43840
rect 21726 43772 21732 43784
rect 21687 43744 21732 43772
rect 21726 43732 21732 43744
rect 21784 43732 21790 43784
rect 22370 43772 22376 43784
rect 22331 43744 22376 43772
rect 22370 43732 22376 43744
rect 22428 43732 22434 43784
rect 23124 43781 23152 43812
rect 24486 43800 24492 43812
rect 24544 43800 24550 43852
rect 25041 43843 25099 43849
rect 25041 43809 25053 43843
rect 25087 43840 25099 43843
rect 25130 43840 25136 43852
rect 25087 43812 25136 43840
rect 25087 43809 25099 43812
rect 25041 43803 25099 43809
rect 25130 43800 25136 43812
rect 25188 43800 25194 43852
rect 25317 43843 25375 43849
rect 25317 43809 25329 43843
rect 25363 43840 25375 43843
rect 25590 43840 25596 43852
rect 25363 43812 25596 43840
rect 25363 43809 25375 43812
rect 25317 43803 25375 43809
rect 25590 43800 25596 43812
rect 25648 43800 25654 43852
rect 26602 43800 26608 43852
rect 26660 43840 26666 43852
rect 26697 43843 26755 43849
rect 26697 43840 26709 43843
rect 26660 43812 26709 43840
rect 26660 43800 26666 43812
rect 26697 43809 26709 43812
rect 26743 43809 26755 43843
rect 27893 43843 27951 43849
rect 27893 43840 27905 43843
rect 26697 43803 26755 43809
rect 26804 43812 27905 43840
rect 23109 43775 23167 43781
rect 23109 43741 23121 43775
rect 23155 43741 23167 43775
rect 23109 43735 23167 43741
rect 23293 43775 23351 43781
rect 23293 43741 23305 43775
rect 23339 43741 23351 43775
rect 23293 43735 23351 43741
rect 23753 43775 23811 43781
rect 23753 43741 23765 43775
rect 23799 43772 23811 43775
rect 23934 43772 23940 43784
rect 23799 43744 23940 43772
rect 23799 43741 23811 43744
rect 23753 43735 23811 43741
rect 19889 43707 19947 43713
rect 19889 43673 19901 43707
rect 19935 43704 19947 43707
rect 20714 43704 20720 43716
rect 19935 43676 20720 43704
rect 19935 43673 19947 43676
rect 19889 43667 19947 43673
rect 20714 43664 20720 43676
rect 20772 43704 20778 43716
rect 20772 43676 21128 43704
rect 20772 43664 20778 43676
rect 21100 43645 21128 43676
rect 23014 43664 23020 43716
rect 23072 43704 23078 43716
rect 23308 43704 23336 43735
rect 23934 43732 23940 43744
rect 23992 43732 23998 43784
rect 24029 43775 24087 43781
rect 24029 43741 24041 43775
rect 24075 43741 24087 43775
rect 24029 43735 24087 43741
rect 23072 43676 23336 43704
rect 24044 43704 24072 43735
rect 24762 43732 24768 43784
rect 24820 43772 24826 43784
rect 26804 43781 26832 43812
rect 27893 43809 27905 43812
rect 27939 43809 27951 43843
rect 27893 43803 27951 43809
rect 28997 43843 29055 43849
rect 28997 43809 29009 43843
rect 29043 43840 29055 43843
rect 29454 43840 29460 43852
rect 29043 43812 29460 43840
rect 29043 43809 29055 43812
rect 28997 43803 29055 43809
rect 29454 43800 29460 43812
rect 29512 43840 29518 43852
rect 29733 43843 29791 43849
rect 29733 43840 29745 43843
rect 29512 43812 29745 43840
rect 29512 43800 29518 43812
rect 29733 43809 29745 43812
rect 29779 43809 29791 43843
rect 29733 43803 29791 43809
rect 32674 43800 32680 43852
rect 32732 43840 32738 43852
rect 34057 43843 34115 43849
rect 34057 43840 34069 43843
rect 32732 43812 34069 43840
rect 32732 43800 32738 43812
rect 34057 43809 34069 43812
rect 34103 43809 34115 43843
rect 34057 43803 34115 43809
rect 24949 43775 25007 43781
rect 24949 43772 24961 43775
rect 24820 43744 24961 43772
rect 24820 43732 24826 43744
rect 24949 43741 24961 43744
rect 24995 43741 25007 43775
rect 24949 43735 25007 43741
rect 26789 43775 26847 43781
rect 26789 43741 26801 43775
rect 26835 43741 26847 43775
rect 26789 43735 26847 43741
rect 26878 43732 26884 43784
rect 26936 43772 26942 43784
rect 27433 43775 27491 43781
rect 27433 43772 27445 43775
rect 26936 43744 27445 43772
rect 26936 43732 26942 43744
rect 27433 43741 27445 43744
rect 27479 43741 27491 43775
rect 28810 43772 28816 43784
rect 28771 43744 28816 43772
rect 27433 43735 27491 43741
rect 28810 43732 28816 43744
rect 28868 43732 28874 43784
rect 30006 43772 30012 43784
rect 29967 43744 30012 43772
rect 30006 43732 30012 43744
rect 30064 43732 30070 43784
rect 32490 43732 32496 43784
rect 32548 43772 32554 43784
rect 32585 43775 32643 43781
rect 32585 43772 32597 43775
rect 32548 43744 32597 43772
rect 32548 43732 32554 43744
rect 32585 43741 32597 43744
rect 32631 43741 32643 43775
rect 32585 43735 32643 43741
rect 33321 43775 33379 43781
rect 33321 43741 33333 43775
rect 33367 43741 33379 43775
rect 33321 43735 33379 43741
rect 33413 43775 33471 43781
rect 33413 43741 33425 43775
rect 33459 43772 33471 43775
rect 33502 43772 33508 43784
rect 33459 43744 33508 43772
rect 33459 43741 33471 43744
rect 33413 43735 33471 43741
rect 25314 43704 25320 43716
rect 24044 43676 25320 43704
rect 23072 43664 23078 43676
rect 25314 43664 25320 43676
rect 25372 43664 25378 43716
rect 32401 43707 32459 43713
rect 32401 43673 32413 43707
rect 32447 43704 32459 43707
rect 32766 43704 32772 43716
rect 32447 43676 32772 43704
rect 32447 43673 32459 43676
rect 32401 43667 32459 43673
rect 32766 43664 32772 43676
rect 32824 43664 32830 43716
rect 33336 43704 33364 43735
rect 33502 43732 33508 43744
rect 33560 43732 33566 43784
rect 33597 43775 33655 43781
rect 33597 43741 33609 43775
rect 33643 43772 33655 43775
rect 33686 43772 33692 43784
rect 33643 43744 33692 43772
rect 33643 43741 33655 43744
rect 33597 43735 33655 43741
rect 33686 43732 33692 43744
rect 33744 43732 33750 43784
rect 34698 43704 34704 43716
rect 33336 43676 34704 43704
rect 34698 43664 34704 43676
rect 34756 43664 34762 43716
rect 35345 43707 35403 43713
rect 35345 43673 35357 43707
rect 35391 43704 35403 43707
rect 35434 43704 35440 43716
rect 35391 43676 35440 43704
rect 35391 43673 35403 43676
rect 35345 43667 35403 43673
rect 35434 43664 35440 43676
rect 35492 43664 35498 43716
rect 35561 43707 35619 43713
rect 35561 43673 35573 43707
rect 35607 43704 35619 43707
rect 35802 43704 35808 43716
rect 35607 43676 35808 43704
rect 35607 43673 35619 43676
rect 35561 43667 35619 43673
rect 35802 43664 35808 43676
rect 35860 43664 35866 43716
rect 21085 43639 21143 43645
rect 21085 43605 21097 43639
rect 21131 43636 21143 43639
rect 21910 43636 21916 43648
rect 21131 43608 21916 43636
rect 21131 43605 21143 43608
rect 21085 43599 21143 43605
rect 21910 43596 21916 43608
rect 21968 43596 21974 43648
rect 23937 43639 23995 43645
rect 23937 43605 23949 43639
rect 23983 43636 23995 43639
rect 24854 43636 24860 43648
rect 23983 43608 24860 43636
rect 23983 43605 23995 43608
rect 23937 43599 23995 43605
rect 24854 43596 24860 43608
rect 24912 43596 24918 43648
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 20530 43392 20536 43444
rect 20588 43432 20594 43444
rect 21177 43435 21235 43441
rect 21177 43432 21189 43435
rect 20588 43404 21189 43432
rect 20588 43392 20594 43404
rect 21177 43401 21189 43404
rect 21223 43401 21235 43435
rect 21177 43395 21235 43401
rect 23566 43392 23572 43444
rect 23624 43432 23630 43444
rect 23845 43435 23903 43441
rect 23845 43432 23857 43435
rect 23624 43404 23857 43432
rect 23624 43392 23630 43404
rect 23845 43401 23857 43404
rect 23891 43401 23903 43435
rect 23845 43395 23903 43401
rect 24489 43435 24547 43441
rect 24489 43401 24501 43435
rect 24535 43432 24547 43435
rect 24854 43432 24860 43444
rect 24535 43404 24860 43432
rect 24535 43401 24547 43404
rect 24489 43395 24547 43401
rect 24854 43392 24860 43404
rect 24912 43392 24918 43444
rect 25590 43432 25596 43444
rect 25551 43404 25596 43432
rect 25590 43392 25596 43404
rect 25648 43392 25654 43444
rect 27417 43435 27475 43441
rect 27417 43401 27429 43435
rect 27463 43432 27475 43435
rect 27522 43432 27528 43444
rect 27463 43404 27528 43432
rect 27463 43401 27475 43404
rect 27417 43395 27475 43401
rect 27522 43392 27528 43404
rect 27580 43392 27586 43444
rect 28166 43432 28172 43444
rect 28127 43404 28172 43432
rect 28166 43392 28172 43404
rect 28224 43392 28230 43444
rect 33778 43432 33784 43444
rect 33739 43404 33784 43432
rect 33778 43392 33784 43404
rect 33836 43392 33842 43444
rect 35069 43435 35127 43441
rect 35069 43401 35081 43435
rect 35115 43432 35127 43435
rect 35434 43432 35440 43444
rect 35115 43404 35440 43432
rect 35115 43401 35127 43404
rect 35069 43395 35127 43401
rect 35434 43392 35440 43404
rect 35492 43392 35498 43444
rect 24673 43367 24731 43373
rect 24673 43333 24685 43367
rect 24719 43364 24731 43367
rect 24762 43364 24768 43376
rect 24719 43336 24768 43364
rect 24719 43333 24731 43336
rect 24673 43327 24731 43333
rect 24762 43324 24768 43336
rect 24820 43324 24826 43376
rect 27614 43364 27620 43376
rect 27575 43336 27620 43364
rect 27614 43324 27620 43336
rect 27672 43324 27678 43376
rect 30098 43364 30104 43376
rect 28276 43336 30104 43364
rect 22462 43296 22468 43308
rect 22423 43268 22468 43296
rect 22462 43256 22468 43268
rect 22520 43256 22526 43308
rect 23293 43299 23351 43305
rect 23293 43265 23305 43299
rect 23339 43296 23351 43299
rect 23382 43296 23388 43308
rect 23339 43268 23388 43296
rect 23339 43265 23351 43268
rect 23293 43259 23351 43265
rect 23382 43256 23388 43268
rect 23440 43256 23446 43308
rect 23753 43299 23811 43305
rect 23753 43265 23765 43299
rect 23799 43296 23811 43299
rect 23842 43296 23848 43308
rect 23799 43268 23848 43296
rect 23799 43265 23811 43268
rect 23753 43259 23811 43265
rect 23842 43256 23848 43268
rect 23900 43256 23906 43308
rect 23937 43299 23995 43305
rect 23937 43265 23949 43299
rect 23983 43296 23995 43299
rect 24026 43296 24032 43308
rect 23983 43268 24032 43296
rect 23983 43265 23995 43268
rect 23937 43259 23995 43265
rect 24026 43256 24032 43268
rect 24084 43256 24090 43308
rect 24857 43299 24915 43305
rect 24857 43265 24869 43299
rect 24903 43296 24915 43299
rect 25130 43296 25136 43308
rect 24903 43268 25136 43296
rect 24903 43265 24915 43268
rect 24857 43259 24915 43265
rect 25130 43256 25136 43268
rect 25188 43256 25194 43308
rect 25314 43256 25320 43308
rect 25372 43296 25378 43308
rect 25501 43299 25559 43305
rect 25501 43296 25513 43299
rect 25372 43268 25513 43296
rect 25372 43256 25378 43268
rect 25501 43265 25513 43268
rect 25547 43265 25559 43299
rect 25774 43296 25780 43308
rect 25687 43268 25780 43296
rect 25501 43259 25559 43265
rect 25774 43256 25780 43268
rect 25832 43296 25838 43308
rect 26329 43299 26387 43305
rect 26329 43296 26341 43299
rect 25832 43268 26341 43296
rect 25832 43256 25838 43268
rect 26329 43265 26341 43268
rect 26375 43296 26387 43299
rect 26786 43296 26792 43308
rect 26375 43268 26792 43296
rect 26375 43265 26387 43268
rect 26329 43259 26387 43265
rect 26786 43256 26792 43268
rect 26844 43296 26850 43308
rect 28276 43305 28304 43336
rect 30098 43324 30104 43336
rect 30156 43324 30162 43376
rect 28261 43299 28319 43305
rect 28261 43296 28273 43299
rect 26844 43268 28273 43296
rect 26844 43256 26850 43268
rect 28261 43265 28273 43268
rect 28307 43265 28319 43299
rect 28261 43259 28319 43265
rect 28994 43256 29000 43308
rect 29052 43296 29058 43308
rect 29365 43299 29423 43305
rect 29365 43296 29377 43299
rect 29052 43268 29377 43296
rect 29052 43256 29058 43268
rect 29365 43265 29377 43268
rect 29411 43265 29423 43299
rect 29365 43259 29423 43265
rect 29638 43256 29644 43308
rect 29696 43296 29702 43308
rect 30009 43299 30067 43305
rect 30009 43296 30021 43299
rect 29696 43268 30021 43296
rect 29696 43256 29702 43268
rect 30009 43265 30021 43268
rect 30055 43265 30067 43299
rect 31294 43296 31300 43308
rect 31255 43268 31300 43296
rect 30009 43259 30067 43265
rect 31294 43256 31300 43268
rect 31352 43256 31358 43308
rect 32398 43256 32404 43308
rect 32456 43296 32462 43308
rect 32953 43299 33011 43305
rect 32953 43296 32965 43299
rect 32456 43268 32965 43296
rect 32456 43256 32462 43268
rect 32953 43265 32965 43268
rect 32999 43265 33011 43299
rect 32953 43259 33011 43265
rect 33134 43256 33140 43308
rect 33192 43296 33198 43308
rect 33597 43299 33655 43305
rect 33597 43296 33609 43299
rect 33192 43268 33609 43296
rect 33192 43256 33198 43268
rect 33597 43265 33609 43268
rect 33643 43265 33655 43299
rect 33597 43259 33655 43265
rect 34514 43256 34520 43308
rect 34572 43296 34578 43308
rect 34885 43299 34943 43305
rect 34885 43296 34897 43299
rect 34572 43268 34897 43296
rect 34572 43256 34578 43268
rect 34885 43265 34897 43268
rect 34931 43296 34943 43299
rect 35529 43299 35587 43305
rect 35529 43296 35541 43299
rect 34931 43268 35541 43296
rect 34931 43265 34943 43268
rect 34885 43259 34943 43265
rect 35529 43265 35541 43268
rect 35575 43265 35587 43299
rect 35529 43259 35587 43265
rect 27890 43188 27896 43240
rect 27948 43228 27954 43240
rect 28721 43231 28779 43237
rect 28721 43228 28733 43231
rect 27948 43200 28733 43228
rect 27948 43188 27954 43200
rect 28721 43197 28733 43200
rect 28767 43197 28779 43231
rect 28721 43191 28779 43197
rect 31662 43188 31668 43240
rect 31720 43228 31726 43240
rect 32309 43231 32367 43237
rect 32309 43228 32321 43231
rect 31720 43200 32321 43228
rect 31720 43188 31726 43200
rect 32309 43197 32321 43200
rect 32355 43197 32367 43231
rect 32309 43191 32367 43197
rect 33318 43188 33324 43240
rect 33376 43228 33382 43240
rect 34241 43231 34299 43237
rect 34241 43228 34253 43231
rect 33376 43200 34253 43228
rect 33376 43188 33382 43200
rect 34241 43197 34253 43200
rect 34287 43197 34299 43231
rect 34241 43191 34299 43197
rect 25498 43120 25504 43172
rect 25556 43160 25562 43172
rect 25777 43163 25835 43169
rect 25777 43160 25789 43163
rect 25556 43132 25789 43160
rect 25556 43120 25562 43132
rect 25777 43129 25789 43132
rect 25823 43129 25835 43163
rect 25777 43123 25835 43129
rect 27249 43163 27307 43169
rect 27249 43129 27261 43163
rect 27295 43160 27307 43163
rect 27338 43160 27344 43172
rect 27295 43132 27344 43160
rect 27295 43129 27307 43132
rect 27249 43123 27307 43129
rect 27338 43120 27344 43132
rect 27396 43120 27402 43172
rect 27430 43092 27436 43104
rect 27391 43064 27436 43092
rect 27430 43052 27436 43064
rect 27488 43052 27494 43104
rect 30650 43092 30656 43104
rect 30611 43064 30656 43092
rect 30650 43052 30656 43064
rect 30708 43052 30714 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 24946 42848 24952 42900
rect 25004 42888 25010 42900
rect 25317 42891 25375 42897
rect 25317 42888 25329 42891
rect 25004 42860 25329 42888
rect 25004 42848 25010 42860
rect 25317 42857 25329 42860
rect 25363 42888 25375 42891
rect 26145 42891 26203 42897
rect 26145 42888 26157 42891
rect 25363 42860 26157 42888
rect 25363 42857 25375 42860
rect 25317 42851 25375 42857
rect 26145 42857 26157 42860
rect 26191 42857 26203 42891
rect 26786 42888 26792 42900
rect 26747 42860 26792 42888
rect 26145 42851 26203 42857
rect 22646 42712 22652 42764
rect 22704 42752 22710 42764
rect 22833 42755 22891 42761
rect 22833 42752 22845 42755
rect 22704 42724 22845 42752
rect 22704 42712 22710 42724
rect 22833 42721 22845 42724
rect 22879 42721 22891 42755
rect 24670 42752 24676 42764
rect 24631 42724 24676 42752
rect 22833 42715 22891 42721
rect 24670 42712 24676 42724
rect 24728 42712 24734 42764
rect 26160 42616 26188 42851
rect 26786 42848 26792 42860
rect 26844 42848 26850 42900
rect 27062 42848 27068 42900
rect 27120 42888 27126 42900
rect 27893 42891 27951 42897
rect 27893 42888 27905 42891
rect 27120 42860 27905 42888
rect 27120 42848 27126 42860
rect 27893 42857 27905 42860
rect 27939 42857 27951 42891
rect 27893 42851 27951 42857
rect 33134 42848 33140 42900
rect 33192 42888 33198 42900
rect 33413 42891 33471 42897
rect 33413 42888 33425 42891
rect 33192 42860 33425 42888
rect 33192 42848 33198 42860
rect 33413 42857 33425 42860
rect 33459 42857 33471 42891
rect 33413 42851 33471 42857
rect 30650 42820 30656 42832
rect 30300 42792 30656 42820
rect 27246 42752 27252 42764
rect 27207 42724 27252 42752
rect 27246 42712 27252 42724
rect 27304 42712 27310 42764
rect 28258 42712 28264 42764
rect 28316 42752 28322 42764
rect 28537 42755 28595 42761
rect 28537 42752 28549 42755
rect 28316 42724 28549 42752
rect 28316 42712 28322 42724
rect 28537 42721 28549 42724
rect 28583 42721 28595 42755
rect 30300 42752 30328 42792
rect 30650 42780 30656 42792
rect 30708 42780 30714 42832
rect 32214 42752 32220 42764
rect 28537 42715 28595 42721
rect 29748 42724 30328 42752
rect 32175 42724 32220 42752
rect 27706 42644 27712 42696
rect 27764 42684 27770 42696
rect 28077 42687 28135 42693
rect 28077 42684 28089 42687
rect 27764 42656 28089 42684
rect 27764 42644 27770 42656
rect 28077 42653 28089 42656
rect 28123 42653 28135 42687
rect 28077 42647 28135 42653
rect 27798 42616 27804 42628
rect 26160 42588 27804 42616
rect 27798 42576 27804 42588
rect 27856 42616 27862 42628
rect 29454 42616 29460 42628
rect 27856 42588 29460 42616
rect 27856 42576 27862 42588
rect 29454 42576 29460 42588
rect 29512 42616 29518 42628
rect 29748 42625 29776 42724
rect 32214 42712 32220 42724
rect 32272 42712 32278 42764
rect 30098 42644 30104 42696
rect 30156 42684 30162 42696
rect 30377 42687 30435 42693
rect 30377 42684 30389 42687
rect 30156 42656 30389 42684
rect 30156 42644 30162 42656
rect 30377 42653 30389 42656
rect 30423 42653 30435 42687
rect 30377 42647 30435 42653
rect 29733 42619 29791 42625
rect 29733 42616 29745 42619
rect 29512 42588 29745 42616
rect 29512 42576 29518 42588
rect 29733 42585 29745 42588
rect 29779 42585 29791 42619
rect 29733 42579 29791 42585
rect 21910 42548 21916 42560
rect 21871 42520 21916 42548
rect 21910 42508 21916 42520
rect 21968 42508 21974 42560
rect 23477 42551 23535 42557
rect 23477 42517 23489 42551
rect 23523 42548 23535 42551
rect 24026 42548 24032 42560
rect 23523 42520 24032 42548
rect 23523 42517 23535 42520
rect 23477 42511 23535 42517
rect 24026 42508 24032 42520
rect 24084 42508 24090 42560
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 24026 42304 24032 42356
rect 24084 42344 24090 42356
rect 24765 42347 24823 42353
rect 24765 42344 24777 42347
rect 24084 42316 24777 42344
rect 24084 42304 24090 42316
rect 24765 42313 24777 42316
rect 24811 42344 24823 42347
rect 25774 42344 25780 42356
rect 24811 42316 25780 42344
rect 24811 42313 24823 42316
rect 24765 42307 24823 42313
rect 25774 42304 25780 42316
rect 25832 42304 25838 42356
rect 27154 42344 27160 42356
rect 27115 42316 27160 42344
rect 27154 42304 27160 42316
rect 27212 42304 27218 42356
rect 27706 42344 27712 42356
rect 27667 42316 27712 42344
rect 27706 42304 27712 42316
rect 27764 42304 27770 42356
rect 28810 42304 28816 42356
rect 28868 42344 28874 42356
rect 28997 42347 29055 42353
rect 28997 42344 29009 42347
rect 28868 42316 29009 42344
rect 28868 42304 28874 42316
rect 28997 42313 29009 42316
rect 29043 42313 29055 42347
rect 29454 42344 29460 42356
rect 29415 42316 29460 42344
rect 28997 42307 29055 42313
rect 29454 42304 29460 42316
rect 29512 42304 29518 42356
rect 28445 42279 28503 42285
rect 28445 42245 28457 42279
rect 28491 42276 28503 42279
rect 30098 42276 30104 42288
rect 28491 42248 30104 42276
rect 28491 42245 28503 42248
rect 28445 42239 28503 42245
rect 30098 42236 30104 42248
rect 30156 42236 30162 42288
rect 23753 42075 23811 42081
rect 23753 42072 23765 42075
rect 22066 42044 23765 42072
rect 21910 41964 21916 42016
rect 21968 42004 21974 42016
rect 22066 42004 22094 42044
rect 23753 42041 23765 42044
rect 23799 42072 23811 42075
rect 25130 42072 25136 42084
rect 23799 42044 25136 42072
rect 23799 42041 23811 42044
rect 23753 42035 23811 42041
rect 25130 42032 25136 42044
rect 25188 42032 25194 42084
rect 21968 41976 22094 42004
rect 21968 41964 21974 41976
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 27798 41800 27804 41812
rect 27759 41772 27804 41800
rect 27798 41760 27804 41772
rect 27856 41760 27862 41812
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 25130 7528 25136 7540
rect 25091 7500 25136 7528
rect 25130 7488 25136 7500
rect 25188 7488 25194 7540
rect 24489 7395 24547 7401
rect 24489 7361 24501 7395
rect 24535 7392 24547 7395
rect 25038 7392 25044 7404
rect 24535 7364 25044 7392
rect 24535 7361 24547 7364
rect 24489 7355 24547 7361
rect 25038 7352 25044 7364
rect 25096 7392 25102 7404
rect 26513 7395 26571 7401
rect 26513 7392 26525 7395
rect 25096 7364 26525 7392
rect 25096 7352 25102 7364
rect 26513 7361 26525 7364
rect 26559 7361 26571 7395
rect 26513 7355 26571 7361
rect 23106 7188 23112 7200
rect 23067 7160 23112 7188
rect 23106 7148 23112 7160
rect 23164 7148 23170 7200
rect 23750 7188 23756 7200
rect 23711 7160 23756 7188
rect 23750 7148 23756 7160
rect 23808 7148 23814 7200
rect 24578 7188 24584 7200
rect 24539 7160 24584 7188
rect 24578 7148 24584 7160
rect 24636 7148 24642 7200
rect 25590 7148 25596 7200
rect 25648 7188 25654 7200
rect 25685 7191 25743 7197
rect 25685 7188 25697 7191
rect 25648 7160 25697 7188
rect 25648 7148 25654 7160
rect 25685 7157 25697 7160
rect 25731 7157 25743 7191
rect 26418 7188 26424 7200
rect 26379 7160 26424 7188
rect 25685 7151 25743 7157
rect 26418 7148 26424 7160
rect 26476 7148 26482 7200
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 25038 6848 25044 6860
rect 23860 6820 25044 6848
rect 21174 6780 21180 6792
rect 21135 6752 21180 6780
rect 21174 6740 21180 6752
rect 21232 6740 21238 6792
rect 21266 6740 21272 6792
rect 21324 6780 21330 6792
rect 23860 6789 23888 6820
rect 25038 6808 25044 6820
rect 25096 6848 25102 6860
rect 25317 6851 25375 6857
rect 25317 6848 25329 6851
rect 25096 6820 25329 6848
rect 25096 6808 25102 6820
rect 25317 6817 25329 6820
rect 25363 6817 25375 6851
rect 25317 6811 25375 6817
rect 22281 6783 22339 6789
rect 22281 6780 22293 6783
rect 21324 6752 22293 6780
rect 21324 6740 21330 6752
rect 22281 6749 22293 6752
rect 22327 6780 22339 6783
rect 22925 6783 22983 6789
rect 22925 6780 22937 6783
rect 22327 6752 22937 6780
rect 22327 6749 22339 6752
rect 22281 6743 22339 6749
rect 22925 6749 22937 6752
rect 22971 6749 22983 6783
rect 22925 6743 22983 6749
rect 23845 6783 23903 6789
rect 23845 6749 23857 6783
rect 23891 6749 23903 6783
rect 25130 6780 25136 6792
rect 23845 6743 23903 6749
rect 24872 6752 25136 6780
rect 24872 6656 24900 6752
rect 25130 6740 25136 6752
rect 25188 6740 25194 6792
rect 26234 6740 26240 6792
rect 26292 6780 26298 6792
rect 26694 6780 26700 6792
rect 26292 6752 26337 6780
rect 26655 6752 26700 6780
rect 26292 6740 26298 6752
rect 26694 6740 26700 6752
rect 26752 6740 26758 6792
rect 27522 6740 27528 6792
rect 27580 6780 27586 6792
rect 27617 6783 27675 6789
rect 27617 6780 27629 6783
rect 27580 6752 27629 6780
rect 27580 6740 27586 6752
rect 27617 6749 27629 6752
rect 27663 6749 27675 6783
rect 27617 6743 27675 6749
rect 27798 6740 27804 6792
rect 27856 6780 27862 6792
rect 28445 6783 28503 6789
rect 28445 6780 28457 6783
rect 27856 6752 28457 6780
rect 27856 6740 27862 6752
rect 28445 6749 28457 6752
rect 28491 6749 28503 6783
rect 28445 6743 28503 6749
rect 22370 6644 22376 6656
rect 22331 6616 22376 6644
rect 22370 6604 22376 6616
rect 22428 6604 22434 6656
rect 23014 6644 23020 6656
rect 22975 6616 23020 6644
rect 23014 6604 23020 6616
rect 23072 6604 23078 6656
rect 23937 6647 23995 6653
rect 23937 6613 23949 6647
rect 23983 6644 23995 6647
rect 24486 6644 24492 6656
rect 23983 6616 24492 6644
rect 23983 6613 23995 6616
rect 23937 6607 23995 6613
rect 24486 6604 24492 6616
rect 24544 6604 24550 6656
rect 24673 6647 24731 6653
rect 24673 6613 24685 6647
rect 24719 6644 24731 6647
rect 24854 6644 24860 6656
rect 24719 6616 24860 6644
rect 24719 6613 24731 6616
rect 24673 6607 24731 6613
rect 24854 6604 24860 6616
rect 24912 6604 24918 6656
rect 27706 6604 27712 6656
rect 27764 6644 27770 6656
rect 28353 6647 28411 6653
rect 28353 6644 28365 6647
rect 27764 6616 28365 6644
rect 27764 6604 27770 6616
rect 28353 6613 28365 6616
rect 28399 6613 28411 6647
rect 28353 6607 28411 6613
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 24486 6372 24492 6384
rect 24447 6344 24492 6372
rect 24486 6332 24492 6344
rect 24544 6332 24550 6384
rect 27706 6372 27712 6384
rect 27667 6344 27712 6372
rect 27706 6332 27712 6344
rect 27764 6332 27770 6384
rect 21266 6304 21272 6316
rect 21227 6276 21272 6304
rect 21266 6264 21272 6276
rect 21324 6264 21330 6316
rect 27522 6304 27528 6316
rect 27483 6276 27528 6304
rect 27522 6264 27528 6276
rect 27580 6264 27586 6316
rect 21361 6239 21419 6245
rect 21361 6205 21373 6239
rect 21407 6236 21419 6239
rect 22278 6236 22284 6248
rect 21407 6208 22284 6236
rect 21407 6205 21419 6208
rect 21361 6199 21419 6205
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 23845 6239 23903 6245
rect 23845 6205 23857 6239
rect 23891 6236 23903 6239
rect 24305 6239 24363 6245
rect 24305 6236 24317 6239
rect 23891 6208 24317 6236
rect 23891 6205 23903 6208
rect 23845 6199 23903 6205
rect 24305 6205 24317 6208
rect 24351 6205 24363 6239
rect 24946 6236 24952 6248
rect 24907 6208 24952 6236
rect 24305 6199 24363 6205
rect 24946 6196 24952 6208
rect 25004 6196 25010 6248
rect 29178 6236 29184 6248
rect 29139 6208 29184 6236
rect 29178 6196 29184 6208
rect 29236 6196 29242 6248
rect 22094 6128 22100 6180
rect 22152 6168 22158 6180
rect 22925 6171 22983 6177
rect 22925 6168 22937 6171
rect 22152 6140 22937 6168
rect 22152 6128 22158 6140
rect 22925 6137 22937 6140
rect 22971 6137 22983 6171
rect 22925 6131 22983 6137
rect 18966 6100 18972 6112
rect 18927 6072 18972 6100
rect 18966 6060 18972 6072
rect 19024 6060 19030 6112
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 19521 6103 19579 6109
rect 19521 6100 19533 6103
rect 19392 6072 19533 6100
rect 19392 6060 19398 6072
rect 19521 6069 19533 6072
rect 19567 6069 19579 6103
rect 20254 6100 20260 6112
rect 20215 6072 20260 6100
rect 19521 6063 19579 6069
rect 20254 6060 20260 6072
rect 20312 6060 20318 6112
rect 22186 6060 22192 6112
rect 22244 6100 22250 6112
rect 22281 6103 22339 6109
rect 22281 6100 22293 6103
rect 22244 6072 22293 6100
rect 22244 6060 22250 6072
rect 22281 6069 22293 6072
rect 22327 6069 22339 6103
rect 22281 6063 22339 6069
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 21266 5788 21272 5840
rect 21324 5828 21330 5840
rect 21324 5800 21496 5828
rect 21324 5788 21330 5800
rect 20162 5760 20168 5772
rect 19996 5732 20168 5760
rect 18598 5652 18604 5704
rect 18656 5692 18662 5704
rect 19996 5701 20024 5732
rect 20162 5720 20168 5732
rect 20220 5760 20226 5772
rect 21468 5769 21496 5800
rect 25038 5788 25044 5840
rect 25096 5828 25102 5840
rect 25096 5800 28120 5828
rect 25096 5788 25102 5800
rect 21453 5763 21511 5769
rect 21453 5760 21465 5763
rect 20220 5732 21465 5760
rect 20220 5720 20226 5732
rect 21453 5729 21465 5732
rect 21499 5729 21511 5763
rect 22186 5760 22192 5772
rect 22147 5732 22192 5760
rect 21453 5723 21511 5729
rect 22186 5720 22192 5732
rect 22244 5720 22250 5772
rect 22370 5760 22376 5772
rect 22331 5732 22376 5760
rect 22370 5720 22376 5732
rect 22428 5720 22434 5772
rect 22922 5760 22928 5772
rect 22883 5732 22928 5760
rect 22922 5720 22928 5732
rect 22980 5720 22986 5772
rect 26234 5720 26240 5772
rect 26292 5760 26298 5772
rect 27617 5763 27675 5769
rect 27617 5760 27629 5763
rect 26292 5732 27629 5760
rect 26292 5720 26298 5732
rect 27617 5729 27629 5732
rect 27663 5729 27675 5763
rect 27617 5723 27675 5729
rect 18693 5695 18751 5701
rect 18693 5692 18705 5695
rect 18656 5664 18705 5692
rect 18656 5652 18662 5664
rect 18693 5661 18705 5664
rect 18739 5661 18751 5695
rect 18693 5655 18751 5661
rect 19981 5695 20039 5701
rect 19981 5661 19993 5695
rect 20027 5661 20039 5695
rect 20806 5692 20812 5704
rect 20767 5664 20812 5692
rect 19981 5655 20039 5661
rect 20806 5652 20812 5664
rect 20864 5652 20870 5704
rect 21269 5695 21327 5701
rect 21269 5661 21281 5695
rect 21315 5692 21327 5695
rect 24854 5692 24860 5704
rect 21315 5664 22232 5692
rect 24767 5664 24860 5692
rect 21315 5661 21327 5664
rect 21269 5655 21327 5661
rect 21284 5624 21312 5655
rect 19444 5596 21312 5624
rect 22204 5624 22232 5664
rect 24854 5652 24860 5664
rect 24912 5652 24918 5704
rect 28092 5701 28120 5800
rect 28077 5695 28135 5701
rect 28077 5661 28089 5695
rect 28123 5661 28135 5695
rect 28077 5655 28135 5661
rect 28905 5695 28963 5701
rect 28905 5661 28917 5695
rect 28951 5692 28963 5695
rect 28994 5692 29000 5704
rect 28951 5664 29000 5692
rect 28951 5661 28963 5664
rect 28905 5655 28963 5661
rect 28994 5652 29000 5664
rect 29052 5652 29058 5704
rect 29917 5695 29975 5701
rect 29917 5692 29929 5695
rect 29564 5664 29929 5692
rect 24872 5624 24900 5652
rect 25130 5624 25136 5636
rect 22204 5596 24900 5624
rect 25091 5596 25136 5624
rect 18966 5516 18972 5568
rect 19024 5556 19030 5568
rect 19444 5565 19472 5596
rect 25130 5584 25136 5596
rect 25188 5584 25194 5636
rect 25777 5627 25835 5633
rect 25777 5593 25789 5627
rect 25823 5624 25835 5627
rect 26602 5624 26608 5636
rect 25823 5596 26608 5624
rect 25823 5593 25835 5596
rect 25777 5587 25835 5593
rect 26602 5584 26608 5596
rect 26660 5584 26666 5636
rect 27433 5627 27491 5633
rect 27433 5593 27445 5627
rect 27479 5624 27491 5627
rect 28169 5627 28227 5633
rect 28169 5624 28181 5627
rect 27479 5596 28181 5624
rect 27479 5593 27491 5596
rect 27433 5587 27491 5593
rect 28169 5593 28181 5596
rect 28215 5593 28227 5627
rect 28169 5587 28227 5593
rect 19429 5559 19487 5565
rect 19429 5556 19441 5559
rect 19024 5528 19441 5556
rect 19024 5516 19030 5528
rect 19429 5525 19441 5528
rect 19475 5525 19487 5559
rect 19429 5519 19487 5525
rect 20073 5559 20131 5565
rect 20073 5525 20085 5559
rect 20119 5556 20131 5559
rect 21726 5556 21732 5568
rect 20119 5528 21732 5556
rect 20119 5525 20131 5528
rect 20073 5519 20131 5525
rect 21726 5516 21732 5528
rect 21784 5516 21790 5568
rect 27798 5516 27804 5568
rect 27856 5556 27862 5568
rect 29564 5556 29592 5664
rect 29917 5661 29929 5664
rect 29963 5661 29975 5695
rect 29917 5655 29975 5661
rect 27856 5528 29592 5556
rect 27856 5516 27862 5528
rect 29638 5516 29644 5568
rect 29696 5556 29702 5568
rect 29825 5559 29883 5565
rect 29825 5556 29837 5559
rect 29696 5528 29837 5556
rect 29696 5516 29702 5528
rect 29825 5525 29837 5528
rect 29871 5525 29883 5559
rect 29825 5519 29883 5525
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 21174 5284 21180 5296
rect 19628 5256 21180 5284
rect 18966 5216 18972 5228
rect 18927 5188 18972 5216
rect 18966 5176 18972 5188
rect 19024 5176 19030 5228
rect 19628 5225 19656 5256
rect 21174 5244 21180 5256
rect 21232 5244 21238 5296
rect 22281 5287 22339 5293
rect 22281 5253 22293 5287
rect 22327 5284 22339 5287
rect 23014 5284 23020 5296
rect 22327 5256 23020 5284
rect 22327 5253 22339 5256
rect 22281 5247 22339 5253
rect 23014 5244 23020 5256
rect 23072 5244 23078 5296
rect 24578 5284 24584 5296
rect 24539 5256 24584 5284
rect 24578 5244 24584 5256
rect 24636 5244 24642 5296
rect 29638 5284 29644 5296
rect 29599 5256 29644 5284
rect 29638 5244 29644 5256
rect 29696 5244 29702 5296
rect 19613 5219 19671 5225
rect 19613 5185 19625 5219
rect 19659 5185 19671 5219
rect 22094 5216 22100 5228
rect 22055 5188 22100 5216
rect 19613 5179 19671 5185
rect 22094 5176 22100 5188
rect 22152 5176 22158 5228
rect 28994 5176 29000 5228
rect 29052 5216 29058 5228
rect 29052 5188 29097 5216
rect 29052 5176 29058 5188
rect 17954 5108 17960 5160
rect 18012 5148 18018 5160
rect 19797 5151 19855 5157
rect 19797 5148 19809 5151
rect 18012 5120 19809 5148
rect 18012 5108 18018 5120
rect 19797 5117 19809 5120
rect 19843 5117 19855 5151
rect 21358 5148 21364 5160
rect 21319 5120 21364 5148
rect 19797 5111 19855 5117
rect 21358 5108 21364 5120
rect 21416 5108 21422 5160
rect 23474 5148 23480 5160
rect 23435 5120 23480 5148
rect 23474 5108 23480 5120
rect 23532 5108 23538 5160
rect 24026 5108 24032 5160
rect 24084 5148 24090 5160
rect 24397 5151 24455 5157
rect 24397 5148 24409 5151
rect 24084 5120 24409 5148
rect 24084 5108 24090 5120
rect 24397 5117 24409 5120
rect 24443 5117 24455 5151
rect 25222 5148 25228 5160
rect 25183 5120 25228 5148
rect 24397 5111 24455 5117
rect 25222 5108 25228 5120
rect 25280 5108 25286 5160
rect 27801 5151 27859 5157
rect 27801 5148 27813 5151
rect 27724 5120 27813 5148
rect 27724 5092 27752 5120
rect 27801 5117 27813 5120
rect 27847 5117 27859 5151
rect 27801 5111 27859 5117
rect 27982 5108 27988 5160
rect 28040 5148 28046 5160
rect 28813 5151 28871 5157
rect 28813 5148 28825 5151
rect 28040 5120 28825 5148
rect 28040 5108 28046 5120
rect 28813 5117 28825 5120
rect 28859 5117 28871 5151
rect 28813 5111 28871 5117
rect 29457 5151 29515 5157
rect 29457 5117 29469 5151
rect 29503 5148 29515 5151
rect 29730 5148 29736 5160
rect 29503 5120 29736 5148
rect 29503 5117 29515 5120
rect 29457 5111 29515 5117
rect 29730 5108 29736 5120
rect 29788 5108 29794 5160
rect 30006 5148 30012 5160
rect 29967 5120 30012 5148
rect 30006 5108 30012 5120
rect 30064 5108 30070 5160
rect 18509 5083 18567 5089
rect 18509 5049 18521 5083
rect 18555 5080 18567 5083
rect 19978 5080 19984 5092
rect 18555 5052 19984 5080
rect 18555 5049 18567 5052
rect 18509 5043 18567 5049
rect 19978 5040 19984 5052
rect 20036 5040 20042 5092
rect 27706 5040 27712 5092
rect 27764 5040 27770 5092
rect 16942 4972 16948 5024
rect 17000 5012 17006 5024
rect 17037 5015 17095 5021
rect 17037 5012 17049 5015
rect 17000 4984 17049 5012
rect 17000 4972 17006 4984
rect 17037 4981 17049 4984
rect 17083 4981 17095 5015
rect 17037 4975 17095 4981
rect 17865 5015 17923 5021
rect 17865 4981 17877 5015
rect 17911 5012 17923 5015
rect 18322 5012 18328 5024
rect 17911 4984 18328 5012
rect 17911 4981 17923 4984
rect 17865 4975 17923 4981
rect 18322 4972 18328 4984
rect 18380 4972 18386 5024
rect 19061 5015 19119 5021
rect 19061 4981 19073 5015
rect 19107 5012 19119 5015
rect 20070 5012 20076 5024
rect 19107 4984 20076 5012
rect 19107 4981 19119 4984
rect 19061 4975 19119 4981
rect 20070 4972 20076 4984
rect 20128 4972 20134 5024
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 23106 4808 23112 4820
rect 22204 4780 23112 4808
rect 20254 4740 20260 4752
rect 19904 4712 20260 4740
rect 17589 4675 17647 4681
rect 17589 4641 17601 4675
rect 17635 4672 17647 4675
rect 19058 4672 19064 4684
rect 17635 4644 19064 4672
rect 17635 4641 17647 4644
rect 17589 4635 17647 4641
rect 19058 4632 19064 4644
rect 19116 4632 19122 4684
rect 19904 4681 19932 4712
rect 20254 4700 20260 4712
rect 20312 4700 20318 4752
rect 19889 4675 19947 4681
rect 19889 4641 19901 4675
rect 19935 4641 19947 4675
rect 20070 4672 20076 4684
rect 20031 4644 20076 4672
rect 19889 4635 19947 4641
rect 20070 4632 20076 4644
rect 20128 4632 20134 4684
rect 21082 4672 21088 4684
rect 21043 4644 21088 4672
rect 21082 4632 21088 4644
rect 21140 4632 21146 4684
rect 22204 4681 22232 4780
rect 23106 4768 23112 4780
rect 23164 4768 23170 4820
rect 27982 4808 27988 4820
rect 27943 4780 27988 4808
rect 27982 4768 27988 4780
rect 28040 4768 28046 4820
rect 29730 4808 29736 4820
rect 29691 4780 29736 4808
rect 29730 4768 29736 4780
rect 29788 4768 29794 4820
rect 22278 4700 22284 4752
rect 22336 4740 22342 4752
rect 22336 4712 22416 4740
rect 22336 4700 22342 4712
rect 22388 4681 22416 4712
rect 22189 4675 22247 4681
rect 22189 4641 22201 4675
rect 22235 4641 22247 4675
rect 22189 4635 22247 4641
rect 22373 4675 22431 4681
rect 22373 4641 22385 4675
rect 22419 4641 22431 4675
rect 23566 4672 23572 4684
rect 23527 4644 23572 4672
rect 22373 4635 22431 4641
rect 23566 4632 23572 4644
rect 23624 4632 23630 4684
rect 25038 4632 25044 4684
rect 25096 4632 25102 4684
rect 25590 4672 25596 4684
rect 25551 4644 25596 4672
rect 25590 4632 25596 4644
rect 25648 4632 25654 4684
rect 26326 4672 26332 4684
rect 26287 4644 26332 4672
rect 26326 4632 26332 4644
rect 26384 4632 26390 4684
rect 30561 4675 30619 4681
rect 30561 4641 30573 4675
rect 30607 4672 30619 4675
rect 31294 4672 31300 4684
rect 30607 4644 31300 4672
rect 30607 4641 30619 4644
rect 30561 4635 30619 4641
rect 31294 4632 31300 4644
rect 31352 4632 31358 4684
rect 15010 4564 15016 4616
rect 15068 4604 15074 4616
rect 15105 4607 15163 4613
rect 15105 4604 15117 4607
rect 15068 4576 15117 4604
rect 15068 4564 15074 4576
rect 15105 4573 15117 4576
rect 15151 4573 15163 4607
rect 15105 4567 15163 4573
rect 15838 4564 15844 4616
rect 15896 4604 15902 4616
rect 15933 4607 15991 4613
rect 15933 4604 15945 4607
rect 15896 4576 15945 4604
rect 15896 4564 15902 4576
rect 15933 4573 15945 4576
rect 15979 4573 15991 4607
rect 15933 4567 15991 4573
rect 16945 4607 17003 4613
rect 16945 4573 16957 4607
rect 16991 4604 17003 4607
rect 17402 4604 17408 4616
rect 16991 4576 17408 4604
rect 16991 4573 17003 4576
rect 16945 4567 17003 4573
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 18046 4604 18052 4616
rect 18007 4576 18052 4604
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 18877 4607 18935 4613
rect 18877 4573 18889 4607
rect 18923 4604 18935 4607
rect 19426 4604 19432 4616
rect 18923 4576 19432 4604
rect 18923 4573 18935 4576
rect 18877 4567 18935 4573
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 24854 4564 24860 4616
rect 24912 4604 24918 4616
rect 24949 4607 25007 4613
rect 24949 4604 24961 4607
rect 24912 4576 24961 4604
rect 24912 4564 24918 4576
rect 24949 4573 24961 4576
rect 24995 4604 25007 4607
rect 25056 4604 25084 4632
rect 24995 4576 25084 4604
rect 24995 4573 25007 4576
rect 24949 4567 25007 4573
rect 27798 4564 27804 4616
rect 27856 4604 27862 4616
rect 27893 4607 27951 4613
rect 27893 4604 27905 4607
rect 27856 4576 27905 4604
rect 27856 4564 27862 4576
rect 27893 4573 27905 4576
rect 27939 4573 27951 4607
rect 27893 4567 27951 4573
rect 28721 4607 28779 4613
rect 28721 4573 28733 4607
rect 28767 4604 28779 4607
rect 28994 4604 29000 4616
rect 28767 4576 29000 4604
rect 28767 4573 28779 4576
rect 28721 4567 28779 4573
rect 25041 4539 25099 4545
rect 25041 4505 25053 4539
rect 25087 4536 25099 4539
rect 25777 4539 25835 4545
rect 25777 4536 25789 4539
rect 25087 4508 25789 4536
rect 25087 4505 25099 4508
rect 25041 4499 25099 4505
rect 25777 4505 25789 4508
rect 25823 4505 25835 4539
rect 27908 4536 27936 4567
rect 28994 4564 29000 4576
rect 29052 4564 29058 4616
rect 31202 4604 31208 4616
rect 31163 4576 31208 4604
rect 31202 4564 31208 4576
rect 31260 4564 31266 4616
rect 31849 4607 31907 4613
rect 31849 4604 31861 4607
rect 31726 4576 31861 4604
rect 31726 4536 31754 4576
rect 31849 4573 31861 4576
rect 31895 4604 31907 4607
rect 32122 4604 32128 4616
rect 31895 4576 32128 4604
rect 31895 4573 31907 4576
rect 31849 4567 31907 4573
rect 32122 4564 32128 4576
rect 32180 4564 32186 4616
rect 32306 4604 32312 4616
rect 32267 4576 32312 4604
rect 32306 4564 32312 4576
rect 32364 4564 32370 4616
rect 27908 4508 31754 4536
rect 25777 4499 25835 4505
rect 31754 4428 31760 4480
rect 31812 4468 31818 4480
rect 31812 4440 31857 4468
rect 31812 4428 31818 4440
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 32122 4156 32128 4208
rect 32180 4196 32186 4208
rect 32180 4168 32536 4196
rect 32180 4156 32186 4168
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 17037 4131 17095 4137
rect 17037 4128 17049 4131
rect 16816 4100 17049 4128
rect 16816 4088 16822 4100
rect 17037 4097 17049 4100
rect 17083 4128 17095 4131
rect 17681 4131 17739 4137
rect 17681 4128 17693 4131
rect 17083 4100 17693 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 17681 4097 17693 4100
rect 17727 4128 17739 4131
rect 18325 4131 18383 4137
rect 18325 4128 18337 4131
rect 17727 4100 18337 4128
rect 17727 4097 17739 4100
rect 17681 4091 17739 4097
rect 18325 4097 18337 4100
rect 18371 4097 18383 4131
rect 18325 4091 18383 4097
rect 15657 4063 15715 4069
rect 15657 4029 15669 4063
rect 15703 4060 15715 4063
rect 17218 4060 17224 4072
rect 15703 4032 17224 4060
rect 15703 4029 15715 4032
rect 15657 4023 15715 4029
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 16301 3995 16359 4001
rect 16301 3961 16313 3995
rect 16347 3992 16359 3995
rect 17678 3992 17684 4004
rect 16347 3964 17684 3992
rect 16347 3961 16359 3964
rect 16301 3955 16359 3961
rect 17678 3952 17684 3964
rect 17736 3952 17742 4004
rect 18340 3992 18368 4091
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 19613 4131 19671 4137
rect 19613 4128 19625 4131
rect 19484 4100 19625 4128
rect 19484 4088 19490 4100
rect 19613 4097 19625 4100
rect 19659 4097 19671 4131
rect 19613 4091 19671 4097
rect 23661 4131 23719 4137
rect 23661 4097 23673 4131
rect 23707 4128 23719 4131
rect 24026 4128 24032 4140
rect 23707 4100 24032 4128
rect 23707 4097 23719 4100
rect 23661 4091 23719 4097
rect 24026 4088 24032 4100
rect 24084 4088 24090 4140
rect 28994 4088 29000 4140
rect 29052 4128 29058 4140
rect 29052 4100 29097 4128
rect 29052 4088 29058 4100
rect 31294 4088 31300 4140
rect 31352 4128 31358 4140
rect 31352 4100 31397 4128
rect 31352 4088 31358 4100
rect 31570 4088 31576 4140
rect 31628 4128 31634 4140
rect 32306 4128 32312 4140
rect 31628 4100 32312 4128
rect 31628 4088 31634 4100
rect 32306 4088 32312 4100
rect 32364 4088 32370 4140
rect 32508 4137 32536 4168
rect 32493 4131 32551 4137
rect 32493 4097 32505 4131
rect 32539 4097 32551 4131
rect 32493 4091 32551 4097
rect 18417 4063 18475 4069
rect 18417 4029 18429 4063
rect 18463 4060 18475 4063
rect 19797 4063 19855 4069
rect 19797 4060 19809 4063
rect 18463 4032 19809 4060
rect 18463 4029 18475 4032
rect 18417 4023 18475 4029
rect 19797 4029 19809 4032
rect 19843 4029 19855 4063
rect 19797 4023 19855 4029
rect 21453 4063 21511 4069
rect 21453 4029 21465 4063
rect 21499 4060 21511 4063
rect 22278 4060 22284 4072
rect 21499 4032 22284 4060
rect 21499 4029 21511 4032
rect 21453 4023 21511 4029
rect 22278 4020 22284 4032
rect 22336 4020 22342 4072
rect 22373 4063 22431 4069
rect 22373 4029 22385 4063
rect 22419 4060 22431 4063
rect 24121 4063 24179 4069
rect 24121 4060 24133 4063
rect 22419 4032 24133 4060
rect 22419 4029 22431 4032
rect 22373 4023 22431 4029
rect 24121 4029 24133 4032
rect 24167 4029 24179 4063
rect 24302 4060 24308 4072
rect 24263 4032 24308 4060
rect 24121 4023 24179 4029
rect 24302 4020 24308 4032
rect 24360 4020 24366 4072
rect 24670 4060 24676 4072
rect 24631 4032 24676 4060
rect 24670 4020 24676 4032
rect 24728 4020 24734 4072
rect 27430 4060 27436 4072
rect 27391 4032 27436 4060
rect 27430 4020 27436 4032
rect 27488 4020 27494 4072
rect 27890 4020 27896 4072
rect 27948 4060 27954 4072
rect 28813 4063 28871 4069
rect 28813 4060 28825 4063
rect 27948 4032 28825 4060
rect 27948 4020 27954 4032
rect 28813 4029 28825 4032
rect 28859 4029 28871 4063
rect 28813 4023 28871 4029
rect 29086 4020 29092 4072
rect 29144 4060 29150 4072
rect 29457 4063 29515 4069
rect 29457 4060 29469 4063
rect 29144 4032 29469 4060
rect 29144 4020 29150 4032
rect 29457 4029 29469 4032
rect 29503 4029 29515 4063
rect 29457 4023 29515 4029
rect 31113 4063 31171 4069
rect 31113 4029 31125 4063
rect 31159 4029 31171 4063
rect 31113 4023 31171 4029
rect 20162 3992 20168 4004
rect 18340 3964 20168 3992
rect 20162 3952 20168 3964
rect 20220 3952 20226 4004
rect 31128 3992 31156 4023
rect 31386 4020 31392 4072
rect 31444 4060 31450 4072
rect 32953 4063 33011 4069
rect 32953 4060 32965 4063
rect 31444 4032 32965 4060
rect 31444 4020 31450 4032
rect 32953 4029 32965 4032
rect 32999 4029 33011 4063
rect 32953 4023 33011 4029
rect 31754 3992 31760 4004
rect 31128 3964 31760 3992
rect 31754 3952 31760 3964
rect 31812 3952 31818 4004
rect 34054 3952 34060 4004
rect 34112 3992 34118 4004
rect 34885 3995 34943 4001
rect 34885 3992 34897 3995
rect 34112 3964 34897 3992
rect 34112 3952 34118 3964
rect 34885 3961 34897 3964
rect 34931 3961 34943 3995
rect 34885 3955 34943 3961
rect 12250 3884 12256 3936
rect 12308 3924 12314 3936
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 12308 3896 12357 3924
rect 12308 3884 12314 3896
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12345 3887 12403 3893
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 13173 3927 13231 3933
rect 13173 3924 13185 3927
rect 13136 3896 13185 3924
rect 13136 3884 13142 3896
rect 13173 3893 13185 3896
rect 13219 3893 13231 3927
rect 13173 3887 13231 3893
rect 13906 3884 13912 3936
rect 13964 3924 13970 3936
rect 14001 3927 14059 3933
rect 14001 3924 14013 3927
rect 13964 3896 14013 3924
rect 13964 3884 13970 3896
rect 14001 3893 14013 3896
rect 14047 3893 14059 3927
rect 14001 3887 14059 3893
rect 15013 3927 15071 3933
rect 15013 3893 15025 3927
rect 15059 3924 15071 3927
rect 15286 3924 15292 3936
rect 15059 3896 15292 3924
rect 15059 3893 15071 3896
rect 15013 3887 15071 3893
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 17129 3927 17187 3933
rect 17129 3893 17141 3927
rect 17175 3924 17187 3927
rect 17494 3924 17500 3936
rect 17175 3896 17500 3924
rect 17175 3893 17187 3896
rect 17129 3887 17187 3893
rect 17494 3884 17500 3896
rect 17552 3884 17558 3936
rect 17770 3924 17776 3936
rect 17731 3896 17776 3924
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 19153 3927 19211 3933
rect 19153 3893 19165 3927
rect 19199 3924 19211 3927
rect 22094 3924 22100 3936
rect 19199 3896 22100 3924
rect 19199 3893 19211 3896
rect 19153 3887 19211 3893
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 23017 3927 23075 3933
rect 23017 3893 23029 3927
rect 23063 3924 23075 3927
rect 24762 3924 24768 3936
rect 23063 3896 24768 3924
rect 23063 3893 23075 3896
rect 23017 3887 23075 3893
rect 24762 3884 24768 3896
rect 24820 3884 24826 3936
rect 25498 3884 25504 3936
rect 25556 3924 25562 3936
rect 26421 3927 26479 3933
rect 26421 3924 26433 3927
rect 25556 3896 26433 3924
rect 25556 3884 25562 3896
rect 26421 3893 26433 3896
rect 26467 3893 26479 3927
rect 26421 3887 26479 3893
rect 31846 3884 31852 3936
rect 31904 3924 31910 3936
rect 32401 3927 32459 3933
rect 32401 3924 32413 3927
rect 31904 3896 32413 3924
rect 31904 3884 31910 3896
rect 32401 3893 32413 3896
rect 32447 3893 32459 3927
rect 32401 3887 32459 3893
rect 32766 3884 32772 3936
rect 32824 3924 32830 3936
rect 33597 3927 33655 3933
rect 33597 3924 33609 3927
rect 32824 3896 33609 3924
rect 32824 3884 32830 3896
rect 33597 3893 33609 3896
rect 33643 3893 33655 3927
rect 33597 3887 33655 3893
rect 33778 3884 33784 3936
rect 33836 3924 33842 3936
rect 34241 3927 34299 3933
rect 34241 3924 34253 3927
rect 33836 3896 34253 3924
rect 33836 3884 33842 3896
rect 34241 3893 34253 3896
rect 34287 3893 34299 3927
rect 34241 3887 34299 3893
rect 35342 3884 35348 3936
rect 35400 3924 35406 3936
rect 35529 3927 35587 3933
rect 35529 3924 35541 3927
rect 35400 3896 35541 3924
rect 35400 3884 35406 3896
rect 35529 3893 35541 3896
rect 35575 3893 35587 3927
rect 35529 3887 35587 3893
rect 47302 3884 47308 3936
rect 47360 3924 47366 3936
rect 47765 3927 47823 3933
rect 47765 3924 47777 3927
rect 47360 3896 47777 3924
rect 47360 3884 47366 3896
rect 47765 3893 47777 3896
rect 47811 3893 47823 3927
rect 47765 3887 47823 3893
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 16853 3723 16911 3729
rect 16853 3689 16865 3723
rect 16899 3720 16911 3723
rect 17954 3720 17960 3732
rect 16899 3692 17960 3720
rect 16899 3689 16911 3692
rect 16853 3683 16911 3689
rect 17954 3680 17960 3692
rect 18012 3680 18018 3732
rect 18785 3723 18843 3729
rect 18785 3689 18797 3723
rect 18831 3720 18843 3723
rect 20254 3720 20260 3732
rect 18831 3692 20260 3720
rect 18831 3689 18843 3692
rect 18785 3683 18843 3689
rect 20254 3680 20260 3692
rect 20312 3680 20318 3732
rect 20349 3723 20407 3729
rect 20349 3689 20361 3723
rect 20395 3720 20407 3723
rect 24302 3720 24308 3732
rect 20395 3692 24308 3720
rect 20395 3689 20407 3692
rect 20349 3683 20407 3689
rect 24302 3680 24308 3692
rect 24360 3680 24366 3732
rect 27890 3720 27896 3732
rect 27851 3692 27896 3720
rect 27890 3680 27896 3692
rect 27948 3680 27954 3732
rect 30742 3680 30748 3732
rect 30800 3720 30806 3732
rect 33321 3723 33379 3729
rect 33321 3720 33333 3723
rect 30800 3692 33333 3720
rect 30800 3680 30806 3692
rect 33321 3689 33333 3692
rect 33367 3689 33379 3723
rect 33321 3683 33379 3689
rect 15013 3655 15071 3661
rect 15013 3621 15025 3655
rect 15059 3652 15071 3655
rect 16390 3652 16396 3664
rect 15059 3624 16396 3652
rect 15059 3621 15071 3624
rect 15013 3615 15071 3621
rect 16390 3612 16396 3624
rect 16448 3612 16454 3664
rect 17126 3612 17132 3664
rect 17184 3652 17190 3664
rect 20530 3652 20536 3664
rect 17184 3624 20536 3652
rect 17184 3612 17190 3624
rect 20530 3612 20536 3624
rect 20588 3612 20594 3664
rect 25130 3652 25136 3664
rect 20732 3624 23980 3652
rect 15657 3587 15715 3593
rect 15657 3553 15669 3587
rect 15703 3584 15715 3587
rect 17589 3587 17647 3593
rect 15703 3556 17540 3584
rect 15703 3553 15715 3556
rect 15657 3547 15715 3553
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 4614 3516 4620 3528
rect 4387 3488 4620 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 4890 3476 4896 3528
rect 4948 3516 4954 3528
rect 4985 3519 5043 3525
rect 4985 3516 4997 3519
rect 4948 3488 4997 3516
rect 4948 3476 4954 3488
rect 4985 3485 4997 3488
rect 5031 3485 5043 3519
rect 4985 3479 5043 3485
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 5813 3519 5871 3525
rect 5813 3516 5825 3519
rect 5776 3488 5825 3516
rect 5776 3476 5782 3488
rect 5813 3485 5825 3488
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 6546 3476 6552 3528
rect 6604 3516 6610 3528
rect 6641 3519 6699 3525
rect 6641 3516 6653 3519
rect 6604 3488 6653 3516
rect 6604 3476 6610 3488
rect 6641 3485 6653 3488
rect 6687 3485 6699 3519
rect 6641 3479 6699 3485
rect 7374 3476 7380 3528
rect 7432 3516 7438 3528
rect 7469 3519 7527 3525
rect 7469 3516 7481 3519
rect 7432 3488 7481 3516
rect 7432 3476 7438 3488
rect 7469 3485 7481 3488
rect 7515 3485 7527 3519
rect 7469 3479 7527 3485
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 8260 3488 8309 3516
rect 8260 3476 8266 3488
rect 8297 3485 8309 3488
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 9088 3488 9137 3516
rect 9088 3476 9094 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9858 3476 9864 3528
rect 9916 3516 9922 3528
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 9916 3488 9965 3516
rect 9916 3476 9922 3488
rect 9953 3485 9965 3488
rect 9999 3485 10011 3519
rect 9953 3479 10011 3485
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 10781 3519 10839 3525
rect 10781 3516 10793 3519
rect 10744 3488 10793 3516
rect 10744 3476 10750 3488
rect 10781 3485 10793 3488
rect 10827 3485 10839 3519
rect 10781 3479 10839 3485
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 11609 3519 11667 3525
rect 11609 3516 11621 3519
rect 11572 3488 11621 3516
rect 11572 3476 11578 3488
rect 11609 3485 11621 3488
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3516 12495 3519
rect 12802 3516 12808 3528
rect 12483 3488 12808 3516
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3516 13139 3519
rect 13630 3516 13636 3528
rect 13127 3488 13636 3516
rect 13127 3485 13139 3488
rect 13081 3479 13139 3485
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3516 13783 3519
rect 14182 3516 14188 3528
rect 13771 3488 14188 3516
rect 13771 3485 13783 3488
rect 13725 3479 13783 3485
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 16114 3516 16120 3528
rect 16027 3488 16120 3516
rect 16114 3476 16120 3488
rect 16172 3516 16178 3528
rect 16758 3516 16764 3528
rect 16172 3488 16764 3516
rect 16172 3476 16178 3488
rect 16758 3476 16764 3488
rect 16816 3476 16822 3528
rect 17512 3516 17540 3556
rect 17589 3553 17601 3587
rect 17635 3584 17647 3587
rect 19242 3584 19248 3596
rect 17635 3556 19248 3584
rect 17635 3553 17647 3556
rect 17589 3547 17647 3553
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 19720 3556 20300 3584
rect 17954 3516 17960 3528
rect 17512 3488 17960 3516
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 18233 3519 18291 3525
rect 18233 3485 18245 3519
rect 18279 3516 18291 3519
rect 18693 3519 18751 3525
rect 18693 3516 18705 3519
rect 18279 3488 18705 3516
rect 18279 3485 18291 3488
rect 18233 3479 18291 3485
rect 18693 3485 18705 3488
rect 18739 3516 18751 3519
rect 19720 3516 19748 3556
rect 20272 3525 20300 3556
rect 18739 3488 19748 3516
rect 19797 3519 19855 3525
rect 18739 3485 18751 3488
rect 18693 3479 18751 3485
rect 19797 3485 19809 3519
rect 19843 3485 19855 3519
rect 19797 3479 19855 3485
rect 20257 3519 20315 3525
rect 20257 3485 20269 3519
rect 20303 3516 20315 3519
rect 20732 3516 20760 3624
rect 20806 3544 20812 3596
rect 20864 3584 20870 3596
rect 21545 3587 21603 3593
rect 21545 3584 21557 3587
rect 20864 3556 21557 3584
rect 20864 3544 20870 3556
rect 21545 3553 21557 3556
rect 21591 3553 21603 3587
rect 21726 3584 21732 3596
rect 21687 3556 21732 3584
rect 21545 3547 21603 3553
rect 21726 3544 21732 3556
rect 21784 3544 21790 3596
rect 22186 3584 22192 3596
rect 22147 3556 22192 3584
rect 22186 3544 22192 3556
rect 22244 3544 22250 3596
rect 20901 3519 20959 3525
rect 20901 3516 20913 3519
rect 20303 3488 20913 3516
rect 20303 3485 20315 3488
rect 20257 3479 20315 3485
rect 20901 3485 20913 3488
rect 20947 3485 20959 3519
rect 20901 3479 20959 3485
rect 18141 3451 18199 3457
rect 18141 3417 18153 3451
rect 18187 3448 18199 3451
rect 19812 3448 19840 3479
rect 22462 3448 22468 3460
rect 18187 3420 19748 3448
rect 19812 3420 22468 3448
rect 18187 3417 18199 3420
rect 18141 3411 18199 3417
rect 16209 3383 16267 3389
rect 16209 3349 16221 3383
rect 16255 3380 16267 3383
rect 16758 3380 16764 3392
rect 16255 3352 16764 3380
rect 16255 3349 16267 3352
rect 16209 3343 16267 3349
rect 16758 3340 16764 3352
rect 16816 3340 16822 3392
rect 19720 3380 19748 3420
rect 22462 3408 22468 3420
rect 22520 3408 22526 3460
rect 23952 3448 23980 3624
rect 24044 3624 25136 3652
rect 24044 3525 24072 3624
rect 25130 3612 25136 3624
rect 25188 3652 25194 3664
rect 25188 3624 26234 3652
rect 25188 3612 25194 3624
rect 25498 3584 25504 3596
rect 25459 3556 25504 3584
rect 25498 3544 25504 3556
rect 25556 3544 25562 3596
rect 26050 3584 26056 3596
rect 26011 3556 26056 3584
rect 26050 3544 26056 3556
rect 26108 3544 26114 3596
rect 26206 3584 26234 3624
rect 30190 3612 30196 3664
rect 30248 3652 30254 3664
rect 30248 3624 31708 3652
rect 30248 3612 30254 3624
rect 26206 3556 27752 3584
rect 24029 3519 24087 3525
rect 24029 3485 24041 3519
rect 24075 3485 24087 3519
rect 24854 3516 24860 3528
rect 24767 3488 24860 3516
rect 24029 3479 24087 3485
rect 24854 3476 24860 3488
rect 24912 3476 24918 3528
rect 27724 3516 27752 3556
rect 31202 3544 31208 3596
rect 31260 3584 31266 3596
rect 31573 3587 31631 3593
rect 31573 3584 31585 3587
rect 31260 3556 31585 3584
rect 31260 3544 31266 3556
rect 31573 3553 31585 3556
rect 31619 3553 31631 3587
rect 31680 3584 31708 3624
rect 31754 3612 31760 3664
rect 31812 3652 31818 3664
rect 31812 3624 32812 3652
rect 31812 3612 31818 3624
rect 31680 3556 32536 3584
rect 31573 3547 31631 3553
rect 27798 3516 27804 3528
rect 27711 3488 27804 3516
rect 27798 3476 27804 3488
rect 27856 3476 27862 3528
rect 28629 3519 28687 3525
rect 28629 3485 28641 3519
rect 28675 3516 28687 3519
rect 28994 3516 29000 3528
rect 28675 3488 29000 3516
rect 28675 3485 28687 3488
rect 28629 3479 28687 3485
rect 28994 3476 29000 3488
rect 29052 3476 29058 3528
rect 32122 3476 32128 3528
rect 32180 3516 32186 3528
rect 32217 3519 32275 3525
rect 32217 3516 32229 3519
rect 32180 3488 32229 3516
rect 32180 3476 32186 3488
rect 32217 3485 32229 3488
rect 32263 3485 32275 3519
rect 32217 3479 32275 3485
rect 24872 3448 24900 3476
rect 23952 3420 24900 3448
rect 24949 3451 25007 3457
rect 24949 3417 24961 3451
rect 24995 3448 25007 3451
rect 25685 3451 25743 3457
rect 25685 3448 25697 3451
rect 24995 3420 25697 3448
rect 24995 3417 25007 3420
rect 24949 3411 25007 3417
rect 25685 3417 25697 3420
rect 25731 3417 25743 3451
rect 25685 3411 25743 3417
rect 28258 3408 28264 3460
rect 28316 3448 28322 3460
rect 29733 3451 29791 3457
rect 29733 3448 29745 3451
rect 28316 3420 29745 3448
rect 28316 3408 28322 3420
rect 29733 3417 29745 3420
rect 29779 3417 29791 3451
rect 29733 3411 29791 3417
rect 31389 3451 31447 3457
rect 31389 3417 31401 3451
rect 31435 3448 31447 3451
rect 32398 3448 32404 3460
rect 31435 3420 32404 3448
rect 31435 3417 31447 3420
rect 31389 3411 31447 3417
rect 32398 3408 32404 3420
rect 32456 3408 32462 3460
rect 32508 3448 32536 3556
rect 32674 3516 32680 3528
rect 32635 3488 32680 3516
rect 32674 3476 32680 3488
rect 32732 3476 32738 3528
rect 32784 3516 32812 3624
rect 33226 3612 33232 3664
rect 33284 3652 33290 3664
rect 34885 3655 34943 3661
rect 34885 3652 34897 3655
rect 33284 3624 34897 3652
rect 33284 3612 33290 3624
rect 34885 3621 34897 3624
rect 34931 3621 34943 3655
rect 34885 3615 34943 3621
rect 35434 3612 35440 3664
rect 35492 3652 35498 3664
rect 36173 3655 36231 3661
rect 36173 3652 36185 3655
rect 35492 3624 36185 3652
rect 35492 3612 35498 3624
rect 36173 3621 36185 3624
rect 36219 3621 36231 3655
rect 36173 3615 36231 3621
rect 37458 3612 37464 3664
rect 37516 3652 37522 3664
rect 38105 3655 38163 3661
rect 38105 3652 38117 3655
rect 37516 3624 38117 3652
rect 37516 3612 37522 3624
rect 38105 3621 38117 3624
rect 38151 3621 38163 3655
rect 38105 3615 38163 3621
rect 40678 3612 40684 3664
rect 40736 3652 40742 3664
rect 41325 3655 41383 3661
rect 41325 3652 41337 3655
rect 40736 3624 41337 3652
rect 40736 3612 40742 3624
rect 41325 3621 41337 3624
rect 41371 3621 41383 3655
rect 41325 3615 41383 3621
rect 46474 3612 46480 3664
rect 46532 3652 46538 3664
rect 47121 3655 47179 3661
rect 47121 3652 47133 3655
rect 46532 3624 47133 3652
rect 46532 3612 46538 3624
rect 47121 3621 47133 3624
rect 47167 3621 47179 3655
rect 47121 3615 47179 3621
rect 34514 3584 34520 3596
rect 33704 3556 34520 3584
rect 33704 3516 33732 3556
rect 34514 3544 34520 3556
rect 34572 3544 34578 3596
rect 34606 3544 34612 3596
rect 34664 3584 34670 3596
rect 35529 3587 35587 3593
rect 35529 3584 35541 3587
rect 34664 3556 35541 3584
rect 34664 3544 34670 3556
rect 35529 3553 35541 3556
rect 35575 3553 35587 3587
rect 35529 3547 35587 3553
rect 35986 3544 35992 3596
rect 36044 3584 36050 3596
rect 36817 3587 36875 3593
rect 36817 3584 36829 3587
rect 36044 3556 36829 3584
rect 36044 3544 36050 3556
rect 36817 3553 36829 3556
rect 36863 3553 36875 3587
rect 36817 3547 36875 3553
rect 41230 3544 41236 3596
rect 41288 3584 41294 3596
rect 41969 3587 42027 3593
rect 41969 3584 41981 3587
rect 41288 3556 41981 3584
rect 41288 3544 41294 3556
rect 41969 3553 41981 3556
rect 42015 3553 42027 3587
rect 41969 3547 42027 3553
rect 47026 3544 47032 3596
rect 47084 3584 47090 3596
rect 47765 3587 47823 3593
rect 47765 3584 47777 3587
rect 47084 3556 47777 3584
rect 47084 3544 47090 3556
rect 47765 3553 47777 3556
rect 47811 3553 47823 3587
rect 47765 3547 47823 3553
rect 32784 3488 33732 3516
rect 33965 3519 34023 3525
rect 33965 3485 33977 3519
rect 34011 3485 34023 3519
rect 33965 3479 34023 3485
rect 33594 3448 33600 3460
rect 32508 3420 33600 3448
rect 33594 3408 33600 3420
rect 33652 3408 33658 3460
rect 20622 3380 20628 3392
rect 19720 3352 20628 3380
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 20993 3383 21051 3389
rect 20993 3349 21005 3383
rect 21039 3380 21051 3383
rect 23842 3380 23848 3392
rect 21039 3352 23848 3380
rect 21039 3349 21051 3352
rect 20993 3343 21051 3349
rect 23842 3340 23848 3352
rect 23900 3340 23906 3392
rect 23937 3383 23995 3389
rect 23937 3349 23949 3383
rect 23983 3380 23995 3383
rect 28810 3380 28816 3392
rect 23983 3352 28816 3380
rect 23983 3349 23995 3352
rect 23937 3343 23995 3349
rect 28810 3340 28816 3352
rect 28868 3340 28874 3392
rect 30466 3340 30472 3392
rect 30524 3380 30530 3392
rect 31754 3380 31760 3392
rect 30524 3352 31760 3380
rect 30524 3340 30530 3352
rect 31754 3340 31760 3352
rect 31812 3340 31818 3392
rect 31938 3340 31944 3392
rect 31996 3380 32002 3392
rect 32125 3383 32183 3389
rect 32125 3380 32137 3383
rect 31996 3352 32137 3380
rect 31996 3340 32002 3352
rect 32125 3349 32137 3352
rect 32171 3349 32183 3383
rect 32125 3343 32183 3349
rect 32214 3340 32220 3392
rect 32272 3380 32278 3392
rect 33980 3380 34008 3479
rect 36538 3476 36544 3528
rect 36596 3516 36602 3528
rect 37461 3519 37519 3525
rect 37461 3516 37473 3519
rect 36596 3488 37473 3516
rect 36596 3476 36602 3488
rect 37461 3485 37473 3488
rect 37507 3485 37519 3519
rect 37461 3479 37519 3485
rect 37918 3476 37924 3528
rect 37976 3516 37982 3528
rect 38749 3519 38807 3525
rect 38749 3516 38761 3519
rect 37976 3488 38761 3516
rect 37976 3476 37982 3488
rect 38749 3485 38761 3488
rect 38795 3485 38807 3519
rect 38749 3479 38807 3485
rect 39298 3476 39304 3528
rect 39356 3516 39362 3528
rect 40037 3519 40095 3525
rect 40037 3516 40049 3519
rect 39356 3488 40049 3516
rect 39356 3476 39362 3488
rect 40037 3485 40049 3488
rect 40083 3485 40095 3519
rect 40037 3479 40095 3485
rect 40126 3476 40132 3528
rect 40184 3516 40190 3528
rect 40681 3519 40739 3525
rect 40681 3516 40693 3519
rect 40184 3488 40693 3516
rect 40184 3476 40190 3488
rect 40681 3485 40693 3488
rect 40727 3485 40739 3519
rect 40681 3479 40739 3485
rect 42610 3476 42616 3528
rect 42668 3516 42674 3528
rect 42705 3519 42763 3525
rect 42705 3516 42717 3519
rect 42668 3488 42717 3516
rect 42668 3476 42674 3488
rect 42705 3485 42717 3488
rect 42751 3485 42763 3519
rect 42705 3479 42763 3485
rect 42886 3476 42892 3528
rect 42944 3516 42950 3528
rect 43349 3519 43407 3525
rect 43349 3516 43361 3519
rect 42944 3488 43361 3516
rect 42944 3476 42950 3488
rect 43349 3485 43361 3488
rect 43395 3485 43407 3519
rect 43349 3479 43407 3485
rect 44542 3476 44548 3528
rect 44600 3516 44606 3528
rect 45189 3519 45247 3525
rect 45189 3516 45201 3519
rect 44600 3488 45201 3516
rect 44600 3476 44606 3488
rect 45189 3485 45201 3488
rect 45235 3485 45247 3519
rect 45189 3479 45247 3485
rect 45370 3476 45376 3528
rect 45428 3516 45434 3528
rect 45833 3519 45891 3525
rect 45833 3516 45845 3519
rect 45428 3488 45845 3516
rect 45428 3476 45434 3488
rect 45833 3485 45845 3488
rect 45879 3485 45891 3519
rect 45833 3479 45891 3485
rect 46198 3476 46204 3528
rect 46256 3516 46262 3528
rect 46477 3519 46535 3525
rect 46477 3516 46489 3519
rect 46256 3488 46489 3516
rect 46256 3476 46262 3488
rect 46477 3485 46489 3488
rect 46523 3485 46535 3519
rect 46477 3479 46535 3485
rect 32272 3352 34008 3380
rect 32272 3340 32278 3352
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 19150 3176 19156 3188
rect 15028 3148 19156 3176
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 14458 3040 14464 3052
rect 13127 3012 14464 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 15028 3049 15056 3148
rect 19150 3136 19156 3148
rect 19208 3136 19214 3188
rect 23750 3176 23756 3188
rect 19628 3148 23756 3176
rect 17494 3108 17500 3120
rect 17455 3080 17500 3108
rect 17494 3068 17500 3080
rect 17552 3068 17558 3120
rect 17770 3068 17776 3120
rect 17828 3108 17834 3120
rect 17828 3080 19472 3108
rect 17828 3068 17834 3080
rect 15013 3043 15071 3049
rect 15013 3009 15025 3043
rect 15059 3009 15071 3043
rect 16114 3040 16120 3052
rect 16075 3012 16120 3040
rect 15013 3003 15071 3009
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 4065 2975 4123 2981
rect 4065 2941 4077 2975
rect 4111 2972 4123 2975
rect 4706 2972 4712 2984
rect 4111 2944 4712 2972
rect 4111 2941 4123 2944
rect 4065 2935 4123 2941
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 5353 2975 5411 2981
rect 5353 2941 5365 2975
rect 5399 2972 5411 2975
rect 5994 2972 6000 2984
rect 5399 2944 6000 2972
rect 5399 2941 5411 2944
rect 5353 2935 5411 2941
rect 5994 2932 6000 2944
rect 6052 2932 6058 2984
rect 14369 2975 14427 2981
rect 14369 2941 14381 2975
rect 14415 2972 14427 2975
rect 16666 2972 16672 2984
rect 14415 2944 16672 2972
rect 14415 2941 14427 2944
rect 14369 2935 14427 2941
rect 16666 2932 16672 2944
rect 16724 2932 16730 2984
rect 17313 2975 17371 2981
rect 17313 2941 17325 2975
rect 17359 2972 17371 2975
rect 18046 2972 18052 2984
rect 17359 2944 18052 2972
rect 17359 2941 17371 2944
rect 17313 2935 17371 2941
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18969 2975 19027 2981
rect 18969 2941 18981 2975
rect 19015 2941 19027 2975
rect 19444 2972 19472 3080
rect 19628 3049 19656 3148
rect 23750 3136 23756 3148
rect 23808 3136 23814 3188
rect 27982 3136 27988 3188
rect 28040 3176 28046 3188
rect 29178 3176 29184 3188
rect 28040 3148 29184 3176
rect 28040 3136 28046 3148
rect 29178 3136 29184 3148
rect 29236 3136 29242 3188
rect 29914 3136 29920 3188
rect 29972 3176 29978 3188
rect 33686 3176 33692 3188
rect 29972 3148 33692 3176
rect 29972 3136 29978 3148
rect 33686 3136 33692 3148
rect 33744 3136 33750 3188
rect 20254 3068 20260 3120
rect 20312 3108 20318 3120
rect 22649 3111 22707 3117
rect 22649 3108 22661 3111
rect 20312 3080 22661 3108
rect 20312 3068 20318 3080
rect 22649 3077 22661 3080
rect 22695 3077 22707 3111
rect 22649 3071 22707 3077
rect 23842 3068 23848 3120
rect 23900 3108 23906 3120
rect 24949 3111 25007 3117
rect 24949 3108 24961 3111
rect 23900 3080 24961 3108
rect 23900 3068 23906 3080
rect 24949 3077 24961 3080
rect 24995 3077 25007 3111
rect 28810 3108 28816 3120
rect 28771 3080 28816 3108
rect 24949 3071 25007 3077
rect 28810 3068 28816 3080
rect 28868 3068 28874 3120
rect 31113 3111 31171 3117
rect 31113 3077 31125 3111
rect 31159 3108 31171 3111
rect 33042 3108 33048 3120
rect 31159 3080 33048 3108
rect 31159 3077 31171 3080
rect 31113 3071 31171 3077
rect 33042 3068 33048 3080
rect 33100 3068 33106 3120
rect 33502 3068 33508 3120
rect 33560 3108 33566 3120
rect 36170 3108 36176 3120
rect 33560 3080 36176 3108
rect 33560 3068 33566 3080
rect 36170 3068 36176 3080
rect 36228 3068 36234 3120
rect 19613 3043 19671 3049
rect 19613 3009 19625 3043
rect 19659 3009 19671 3043
rect 22462 3040 22468 3052
rect 22423 3012 22468 3040
rect 19613 3003 19671 3009
rect 22462 3000 22468 3012
rect 22520 3000 22526 3052
rect 24762 3040 24768 3052
rect 24723 3012 24768 3040
rect 24762 3000 24768 3012
rect 24820 3000 24826 3052
rect 28994 3000 29000 3052
rect 29052 3040 29058 3052
rect 29052 3012 29097 3040
rect 29052 3000 29058 3012
rect 32858 3000 32864 3052
rect 32916 3040 32922 3052
rect 33594 3040 33600 3052
rect 32916 3012 33088 3040
rect 33555 3012 33600 3040
rect 32916 3000 32922 3012
rect 19797 2975 19855 2981
rect 19797 2972 19809 2975
rect 19444 2944 19809 2972
rect 18969 2935 19027 2941
rect 19797 2941 19809 2944
rect 19843 2941 19855 2975
rect 19797 2935 19855 2941
rect 21453 2975 21511 2981
rect 21453 2941 21465 2975
rect 21499 2972 21511 2975
rect 23842 2972 23848 2984
rect 21499 2944 23848 2972
rect 21499 2941 21511 2944
rect 21453 2935 21511 2941
rect 12437 2907 12495 2913
rect 12437 2873 12449 2907
rect 12483 2904 12495 2907
rect 13354 2904 13360 2916
rect 12483 2876 13360 2904
rect 12483 2873 12495 2876
rect 12437 2867 12495 2873
rect 13354 2864 13360 2876
rect 13412 2864 13418 2916
rect 15657 2907 15715 2913
rect 15657 2873 15669 2907
rect 15703 2904 15715 2907
rect 17126 2904 17132 2916
rect 15703 2876 17132 2904
rect 15703 2873 15715 2876
rect 15657 2867 15715 2873
rect 17126 2864 17132 2876
rect 17184 2864 17190 2916
rect 3421 2839 3479 2845
rect 3421 2805 3433 2839
rect 3467 2836 3479 2839
rect 3510 2836 3516 2848
rect 3467 2808 3516 2836
rect 3467 2805 3479 2808
rect 3421 2799 3479 2805
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 4709 2839 4767 2845
rect 4709 2805 4721 2839
rect 4755 2836 4767 2839
rect 5166 2836 5172 2848
rect 4755 2808 5172 2836
rect 4755 2805 4767 2808
rect 4709 2799 4767 2805
rect 5166 2796 5172 2808
rect 5224 2796 5230 2848
rect 5997 2839 6055 2845
rect 5997 2805 6009 2839
rect 6043 2836 6055 2839
rect 6270 2836 6276 2848
rect 6043 2808 6276 2836
rect 6043 2805 6055 2808
rect 5997 2799 6055 2805
rect 6270 2796 6276 2808
rect 6328 2796 6334 2848
rect 7285 2839 7343 2845
rect 7285 2805 7297 2839
rect 7331 2836 7343 2839
rect 7650 2836 7656 2848
rect 7331 2808 7656 2836
rect 7331 2805 7343 2808
rect 7285 2799 7343 2805
rect 7650 2796 7656 2808
rect 7708 2796 7714 2848
rect 7929 2839 7987 2845
rect 7929 2805 7941 2839
rect 7975 2836 7987 2839
rect 8478 2836 8484 2848
rect 7975 2808 8484 2836
rect 7975 2805 7987 2808
rect 7929 2799 7987 2805
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 8573 2839 8631 2845
rect 8573 2805 8585 2839
rect 8619 2836 8631 2839
rect 8754 2836 8760 2848
rect 8619 2808 8760 2836
rect 8619 2805 8631 2808
rect 8573 2799 8631 2805
rect 8754 2796 8760 2808
rect 8812 2796 8818 2848
rect 9217 2839 9275 2845
rect 9217 2805 9229 2839
rect 9263 2836 9275 2839
rect 9582 2836 9588 2848
rect 9263 2808 9588 2836
rect 9263 2805 9275 2808
rect 9217 2799 9275 2805
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 9861 2839 9919 2845
rect 9861 2805 9873 2839
rect 9907 2836 9919 2839
rect 10410 2836 10416 2848
rect 9907 2808 10416 2836
rect 9907 2805 9919 2808
rect 9861 2799 9919 2805
rect 10410 2796 10416 2808
rect 10468 2796 10474 2848
rect 10505 2839 10563 2845
rect 10505 2805 10517 2839
rect 10551 2836 10563 2839
rect 10962 2836 10968 2848
rect 10551 2808 10968 2836
rect 10551 2805 10563 2808
rect 10505 2799 10563 2805
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2836 11207 2839
rect 11790 2836 11796 2848
rect 11195 2808 11796 2836
rect 11195 2805 11207 2808
rect 11149 2799 11207 2805
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 13725 2839 13783 2845
rect 13725 2805 13737 2839
rect 13771 2836 13783 2839
rect 16114 2836 16120 2848
rect 13771 2808 16120 2836
rect 13771 2805 13783 2808
rect 13725 2799 13783 2805
rect 16114 2796 16120 2808
rect 16172 2796 16178 2848
rect 16209 2839 16267 2845
rect 16209 2805 16221 2839
rect 16255 2836 16267 2839
rect 17862 2836 17868 2848
rect 16255 2808 17868 2836
rect 16255 2805 16267 2808
rect 16209 2799 16267 2805
rect 17862 2796 17868 2808
rect 17920 2796 17926 2848
rect 17954 2796 17960 2848
rect 18012 2836 18018 2848
rect 18874 2836 18880 2848
rect 18012 2808 18880 2836
rect 18012 2796 18018 2808
rect 18874 2796 18880 2808
rect 18932 2796 18938 2848
rect 18984 2836 19012 2935
rect 23842 2932 23848 2944
rect 23900 2932 23906 2984
rect 24305 2975 24363 2981
rect 24305 2941 24317 2975
rect 24351 2972 24363 2975
rect 24394 2972 24400 2984
rect 24351 2944 24400 2972
rect 24351 2941 24363 2944
rect 24305 2935 24363 2941
rect 24394 2932 24400 2944
rect 24452 2932 24458 2984
rect 25498 2972 25504 2984
rect 25459 2944 25504 2972
rect 25498 2932 25504 2944
rect 25556 2932 25562 2984
rect 26878 2932 26884 2984
rect 26936 2972 26942 2984
rect 27157 2975 27215 2981
rect 27157 2972 27169 2975
rect 26936 2944 27169 2972
rect 26936 2932 26942 2944
rect 27157 2941 27169 2944
rect 27203 2941 27215 2975
rect 27157 2935 27215 2941
rect 28534 2932 28540 2984
rect 28592 2972 28598 2984
rect 29457 2975 29515 2981
rect 29457 2972 29469 2975
rect 28592 2944 29469 2972
rect 28592 2932 28598 2944
rect 29457 2941 29469 2944
rect 29503 2941 29515 2975
rect 29457 2935 29515 2941
rect 31297 2975 31355 2981
rect 31297 2941 31309 2975
rect 31343 2972 31355 2975
rect 32953 2975 33011 2981
rect 32953 2972 32965 2975
rect 31343 2944 32965 2972
rect 31343 2941 31355 2944
rect 31297 2935 31355 2941
rect 32953 2941 32965 2944
rect 32999 2941 33011 2975
rect 33060 2972 33088 3012
rect 33594 3000 33600 3012
rect 33652 3000 33658 3052
rect 35529 3043 35587 3049
rect 35529 3040 35541 3043
rect 33704 3012 35541 3040
rect 33704 2972 33732 3012
rect 35529 3009 35541 3012
rect 35575 3009 35587 3043
rect 35529 3003 35587 3009
rect 35710 3000 35716 3052
rect 35768 3040 35774 3052
rect 37461 3043 37519 3049
rect 37461 3040 37473 3043
rect 35768 3012 37473 3040
rect 35768 3000 35774 3012
rect 37461 3009 37473 3012
rect 37507 3009 37519 3043
rect 37461 3003 37519 3009
rect 33060 2944 33732 2972
rect 32953 2935 33011 2941
rect 34790 2932 34796 2984
rect 34848 2972 34854 2984
rect 37366 2972 37372 2984
rect 34848 2944 37372 2972
rect 34848 2932 34854 2944
rect 37366 2932 37372 2944
rect 37424 2932 37430 2984
rect 37642 2932 37648 2984
rect 37700 2972 37706 2984
rect 38749 2975 38807 2981
rect 38749 2972 38761 2975
rect 37700 2944 38761 2972
rect 37700 2932 37706 2944
rect 38749 2941 38761 2944
rect 38795 2941 38807 2975
rect 38749 2935 38807 2941
rect 39850 2932 39856 2984
rect 39908 2972 39914 2984
rect 40681 2975 40739 2981
rect 40681 2972 40693 2975
rect 39908 2944 40693 2972
rect 39908 2932 39914 2944
rect 40681 2941 40693 2944
rect 40727 2941 40739 2975
rect 40681 2935 40739 2941
rect 42334 2932 42340 2984
rect 42392 2972 42398 2984
rect 43257 2975 43315 2981
rect 43257 2972 43269 2975
rect 42392 2944 43269 2972
rect 42392 2932 42398 2944
rect 43257 2941 43269 2944
rect 43303 2941 43315 2975
rect 43257 2935 43315 2941
rect 44266 2932 44272 2984
rect 44324 2972 44330 2984
rect 45189 2975 45247 2981
rect 45189 2972 45201 2975
rect 44324 2944 45201 2972
rect 44324 2932 44330 2944
rect 45189 2941 45201 2944
rect 45235 2941 45247 2975
rect 45189 2935 45247 2941
rect 31018 2864 31024 2916
rect 31076 2904 31082 2916
rect 34241 2907 34299 2913
rect 34241 2904 34253 2907
rect 31076 2876 34253 2904
rect 31076 2864 31082 2876
rect 34241 2873 34253 2876
rect 34287 2873 34299 2907
rect 34241 2867 34299 2873
rect 34330 2864 34336 2916
rect 34388 2904 34394 2916
rect 36173 2907 36231 2913
rect 36173 2904 36185 2907
rect 34388 2876 36185 2904
rect 34388 2864 34394 2876
rect 36173 2873 36185 2876
rect 36219 2873 36231 2907
rect 36173 2867 36231 2873
rect 36814 2864 36820 2916
rect 36872 2904 36878 2916
rect 38105 2907 38163 2913
rect 38105 2904 38117 2907
rect 36872 2876 38117 2904
rect 36872 2864 36878 2876
rect 38105 2873 38117 2876
rect 38151 2873 38163 2907
rect 38105 2867 38163 2873
rect 38470 2864 38476 2916
rect 38528 2904 38534 2916
rect 39393 2907 39451 2913
rect 39393 2904 39405 2907
rect 38528 2876 39405 2904
rect 38528 2864 38534 2876
rect 39393 2873 39405 2876
rect 39439 2873 39451 2907
rect 39393 2867 39451 2873
rect 40402 2864 40408 2916
rect 40460 2904 40466 2916
rect 41325 2907 41383 2913
rect 41325 2904 41337 2907
rect 40460 2876 41337 2904
rect 40460 2864 40466 2876
rect 41325 2873 41337 2876
rect 41371 2873 41383 2907
rect 41325 2867 41383 2873
rect 43162 2864 43168 2916
rect 43220 2904 43226 2916
rect 43901 2907 43959 2913
rect 43901 2904 43913 2907
rect 43220 2876 43913 2904
rect 43220 2864 43226 2876
rect 43901 2873 43913 2876
rect 43947 2873 43959 2907
rect 43901 2867 43959 2873
rect 45094 2864 45100 2916
rect 45152 2904 45158 2916
rect 45833 2907 45891 2913
rect 45833 2904 45845 2907
rect 45152 2876 45845 2904
rect 45152 2864 45158 2876
rect 45833 2873 45845 2876
rect 45879 2873 45891 2907
rect 45833 2867 45891 2873
rect 21634 2836 21640 2848
rect 18984 2808 21640 2836
rect 21634 2796 21640 2808
rect 21692 2796 21698 2848
rect 28810 2796 28816 2848
rect 28868 2836 28874 2848
rect 30006 2836 30012 2848
rect 28868 2808 30012 2836
rect 28868 2796 28874 2808
rect 30006 2796 30012 2808
rect 30064 2796 30070 2848
rect 30374 2796 30380 2848
rect 30432 2836 30438 2848
rect 32309 2839 32367 2845
rect 32309 2836 32321 2839
rect 30432 2808 32321 2836
rect 30432 2796 30438 2808
rect 32309 2805 32321 2808
rect 32355 2805 32367 2839
rect 32309 2799 32367 2805
rect 32490 2796 32496 2848
rect 32548 2836 32554 2848
rect 34885 2839 34943 2845
rect 34885 2836 34897 2839
rect 32548 2808 34897 2836
rect 32548 2796 32554 2808
rect 34885 2805 34897 2808
rect 34931 2805 34943 2839
rect 34885 2799 34943 2805
rect 38746 2796 38752 2848
rect 38804 2836 38810 2848
rect 40037 2839 40095 2845
rect 40037 2836 40049 2839
rect 38804 2808 40049 2836
rect 38804 2796 38810 2808
rect 40037 2805 40049 2808
rect 40083 2805 40095 2839
rect 40037 2799 40095 2805
rect 41782 2796 41788 2848
rect 41840 2836 41846 2848
rect 42613 2839 42671 2845
rect 42613 2836 42625 2839
rect 41840 2808 42625 2836
rect 41840 2796 41846 2808
rect 42613 2805 42625 2808
rect 42659 2805 42671 2839
rect 42613 2799 42671 2805
rect 43714 2796 43720 2848
rect 43772 2836 43778 2848
rect 44545 2839 44603 2845
rect 44545 2836 44557 2839
rect 43772 2808 44557 2836
rect 43772 2796 43778 2808
rect 44545 2805 44557 2808
rect 44591 2805 44603 2839
rect 44545 2799 44603 2805
rect 45646 2796 45652 2848
rect 45704 2836 45710 2848
rect 46477 2839 46535 2845
rect 46477 2836 46489 2839
rect 45704 2808 46489 2836
rect 45704 2796 45710 2808
rect 46477 2805 46489 2808
rect 46523 2805 46535 2839
rect 46477 2799 46535 2805
rect 46750 2796 46756 2848
rect 46808 2836 46814 2848
rect 47765 2839 47823 2845
rect 47765 2836 47777 2839
rect 46808 2808 47777 2836
rect 46808 2796 46814 2808
rect 47765 2805 47777 2808
rect 47811 2805 47823 2839
rect 47765 2799 47823 2805
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 13725 2635 13783 2641
rect 13725 2601 13737 2635
rect 13771 2632 13783 2635
rect 18046 2632 18052 2644
rect 13771 2604 18052 2632
rect 13771 2601 13783 2604
rect 13725 2595 13783 2601
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 32398 2632 32404 2644
rect 32359 2604 32404 2632
rect 32398 2592 32404 2604
rect 32456 2592 32462 2644
rect 33042 2632 33048 2644
rect 33003 2604 33048 2632
rect 33042 2592 33048 2604
rect 33100 2592 33106 2644
rect 33594 2632 33600 2644
rect 33555 2604 33600 2632
rect 33594 2592 33600 2604
rect 33652 2592 33658 2644
rect 34514 2592 34520 2644
rect 34572 2632 34578 2644
rect 34885 2635 34943 2641
rect 34885 2632 34897 2635
rect 34572 2604 34897 2632
rect 34572 2592 34578 2604
rect 34885 2601 34897 2604
rect 34931 2601 34943 2635
rect 36170 2632 36176 2644
rect 36131 2604 36176 2632
rect 34885 2595 34943 2601
rect 36170 2592 36176 2604
rect 36228 2592 36234 2644
rect 37366 2592 37372 2644
rect 37424 2632 37430 2644
rect 37461 2635 37519 2641
rect 37461 2632 37473 2635
rect 37424 2604 37473 2632
rect 37424 2592 37430 2604
rect 37461 2601 37473 2604
rect 37507 2601 37519 2635
rect 37461 2595 37519 2601
rect 5353 2567 5411 2573
rect 5353 2533 5365 2567
rect 5399 2564 5411 2567
rect 6822 2564 6828 2576
rect 5399 2536 6828 2564
rect 5399 2533 5411 2536
rect 5353 2527 5411 2533
rect 6822 2524 6828 2536
rect 6880 2524 6886 2576
rect 7285 2567 7343 2573
rect 7285 2533 7297 2567
rect 7331 2564 7343 2567
rect 7926 2564 7932 2576
rect 7331 2536 7932 2564
rect 7331 2533 7343 2536
rect 7285 2527 7343 2533
rect 7926 2524 7932 2536
rect 7984 2524 7990 2576
rect 9861 2567 9919 2573
rect 9861 2533 9873 2567
rect 9907 2564 9919 2567
rect 11238 2564 11244 2576
rect 9907 2536 11244 2564
rect 9907 2533 9919 2536
rect 9861 2527 9919 2533
rect 11238 2524 11244 2536
rect 11296 2524 11302 2576
rect 12437 2567 12495 2573
rect 12437 2533 12449 2567
rect 12483 2564 12495 2567
rect 14734 2564 14740 2576
rect 12483 2536 14740 2564
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 14734 2524 14740 2536
rect 14792 2524 14798 2576
rect 31938 2564 31944 2576
rect 28828 2536 31944 2564
rect 4709 2499 4767 2505
rect 4709 2465 4721 2499
rect 4755 2496 4767 2499
rect 5442 2496 5448 2508
rect 4755 2468 5448 2496
rect 4755 2465 4767 2468
rect 4709 2459 4767 2465
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 10134 2496 10140 2508
rect 8619 2468 10140 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2496 11207 2499
rect 12526 2496 12532 2508
rect 11195 2468 12532 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 12526 2456 12532 2468
rect 12584 2456 12590 2508
rect 13081 2499 13139 2505
rect 13081 2465 13093 2499
rect 13127 2496 13139 2499
rect 15470 2496 15476 2508
rect 13127 2468 15476 2496
rect 13127 2465 13139 2468
rect 13081 2459 13139 2465
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 16758 2456 16764 2508
rect 16816 2496 16822 2508
rect 17221 2499 17279 2505
rect 17221 2496 17233 2499
rect 16816 2468 17233 2496
rect 16816 2456 16822 2468
rect 17221 2465 17233 2468
rect 17267 2465 17279 2499
rect 17221 2459 17279 2465
rect 17862 2456 17868 2508
rect 17920 2496 17926 2508
rect 19797 2499 19855 2505
rect 19797 2496 19809 2499
rect 17920 2468 19809 2496
rect 17920 2456 17926 2468
rect 19797 2465 19809 2468
rect 19843 2465 19855 2499
rect 19797 2459 19855 2465
rect 21453 2499 21511 2505
rect 21453 2465 21465 2499
rect 21499 2496 21511 2499
rect 22738 2496 22744 2508
rect 21499 2468 22744 2496
rect 21499 2465 21511 2468
rect 21453 2459 21511 2465
rect 22738 2456 22744 2468
rect 22796 2456 22802 2508
rect 25774 2496 25780 2508
rect 25735 2468 25780 2496
rect 25774 2456 25780 2468
rect 25832 2456 25838 2508
rect 26418 2496 26424 2508
rect 26379 2468 26424 2496
rect 26418 2456 26424 2468
rect 26476 2456 26482 2508
rect 26605 2499 26663 2505
rect 26605 2465 26617 2499
rect 26651 2496 26663 2499
rect 26694 2496 26700 2508
rect 26651 2468 26700 2496
rect 26651 2465 26663 2468
rect 26605 2459 26663 2465
rect 26694 2456 26700 2468
rect 26752 2456 26758 2508
rect 28828 2505 28856 2536
rect 31938 2524 31944 2536
rect 31996 2524 32002 2576
rect 38194 2524 38200 2576
rect 38252 2564 38258 2576
rect 40037 2567 40095 2573
rect 40037 2564 40049 2567
rect 38252 2536 40049 2564
rect 38252 2524 38258 2536
rect 40037 2533 40049 2536
rect 40083 2533 40095 2567
rect 40037 2527 40095 2533
rect 42058 2524 42064 2576
rect 42116 2564 42122 2576
rect 43901 2567 43959 2573
rect 43901 2564 43913 2567
rect 42116 2536 43913 2564
rect 42116 2524 42122 2536
rect 43901 2533 43913 2536
rect 43947 2533 43959 2567
rect 43901 2527 43959 2533
rect 44818 2524 44824 2576
rect 44876 2564 44882 2576
rect 46477 2567 46535 2573
rect 46477 2564 46489 2567
rect 44876 2536 46489 2564
rect 44876 2524 44882 2536
rect 46477 2533 46489 2536
rect 46523 2533 46535 2567
rect 46477 2527 46535 2533
rect 28813 2499 28871 2505
rect 28813 2465 28825 2499
rect 28859 2465 28871 2499
rect 28813 2459 28871 2465
rect 28997 2499 29055 2505
rect 28997 2465 29009 2499
rect 29043 2496 29055 2499
rect 30374 2496 30380 2508
rect 29043 2468 30380 2496
rect 29043 2465 29055 2468
rect 28997 2459 29055 2465
rect 30374 2456 30380 2468
rect 30432 2456 30438 2508
rect 31573 2499 31631 2505
rect 31573 2465 31585 2499
rect 31619 2496 31631 2499
rect 32674 2496 32680 2508
rect 31619 2468 32680 2496
rect 31619 2465 31631 2468
rect 31573 2459 31631 2465
rect 32674 2456 32680 2468
rect 32732 2456 32738 2508
rect 37090 2456 37096 2508
rect 37148 2496 37154 2508
rect 38749 2499 38807 2505
rect 38749 2496 38761 2499
rect 37148 2468 38761 2496
rect 37148 2456 37154 2468
rect 38749 2465 38761 2468
rect 38795 2465 38807 2499
rect 38749 2459 38807 2465
rect 39022 2456 39028 2508
rect 39080 2496 39086 2508
rect 40681 2499 40739 2505
rect 40681 2496 40693 2499
rect 39080 2468 40693 2496
rect 39080 2456 39086 2468
rect 40681 2465 40693 2468
rect 40727 2465 40739 2499
rect 40681 2459 40739 2465
rect 40954 2456 40960 2508
rect 41012 2496 41018 2508
rect 42613 2499 42671 2505
rect 42613 2496 42625 2499
rect 41012 2468 42625 2496
rect 41012 2456 41018 2468
rect 42613 2465 42625 2468
rect 42659 2465 42671 2499
rect 42613 2459 42671 2465
rect 43438 2456 43444 2508
rect 43496 2496 43502 2508
rect 45189 2499 45247 2505
rect 45189 2496 45201 2499
rect 43496 2468 45201 2496
rect 43496 2456 43502 2468
rect 45189 2465 45201 2468
rect 45235 2465 45247 2499
rect 45189 2459 45247 2465
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2590 2428 2596 2440
rect 2179 2400 2596 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 3142 2428 3148 2440
rect 2823 2400 3148 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 3142 2388 3148 2400
rect 3200 2388 3206 2440
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 3878 2428 3884 2440
rect 3467 2400 3884 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 3878 2388 3884 2400
rect 3936 2388 3942 2440
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 7098 2428 7104 2440
rect 6043 2400 7104 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 12066 2428 12072 2440
rect 10551 2400 12072 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 7944 2360 7972 2391
rect 12066 2388 12072 2400
rect 12124 2388 12130 2440
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2428 15071 2431
rect 15562 2428 15568 2440
rect 15059 2400 15568 2428
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2397 15715 2431
rect 15657 2391 15715 2397
rect 16301 2431 16359 2437
rect 16301 2397 16313 2431
rect 16347 2428 16359 2431
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 16347 2400 17049 2428
rect 16347 2397 16359 2400
rect 16301 2391 16359 2397
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 9306 2360 9312 2372
rect 7944 2332 9312 2360
rect 9306 2320 9312 2332
rect 9364 2320 9370 2372
rect 15672 2292 15700 2391
rect 19242 2388 19248 2440
rect 19300 2428 19306 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19300 2400 19625 2428
rect 19300 2388 19306 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 22094 2388 22100 2440
rect 22152 2428 22158 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 22152 2400 22201 2428
rect 22152 2388 22158 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 32122 2388 32128 2440
rect 32180 2428 32186 2440
rect 32493 2431 32551 2437
rect 32493 2428 32505 2431
rect 32180 2400 32505 2428
rect 32180 2388 32186 2400
rect 32493 2397 32505 2400
rect 32539 2428 32551 2431
rect 32953 2431 33011 2437
rect 32953 2428 32965 2431
rect 32539 2400 32965 2428
rect 32539 2397 32551 2400
rect 32493 2391 32551 2397
rect 32953 2397 32965 2400
rect 32999 2397 33011 2431
rect 32953 2391 33011 2397
rect 35529 2431 35587 2437
rect 35529 2397 35541 2431
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 18877 2363 18935 2369
rect 18877 2329 18889 2363
rect 18923 2329 18935 2363
rect 18877 2323 18935 2329
rect 18782 2292 18788 2304
rect 15672 2264 18788 2292
rect 18782 2252 18788 2264
rect 18840 2252 18846 2304
rect 18892 2292 18920 2323
rect 20622 2320 20628 2372
rect 20680 2360 20686 2372
rect 22373 2363 22431 2369
rect 22373 2360 22385 2363
rect 20680 2332 22385 2360
rect 20680 2320 20686 2332
rect 22373 2329 22385 2332
rect 22419 2329 22431 2363
rect 22373 2323 22431 2329
rect 24029 2363 24087 2369
rect 24029 2329 24041 2363
rect 24075 2360 24087 2363
rect 24118 2360 24124 2372
rect 24075 2332 24124 2360
rect 24075 2329 24087 2332
rect 24029 2323 24087 2329
rect 24118 2320 24124 2332
rect 24176 2320 24182 2372
rect 27154 2360 27160 2372
rect 27115 2332 27160 2360
rect 27154 2320 27160 2332
rect 27212 2320 27218 2372
rect 29362 2320 29368 2372
rect 29420 2360 29426 2372
rect 29733 2363 29791 2369
rect 29733 2360 29745 2363
rect 29420 2332 29745 2360
rect 29420 2320 29426 2332
rect 29733 2329 29745 2332
rect 29779 2329 29791 2363
rect 29733 2323 29791 2329
rect 31389 2363 31447 2369
rect 31389 2329 31401 2363
rect 31435 2360 31447 2363
rect 31846 2360 31852 2372
rect 31435 2332 31852 2360
rect 31435 2329 31447 2332
rect 31389 2323 31447 2329
rect 31846 2320 31852 2332
rect 31904 2320 31910 2372
rect 31938 2320 31944 2372
rect 31996 2360 32002 2372
rect 35544 2360 35572 2391
rect 36262 2388 36268 2440
rect 36320 2428 36326 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 36320 2400 38117 2428
rect 36320 2388 36326 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 39574 2388 39580 2440
rect 39632 2428 39638 2440
rect 41325 2431 41383 2437
rect 41325 2428 41337 2431
rect 39632 2400 41337 2428
rect 39632 2388 39638 2400
rect 41325 2397 41337 2400
rect 41371 2397 41383 2431
rect 41325 2391 41383 2397
rect 41506 2388 41512 2440
rect 41564 2428 41570 2440
rect 43257 2431 43315 2437
rect 43257 2428 43269 2431
rect 41564 2400 43269 2428
rect 41564 2388 41570 2400
rect 43257 2397 43269 2400
rect 43303 2397 43315 2431
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 43257 2391 43315 2397
rect 45526 2400 45845 2428
rect 31996 2332 35572 2360
rect 31996 2320 32002 2332
rect 43990 2320 43996 2372
rect 44048 2360 44054 2372
rect 45526 2360 45554 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 45922 2388 45928 2440
rect 45980 2428 45986 2440
rect 47765 2431 47823 2437
rect 47765 2428 47777 2431
rect 45980 2400 47777 2428
rect 45980 2388 45986 2400
rect 47765 2397 47777 2400
rect 47811 2397 47823 2431
rect 47765 2391 47823 2397
rect 44048 2332 45554 2360
rect 44048 2320 44054 2332
rect 21910 2292 21916 2304
rect 18892 2264 21916 2292
rect 21910 2252 21916 2264
rect 21968 2252 21974 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 18782 2048 18788 2100
rect 18840 2088 18846 2100
rect 20806 2088 20812 2100
rect 18840 2060 20812 2088
rect 18840 2048 18846 2060
rect 20806 2048 20812 2060
rect 20864 2048 20870 2100
rect 15562 1980 15568 2032
rect 15620 2020 15626 2032
rect 20254 2020 20260 2032
rect 15620 1992 20260 2020
rect 15620 1980 15626 1992
rect 20254 1980 20260 1992
rect 20312 1980 20318 2032
rect 19058 1912 19064 1964
rect 19116 1952 19122 1964
rect 19702 1952 19708 1964
rect 19116 1924 19708 1952
rect 19116 1912 19122 1924
rect 19702 1912 19708 1924
rect 19760 1912 19766 1964
<< via1 >>
rect 10968 47812 11020 47864
rect 20720 47812 20772 47864
rect 15384 47744 15436 47796
rect 23388 47744 23440 47796
rect 18880 47608 18932 47660
rect 20904 47608 20956 47660
rect 23664 47608 23716 47660
rect 25688 47608 25740 47660
rect 14556 47540 14608 47592
rect 20352 47540 20404 47592
rect 13176 47472 13228 47524
rect 21456 47472 21508 47524
rect 23756 47472 23808 47524
rect 30288 47472 30340 47524
rect 37832 47472 37884 47524
rect 38384 47472 38436 47524
rect 11704 47404 11756 47456
rect 17776 47404 17828 47456
rect 18144 47404 18196 47456
rect 24032 47404 24084 47456
rect 29828 47404 29880 47456
rect 30012 47404 30064 47456
rect 43444 47404 43496 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 5080 47200 5132 47252
rect 7288 47243 7340 47252
rect 7288 47209 7297 47243
rect 7297 47209 7331 47243
rect 7331 47209 7340 47243
rect 7288 47200 7340 47209
rect 7932 47243 7984 47252
rect 7932 47209 7941 47243
rect 7941 47209 7975 47243
rect 7975 47209 7984 47243
rect 7932 47200 7984 47209
rect 8392 47243 8444 47252
rect 8392 47209 8401 47243
rect 8401 47209 8435 47243
rect 8435 47209 8444 47243
rect 8392 47200 8444 47209
rect 9680 47243 9732 47252
rect 9680 47209 9689 47243
rect 9689 47209 9723 47243
rect 9723 47209 9732 47243
rect 9680 47200 9732 47209
rect 10784 47243 10836 47252
rect 10784 47209 10793 47243
rect 10793 47209 10827 47243
rect 10827 47209 10836 47243
rect 10784 47200 10836 47209
rect 11888 47243 11940 47252
rect 11888 47209 11897 47243
rect 11897 47209 11931 47243
rect 11931 47209 11940 47243
rect 11888 47200 11940 47209
rect 12992 47243 13044 47252
rect 12992 47209 13001 47243
rect 13001 47209 13035 47243
rect 13035 47209 13044 47243
rect 12992 47200 13044 47209
rect 13912 47200 13964 47252
rect 15200 47243 15252 47252
rect 15200 47209 15209 47243
rect 15209 47209 15243 47243
rect 15243 47209 15252 47243
rect 15200 47200 15252 47209
rect 16120 47243 16172 47252
rect 16120 47209 16129 47243
rect 16129 47209 16163 47243
rect 16163 47209 16172 47243
rect 16120 47200 16172 47209
rect 17224 47243 17276 47252
rect 17224 47209 17233 47243
rect 17233 47209 17267 47243
rect 17267 47209 17276 47243
rect 17224 47200 17276 47209
rect 19432 47200 19484 47252
rect 22744 47200 22796 47252
rect 23388 47243 23440 47252
rect 23388 47209 23397 47243
rect 23397 47209 23431 47243
rect 23431 47209 23440 47243
rect 23388 47200 23440 47209
rect 23848 47200 23900 47252
rect 26056 47200 26108 47252
rect 35440 47200 35492 47252
rect 43444 47243 43496 47252
rect 43444 47209 43453 47243
rect 43453 47209 43487 47243
rect 43487 47209 43496 47243
rect 43444 47200 43496 47209
rect 44272 47243 44324 47252
rect 44272 47209 44281 47243
rect 44281 47209 44315 47243
rect 44315 47209 44324 47243
rect 44272 47200 44324 47209
rect 45928 47200 45980 47252
rect 4068 47107 4120 47116
rect 4068 47073 4077 47107
rect 4077 47073 4111 47107
rect 4111 47073 4120 47107
rect 4068 47064 4120 47073
rect 11704 47064 11756 47116
rect 5632 47039 5684 47048
rect 5632 47005 5641 47039
rect 5641 47005 5675 47039
rect 5675 47005 5684 47039
rect 5632 46996 5684 47005
rect 9864 47039 9916 47048
rect 9864 47005 9873 47039
rect 9873 47005 9907 47039
rect 9907 47005 9916 47039
rect 9864 46996 9916 47005
rect 10968 47039 11020 47048
rect 10968 47005 10977 47039
rect 10977 47005 11011 47039
rect 11011 47005 11020 47039
rect 10968 46996 11020 47005
rect 13176 47039 13228 47048
rect 13176 47005 13185 47039
rect 13185 47005 13219 47039
rect 13219 47005 13228 47039
rect 13176 46996 13228 47005
rect 14556 47039 14608 47048
rect 14556 47005 14565 47039
rect 14565 47005 14599 47039
rect 14599 47005 14608 47039
rect 14556 46996 14608 47005
rect 15384 47039 15436 47048
rect 15384 47005 15393 47039
rect 15393 47005 15427 47039
rect 15427 47005 15436 47039
rect 15384 46996 15436 47005
rect 18052 47064 18104 47116
rect 18144 47039 18196 47048
rect 18144 47005 18153 47039
rect 18153 47005 18187 47039
rect 18187 47005 18196 47039
rect 18144 46996 18196 47005
rect 18328 47064 18380 47116
rect 18880 47039 18932 47048
rect 18880 47005 18889 47039
rect 18889 47005 18923 47039
rect 18923 47005 18932 47039
rect 18880 46996 18932 47005
rect 19340 47064 19392 47116
rect 26792 47132 26844 47184
rect 35992 47132 36044 47184
rect 21640 47064 21692 47116
rect 23204 47064 23256 47116
rect 23848 47107 23900 47116
rect 23848 47073 23857 47107
rect 23857 47073 23891 47107
rect 23891 47073 23900 47107
rect 23848 47064 23900 47073
rect 20260 46996 20312 47048
rect 21088 46996 21140 47048
rect 18696 46860 18748 46912
rect 19432 46860 19484 46912
rect 20444 46928 20496 46980
rect 22100 46996 22152 47048
rect 23296 46996 23348 47048
rect 23572 47039 23624 47048
rect 23572 47005 23581 47039
rect 23581 47005 23615 47039
rect 23615 47005 23624 47039
rect 23572 46996 23624 47005
rect 23756 47039 23808 47048
rect 23756 47005 23765 47039
rect 23765 47005 23799 47039
rect 23799 47005 23808 47039
rect 23756 46996 23808 47005
rect 24032 47039 24084 47048
rect 24032 47005 24041 47039
rect 24041 47005 24075 47039
rect 24075 47005 24084 47039
rect 24032 46996 24084 47005
rect 31760 47064 31812 47116
rect 31944 47064 31996 47116
rect 33232 47064 33284 47116
rect 33968 47107 34020 47116
rect 33968 47073 33977 47107
rect 33977 47073 34011 47107
rect 34011 47073 34020 47107
rect 33968 47064 34020 47073
rect 34152 47064 34204 47116
rect 37556 47064 37608 47116
rect 37832 47107 37884 47116
rect 37832 47073 37841 47107
rect 37841 47073 37875 47107
rect 37875 47073 37884 47107
rect 37832 47064 37884 47073
rect 25688 47039 25740 47048
rect 25688 47005 25697 47039
rect 25697 47005 25731 47039
rect 25731 47005 25740 47039
rect 25688 46996 25740 47005
rect 25872 47039 25924 47048
rect 25872 47005 25881 47039
rect 25881 47005 25915 47039
rect 25915 47005 25924 47039
rect 25872 46996 25924 47005
rect 26148 46996 26200 47048
rect 26424 46996 26476 47048
rect 27160 47039 27212 47048
rect 27160 47005 27169 47039
rect 27169 47005 27203 47039
rect 27203 47005 27212 47039
rect 27160 46996 27212 47005
rect 27620 46996 27672 47048
rect 29368 46996 29420 47048
rect 29736 46996 29788 47048
rect 29920 46996 29972 47048
rect 32220 46996 32272 47048
rect 33784 47039 33836 47048
rect 33784 47005 33793 47039
rect 33793 47005 33827 47039
rect 33827 47005 33836 47039
rect 33784 46996 33836 47005
rect 36084 46996 36136 47048
rect 37648 47039 37700 47048
rect 21916 46860 21968 46912
rect 24676 46928 24728 46980
rect 29184 46971 29236 46980
rect 22928 46860 22980 46912
rect 25504 46903 25556 46912
rect 25504 46869 25513 46903
rect 25513 46869 25547 46903
rect 25547 46869 25556 46903
rect 25504 46860 25556 46869
rect 29184 46937 29193 46971
rect 29193 46937 29227 46971
rect 29227 46937 29236 46971
rect 29184 46928 29236 46937
rect 31668 46928 31720 46980
rect 31852 46928 31904 46980
rect 30840 46860 30892 46912
rect 32220 46860 32272 46912
rect 33324 46860 33376 46912
rect 35348 46860 35400 46912
rect 37648 47005 37657 47039
rect 37657 47005 37691 47039
rect 37691 47005 37700 47039
rect 37648 46996 37700 47005
rect 37280 46928 37332 46980
rect 37372 46928 37424 46980
rect 40040 47107 40092 47116
rect 40040 47073 40049 47107
rect 40049 47073 40083 47107
rect 40083 47073 40092 47107
rect 40040 47064 40092 47073
rect 41604 47064 41656 47116
rect 38844 46996 38896 47048
rect 40224 46996 40276 47048
rect 41972 46971 42024 46980
rect 41972 46937 41981 46971
rect 41981 46937 42015 46971
rect 42015 46937 42024 46971
rect 41972 46928 42024 46937
rect 42984 46996 43036 47048
rect 43812 46996 43864 47048
rect 44180 46996 44232 47048
rect 45192 46996 45244 47048
rect 36636 46860 36688 46912
rect 36912 46860 36964 46912
rect 37464 46903 37516 46912
rect 37464 46869 37473 46903
rect 37473 46869 37507 46903
rect 37507 46869 37516 46903
rect 37464 46860 37516 46869
rect 38660 46860 38712 46912
rect 42156 46860 42208 46912
rect 43260 46928 43312 46980
rect 44824 46860 44876 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 4068 46656 4120 46708
rect 18420 46699 18472 46708
rect 18420 46665 18429 46699
rect 18429 46665 18463 46699
rect 18463 46665 18472 46699
rect 18420 46656 18472 46665
rect 20536 46656 20588 46708
rect 22100 46656 22152 46708
rect 23848 46699 23900 46708
rect 23848 46665 23857 46699
rect 23857 46665 23891 46699
rect 23891 46665 23900 46699
rect 23848 46656 23900 46665
rect 25688 46656 25740 46708
rect 25964 46656 26016 46708
rect 30104 46656 30156 46708
rect 4804 46563 4856 46572
rect 4804 46529 4813 46563
rect 4813 46529 4847 46563
rect 4847 46529 4856 46563
rect 4804 46520 4856 46529
rect 6000 46563 6052 46572
rect 6000 46529 6009 46563
rect 6009 46529 6043 46563
rect 6043 46529 6052 46563
rect 6000 46520 6052 46529
rect 5632 46452 5684 46504
rect 7012 46563 7064 46572
rect 7012 46529 7021 46563
rect 7021 46529 7055 46563
rect 7055 46529 7064 46563
rect 7012 46520 7064 46529
rect 9220 46563 9272 46572
rect 9220 46529 9229 46563
rect 9229 46529 9263 46563
rect 9263 46529 9272 46563
rect 9220 46520 9272 46529
rect 10324 46563 10376 46572
rect 10324 46529 10333 46563
rect 10333 46529 10367 46563
rect 10367 46529 10376 46563
rect 10324 46520 10376 46529
rect 11336 46520 11388 46572
rect 12532 46563 12584 46572
rect 12532 46529 12541 46563
rect 12541 46529 12575 46563
rect 12575 46529 12584 46563
rect 12532 46520 12584 46529
rect 13636 46563 13688 46572
rect 13636 46529 13645 46563
rect 13645 46529 13679 46563
rect 13679 46529 13688 46563
rect 13636 46520 13688 46529
rect 14740 46563 14792 46572
rect 14740 46529 14749 46563
rect 14749 46529 14783 46563
rect 14783 46529 14792 46563
rect 14740 46520 14792 46529
rect 15844 46563 15896 46572
rect 15844 46529 15853 46563
rect 15853 46529 15887 46563
rect 15887 46529 15896 46563
rect 15844 46520 15896 46529
rect 17960 46520 18012 46572
rect 19340 46563 19392 46572
rect 19340 46529 19349 46563
rect 19349 46529 19383 46563
rect 19383 46529 19392 46563
rect 19340 46520 19392 46529
rect 20260 46520 20312 46572
rect 20720 46520 20772 46572
rect 19524 46452 19576 46504
rect 19800 46495 19852 46504
rect 19800 46461 19809 46495
rect 19809 46461 19843 46495
rect 19843 46461 19852 46495
rect 19800 46452 19852 46461
rect 18696 46384 18748 46436
rect 21548 46520 21600 46572
rect 22284 46520 22336 46572
rect 22836 46588 22888 46640
rect 23296 46588 23348 46640
rect 24860 46588 24912 46640
rect 25228 46631 25280 46640
rect 25228 46597 25237 46631
rect 25237 46597 25271 46631
rect 25271 46597 25280 46631
rect 25228 46588 25280 46597
rect 22744 46563 22796 46572
rect 22744 46529 22753 46563
rect 22753 46529 22787 46563
rect 22787 46529 22796 46563
rect 22744 46520 22796 46529
rect 23664 46520 23716 46572
rect 24032 46563 24084 46572
rect 24032 46529 24041 46563
rect 24041 46529 24075 46563
rect 24075 46529 24084 46563
rect 24032 46520 24084 46529
rect 24216 46563 24268 46572
rect 24216 46529 24225 46563
rect 24225 46529 24259 46563
rect 24259 46529 24268 46563
rect 24216 46520 24268 46529
rect 24492 46520 24544 46572
rect 24676 46520 24728 46572
rect 24768 46520 24820 46572
rect 28080 46588 28132 46640
rect 29092 46588 29144 46640
rect 25872 46520 25924 46572
rect 26148 46520 26200 46572
rect 22928 46452 22980 46504
rect 23020 46452 23072 46504
rect 24308 46495 24360 46504
rect 24308 46461 24317 46495
rect 24317 46461 24351 46495
rect 24351 46461 24360 46495
rect 24308 46452 24360 46461
rect 20260 46384 20312 46436
rect 24952 46384 25004 46436
rect 25228 46452 25280 46504
rect 27068 46520 27120 46572
rect 26424 46495 26476 46504
rect 26424 46461 26433 46495
rect 26433 46461 26467 46495
rect 26467 46461 26476 46495
rect 26424 46452 26476 46461
rect 28172 46520 28224 46572
rect 28448 46563 28500 46572
rect 28448 46529 28457 46563
rect 28457 46529 28491 46563
rect 28491 46529 28500 46563
rect 28448 46520 28500 46529
rect 28540 46563 28592 46572
rect 28540 46529 28549 46563
rect 28549 46529 28583 46563
rect 28583 46529 28592 46563
rect 29368 46563 29420 46572
rect 28540 46520 28592 46529
rect 29368 46529 29377 46563
rect 29377 46529 29411 46563
rect 29411 46529 29420 46563
rect 29368 46520 29420 46529
rect 29828 46588 29880 46640
rect 30656 46563 30708 46572
rect 29184 46495 29236 46504
rect 29184 46461 29193 46495
rect 29193 46461 29227 46495
rect 29227 46461 29236 46495
rect 29184 46452 29236 46461
rect 30656 46529 30665 46563
rect 30665 46529 30699 46563
rect 30699 46529 30708 46563
rect 30656 46520 30708 46529
rect 30748 46520 30800 46572
rect 31852 46588 31904 46640
rect 33784 46656 33836 46708
rect 34060 46656 34112 46708
rect 34796 46656 34848 46708
rect 33784 46520 33836 46572
rect 34152 46563 34204 46572
rect 34152 46529 34158 46563
rect 34158 46529 34192 46563
rect 34192 46529 34204 46563
rect 34152 46520 34204 46529
rect 37372 46588 37424 46640
rect 31668 46452 31720 46504
rect 31852 46452 31904 46504
rect 32036 46452 32088 46504
rect 32588 46495 32640 46504
rect 32588 46461 32597 46495
rect 32597 46461 32631 46495
rect 32631 46461 32640 46495
rect 32588 46452 32640 46461
rect 33508 46452 33560 46504
rect 35532 46452 35584 46504
rect 36268 46520 36320 46572
rect 36452 46495 36504 46504
rect 36452 46461 36461 46495
rect 36461 46461 36495 46495
rect 36495 46461 36504 46495
rect 36452 46452 36504 46461
rect 37464 46520 37516 46572
rect 38108 46520 38160 46572
rect 38476 46452 38528 46504
rect 38844 46520 38896 46572
rect 39120 46563 39172 46572
rect 39120 46529 39129 46563
rect 39129 46529 39163 46563
rect 39163 46529 39172 46563
rect 39120 46520 39172 46529
rect 40868 46563 40920 46572
rect 40868 46529 40877 46563
rect 40877 46529 40911 46563
rect 40911 46529 40920 46563
rect 40868 46520 40920 46529
rect 42616 46520 42668 46572
rect 43352 46520 43404 46572
rect 44456 46520 44508 46572
rect 45836 46563 45888 46572
rect 45836 46529 45845 46563
rect 45845 46529 45879 46563
rect 45879 46529 45888 46563
rect 45836 46520 45888 46529
rect 43720 46452 43772 46504
rect 18788 46316 18840 46368
rect 20076 46316 20128 46368
rect 20904 46359 20956 46368
rect 20904 46325 20913 46359
rect 20913 46325 20947 46359
rect 20947 46325 20956 46359
rect 20904 46316 20956 46325
rect 21456 46359 21508 46368
rect 21456 46325 21465 46359
rect 21465 46325 21499 46359
rect 21499 46325 21508 46359
rect 21456 46316 21508 46325
rect 23756 46316 23808 46368
rect 25136 46316 25188 46368
rect 30472 46384 30524 46436
rect 37096 46384 37148 46436
rect 38752 46384 38804 46436
rect 41512 46384 41564 46436
rect 27344 46316 27396 46368
rect 27804 46316 27856 46368
rect 31852 46316 31904 46368
rect 32036 46316 32088 46368
rect 34336 46316 34388 46368
rect 34796 46316 34848 46368
rect 35532 46316 35584 46368
rect 35992 46316 36044 46368
rect 37556 46316 37608 46368
rect 37924 46316 37976 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 5908 46155 5960 46164
rect 5908 46121 5917 46155
rect 5917 46121 5951 46155
rect 5951 46121 5960 46155
rect 5908 46112 5960 46121
rect 16948 46155 17000 46164
rect 16948 46121 16957 46155
rect 16957 46121 16991 46155
rect 16991 46121 17000 46155
rect 16948 46112 17000 46121
rect 18052 46155 18104 46164
rect 18052 46121 18061 46155
rect 18061 46121 18095 46155
rect 18095 46121 18104 46155
rect 18052 46112 18104 46121
rect 18696 46155 18748 46164
rect 18696 46121 18705 46155
rect 18705 46121 18739 46155
rect 18739 46121 18748 46155
rect 18696 46112 18748 46121
rect 18788 46112 18840 46164
rect 21272 46112 21324 46164
rect 22744 46155 22796 46164
rect 22744 46121 22753 46155
rect 22753 46121 22787 46155
rect 22787 46121 22796 46155
rect 22744 46112 22796 46121
rect 22836 46112 22888 46164
rect 24952 46155 25004 46164
rect 20720 46044 20772 46096
rect 22652 46044 22704 46096
rect 23940 46044 23992 46096
rect 24952 46121 24961 46155
rect 24961 46121 24995 46155
rect 24995 46121 25004 46155
rect 24952 46112 25004 46121
rect 27344 46112 27396 46164
rect 28540 46112 28592 46164
rect 25136 46044 25188 46096
rect 25228 46044 25280 46096
rect 20444 45976 20496 46028
rect 19800 45951 19852 45960
rect 19800 45917 19809 45951
rect 19809 45917 19843 45951
rect 19843 45917 19852 45951
rect 19800 45908 19852 45917
rect 19984 45951 20036 45960
rect 19984 45917 19993 45951
rect 19993 45917 20027 45951
rect 20027 45917 20036 45951
rect 23112 45976 23164 46028
rect 23664 46019 23716 46028
rect 23664 45985 23673 46019
rect 23673 45985 23707 46019
rect 23707 45985 23716 46019
rect 23664 45976 23716 45985
rect 19984 45908 20036 45917
rect 21364 45951 21416 45960
rect 21364 45917 21373 45951
rect 21373 45917 21407 45951
rect 21407 45917 21416 45951
rect 21364 45908 21416 45917
rect 21548 45951 21600 45960
rect 21548 45917 21557 45951
rect 21557 45917 21591 45951
rect 21591 45917 21600 45951
rect 24768 45976 24820 46028
rect 25872 46044 25924 46096
rect 21548 45908 21600 45917
rect 9864 45772 9916 45824
rect 20260 45772 20312 45824
rect 22560 45840 22612 45892
rect 23112 45883 23164 45892
rect 23112 45849 23121 45883
rect 23121 45849 23155 45883
rect 23155 45849 23164 45883
rect 23112 45840 23164 45849
rect 25504 45976 25556 46028
rect 25136 45951 25188 45960
rect 25136 45917 25145 45951
rect 25145 45917 25179 45951
rect 25179 45917 25188 45951
rect 25136 45908 25188 45917
rect 26056 45908 26108 45960
rect 26700 45951 26752 45960
rect 26700 45917 26709 45951
rect 26709 45917 26743 45951
rect 26743 45917 26752 45951
rect 26700 45908 26752 45917
rect 26792 45951 26844 45960
rect 26792 45917 26801 45951
rect 26801 45917 26835 45951
rect 26835 45917 26844 45951
rect 28172 46044 28224 46096
rect 28448 46044 28500 46096
rect 29184 46112 29236 46164
rect 28724 46019 28776 46028
rect 28724 45985 28733 46019
rect 28733 45985 28767 46019
rect 28767 45985 28776 46019
rect 28724 45976 28776 45985
rect 29828 46044 29880 46096
rect 30288 46087 30340 46096
rect 30288 46053 30297 46087
rect 30297 46053 30331 46087
rect 30331 46053 30340 46087
rect 30288 46044 30340 46053
rect 32588 46112 32640 46164
rect 31760 46044 31812 46096
rect 32036 46044 32088 46096
rect 32956 46087 33008 46096
rect 32956 46053 32965 46087
rect 32965 46053 32999 46087
rect 32999 46053 33008 46087
rect 32956 46044 33008 46053
rect 32128 45976 32180 46028
rect 37924 46112 37976 46164
rect 38108 46155 38160 46164
rect 38108 46121 38117 46155
rect 38117 46121 38151 46155
rect 38151 46121 38160 46155
rect 38108 46112 38160 46121
rect 38384 46112 38436 46164
rect 33232 46044 33284 46096
rect 33324 46044 33376 46096
rect 33784 46044 33836 46096
rect 34980 46019 35032 46028
rect 34980 45985 34989 46019
rect 34989 45985 35023 46019
rect 35023 45985 35032 46019
rect 34980 45976 35032 45985
rect 35440 45976 35492 46028
rect 35532 45976 35584 46028
rect 26792 45908 26844 45917
rect 21548 45772 21600 45824
rect 21732 45815 21784 45824
rect 21732 45781 21741 45815
rect 21741 45781 21775 45815
rect 21775 45781 21784 45815
rect 21732 45772 21784 45781
rect 24032 45772 24084 45824
rect 27344 45772 27396 45824
rect 28356 45908 28408 45960
rect 27988 45840 28040 45892
rect 30012 45908 30064 45960
rect 30472 45951 30524 45960
rect 30472 45917 30481 45951
rect 30481 45917 30515 45951
rect 30515 45917 30524 45951
rect 30472 45908 30524 45917
rect 30748 45951 30800 45960
rect 30748 45917 30757 45951
rect 30757 45917 30791 45951
rect 30791 45917 30800 45951
rect 30748 45908 30800 45917
rect 31760 45951 31812 45960
rect 31760 45917 31769 45951
rect 31769 45917 31803 45951
rect 31803 45917 31812 45951
rect 31760 45908 31812 45917
rect 32956 45908 33008 45960
rect 34060 45908 34112 45960
rect 34520 45908 34572 45960
rect 35808 45976 35860 46028
rect 36544 46019 36596 46028
rect 30656 45883 30708 45892
rect 30656 45849 30665 45883
rect 30665 45849 30699 45883
rect 30699 45849 30708 45883
rect 30656 45840 30708 45849
rect 33508 45840 33560 45892
rect 34612 45840 34664 45892
rect 35716 45951 35768 45960
rect 35716 45917 35725 45951
rect 35725 45917 35759 45951
rect 35759 45917 35768 45951
rect 36544 45985 36553 46019
rect 36553 45985 36587 46019
rect 36587 45985 36596 46019
rect 36544 45976 36596 45985
rect 38292 46044 38344 46096
rect 38476 46087 38528 46096
rect 38476 46053 38485 46087
rect 38485 46053 38519 46087
rect 38519 46053 38528 46087
rect 38476 46044 38528 46053
rect 38568 46044 38620 46096
rect 35716 45908 35768 45917
rect 35992 45951 36044 45960
rect 35992 45917 36001 45951
rect 36001 45917 36035 45951
rect 36035 45917 36044 45951
rect 35992 45908 36044 45917
rect 36452 45908 36504 45960
rect 37372 45908 37424 45960
rect 38016 45908 38068 45960
rect 38936 46112 38988 46164
rect 41144 46112 41196 46164
rect 42248 46112 42300 46164
rect 43260 46155 43312 46164
rect 43260 46121 43269 46155
rect 43269 46121 43303 46155
rect 43303 46121 43312 46155
rect 43260 46112 43312 46121
rect 43812 46155 43864 46164
rect 43812 46121 43821 46155
rect 43821 46121 43855 46155
rect 43855 46121 43864 46155
rect 43812 46112 43864 46121
rect 44180 46112 44232 46164
rect 45192 46155 45244 46164
rect 45192 46121 45201 46155
rect 45201 46121 45235 46155
rect 45235 46121 45244 46155
rect 45192 46112 45244 46121
rect 40316 46044 40368 46096
rect 38844 45908 38896 45960
rect 28724 45772 28776 45824
rect 31392 45772 31444 45824
rect 31944 45772 31996 45824
rect 33968 45815 34020 45824
rect 33968 45781 33977 45815
rect 33977 45781 34011 45815
rect 34011 45781 34020 45815
rect 33968 45772 34020 45781
rect 35716 45772 35768 45824
rect 36728 45840 36780 45892
rect 39212 45840 39264 45892
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 23112 45611 23164 45620
rect 17776 45543 17828 45552
rect 17776 45509 17785 45543
rect 17785 45509 17819 45543
rect 17819 45509 17828 45543
rect 17776 45500 17828 45509
rect 20536 45500 20588 45552
rect 23112 45577 23121 45611
rect 23121 45577 23155 45611
rect 23155 45577 23164 45611
rect 23112 45568 23164 45577
rect 24032 45568 24084 45620
rect 20812 45500 20864 45552
rect 19064 45432 19116 45484
rect 22376 45432 22428 45484
rect 23756 45432 23808 45484
rect 20168 45364 20220 45416
rect 19432 45296 19484 45348
rect 21364 45364 21416 45416
rect 21916 45364 21968 45416
rect 23296 45407 23348 45416
rect 23296 45373 23305 45407
rect 23305 45373 23339 45407
rect 23339 45373 23348 45407
rect 23296 45364 23348 45373
rect 23480 45407 23532 45416
rect 23480 45373 23489 45407
rect 23489 45373 23523 45407
rect 23523 45373 23532 45407
rect 23480 45364 23532 45373
rect 25320 45500 25372 45552
rect 26056 45568 26108 45620
rect 26240 45611 26292 45620
rect 26240 45577 26249 45611
rect 26249 45577 26283 45611
rect 26283 45577 26292 45611
rect 26240 45568 26292 45577
rect 27344 45568 27396 45620
rect 28080 45611 28132 45620
rect 28080 45577 28089 45611
rect 28089 45577 28123 45611
rect 28123 45577 28132 45611
rect 28080 45568 28132 45577
rect 30748 45611 30800 45620
rect 30748 45577 30757 45611
rect 30757 45577 30791 45611
rect 30791 45577 30800 45611
rect 30748 45568 30800 45577
rect 21272 45296 21324 45348
rect 22100 45296 22152 45348
rect 24860 45432 24912 45484
rect 25780 45475 25832 45484
rect 25780 45441 25797 45475
rect 25797 45441 25832 45475
rect 25780 45432 25832 45441
rect 31392 45500 31444 45552
rect 31944 45500 31996 45552
rect 34612 45568 34664 45620
rect 33416 45543 33468 45552
rect 27620 45475 27672 45484
rect 25504 45364 25556 45416
rect 27620 45441 27629 45475
rect 27629 45441 27663 45475
rect 27663 45441 27672 45475
rect 27620 45432 27672 45441
rect 28448 45475 28500 45484
rect 28448 45441 28457 45475
rect 28457 45441 28491 45475
rect 28491 45441 28500 45475
rect 28448 45432 28500 45441
rect 29276 45475 29328 45484
rect 29276 45441 29285 45475
rect 29285 45441 29319 45475
rect 29319 45441 29328 45475
rect 29276 45432 29328 45441
rect 29552 45475 29604 45484
rect 29552 45441 29561 45475
rect 29561 45441 29595 45475
rect 29595 45441 29604 45475
rect 29552 45432 29604 45441
rect 32312 45475 32364 45484
rect 19984 45271 20036 45280
rect 19984 45237 19993 45271
rect 19993 45237 20027 45271
rect 20027 45237 20036 45271
rect 19984 45228 20036 45237
rect 20352 45228 20404 45280
rect 21088 45271 21140 45280
rect 21088 45237 21097 45271
rect 21097 45237 21131 45271
rect 21131 45237 21140 45271
rect 21088 45228 21140 45237
rect 22376 45271 22428 45280
rect 22376 45237 22385 45271
rect 22385 45237 22419 45271
rect 22419 45237 22428 45271
rect 22376 45228 22428 45237
rect 24308 45271 24360 45280
rect 24308 45237 24317 45271
rect 24317 45237 24351 45271
rect 24351 45237 24360 45271
rect 24308 45228 24360 45237
rect 24768 45228 24820 45280
rect 28724 45364 28776 45416
rect 27620 45296 27672 45348
rect 28356 45296 28408 45348
rect 28632 45296 28684 45348
rect 29920 45364 29972 45416
rect 30472 45407 30524 45416
rect 30472 45373 30481 45407
rect 30481 45373 30515 45407
rect 30515 45373 30524 45407
rect 30472 45364 30524 45373
rect 32312 45441 32321 45475
rect 32321 45441 32355 45475
rect 32355 45441 32364 45475
rect 32312 45432 32364 45441
rect 32588 45475 32640 45484
rect 31852 45296 31904 45348
rect 32588 45441 32597 45475
rect 32597 45441 32631 45475
rect 32631 45441 32640 45475
rect 32588 45432 32640 45441
rect 33416 45509 33425 45543
rect 33425 45509 33459 45543
rect 33459 45509 33468 45543
rect 33416 45500 33468 45509
rect 33784 45543 33836 45552
rect 32956 45432 33008 45484
rect 33784 45509 33793 45543
rect 33793 45509 33827 45543
rect 33827 45509 33836 45543
rect 33784 45500 33836 45509
rect 33968 45500 34020 45552
rect 34336 45500 34388 45552
rect 35532 45568 35584 45620
rect 36268 45568 36320 45620
rect 36360 45568 36412 45620
rect 38108 45568 38160 45620
rect 38200 45568 38252 45620
rect 35716 45500 35768 45552
rect 35440 45475 35492 45484
rect 33600 45296 33652 45348
rect 35440 45441 35449 45475
rect 35449 45441 35483 45475
rect 35483 45441 35492 45475
rect 35440 45432 35492 45441
rect 35808 45432 35860 45484
rect 35992 45475 36044 45484
rect 35992 45441 36001 45475
rect 36001 45441 36035 45475
rect 36035 45441 36044 45475
rect 35992 45432 36044 45441
rect 36176 45432 36228 45484
rect 37372 45432 37424 45484
rect 38568 45500 38620 45552
rect 34060 45407 34112 45416
rect 34060 45373 34069 45407
rect 34069 45373 34103 45407
rect 34103 45373 34112 45407
rect 34060 45364 34112 45373
rect 37464 45407 37516 45416
rect 37464 45373 37473 45407
rect 37473 45373 37507 45407
rect 37507 45373 37516 45407
rect 37464 45364 37516 45373
rect 37556 45364 37608 45416
rect 39304 45568 39356 45620
rect 39212 45407 39264 45416
rect 36544 45296 36596 45348
rect 39212 45373 39221 45407
rect 39221 45373 39255 45407
rect 39255 45373 39264 45407
rect 39212 45364 39264 45373
rect 40408 45432 40460 45484
rect 41604 45364 41656 45416
rect 29460 45228 29512 45280
rect 31760 45228 31812 45280
rect 35348 45228 35400 45280
rect 35716 45228 35768 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19340 45024 19392 45076
rect 22560 45067 22612 45076
rect 22560 45033 22569 45067
rect 22569 45033 22603 45067
rect 22603 45033 22612 45067
rect 22560 45024 22612 45033
rect 22744 45024 22796 45076
rect 20260 44956 20312 45008
rect 21272 44956 21324 45008
rect 23756 45024 23808 45076
rect 25964 45067 26016 45076
rect 25964 45033 25973 45067
rect 25973 45033 26007 45067
rect 26007 45033 26016 45067
rect 25964 45024 26016 45033
rect 26424 45024 26476 45076
rect 29092 45024 29144 45076
rect 30472 45024 30524 45076
rect 31944 45024 31996 45076
rect 32588 45024 32640 45076
rect 33508 45024 33560 45076
rect 33784 45024 33836 45076
rect 26240 44956 26292 45008
rect 29368 44956 29420 45008
rect 20536 44931 20588 44940
rect 20536 44897 20545 44931
rect 20545 44897 20579 44931
rect 20579 44897 20588 44931
rect 21640 44931 21692 44940
rect 20536 44888 20588 44897
rect 20076 44863 20128 44872
rect 20076 44829 20085 44863
rect 20085 44829 20119 44863
rect 20119 44829 20128 44863
rect 20076 44820 20128 44829
rect 20812 44820 20864 44872
rect 21640 44897 21649 44931
rect 21649 44897 21683 44931
rect 21683 44897 21692 44931
rect 21640 44888 21692 44897
rect 23664 44888 23716 44940
rect 22744 44863 22796 44872
rect 22744 44829 22753 44863
rect 22753 44829 22787 44863
rect 22787 44829 22796 44863
rect 22744 44820 22796 44829
rect 23296 44820 23348 44872
rect 23480 44820 23532 44872
rect 24584 44863 24636 44872
rect 24584 44829 24593 44863
rect 24593 44829 24627 44863
rect 24627 44829 24636 44863
rect 24584 44820 24636 44829
rect 24860 44863 24912 44872
rect 24860 44829 24869 44863
rect 24869 44829 24903 44863
rect 24903 44829 24912 44863
rect 24860 44820 24912 44829
rect 25320 44820 25372 44872
rect 25872 44863 25924 44872
rect 25872 44829 25881 44863
rect 25881 44829 25915 44863
rect 25915 44829 25924 44863
rect 25872 44820 25924 44829
rect 27620 44888 27672 44940
rect 19984 44684 20036 44736
rect 20812 44684 20864 44736
rect 23296 44727 23348 44736
rect 23296 44693 23305 44727
rect 23305 44693 23339 44727
rect 23339 44693 23348 44727
rect 23296 44684 23348 44693
rect 24308 44684 24360 44736
rect 27528 44820 27580 44872
rect 27804 44820 27856 44872
rect 28540 44820 28592 44872
rect 28724 44863 28776 44872
rect 28724 44829 28733 44863
rect 28733 44829 28767 44863
rect 28767 44829 28776 44863
rect 28724 44820 28776 44829
rect 29552 44820 29604 44872
rect 28448 44752 28500 44804
rect 26608 44684 26660 44736
rect 26884 44727 26936 44736
rect 26884 44693 26893 44727
rect 26893 44693 26927 44727
rect 26927 44693 26936 44727
rect 26884 44684 26936 44693
rect 27436 44684 27488 44736
rect 28080 44684 28132 44736
rect 29828 44820 29880 44872
rect 30104 44863 30156 44872
rect 30104 44829 30113 44863
rect 30113 44829 30147 44863
rect 30147 44829 30156 44863
rect 32036 44956 32088 45008
rect 33232 44956 33284 45008
rect 31852 44888 31904 44940
rect 32496 44888 32548 44940
rect 37648 45024 37700 45076
rect 38660 45024 38712 45076
rect 40040 45067 40092 45076
rect 40040 45033 40049 45067
rect 40049 45033 40083 45067
rect 40083 45033 40092 45067
rect 40040 45024 40092 45033
rect 40868 45024 40920 45076
rect 34612 44956 34664 45008
rect 35348 44956 35400 45008
rect 30104 44820 30156 44829
rect 31668 44820 31720 44872
rect 32772 44863 32824 44872
rect 32772 44829 32781 44863
rect 32781 44829 32815 44863
rect 32815 44829 32824 44863
rect 32772 44820 32824 44829
rect 35072 44863 35124 44872
rect 32128 44752 32180 44804
rect 35072 44829 35081 44863
rect 35081 44829 35115 44863
rect 35115 44829 35124 44863
rect 35072 44820 35124 44829
rect 36268 44888 36320 44940
rect 37464 44931 37516 44940
rect 37464 44897 37473 44931
rect 37473 44897 37507 44931
rect 37507 44897 37516 44931
rect 37464 44888 37516 44897
rect 38752 44888 38804 44940
rect 34152 44752 34204 44804
rect 30012 44684 30064 44736
rect 34612 44684 34664 44736
rect 34980 44752 35032 44804
rect 37372 44863 37424 44872
rect 35624 44752 35676 44804
rect 37372 44829 37381 44863
rect 37381 44829 37415 44863
rect 37415 44829 37424 44863
rect 37372 44820 37424 44829
rect 38016 44820 38068 44872
rect 38108 44820 38160 44872
rect 35808 44684 35860 44736
rect 36912 44752 36964 44804
rect 37924 44752 37976 44804
rect 38292 44752 38344 44804
rect 36820 44684 36872 44736
rect 38476 44684 38528 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 20260 44523 20312 44532
rect 20260 44489 20269 44523
rect 20269 44489 20303 44523
rect 20303 44489 20312 44523
rect 20260 44480 20312 44489
rect 19432 44412 19484 44464
rect 23848 44480 23900 44532
rect 24216 44480 24268 44532
rect 25780 44480 25832 44532
rect 25872 44480 25924 44532
rect 25136 44412 25188 44464
rect 25964 44412 26016 44464
rect 26884 44412 26936 44464
rect 28540 44480 28592 44532
rect 32312 44523 32364 44532
rect 32312 44489 32321 44523
rect 32321 44489 32355 44523
rect 32355 44489 32364 44523
rect 32312 44480 32364 44489
rect 33600 44480 33652 44532
rect 34612 44480 34664 44532
rect 34980 44480 35032 44532
rect 20812 44387 20864 44396
rect 20812 44353 20821 44387
rect 20821 44353 20855 44387
rect 20855 44353 20864 44387
rect 20812 44344 20864 44353
rect 22652 44344 22704 44396
rect 23756 44344 23808 44396
rect 23296 44319 23348 44328
rect 23296 44285 23305 44319
rect 23305 44285 23339 44319
rect 23339 44285 23348 44319
rect 23296 44276 23348 44285
rect 24768 44387 24820 44396
rect 24768 44353 24777 44387
rect 24777 44353 24811 44387
rect 24811 44353 24820 44387
rect 25320 44387 25372 44396
rect 24768 44344 24820 44353
rect 25320 44353 25329 44387
rect 25329 44353 25363 44387
rect 25363 44353 25372 44387
rect 25320 44344 25372 44353
rect 25596 44344 25648 44396
rect 26608 44387 26660 44396
rect 26608 44353 26617 44387
rect 26617 44353 26651 44387
rect 26651 44353 26660 44387
rect 27804 44387 27856 44396
rect 26608 44344 26660 44353
rect 27804 44353 27813 44387
rect 27813 44353 27847 44387
rect 27847 44353 27856 44387
rect 27804 44344 27856 44353
rect 28080 44412 28132 44464
rect 29460 44412 29512 44464
rect 29736 44412 29788 44464
rect 34796 44412 34848 44464
rect 35440 44480 35492 44532
rect 35716 44412 35768 44464
rect 36912 44480 36964 44532
rect 37464 44523 37516 44532
rect 37464 44489 37473 44523
rect 37473 44489 37507 44523
rect 37507 44489 37516 44523
rect 37464 44480 37516 44489
rect 38108 44480 38160 44532
rect 29276 44344 29328 44396
rect 32496 44387 32548 44396
rect 32496 44353 32505 44387
rect 32505 44353 32539 44387
rect 32539 44353 32548 44387
rect 32496 44344 32548 44353
rect 27344 44276 27396 44328
rect 29184 44319 29236 44328
rect 29184 44285 29193 44319
rect 29193 44285 29227 44319
rect 29227 44285 29236 44319
rect 29184 44276 29236 44285
rect 30196 44319 30248 44328
rect 30196 44285 30205 44319
rect 30205 44285 30239 44319
rect 30239 44285 30248 44319
rect 30196 44276 30248 44285
rect 31576 44319 31628 44328
rect 19984 44140 20036 44192
rect 20720 44140 20772 44192
rect 23940 44140 23992 44192
rect 24584 44140 24636 44192
rect 25136 44208 25188 44260
rect 29092 44208 29144 44260
rect 31576 44285 31585 44319
rect 31585 44285 31619 44319
rect 31619 44285 31628 44319
rect 31576 44276 31628 44285
rect 32772 44276 32824 44328
rect 34612 44319 34664 44328
rect 34612 44285 34621 44319
rect 34621 44285 34655 44319
rect 34655 44285 34664 44319
rect 34612 44276 34664 44285
rect 35348 44344 35400 44396
rect 36268 44344 36320 44396
rect 36912 44344 36964 44396
rect 36084 44208 36136 44260
rect 38568 44344 38620 44396
rect 37924 44319 37976 44328
rect 37924 44285 37933 44319
rect 37933 44285 37967 44319
rect 37967 44285 37976 44319
rect 37924 44276 37976 44285
rect 38476 44208 38528 44260
rect 25412 44140 25464 44192
rect 27528 44140 27580 44192
rect 35072 44140 35124 44192
rect 35716 44140 35768 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 20536 43936 20588 43988
rect 21088 43936 21140 43988
rect 23204 43936 23256 43988
rect 23756 43979 23808 43988
rect 23756 43945 23765 43979
rect 23765 43945 23799 43979
rect 23799 43945 23808 43979
rect 23756 43936 23808 43945
rect 25044 43936 25096 43988
rect 26700 43936 26752 43988
rect 27344 43936 27396 43988
rect 29184 43936 29236 43988
rect 31576 43936 31628 43988
rect 32588 43936 32640 43988
rect 34060 43936 34112 43988
rect 35440 43936 35492 43988
rect 35716 43979 35768 43988
rect 35716 43945 35725 43979
rect 35725 43945 35759 43979
rect 35759 43945 35768 43979
rect 35716 43936 35768 43945
rect 35900 43936 35952 43988
rect 36636 43936 36688 43988
rect 20904 43868 20956 43920
rect 29920 43868 29972 43920
rect 30564 43868 30616 43920
rect 21732 43775 21784 43784
rect 21732 43741 21741 43775
rect 21741 43741 21775 43775
rect 21775 43741 21784 43775
rect 21732 43732 21784 43741
rect 22376 43775 22428 43784
rect 22376 43741 22385 43775
rect 22385 43741 22419 43775
rect 22419 43741 22428 43775
rect 22376 43732 22428 43741
rect 24492 43800 24544 43852
rect 25136 43800 25188 43852
rect 25596 43800 25648 43852
rect 26608 43800 26660 43852
rect 20720 43664 20772 43716
rect 23020 43664 23072 43716
rect 23940 43732 23992 43784
rect 24768 43732 24820 43784
rect 29460 43800 29512 43852
rect 32680 43800 32732 43852
rect 26884 43732 26936 43784
rect 28816 43775 28868 43784
rect 28816 43741 28825 43775
rect 28825 43741 28859 43775
rect 28859 43741 28868 43775
rect 28816 43732 28868 43741
rect 30012 43775 30064 43784
rect 30012 43741 30021 43775
rect 30021 43741 30055 43775
rect 30055 43741 30064 43775
rect 30012 43732 30064 43741
rect 32496 43732 32548 43784
rect 25320 43664 25372 43716
rect 32772 43664 32824 43716
rect 33508 43732 33560 43784
rect 33692 43732 33744 43784
rect 34704 43664 34756 43716
rect 35440 43664 35492 43716
rect 35808 43664 35860 43716
rect 21916 43596 21968 43648
rect 24860 43596 24912 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 20536 43392 20588 43444
rect 23572 43392 23624 43444
rect 24860 43392 24912 43444
rect 25596 43435 25648 43444
rect 25596 43401 25605 43435
rect 25605 43401 25639 43435
rect 25639 43401 25648 43435
rect 25596 43392 25648 43401
rect 27528 43392 27580 43444
rect 28172 43435 28224 43444
rect 28172 43401 28181 43435
rect 28181 43401 28215 43435
rect 28215 43401 28224 43435
rect 28172 43392 28224 43401
rect 33784 43435 33836 43444
rect 33784 43401 33793 43435
rect 33793 43401 33827 43435
rect 33827 43401 33836 43435
rect 33784 43392 33836 43401
rect 35440 43392 35492 43444
rect 24768 43324 24820 43376
rect 27620 43367 27672 43376
rect 27620 43333 27629 43367
rect 27629 43333 27663 43367
rect 27663 43333 27672 43367
rect 27620 43324 27672 43333
rect 22468 43299 22520 43308
rect 22468 43265 22477 43299
rect 22477 43265 22511 43299
rect 22511 43265 22520 43299
rect 22468 43256 22520 43265
rect 23388 43256 23440 43308
rect 23848 43256 23900 43308
rect 24032 43256 24084 43308
rect 25136 43256 25188 43308
rect 25320 43256 25372 43308
rect 25780 43299 25832 43308
rect 25780 43265 25789 43299
rect 25789 43265 25823 43299
rect 25823 43265 25832 43299
rect 25780 43256 25832 43265
rect 26792 43256 26844 43308
rect 30104 43324 30156 43376
rect 29000 43256 29052 43308
rect 29644 43256 29696 43308
rect 31300 43299 31352 43308
rect 31300 43265 31309 43299
rect 31309 43265 31343 43299
rect 31343 43265 31352 43299
rect 31300 43256 31352 43265
rect 32404 43256 32456 43308
rect 33140 43256 33192 43308
rect 34520 43256 34572 43308
rect 27896 43188 27948 43240
rect 31668 43188 31720 43240
rect 33324 43188 33376 43240
rect 25504 43120 25556 43172
rect 27344 43120 27396 43172
rect 27436 43095 27488 43104
rect 27436 43061 27445 43095
rect 27445 43061 27479 43095
rect 27479 43061 27488 43095
rect 27436 43052 27488 43061
rect 30656 43095 30708 43104
rect 30656 43061 30665 43095
rect 30665 43061 30699 43095
rect 30699 43061 30708 43095
rect 30656 43052 30708 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 24952 42848 25004 42900
rect 26792 42891 26844 42900
rect 22652 42712 22704 42764
rect 24676 42755 24728 42764
rect 24676 42721 24685 42755
rect 24685 42721 24719 42755
rect 24719 42721 24728 42755
rect 24676 42712 24728 42721
rect 26792 42857 26801 42891
rect 26801 42857 26835 42891
rect 26835 42857 26844 42891
rect 26792 42848 26844 42857
rect 27068 42848 27120 42900
rect 33140 42848 33192 42900
rect 27252 42755 27304 42764
rect 27252 42721 27261 42755
rect 27261 42721 27295 42755
rect 27295 42721 27304 42755
rect 27252 42712 27304 42721
rect 28264 42712 28316 42764
rect 30656 42780 30708 42832
rect 32220 42755 32272 42764
rect 27712 42644 27764 42696
rect 27804 42576 27856 42628
rect 29460 42576 29512 42628
rect 32220 42721 32229 42755
rect 32229 42721 32263 42755
rect 32263 42721 32272 42755
rect 32220 42712 32272 42721
rect 30104 42644 30156 42696
rect 21916 42551 21968 42560
rect 21916 42517 21925 42551
rect 21925 42517 21959 42551
rect 21959 42517 21968 42551
rect 21916 42508 21968 42517
rect 24032 42551 24084 42560
rect 24032 42517 24041 42551
rect 24041 42517 24075 42551
rect 24075 42517 24084 42551
rect 24032 42508 24084 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 24032 42304 24084 42356
rect 25780 42304 25832 42356
rect 27160 42347 27212 42356
rect 27160 42313 27169 42347
rect 27169 42313 27203 42347
rect 27203 42313 27212 42347
rect 27160 42304 27212 42313
rect 27712 42347 27764 42356
rect 27712 42313 27721 42347
rect 27721 42313 27755 42347
rect 27755 42313 27764 42347
rect 27712 42304 27764 42313
rect 28816 42304 28868 42356
rect 29460 42347 29512 42356
rect 29460 42313 29469 42347
rect 29469 42313 29503 42347
rect 29503 42313 29512 42347
rect 29460 42304 29512 42313
rect 30104 42236 30156 42288
rect 21916 41964 21968 42016
rect 25136 42032 25188 42084
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 27804 41803 27856 41812
rect 27804 41769 27813 41803
rect 27813 41769 27847 41803
rect 27847 41769 27856 41803
rect 27804 41760 27856 41769
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 25136 7531 25188 7540
rect 25136 7497 25145 7531
rect 25145 7497 25179 7531
rect 25179 7497 25188 7531
rect 25136 7488 25188 7497
rect 25044 7352 25096 7404
rect 23112 7191 23164 7200
rect 23112 7157 23121 7191
rect 23121 7157 23155 7191
rect 23155 7157 23164 7191
rect 23112 7148 23164 7157
rect 23756 7191 23808 7200
rect 23756 7157 23765 7191
rect 23765 7157 23799 7191
rect 23799 7157 23808 7191
rect 23756 7148 23808 7157
rect 24584 7191 24636 7200
rect 24584 7157 24593 7191
rect 24593 7157 24627 7191
rect 24627 7157 24636 7191
rect 24584 7148 24636 7157
rect 25596 7148 25648 7200
rect 26424 7191 26476 7200
rect 26424 7157 26433 7191
rect 26433 7157 26467 7191
rect 26467 7157 26476 7191
rect 26424 7148 26476 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 21180 6783 21232 6792
rect 21180 6749 21189 6783
rect 21189 6749 21223 6783
rect 21223 6749 21232 6783
rect 21180 6740 21232 6749
rect 21272 6740 21324 6792
rect 25044 6808 25096 6860
rect 25136 6783 25188 6792
rect 25136 6749 25145 6783
rect 25145 6749 25179 6783
rect 25179 6749 25188 6783
rect 25136 6740 25188 6749
rect 26240 6783 26292 6792
rect 26240 6749 26249 6783
rect 26249 6749 26283 6783
rect 26283 6749 26292 6783
rect 26700 6783 26752 6792
rect 26240 6740 26292 6749
rect 26700 6749 26709 6783
rect 26709 6749 26743 6783
rect 26743 6749 26752 6783
rect 26700 6740 26752 6749
rect 27528 6740 27580 6792
rect 27804 6740 27856 6792
rect 22376 6647 22428 6656
rect 22376 6613 22385 6647
rect 22385 6613 22419 6647
rect 22419 6613 22428 6647
rect 22376 6604 22428 6613
rect 23020 6647 23072 6656
rect 23020 6613 23029 6647
rect 23029 6613 23063 6647
rect 23063 6613 23072 6647
rect 23020 6604 23072 6613
rect 24492 6604 24544 6656
rect 24860 6604 24912 6656
rect 27712 6604 27764 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 24492 6375 24544 6384
rect 24492 6341 24501 6375
rect 24501 6341 24535 6375
rect 24535 6341 24544 6375
rect 24492 6332 24544 6341
rect 27712 6375 27764 6384
rect 27712 6341 27721 6375
rect 27721 6341 27755 6375
rect 27755 6341 27764 6375
rect 27712 6332 27764 6341
rect 21272 6307 21324 6316
rect 21272 6273 21281 6307
rect 21281 6273 21315 6307
rect 21315 6273 21324 6307
rect 21272 6264 21324 6273
rect 27528 6307 27580 6316
rect 27528 6273 27537 6307
rect 27537 6273 27571 6307
rect 27571 6273 27580 6307
rect 27528 6264 27580 6273
rect 22284 6196 22336 6248
rect 24952 6239 25004 6248
rect 24952 6205 24961 6239
rect 24961 6205 24995 6239
rect 24995 6205 25004 6239
rect 24952 6196 25004 6205
rect 29184 6239 29236 6248
rect 29184 6205 29193 6239
rect 29193 6205 29227 6239
rect 29227 6205 29236 6239
rect 29184 6196 29236 6205
rect 22100 6128 22152 6180
rect 18972 6103 19024 6112
rect 18972 6069 18981 6103
rect 18981 6069 19015 6103
rect 19015 6069 19024 6103
rect 18972 6060 19024 6069
rect 19340 6060 19392 6112
rect 20260 6103 20312 6112
rect 20260 6069 20269 6103
rect 20269 6069 20303 6103
rect 20303 6069 20312 6103
rect 20260 6060 20312 6069
rect 22192 6060 22244 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 21272 5788 21324 5840
rect 18604 5652 18656 5704
rect 20168 5720 20220 5772
rect 25044 5788 25096 5840
rect 22192 5763 22244 5772
rect 22192 5729 22201 5763
rect 22201 5729 22235 5763
rect 22235 5729 22244 5763
rect 22192 5720 22244 5729
rect 22376 5763 22428 5772
rect 22376 5729 22385 5763
rect 22385 5729 22419 5763
rect 22419 5729 22428 5763
rect 22376 5720 22428 5729
rect 22928 5763 22980 5772
rect 22928 5729 22937 5763
rect 22937 5729 22971 5763
rect 22971 5729 22980 5763
rect 22928 5720 22980 5729
rect 26240 5720 26292 5772
rect 20812 5695 20864 5704
rect 20812 5661 20821 5695
rect 20821 5661 20855 5695
rect 20855 5661 20864 5695
rect 20812 5652 20864 5661
rect 24860 5695 24912 5704
rect 24860 5661 24869 5695
rect 24869 5661 24903 5695
rect 24903 5661 24912 5695
rect 24860 5652 24912 5661
rect 29000 5652 29052 5704
rect 25136 5627 25188 5636
rect 18972 5516 19024 5568
rect 25136 5593 25145 5627
rect 25145 5593 25179 5627
rect 25179 5593 25188 5627
rect 25136 5584 25188 5593
rect 26608 5584 26660 5636
rect 21732 5516 21784 5568
rect 27804 5516 27856 5568
rect 29644 5516 29696 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 18972 5219 19024 5228
rect 18972 5185 18981 5219
rect 18981 5185 19015 5219
rect 19015 5185 19024 5219
rect 18972 5176 19024 5185
rect 21180 5244 21232 5296
rect 23020 5244 23072 5296
rect 24584 5287 24636 5296
rect 24584 5253 24593 5287
rect 24593 5253 24627 5287
rect 24627 5253 24636 5287
rect 24584 5244 24636 5253
rect 29644 5287 29696 5296
rect 29644 5253 29653 5287
rect 29653 5253 29687 5287
rect 29687 5253 29696 5287
rect 29644 5244 29696 5253
rect 22100 5219 22152 5228
rect 22100 5185 22109 5219
rect 22109 5185 22143 5219
rect 22143 5185 22152 5219
rect 22100 5176 22152 5185
rect 29000 5219 29052 5228
rect 29000 5185 29009 5219
rect 29009 5185 29043 5219
rect 29043 5185 29052 5219
rect 29000 5176 29052 5185
rect 17960 5108 18012 5160
rect 21364 5151 21416 5160
rect 21364 5117 21373 5151
rect 21373 5117 21407 5151
rect 21407 5117 21416 5151
rect 21364 5108 21416 5117
rect 23480 5151 23532 5160
rect 23480 5117 23489 5151
rect 23489 5117 23523 5151
rect 23523 5117 23532 5151
rect 23480 5108 23532 5117
rect 24032 5108 24084 5160
rect 25228 5151 25280 5160
rect 25228 5117 25237 5151
rect 25237 5117 25271 5151
rect 25271 5117 25280 5151
rect 25228 5108 25280 5117
rect 27988 5108 28040 5160
rect 29736 5108 29788 5160
rect 30012 5151 30064 5160
rect 30012 5117 30021 5151
rect 30021 5117 30055 5151
rect 30055 5117 30064 5151
rect 30012 5108 30064 5117
rect 19984 5040 20036 5092
rect 27712 5040 27764 5092
rect 16948 4972 17000 5024
rect 18328 4972 18380 5024
rect 20076 4972 20128 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19064 4632 19116 4684
rect 20260 4700 20312 4752
rect 20076 4675 20128 4684
rect 20076 4641 20085 4675
rect 20085 4641 20119 4675
rect 20119 4641 20128 4675
rect 20076 4632 20128 4641
rect 21088 4675 21140 4684
rect 21088 4641 21097 4675
rect 21097 4641 21131 4675
rect 21131 4641 21140 4675
rect 21088 4632 21140 4641
rect 23112 4768 23164 4820
rect 27988 4811 28040 4820
rect 27988 4777 27997 4811
rect 27997 4777 28031 4811
rect 28031 4777 28040 4811
rect 27988 4768 28040 4777
rect 29736 4811 29788 4820
rect 29736 4777 29745 4811
rect 29745 4777 29779 4811
rect 29779 4777 29788 4811
rect 29736 4768 29788 4777
rect 22284 4700 22336 4752
rect 23572 4675 23624 4684
rect 23572 4641 23581 4675
rect 23581 4641 23615 4675
rect 23615 4641 23624 4675
rect 23572 4632 23624 4641
rect 25044 4632 25096 4684
rect 25596 4675 25648 4684
rect 25596 4641 25605 4675
rect 25605 4641 25639 4675
rect 25639 4641 25648 4675
rect 25596 4632 25648 4641
rect 26332 4675 26384 4684
rect 26332 4641 26341 4675
rect 26341 4641 26375 4675
rect 26375 4641 26384 4675
rect 26332 4632 26384 4641
rect 31300 4632 31352 4684
rect 15016 4564 15068 4616
rect 15844 4564 15896 4616
rect 17408 4564 17460 4616
rect 18052 4607 18104 4616
rect 18052 4573 18061 4607
rect 18061 4573 18095 4607
rect 18095 4573 18104 4607
rect 18052 4564 18104 4573
rect 19432 4564 19484 4616
rect 24860 4564 24912 4616
rect 27804 4564 27856 4616
rect 29000 4564 29052 4616
rect 31208 4607 31260 4616
rect 31208 4573 31217 4607
rect 31217 4573 31251 4607
rect 31251 4573 31260 4607
rect 31208 4564 31260 4573
rect 32128 4564 32180 4616
rect 32312 4607 32364 4616
rect 32312 4573 32321 4607
rect 32321 4573 32355 4607
rect 32355 4573 32364 4607
rect 32312 4564 32364 4573
rect 31760 4471 31812 4480
rect 31760 4437 31769 4471
rect 31769 4437 31803 4471
rect 31803 4437 31812 4471
rect 31760 4428 31812 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 32128 4156 32180 4208
rect 16764 4088 16816 4140
rect 17224 4020 17276 4072
rect 17684 3952 17736 4004
rect 19432 4088 19484 4140
rect 24032 4088 24084 4140
rect 29000 4131 29052 4140
rect 29000 4097 29009 4131
rect 29009 4097 29043 4131
rect 29043 4097 29052 4131
rect 29000 4088 29052 4097
rect 31300 4131 31352 4140
rect 31300 4097 31309 4131
rect 31309 4097 31343 4131
rect 31343 4097 31352 4131
rect 31300 4088 31352 4097
rect 31576 4088 31628 4140
rect 32312 4088 32364 4140
rect 22284 4020 22336 4072
rect 24308 4063 24360 4072
rect 24308 4029 24317 4063
rect 24317 4029 24351 4063
rect 24351 4029 24360 4063
rect 24308 4020 24360 4029
rect 24676 4063 24728 4072
rect 24676 4029 24685 4063
rect 24685 4029 24719 4063
rect 24719 4029 24728 4063
rect 24676 4020 24728 4029
rect 27436 4063 27488 4072
rect 27436 4029 27445 4063
rect 27445 4029 27479 4063
rect 27479 4029 27488 4063
rect 27436 4020 27488 4029
rect 27896 4020 27948 4072
rect 29092 4020 29144 4072
rect 20168 3952 20220 4004
rect 31392 4020 31444 4072
rect 31760 3952 31812 4004
rect 34060 3952 34112 4004
rect 12256 3884 12308 3936
rect 13084 3884 13136 3936
rect 13912 3884 13964 3936
rect 15292 3884 15344 3936
rect 17500 3884 17552 3936
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 22100 3884 22152 3936
rect 24768 3884 24820 3936
rect 25504 3884 25556 3936
rect 31852 3884 31904 3936
rect 32772 3884 32824 3936
rect 33784 3884 33836 3936
rect 35348 3884 35400 3936
rect 47308 3884 47360 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 17960 3680 18012 3732
rect 20260 3680 20312 3732
rect 24308 3680 24360 3732
rect 27896 3723 27948 3732
rect 27896 3689 27905 3723
rect 27905 3689 27939 3723
rect 27939 3689 27948 3723
rect 27896 3680 27948 3689
rect 30748 3680 30800 3732
rect 16396 3612 16448 3664
rect 17132 3612 17184 3664
rect 20536 3612 20588 3664
rect 4620 3476 4672 3528
rect 4896 3476 4948 3528
rect 5724 3476 5776 3528
rect 6552 3476 6604 3528
rect 7380 3476 7432 3528
rect 8208 3476 8260 3528
rect 9036 3476 9088 3528
rect 9864 3476 9916 3528
rect 10692 3476 10744 3528
rect 11520 3476 11572 3528
rect 12808 3476 12860 3528
rect 13636 3476 13688 3528
rect 14188 3476 14240 3528
rect 16120 3519 16172 3528
rect 16120 3485 16129 3519
rect 16129 3485 16163 3519
rect 16163 3485 16172 3519
rect 16764 3519 16816 3528
rect 16120 3476 16172 3485
rect 16764 3485 16773 3519
rect 16773 3485 16807 3519
rect 16807 3485 16816 3519
rect 16764 3476 16816 3485
rect 19248 3544 19300 3596
rect 17960 3476 18012 3528
rect 20812 3544 20864 3596
rect 21732 3587 21784 3596
rect 21732 3553 21741 3587
rect 21741 3553 21775 3587
rect 21775 3553 21784 3587
rect 21732 3544 21784 3553
rect 22192 3587 22244 3596
rect 22192 3553 22201 3587
rect 22201 3553 22235 3587
rect 22235 3553 22244 3587
rect 22192 3544 22244 3553
rect 16764 3340 16816 3392
rect 22468 3408 22520 3460
rect 25136 3612 25188 3664
rect 25504 3587 25556 3596
rect 25504 3553 25513 3587
rect 25513 3553 25547 3587
rect 25547 3553 25556 3587
rect 25504 3544 25556 3553
rect 26056 3587 26108 3596
rect 26056 3553 26065 3587
rect 26065 3553 26099 3587
rect 26099 3553 26108 3587
rect 26056 3544 26108 3553
rect 30196 3612 30248 3664
rect 24860 3519 24912 3528
rect 24860 3485 24869 3519
rect 24869 3485 24903 3519
rect 24903 3485 24912 3519
rect 24860 3476 24912 3485
rect 31208 3544 31260 3596
rect 31760 3612 31812 3664
rect 27804 3519 27856 3528
rect 27804 3485 27813 3519
rect 27813 3485 27847 3519
rect 27847 3485 27856 3519
rect 27804 3476 27856 3485
rect 29000 3476 29052 3528
rect 32128 3476 32180 3528
rect 28264 3408 28316 3460
rect 32404 3408 32456 3460
rect 32680 3519 32732 3528
rect 32680 3485 32689 3519
rect 32689 3485 32723 3519
rect 32723 3485 32732 3519
rect 32680 3476 32732 3485
rect 33232 3612 33284 3664
rect 35440 3612 35492 3664
rect 37464 3612 37516 3664
rect 40684 3612 40736 3664
rect 46480 3612 46532 3664
rect 34520 3544 34572 3596
rect 34612 3544 34664 3596
rect 35992 3544 36044 3596
rect 41236 3544 41288 3596
rect 47032 3544 47084 3596
rect 33600 3408 33652 3460
rect 20628 3340 20680 3392
rect 23848 3340 23900 3392
rect 28816 3340 28868 3392
rect 30472 3340 30524 3392
rect 31760 3340 31812 3392
rect 31944 3340 31996 3392
rect 32220 3340 32272 3392
rect 36544 3476 36596 3528
rect 37924 3476 37976 3528
rect 39304 3476 39356 3528
rect 40132 3476 40184 3528
rect 42616 3476 42668 3528
rect 42892 3476 42944 3528
rect 44548 3476 44600 3528
rect 45376 3476 45428 3528
rect 46204 3476 46256 3528
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 14464 3000 14516 3052
rect 19156 3136 19208 3188
rect 17500 3111 17552 3120
rect 17500 3077 17509 3111
rect 17509 3077 17543 3111
rect 17543 3077 17552 3111
rect 17500 3068 17552 3077
rect 17776 3068 17828 3120
rect 16120 3043 16172 3052
rect 16120 3009 16129 3043
rect 16129 3009 16163 3043
rect 16163 3009 16172 3043
rect 16120 3000 16172 3009
rect 4712 2932 4764 2984
rect 6000 2932 6052 2984
rect 16672 2932 16724 2984
rect 18052 2932 18104 2984
rect 23756 3136 23808 3188
rect 27988 3136 28040 3188
rect 29184 3136 29236 3188
rect 29920 3136 29972 3188
rect 33692 3136 33744 3188
rect 20260 3068 20312 3120
rect 23848 3068 23900 3120
rect 28816 3111 28868 3120
rect 28816 3077 28825 3111
rect 28825 3077 28859 3111
rect 28859 3077 28868 3111
rect 28816 3068 28868 3077
rect 33048 3068 33100 3120
rect 33508 3068 33560 3120
rect 36176 3068 36228 3120
rect 22468 3043 22520 3052
rect 22468 3009 22477 3043
rect 22477 3009 22511 3043
rect 22511 3009 22520 3043
rect 22468 3000 22520 3009
rect 24768 3043 24820 3052
rect 24768 3009 24777 3043
rect 24777 3009 24811 3043
rect 24811 3009 24820 3043
rect 24768 3000 24820 3009
rect 29000 3043 29052 3052
rect 29000 3009 29009 3043
rect 29009 3009 29043 3043
rect 29043 3009 29052 3043
rect 29000 3000 29052 3009
rect 32864 3000 32916 3052
rect 33600 3043 33652 3052
rect 13360 2864 13412 2916
rect 17132 2864 17184 2916
rect 3516 2796 3568 2848
rect 5172 2796 5224 2848
rect 6276 2796 6328 2848
rect 7656 2796 7708 2848
rect 8484 2796 8536 2848
rect 8760 2796 8812 2848
rect 9588 2796 9640 2848
rect 10416 2796 10468 2848
rect 10968 2796 11020 2848
rect 11796 2796 11848 2848
rect 16120 2796 16172 2848
rect 17868 2796 17920 2848
rect 17960 2796 18012 2848
rect 18880 2796 18932 2848
rect 23848 2932 23900 2984
rect 24400 2932 24452 2984
rect 25504 2975 25556 2984
rect 25504 2941 25513 2975
rect 25513 2941 25547 2975
rect 25547 2941 25556 2975
rect 25504 2932 25556 2941
rect 26884 2932 26936 2984
rect 28540 2932 28592 2984
rect 33600 3009 33609 3043
rect 33609 3009 33643 3043
rect 33643 3009 33652 3043
rect 33600 3000 33652 3009
rect 35716 3000 35768 3052
rect 34796 2932 34848 2984
rect 37372 2932 37424 2984
rect 37648 2932 37700 2984
rect 39856 2932 39908 2984
rect 42340 2932 42392 2984
rect 44272 2932 44324 2984
rect 31024 2864 31076 2916
rect 34336 2864 34388 2916
rect 36820 2864 36872 2916
rect 38476 2864 38528 2916
rect 40408 2864 40460 2916
rect 43168 2864 43220 2916
rect 45100 2864 45152 2916
rect 21640 2796 21692 2848
rect 28816 2796 28868 2848
rect 30012 2796 30064 2848
rect 30380 2796 30432 2848
rect 32496 2796 32548 2848
rect 38752 2796 38804 2848
rect 41788 2796 41840 2848
rect 43720 2796 43772 2848
rect 45652 2796 45704 2848
rect 46756 2796 46808 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 18052 2592 18104 2644
rect 32404 2635 32456 2644
rect 32404 2601 32413 2635
rect 32413 2601 32447 2635
rect 32447 2601 32456 2635
rect 32404 2592 32456 2601
rect 33048 2635 33100 2644
rect 33048 2601 33057 2635
rect 33057 2601 33091 2635
rect 33091 2601 33100 2635
rect 33048 2592 33100 2601
rect 33600 2635 33652 2644
rect 33600 2601 33609 2635
rect 33609 2601 33643 2635
rect 33643 2601 33652 2635
rect 33600 2592 33652 2601
rect 34520 2592 34572 2644
rect 36176 2635 36228 2644
rect 36176 2601 36185 2635
rect 36185 2601 36219 2635
rect 36219 2601 36228 2635
rect 36176 2592 36228 2601
rect 37372 2592 37424 2644
rect 6828 2524 6880 2576
rect 7932 2524 7984 2576
rect 11244 2524 11296 2576
rect 14740 2524 14792 2576
rect 5448 2456 5500 2508
rect 10140 2456 10192 2508
rect 12532 2456 12584 2508
rect 15476 2456 15528 2508
rect 16764 2456 16816 2508
rect 17868 2456 17920 2508
rect 22744 2456 22796 2508
rect 25780 2499 25832 2508
rect 25780 2465 25789 2499
rect 25789 2465 25823 2499
rect 25823 2465 25832 2499
rect 25780 2456 25832 2465
rect 26424 2499 26476 2508
rect 26424 2465 26433 2499
rect 26433 2465 26467 2499
rect 26467 2465 26476 2499
rect 26424 2456 26476 2465
rect 26700 2456 26752 2508
rect 31944 2524 31996 2576
rect 38200 2524 38252 2576
rect 42064 2524 42116 2576
rect 44824 2524 44876 2576
rect 30380 2456 30432 2508
rect 32680 2456 32732 2508
rect 37096 2456 37148 2508
rect 39028 2456 39080 2508
rect 40960 2456 41012 2508
rect 43444 2456 43496 2508
rect 2596 2388 2648 2440
rect 3148 2388 3200 2440
rect 3884 2388 3936 2440
rect 7104 2388 7156 2440
rect 12072 2388 12124 2440
rect 15568 2388 15620 2440
rect 9312 2320 9364 2372
rect 19248 2388 19300 2440
rect 22100 2388 22152 2440
rect 32128 2388 32180 2440
rect 18788 2252 18840 2304
rect 20628 2320 20680 2372
rect 24124 2320 24176 2372
rect 27160 2363 27212 2372
rect 27160 2329 27169 2363
rect 27169 2329 27203 2363
rect 27203 2329 27212 2363
rect 27160 2320 27212 2329
rect 29368 2320 29420 2372
rect 31852 2320 31904 2372
rect 31944 2320 31996 2372
rect 36268 2388 36320 2440
rect 39580 2388 39632 2440
rect 41512 2388 41564 2440
rect 43996 2320 44048 2372
rect 45928 2388 45980 2440
rect 21916 2252 21968 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 18788 2048 18840 2100
rect 20812 2048 20864 2100
rect 15568 1980 15620 2032
rect 20260 1980 20312 2032
rect 19064 1912 19116 1964
rect 19708 1912 19760 1964
<< metal2 >>
rect 3974 49314 4030 50000
rect 3974 49286 4108 49314
rect 3974 49200 4030 49286
rect 4080 47122 4108 49286
rect 4342 49200 4398 50000
rect 4710 49314 4766 50000
rect 4710 49286 4844 49314
rect 4710 49200 4766 49286
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4068 47116 4120 47122
rect 4068 47058 4120 47064
rect 4080 46714 4108 47058
rect 4068 46708 4120 46714
rect 4068 46650 4120 46656
rect 4816 46578 4844 49286
rect 5078 49200 5134 50000
rect 5446 49200 5502 50000
rect 5814 49314 5870 50000
rect 6182 49314 6238 50000
rect 5814 49286 5948 49314
rect 5814 49200 5870 49286
rect 5092 47258 5120 49200
rect 5080 47252 5132 47258
rect 5080 47194 5132 47200
rect 5632 47048 5684 47054
rect 5632 46990 5684 46996
rect 4804 46572 4856 46578
rect 4804 46514 4856 46520
rect 5644 46510 5672 46990
rect 5632 46504 5684 46510
rect 5632 46446 5684 46452
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 5920 46170 5948 49286
rect 6012 49286 6238 49314
rect 6012 46578 6040 49286
rect 6182 49200 6238 49286
rect 6550 49200 6606 50000
rect 6918 49314 6974 50000
rect 6918 49286 7052 49314
rect 6918 49200 6974 49286
rect 7024 46578 7052 49286
rect 7286 49200 7342 50000
rect 7654 49200 7710 50000
rect 8022 49314 8078 50000
rect 7944 49286 8078 49314
rect 7300 47258 7328 49200
rect 7944 47258 7972 49286
rect 8022 49200 8078 49286
rect 8390 49200 8446 50000
rect 8758 49200 8814 50000
rect 9126 49314 9182 50000
rect 9494 49314 9550 50000
rect 9126 49286 9260 49314
rect 9126 49200 9182 49286
rect 8404 47258 8432 49200
rect 7288 47252 7340 47258
rect 7288 47194 7340 47200
rect 7932 47252 7984 47258
rect 7932 47194 7984 47200
rect 8392 47252 8444 47258
rect 8392 47194 8444 47200
rect 9232 46578 9260 49286
rect 9494 49286 9628 49314
rect 9494 49200 9550 49286
rect 9600 48090 9628 49286
rect 9862 49200 9918 50000
rect 10230 49314 10286 50000
rect 10598 49314 10654 50000
rect 10230 49286 10364 49314
rect 10230 49200 10286 49286
rect 9600 48062 9720 48090
rect 9692 47258 9720 48062
rect 9680 47252 9732 47258
rect 9680 47194 9732 47200
rect 9864 47048 9916 47054
rect 9864 46990 9916 46996
rect 6000 46572 6052 46578
rect 6000 46514 6052 46520
rect 7012 46572 7064 46578
rect 7012 46514 7064 46520
rect 9220 46572 9272 46578
rect 9220 46514 9272 46520
rect 5908 46164 5960 46170
rect 5908 46106 5960 46112
rect 9876 45830 9904 46990
rect 10336 46578 10364 49286
rect 10598 49286 10824 49314
rect 10598 49200 10654 49286
rect 10796 47258 10824 49286
rect 10966 49200 11022 50000
rect 11334 49200 11390 50000
rect 11702 49314 11758 50000
rect 11702 49286 11928 49314
rect 11702 49200 11758 49286
rect 10968 47864 11020 47870
rect 10968 47806 11020 47812
rect 10784 47252 10836 47258
rect 10784 47194 10836 47200
rect 10980 47054 11008 47806
rect 10968 47048 11020 47054
rect 10968 46990 11020 46996
rect 11348 46578 11376 49200
rect 11704 47456 11756 47462
rect 11704 47398 11756 47404
rect 11716 47122 11744 47398
rect 11900 47258 11928 49286
rect 12070 49200 12126 50000
rect 12438 49314 12494 50000
rect 12806 49314 12862 50000
rect 12438 49286 12572 49314
rect 12438 49200 12494 49286
rect 11888 47252 11940 47258
rect 11888 47194 11940 47200
rect 11704 47116 11756 47122
rect 11704 47058 11756 47064
rect 12544 46578 12572 49286
rect 12806 49286 13032 49314
rect 12806 49200 12862 49286
rect 13004 47258 13032 49286
rect 13174 49200 13230 50000
rect 13542 49314 13598 50000
rect 13542 49286 13676 49314
rect 13542 49200 13598 49286
rect 13176 47524 13228 47530
rect 13176 47466 13228 47472
rect 12992 47252 13044 47258
rect 12992 47194 13044 47200
rect 13188 47054 13216 47466
rect 13176 47048 13228 47054
rect 13176 46990 13228 46996
rect 13648 46578 13676 49286
rect 13910 49200 13966 50000
rect 14278 49200 14334 50000
rect 14646 49314 14702 50000
rect 15014 49314 15070 50000
rect 14646 49286 14780 49314
rect 14646 49200 14702 49286
rect 13924 47258 13952 49200
rect 14556 47592 14608 47598
rect 14556 47534 14608 47540
rect 13912 47252 13964 47258
rect 13912 47194 13964 47200
rect 14568 47054 14596 47534
rect 14556 47048 14608 47054
rect 14556 46990 14608 46996
rect 14752 46578 14780 49286
rect 15014 49286 15148 49314
rect 15014 49200 15070 49286
rect 15120 48090 15148 49286
rect 15382 49200 15438 50000
rect 15750 49314 15806 50000
rect 15750 49286 15884 49314
rect 15750 49200 15806 49286
rect 15120 48062 15240 48090
rect 15212 47258 15240 48062
rect 15384 47796 15436 47802
rect 15384 47738 15436 47744
rect 15200 47252 15252 47258
rect 15200 47194 15252 47200
rect 15396 47054 15424 47738
rect 15384 47048 15436 47054
rect 15384 46990 15436 46996
rect 15856 46578 15884 49286
rect 16118 49200 16174 50000
rect 16486 49200 16542 50000
rect 16854 49314 16910 50000
rect 16854 49286 16988 49314
rect 16854 49200 16910 49286
rect 16132 47258 16160 49200
rect 16120 47252 16172 47258
rect 16120 47194 16172 47200
rect 10324 46572 10376 46578
rect 10324 46514 10376 46520
rect 11336 46572 11388 46578
rect 11336 46514 11388 46520
rect 12532 46572 12584 46578
rect 12532 46514 12584 46520
rect 13636 46572 13688 46578
rect 13636 46514 13688 46520
rect 14740 46572 14792 46578
rect 14740 46514 14792 46520
rect 15844 46572 15896 46578
rect 15844 46514 15896 46520
rect 16960 46170 16988 49286
rect 17222 49200 17278 50000
rect 17590 49200 17646 50000
rect 17958 49200 18014 50000
rect 18326 49314 18382 50000
rect 18326 49286 18460 49314
rect 18326 49200 18382 49286
rect 17236 47258 17264 49200
rect 17776 47456 17828 47462
rect 17776 47398 17828 47404
rect 17224 47252 17276 47258
rect 17224 47194 17276 47200
rect 16948 46164 17000 46170
rect 16948 46106 17000 46112
rect 9864 45824 9916 45830
rect 9864 45766 9916 45772
rect 17788 45558 17816 47398
rect 17972 46578 18000 49200
rect 18144 47456 18196 47462
rect 18144 47398 18196 47404
rect 18052 47116 18104 47122
rect 18052 47058 18104 47064
rect 18064 46866 18092 47058
rect 18156 47054 18184 47398
rect 18328 47116 18380 47122
rect 18328 47058 18380 47064
rect 18144 47048 18196 47054
rect 18144 46990 18196 46996
rect 18340 46866 18368 47058
rect 18064 46838 18368 46866
rect 17960 46572 18012 46578
rect 17960 46514 18012 46520
rect 18064 46170 18092 46838
rect 18432 46714 18460 49286
rect 18694 49200 18750 50000
rect 19062 49200 19118 50000
rect 19430 49200 19486 50000
rect 19798 49200 19854 50000
rect 20166 49200 20222 50000
rect 20534 49200 20590 50000
rect 20902 49200 20958 50000
rect 21270 49200 21326 50000
rect 21638 49200 21694 50000
rect 22006 49200 22062 50000
rect 22374 49200 22430 50000
rect 22742 49200 22798 50000
rect 23110 49200 23166 50000
rect 23478 49200 23534 50000
rect 23846 49200 23902 50000
rect 24214 49314 24270 50000
rect 23952 49286 24270 49314
rect 18880 47660 18932 47666
rect 18880 47602 18932 47608
rect 18892 47054 18920 47602
rect 18880 47048 18932 47054
rect 18880 46990 18932 46996
rect 18696 46912 18748 46918
rect 18696 46854 18748 46860
rect 18420 46708 18472 46714
rect 18420 46650 18472 46656
rect 18708 46442 18736 46854
rect 18696 46436 18748 46442
rect 18696 46378 18748 46384
rect 18708 46170 18736 46378
rect 18788 46368 18840 46374
rect 18788 46310 18840 46316
rect 18800 46170 18828 46310
rect 18052 46164 18104 46170
rect 18052 46106 18104 46112
rect 18696 46164 18748 46170
rect 18696 46106 18748 46112
rect 18788 46164 18840 46170
rect 18788 46106 18840 46112
rect 17776 45552 17828 45558
rect 17776 45494 17828 45500
rect 19076 45490 19104 49200
rect 19444 47258 19472 49200
rect 19432 47252 19484 47258
rect 19432 47194 19484 47200
rect 19340 47116 19392 47122
rect 19340 47058 19392 47064
rect 19352 46578 19380 47058
rect 19432 46912 19484 46918
rect 19432 46854 19484 46860
rect 19340 46572 19392 46578
rect 19340 46514 19392 46520
rect 19064 45484 19116 45490
rect 19064 45426 19116 45432
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 19352 45082 19380 46514
rect 19444 46073 19472 46854
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19524 46504 19576 46510
rect 19524 46446 19576 46452
rect 19800 46504 19852 46510
rect 19852 46452 20024 46458
rect 19800 46446 20024 46452
rect 19430 46064 19486 46073
rect 19430 45999 19486 46008
rect 19536 45914 19564 46446
rect 19812 46430 20024 46446
rect 19798 46064 19854 46073
rect 19798 45999 19854 46008
rect 19812 45966 19840 45999
rect 19996 45966 20024 46430
rect 20076 46368 20128 46374
rect 20076 46310 20128 46316
rect 19444 45886 19564 45914
rect 19800 45960 19852 45966
rect 19800 45902 19852 45908
rect 19984 45960 20036 45966
rect 19984 45902 20036 45908
rect 19444 45354 19472 45886
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19432 45348 19484 45354
rect 19432 45290 19484 45296
rect 19340 45076 19392 45082
rect 19340 45018 19392 45024
rect 19444 44470 19472 45290
rect 19996 45286 20024 45902
rect 19984 45280 20036 45286
rect 19984 45222 20036 45228
rect 19996 44742 20024 45222
rect 20088 44878 20116 46310
rect 20180 45422 20208 49200
rect 20352 47592 20404 47598
rect 20352 47534 20404 47540
rect 20260 47048 20312 47054
rect 20260 46990 20312 46996
rect 20272 46578 20300 46990
rect 20260 46572 20312 46578
rect 20260 46514 20312 46520
rect 20272 46442 20300 46514
rect 20260 46436 20312 46442
rect 20260 46378 20312 46384
rect 20260 45824 20312 45830
rect 20260 45766 20312 45772
rect 20168 45416 20220 45422
rect 20168 45358 20220 45364
rect 20272 45014 20300 45766
rect 20364 45286 20392 47534
rect 20444 46980 20496 46986
rect 20444 46922 20496 46928
rect 20456 46034 20484 46922
rect 20548 46714 20576 49200
rect 20720 47864 20772 47870
rect 20720 47806 20772 47812
rect 20536 46708 20588 46714
rect 20536 46650 20588 46656
rect 20732 46578 20760 47806
rect 20904 47660 20956 47666
rect 20904 47602 20956 47608
rect 20720 46572 20772 46578
rect 20720 46514 20772 46520
rect 20732 46102 20760 46514
rect 20916 46374 20944 47602
rect 21088 47048 21140 47054
rect 21088 46990 21140 46996
rect 20904 46368 20956 46374
rect 20904 46310 20956 46316
rect 20720 46096 20772 46102
rect 20720 46038 20772 46044
rect 20444 46028 20496 46034
rect 20444 45970 20496 45976
rect 20536 45552 20588 45558
rect 20812 45552 20864 45558
rect 20536 45494 20588 45500
rect 20810 45520 20812 45529
rect 20864 45520 20866 45529
rect 20352 45280 20404 45286
rect 20352 45222 20404 45228
rect 20260 45008 20312 45014
rect 20260 44950 20312 44956
rect 20076 44872 20128 44878
rect 20076 44814 20128 44820
rect 19984 44736 20036 44742
rect 19984 44678 20036 44684
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19432 44464 19484 44470
rect 19432 44406 19484 44412
rect 19996 44198 20024 44678
rect 20272 44538 20300 44950
rect 20548 44946 20576 45494
rect 20810 45455 20866 45464
rect 20536 44940 20588 44946
rect 20536 44882 20588 44888
rect 20260 44532 20312 44538
rect 20260 44474 20312 44480
rect 19984 44192 20036 44198
rect 19984 44134 20036 44140
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 20548 43994 20576 44882
rect 20824 44878 20852 45455
rect 20812 44872 20864 44878
rect 20812 44814 20864 44820
rect 20812 44736 20864 44742
rect 20812 44678 20864 44684
rect 20824 44402 20852 44678
rect 20812 44396 20864 44402
rect 20812 44338 20864 44344
rect 20720 44192 20772 44198
rect 20720 44134 20772 44140
rect 20536 43988 20588 43994
rect 20536 43930 20588 43936
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 20548 43450 20576 43930
rect 20732 43722 20760 44134
rect 20916 43926 20944 46310
rect 21100 45286 21128 46990
rect 21284 46170 21312 49200
rect 21456 47524 21508 47530
rect 21456 47466 21508 47472
rect 21468 46374 21496 47466
rect 21652 47122 21680 49200
rect 21640 47116 21692 47122
rect 21640 47058 21692 47064
rect 22100 47048 22152 47054
rect 22100 46990 22152 46996
rect 21916 46912 21968 46918
rect 21916 46854 21968 46860
rect 21548 46572 21600 46578
rect 21548 46514 21600 46520
rect 21456 46368 21508 46374
rect 21456 46310 21508 46316
rect 21272 46164 21324 46170
rect 21272 46106 21324 46112
rect 21560 45966 21588 46514
rect 21364 45960 21416 45966
rect 21364 45902 21416 45908
rect 21548 45960 21600 45966
rect 21548 45902 21600 45908
rect 21376 45422 21404 45902
rect 21548 45824 21600 45830
rect 21732 45824 21784 45830
rect 21600 45784 21680 45812
rect 21548 45766 21600 45772
rect 21364 45416 21416 45422
rect 21364 45358 21416 45364
rect 21272 45348 21324 45354
rect 21272 45290 21324 45296
rect 21088 45280 21140 45286
rect 21088 45222 21140 45228
rect 21100 43994 21128 45222
rect 21284 45014 21312 45290
rect 21272 45008 21324 45014
rect 21652 44985 21680 45784
rect 21732 45766 21784 45772
rect 21272 44950 21324 44956
rect 21638 44976 21694 44985
rect 21638 44911 21640 44920
rect 21692 44911 21694 44920
rect 21640 44882 21692 44888
rect 21088 43988 21140 43994
rect 21088 43930 21140 43936
rect 20904 43920 20956 43926
rect 20904 43862 20956 43868
rect 21744 43790 21772 45766
rect 21928 45422 21956 46854
rect 22112 46714 22140 46990
rect 22100 46708 22152 46714
rect 22100 46650 22152 46656
rect 22112 45554 22140 46650
rect 22284 46572 22336 46578
rect 22284 46514 22336 46520
rect 22296 45642 22324 46514
rect 22388 46186 22416 49200
rect 22756 47258 22784 49200
rect 23388 47796 23440 47802
rect 23388 47738 23440 47744
rect 23400 47258 23428 47738
rect 22744 47252 22796 47258
rect 22744 47194 22796 47200
rect 23388 47252 23440 47258
rect 23388 47194 23440 47200
rect 23204 47116 23256 47122
rect 23204 47058 23256 47064
rect 22928 46912 22980 46918
rect 22928 46854 22980 46860
rect 22836 46640 22888 46646
rect 22836 46582 22888 46588
rect 22744 46572 22796 46578
rect 22744 46514 22796 46520
rect 22388 46158 22508 46186
rect 22756 46170 22784 46514
rect 22848 46170 22876 46582
rect 22940 46510 22968 46854
rect 22928 46504 22980 46510
rect 22928 46446 22980 46452
rect 23020 46504 23072 46510
rect 23020 46446 23072 46452
rect 22020 45526 22140 45554
rect 22204 45614 22324 45642
rect 22374 45656 22430 45665
rect 21916 45416 21968 45422
rect 22020 45393 22048 45526
rect 21916 45358 21968 45364
rect 22006 45384 22062 45393
rect 21732 43784 21784 43790
rect 21732 43726 21784 43732
rect 20720 43716 20772 43722
rect 20720 43658 20772 43664
rect 21928 43654 21956 45358
rect 22204 45370 22232 45614
rect 22374 45591 22430 45600
rect 22388 45490 22416 45591
rect 22376 45484 22428 45490
rect 22376 45426 22428 45432
rect 22112 45354 22232 45370
rect 22006 45319 22062 45328
rect 22100 45348 22232 45354
rect 22152 45342 22232 45348
rect 22100 45290 22152 45296
rect 22376 45280 22428 45286
rect 22376 45222 22428 45228
rect 22388 43790 22416 45222
rect 22376 43784 22428 43790
rect 22376 43726 22428 43732
rect 21916 43648 21968 43654
rect 21916 43590 21968 43596
rect 20536 43444 20588 43450
rect 20536 43386 20588 43392
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 21928 42566 21956 43590
rect 22480 43314 22508 46158
rect 22744 46164 22796 46170
rect 22744 46106 22796 46112
rect 22836 46164 22888 46170
rect 22836 46106 22888 46112
rect 22652 46096 22704 46102
rect 22652 46038 22704 46044
rect 22560 45892 22612 45898
rect 22560 45834 22612 45840
rect 22572 45082 22600 45834
rect 22560 45076 22612 45082
rect 22560 45018 22612 45024
rect 22664 44402 22692 46038
rect 22744 45076 22796 45082
rect 22744 45018 22796 45024
rect 22756 44878 22784 45018
rect 22744 44872 22796 44878
rect 22744 44814 22796 44820
rect 22652 44396 22704 44402
rect 22652 44338 22704 44344
rect 22468 43308 22520 43314
rect 22468 43250 22520 43256
rect 22664 42770 22692 44338
rect 23032 43722 23060 46446
rect 23112 46028 23164 46034
rect 23112 45970 23164 45976
rect 23124 45898 23152 45970
rect 23112 45892 23164 45898
rect 23112 45834 23164 45840
rect 23124 45626 23152 45834
rect 23112 45620 23164 45626
rect 23112 45562 23164 45568
rect 23216 43994 23244 47058
rect 23296 47048 23348 47054
rect 23296 46990 23348 46996
rect 23308 46646 23336 46990
rect 23296 46640 23348 46646
rect 23296 46582 23348 46588
rect 23492 45554 23520 49200
rect 23664 47660 23716 47666
rect 23664 47602 23716 47608
rect 23572 47048 23624 47054
rect 23572 46990 23624 46996
rect 23400 45526 23520 45554
rect 23296 45416 23348 45422
rect 23296 45358 23348 45364
rect 23308 44878 23336 45358
rect 23296 44872 23348 44878
rect 23296 44814 23348 44820
rect 23296 44736 23348 44742
rect 23296 44678 23348 44684
rect 23308 44334 23336 44678
rect 23296 44328 23348 44334
rect 23296 44270 23348 44276
rect 23204 43988 23256 43994
rect 23204 43930 23256 43936
rect 23020 43716 23072 43722
rect 23020 43658 23072 43664
rect 23400 43314 23428 45526
rect 23480 45416 23532 45422
rect 23480 45358 23532 45364
rect 23492 45257 23520 45358
rect 23478 45248 23534 45257
rect 23478 45183 23534 45192
rect 23492 44878 23520 45183
rect 23480 44872 23532 44878
rect 23480 44814 23532 44820
rect 23584 43450 23612 46990
rect 23676 46578 23704 47602
rect 23756 47524 23808 47530
rect 23756 47466 23808 47472
rect 23768 47054 23796 47466
rect 23860 47258 23888 49200
rect 23848 47252 23900 47258
rect 23848 47194 23900 47200
rect 23848 47116 23900 47122
rect 23848 47058 23900 47064
rect 23756 47048 23808 47054
rect 23756 46990 23808 46996
rect 23860 46714 23888 47058
rect 23848 46708 23900 46714
rect 23848 46650 23900 46656
rect 23664 46572 23716 46578
rect 23664 46514 23716 46520
rect 23756 46368 23808 46374
rect 23756 46310 23808 46316
rect 23664 46028 23716 46034
rect 23664 45970 23716 45976
rect 23676 44946 23704 45970
rect 23768 45490 23796 46310
rect 23952 46102 23980 49286
rect 24214 49200 24270 49286
rect 24582 49200 24638 50000
rect 24950 49200 25006 50000
rect 25318 49200 25374 50000
rect 25686 49200 25742 50000
rect 26054 49200 26110 50000
rect 26422 49200 26478 50000
rect 26790 49200 26846 50000
rect 27158 49314 27214 50000
rect 27158 49286 27292 49314
rect 27158 49200 27214 49286
rect 24032 47456 24084 47462
rect 24032 47398 24084 47404
rect 24044 47054 24072 47398
rect 24032 47048 24084 47054
rect 24032 46990 24084 46996
rect 24032 46572 24084 46578
rect 24032 46514 24084 46520
rect 24216 46572 24268 46578
rect 24216 46514 24268 46520
rect 24492 46572 24544 46578
rect 24492 46514 24544 46520
rect 23940 46096 23992 46102
rect 23940 46038 23992 46044
rect 24044 45830 24072 46514
rect 24032 45824 24084 45830
rect 24032 45766 24084 45772
rect 24044 45626 24072 45766
rect 24032 45620 24084 45626
rect 24032 45562 24084 45568
rect 23756 45484 23808 45490
rect 23756 45426 23808 45432
rect 23768 45082 23796 45426
rect 23756 45076 23808 45082
rect 23756 45018 23808 45024
rect 23664 44940 23716 44946
rect 23664 44882 23716 44888
rect 24228 44538 24256 46514
rect 24308 46504 24360 46510
rect 24306 46472 24308 46481
rect 24360 46472 24362 46481
rect 24306 46407 24362 46416
rect 24308 45280 24360 45286
rect 24308 45222 24360 45228
rect 24320 44742 24348 45222
rect 24308 44736 24360 44742
rect 24308 44678 24360 44684
rect 23848 44532 23900 44538
rect 23848 44474 23900 44480
rect 24216 44532 24268 44538
rect 24216 44474 24268 44480
rect 23756 44396 23808 44402
rect 23756 44338 23808 44344
rect 23768 43994 23796 44338
rect 23756 43988 23808 43994
rect 23756 43930 23808 43936
rect 23572 43444 23624 43450
rect 23572 43386 23624 43392
rect 23860 43314 23888 44474
rect 23940 44192 23992 44198
rect 23940 44134 23992 44140
rect 23952 43790 23980 44134
rect 24504 43858 24532 46514
rect 24596 45948 24624 49200
rect 24676 46980 24728 46986
rect 24676 46922 24728 46928
rect 24688 46578 24716 46922
rect 24860 46640 24912 46646
rect 24858 46608 24860 46617
rect 24912 46608 24914 46617
rect 24676 46572 24728 46578
rect 24676 46514 24728 46520
rect 24768 46572 24820 46578
rect 24964 46594 24992 49200
rect 25228 46640 25280 46646
rect 24964 46566 25084 46594
rect 25228 46582 25280 46588
rect 24858 46543 24914 46552
rect 24768 46514 24820 46520
rect 24780 46034 24808 46514
rect 24768 46028 24820 46034
rect 24768 45970 24820 45976
rect 24596 45920 24716 45948
rect 24584 44872 24636 44878
rect 24584 44814 24636 44820
rect 24596 44198 24624 44814
rect 24584 44192 24636 44198
rect 24584 44134 24636 44140
rect 24492 43852 24544 43858
rect 24492 43794 24544 43800
rect 23940 43784 23992 43790
rect 23940 43726 23992 43732
rect 23388 43308 23440 43314
rect 23388 43250 23440 43256
rect 23848 43308 23900 43314
rect 23848 43250 23900 43256
rect 24032 43308 24084 43314
rect 24032 43250 24084 43256
rect 22652 42764 22704 42770
rect 22652 42706 22704 42712
rect 24044 42566 24072 43250
rect 24688 42770 24716 45920
rect 24872 45490 24900 46543
rect 24952 46436 25004 46442
rect 24952 46378 25004 46384
rect 24964 46170 24992 46378
rect 24952 46164 25004 46170
rect 24952 46106 25004 46112
rect 24860 45484 24912 45490
rect 24912 45444 24992 45472
rect 24860 45426 24912 45432
rect 24768 45280 24820 45286
rect 24768 45222 24820 45228
rect 24780 44402 24808 45222
rect 24860 44872 24912 44878
rect 24860 44814 24912 44820
rect 24768 44396 24820 44402
rect 24768 44338 24820 44344
rect 24780 43790 24808 44338
rect 24768 43784 24820 43790
rect 24768 43726 24820 43732
rect 24780 43382 24808 43726
rect 24872 43654 24900 44814
rect 24860 43648 24912 43654
rect 24860 43590 24912 43596
rect 24872 43450 24900 43590
rect 24860 43444 24912 43450
rect 24860 43386 24912 43392
rect 24768 43376 24820 43382
rect 24768 43318 24820 43324
rect 24964 42906 24992 45444
rect 25056 43994 25084 46566
rect 25240 46510 25268 46582
rect 25228 46504 25280 46510
rect 25228 46446 25280 46452
rect 25136 46368 25188 46374
rect 25136 46310 25188 46316
rect 25148 46102 25176 46310
rect 25240 46102 25268 46446
rect 25136 46096 25188 46102
rect 25136 46038 25188 46044
rect 25228 46096 25280 46102
rect 25228 46038 25280 46044
rect 25136 45960 25188 45966
rect 25136 45902 25188 45908
rect 25148 44470 25176 45902
rect 25332 45558 25360 49200
rect 25700 47666 25728 49200
rect 25688 47660 25740 47666
rect 25688 47602 25740 47608
rect 26068 47258 26096 49200
rect 26056 47252 26108 47258
rect 26056 47194 26108 47200
rect 26436 47054 26464 49200
rect 26804 47190 26832 49200
rect 26792 47184 26844 47190
rect 26792 47126 26844 47132
rect 25688 47048 25740 47054
rect 25688 46990 25740 46996
rect 25872 47048 25924 47054
rect 25872 46990 25924 46996
rect 26148 47048 26200 47054
rect 26148 46990 26200 46996
rect 26424 47048 26476 47054
rect 26424 46990 26476 46996
rect 27160 47048 27212 47054
rect 27160 46990 27212 46996
rect 25504 46912 25556 46918
rect 25504 46854 25556 46860
rect 25516 46034 25544 46854
rect 25700 46714 25728 46990
rect 25688 46708 25740 46714
rect 25884 46696 25912 46990
rect 25964 46708 26016 46714
rect 25884 46668 25964 46696
rect 25688 46650 25740 46656
rect 25964 46650 26016 46656
rect 25872 46572 25924 46578
rect 25872 46514 25924 46520
rect 25884 46102 25912 46514
rect 25872 46096 25924 46102
rect 25872 46038 25924 46044
rect 25504 46028 25556 46034
rect 25504 45970 25556 45976
rect 25320 45552 25372 45558
rect 25372 45512 25452 45540
rect 25320 45494 25372 45500
rect 25320 44872 25372 44878
rect 25320 44814 25372 44820
rect 25136 44464 25188 44470
rect 25136 44406 25188 44412
rect 25332 44402 25360 44814
rect 25320 44396 25372 44402
rect 25320 44338 25372 44344
rect 25136 44260 25188 44266
rect 25136 44202 25188 44208
rect 25044 43988 25096 43994
rect 25044 43930 25096 43936
rect 25148 43858 25176 44202
rect 25136 43852 25188 43858
rect 25136 43794 25188 43800
rect 25148 43314 25176 43794
rect 25332 43722 25360 44338
rect 25424 44198 25452 45512
rect 25780 45484 25832 45490
rect 25780 45426 25832 45432
rect 25504 45416 25556 45422
rect 25504 45358 25556 45364
rect 25412 44192 25464 44198
rect 25412 44134 25464 44140
rect 25320 43716 25372 43722
rect 25320 43658 25372 43664
rect 25332 43314 25360 43658
rect 25136 43308 25188 43314
rect 25136 43250 25188 43256
rect 25320 43308 25372 43314
rect 25320 43250 25372 43256
rect 25516 43178 25544 45358
rect 25792 44538 25820 45426
rect 25884 44878 25912 46038
rect 25976 45082 26004 46650
rect 26160 46578 26188 46990
rect 26422 46608 26478 46617
rect 26148 46572 26200 46578
rect 26422 46543 26478 46552
rect 27068 46572 27120 46578
rect 26148 46514 26200 46520
rect 26436 46510 26464 46543
rect 27068 46514 27120 46520
rect 26424 46504 26476 46510
rect 26424 46446 26476 46452
rect 26068 45966 26096 45997
rect 26056 45960 26108 45966
rect 26054 45928 26056 45937
rect 26700 45960 26752 45966
rect 26108 45928 26110 45937
rect 26792 45960 26844 45966
rect 26700 45902 26752 45908
rect 26790 45928 26792 45937
rect 26844 45928 26846 45937
rect 26054 45863 26110 45872
rect 26068 45626 26096 45863
rect 26238 45656 26294 45665
rect 26056 45620 26108 45626
rect 26238 45591 26240 45600
rect 26056 45562 26108 45568
rect 26292 45591 26294 45600
rect 26240 45562 26292 45568
rect 26238 45248 26294 45257
rect 26238 45183 26294 45192
rect 25964 45076 26016 45082
rect 25964 45018 26016 45024
rect 25872 44872 25924 44878
rect 25872 44814 25924 44820
rect 25884 44538 25912 44814
rect 25780 44532 25832 44538
rect 25780 44474 25832 44480
rect 25872 44532 25924 44538
rect 25872 44474 25924 44480
rect 25976 44470 26004 45018
rect 26252 45014 26280 45183
rect 26424 45076 26476 45082
rect 26424 45018 26476 45024
rect 26240 45008 26292 45014
rect 26436 44985 26464 45018
rect 26240 44950 26292 44956
rect 26422 44976 26478 44985
rect 26422 44911 26478 44920
rect 26608 44736 26660 44742
rect 26608 44678 26660 44684
rect 25964 44464 26016 44470
rect 25964 44406 26016 44412
rect 26620 44402 26648 44678
rect 25596 44396 25648 44402
rect 25596 44338 25648 44344
rect 26608 44396 26660 44402
rect 26608 44338 26660 44344
rect 25608 43858 25636 44338
rect 26620 43858 26648 44338
rect 26712 43994 26740 45902
rect 26790 45863 26846 45872
rect 26884 44736 26936 44742
rect 26884 44678 26936 44684
rect 26896 44470 26924 44678
rect 26884 44464 26936 44470
rect 26884 44406 26936 44412
rect 26700 43988 26752 43994
rect 26700 43930 26752 43936
rect 25596 43852 25648 43858
rect 25596 43794 25648 43800
rect 26608 43852 26660 43858
rect 26608 43794 26660 43800
rect 25608 43450 25636 43794
rect 26896 43790 26924 44406
rect 26884 43784 26936 43790
rect 26884 43726 26936 43732
rect 25596 43444 25648 43450
rect 25596 43386 25648 43392
rect 25780 43308 25832 43314
rect 25780 43250 25832 43256
rect 26792 43308 26844 43314
rect 26792 43250 26844 43256
rect 25504 43172 25556 43178
rect 25504 43114 25556 43120
rect 24952 42900 25004 42906
rect 24952 42842 25004 42848
rect 24676 42764 24728 42770
rect 24676 42706 24728 42712
rect 21916 42560 21968 42566
rect 21916 42502 21968 42508
rect 24032 42560 24084 42566
rect 24032 42502 24084 42508
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 21928 42022 21956 42502
rect 24044 42362 24072 42502
rect 25792 42362 25820 43250
rect 26804 42906 26832 43250
rect 27080 42906 27108 46514
rect 26792 42900 26844 42906
rect 26792 42842 26844 42848
rect 27068 42900 27120 42906
rect 27068 42842 27120 42848
rect 27172 42362 27200 46990
rect 27264 42770 27292 49286
rect 27526 49200 27582 50000
rect 27894 49200 27950 50000
rect 28262 49200 28318 50000
rect 28630 49314 28686 50000
rect 28630 49286 28856 49314
rect 28630 49200 28686 49286
rect 27342 46608 27398 46617
rect 27342 46543 27398 46552
rect 27356 46374 27384 46543
rect 27344 46368 27396 46374
rect 27344 46310 27396 46316
rect 27356 46170 27384 46310
rect 27344 46164 27396 46170
rect 27344 46106 27396 46112
rect 27356 45830 27384 46106
rect 27344 45824 27396 45830
rect 27344 45766 27396 45772
rect 27356 45626 27384 45766
rect 27540 45665 27568 49200
rect 27620 47048 27672 47054
rect 27620 46990 27672 46996
rect 27526 45656 27582 45665
rect 27344 45620 27396 45626
rect 27526 45591 27582 45600
rect 27344 45562 27396 45568
rect 27632 45490 27660 46990
rect 27802 46472 27858 46481
rect 27802 46407 27858 46416
rect 27816 46374 27844 46407
rect 27804 46368 27856 46374
rect 27804 46310 27856 46316
rect 27620 45484 27672 45490
rect 27620 45426 27672 45432
rect 27620 45348 27672 45354
rect 27620 45290 27672 45296
rect 27632 44946 27660 45290
rect 27620 44940 27672 44946
rect 27620 44882 27672 44888
rect 27528 44872 27580 44878
rect 27528 44814 27580 44820
rect 27436 44736 27488 44742
rect 27436 44678 27488 44684
rect 27344 44328 27396 44334
rect 27344 44270 27396 44276
rect 27356 43994 27384 44270
rect 27344 43988 27396 43994
rect 27344 43930 27396 43936
rect 27356 43178 27384 43930
rect 27344 43172 27396 43178
rect 27344 43114 27396 43120
rect 27448 43110 27476 44678
rect 27540 44198 27568 44814
rect 27528 44192 27580 44198
rect 27528 44134 27580 44140
rect 27540 43450 27568 44134
rect 27528 43444 27580 43450
rect 27528 43386 27580 43392
rect 27632 43382 27660 44882
rect 27804 44872 27856 44878
rect 27804 44814 27856 44820
rect 27816 44402 27844 44814
rect 27804 44396 27856 44402
rect 27804 44338 27856 44344
rect 27620 43376 27672 43382
rect 27620 43318 27672 43324
rect 27908 43246 27936 49200
rect 28080 46640 28132 46646
rect 28080 46582 28132 46588
rect 27986 45928 28042 45937
rect 27986 45863 27988 45872
rect 28040 45863 28042 45872
rect 27988 45834 28040 45840
rect 28092 45626 28120 46582
rect 28172 46572 28224 46578
rect 28172 46514 28224 46520
rect 28184 46102 28212 46514
rect 28172 46096 28224 46102
rect 28172 46038 28224 46044
rect 28080 45620 28132 45626
rect 28080 45562 28132 45568
rect 28080 44736 28132 44742
rect 28080 44678 28132 44684
rect 28092 44470 28120 44678
rect 28080 44464 28132 44470
rect 28080 44406 28132 44412
rect 28184 43450 28212 46038
rect 28172 43444 28224 43450
rect 28172 43386 28224 43392
rect 27896 43240 27948 43246
rect 27896 43182 27948 43188
rect 27436 43104 27488 43110
rect 27436 43046 27488 43052
rect 28276 42770 28304 49200
rect 28448 46572 28500 46578
rect 28448 46514 28500 46520
rect 28540 46572 28592 46578
rect 28540 46514 28592 46520
rect 28460 46102 28488 46514
rect 28552 46170 28580 46514
rect 28540 46164 28592 46170
rect 28540 46106 28592 46112
rect 28448 46096 28500 46102
rect 28448 46038 28500 46044
rect 28356 45960 28408 45966
rect 28356 45902 28408 45908
rect 28368 45354 28396 45902
rect 28460 45490 28488 46038
rect 28724 46028 28776 46034
rect 28724 45970 28776 45976
rect 28736 45830 28764 45970
rect 28724 45824 28776 45830
rect 28644 45784 28724 45812
rect 28448 45484 28500 45490
rect 28448 45426 28500 45432
rect 28356 45348 28408 45354
rect 28356 45290 28408 45296
rect 28460 44810 28488 45426
rect 28644 45354 28672 45784
rect 28724 45766 28776 45772
rect 28724 45416 28776 45422
rect 28724 45358 28776 45364
rect 28632 45348 28684 45354
rect 28632 45290 28684 45296
rect 28540 44872 28592 44878
rect 28644 44860 28672 45290
rect 28736 44878 28764 45358
rect 28592 44832 28672 44860
rect 28724 44872 28776 44878
rect 28540 44814 28592 44820
rect 28724 44814 28776 44820
rect 28448 44804 28500 44810
rect 28448 44746 28500 44752
rect 28552 44538 28580 44814
rect 28540 44532 28592 44538
rect 28540 44474 28592 44480
rect 28828 43790 28856 49286
rect 28998 49200 29054 50000
rect 29366 49314 29422 50000
rect 29366 49286 29684 49314
rect 29366 49200 29422 49286
rect 28816 43784 28868 43790
rect 28816 43726 28868 43732
rect 27252 42764 27304 42770
rect 27252 42706 27304 42712
rect 28264 42764 28316 42770
rect 28264 42706 28316 42712
rect 27712 42696 27764 42702
rect 27712 42638 27764 42644
rect 27724 42401 27752 42638
rect 27804 42628 27856 42634
rect 27804 42570 27856 42576
rect 27710 42392 27766 42401
rect 24032 42356 24084 42362
rect 24032 42298 24084 42304
rect 25780 42356 25832 42362
rect 25780 42298 25832 42304
rect 27160 42356 27212 42362
rect 27710 42327 27712 42336
rect 27160 42298 27212 42304
rect 27764 42327 27766 42336
rect 27712 42298 27764 42304
rect 25136 42084 25188 42090
rect 25136 42026 25188 42032
rect 21916 42016 21968 42022
rect 21916 41958 21968 41964
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 25148 7546 25176 42026
rect 27816 41818 27844 42570
rect 28828 42362 28856 43726
rect 29012 43314 29040 49200
rect 29368 47048 29420 47054
rect 29368 46990 29420 46996
rect 29184 46980 29236 46986
rect 29184 46922 29236 46928
rect 29092 46640 29144 46646
rect 29092 46582 29144 46588
rect 29104 45082 29132 46582
rect 29196 46510 29224 46922
rect 29380 46578 29408 46990
rect 29368 46572 29420 46578
rect 29368 46514 29420 46520
rect 29184 46504 29236 46510
rect 29184 46446 29236 46452
rect 29196 46170 29224 46446
rect 29184 46164 29236 46170
rect 29184 46106 29236 46112
rect 29276 45484 29328 45490
rect 29276 45426 29328 45432
rect 29092 45076 29144 45082
rect 29092 45018 29144 45024
rect 29104 44266 29132 45018
rect 29288 44402 29316 45426
rect 29380 45014 29408 46514
rect 29552 45484 29604 45490
rect 29552 45426 29604 45432
rect 29460 45280 29512 45286
rect 29460 45222 29512 45228
rect 29368 45008 29420 45014
rect 29368 44950 29420 44956
rect 29472 44470 29500 45222
rect 29564 44878 29592 45426
rect 29552 44872 29604 44878
rect 29552 44814 29604 44820
rect 29460 44464 29512 44470
rect 29460 44406 29512 44412
rect 29276 44396 29328 44402
rect 29276 44338 29328 44344
rect 29184 44328 29236 44334
rect 29184 44270 29236 44276
rect 29092 44260 29144 44266
rect 29092 44202 29144 44208
rect 29196 43994 29224 44270
rect 29184 43988 29236 43994
rect 29184 43930 29236 43936
rect 29472 43858 29500 44406
rect 29460 43852 29512 43858
rect 29460 43794 29512 43800
rect 29656 43314 29684 49286
rect 29734 49200 29790 50000
rect 30102 49200 30158 50000
rect 30470 49200 30526 50000
rect 30838 49200 30894 50000
rect 31206 49314 31262 50000
rect 31206 49286 31340 49314
rect 31206 49200 31262 49286
rect 29748 47054 29776 49200
rect 29828 47456 29880 47462
rect 29828 47398 29880 47404
rect 30012 47456 30064 47462
rect 30012 47398 30064 47404
rect 29736 47048 29788 47054
rect 29736 46990 29788 46996
rect 29748 44470 29776 46990
rect 29840 46646 29868 47398
rect 29920 47048 29972 47054
rect 29920 46990 29972 46996
rect 29828 46640 29880 46646
rect 29828 46582 29880 46588
rect 29828 46096 29880 46102
rect 29828 46038 29880 46044
rect 29840 45937 29868 46038
rect 29826 45928 29882 45937
rect 29826 45863 29882 45872
rect 29840 44878 29868 45863
rect 29932 45422 29960 46990
rect 30024 45966 30052 47398
rect 30116 46714 30144 49200
rect 30288 47524 30340 47530
rect 30288 47466 30340 47472
rect 30104 46708 30156 46714
rect 30104 46650 30156 46656
rect 30300 46102 30328 47466
rect 30484 46594 30512 49200
rect 30852 46918 30880 49200
rect 30840 46912 30892 46918
rect 30840 46854 30892 46860
rect 30654 46608 30710 46617
rect 30484 46566 30604 46594
rect 30472 46436 30524 46442
rect 30472 46378 30524 46384
rect 30288 46096 30340 46102
rect 30288 46038 30340 46044
rect 30484 45966 30512 46378
rect 30012 45960 30064 45966
rect 30012 45902 30064 45908
rect 30472 45960 30524 45966
rect 30472 45902 30524 45908
rect 29920 45416 29972 45422
rect 29920 45358 29972 45364
rect 29828 44872 29880 44878
rect 29828 44814 29880 44820
rect 29736 44464 29788 44470
rect 29736 44406 29788 44412
rect 29932 43926 29960 45358
rect 30024 44860 30052 45902
rect 30472 45416 30524 45422
rect 30472 45358 30524 45364
rect 30484 45082 30512 45358
rect 30472 45076 30524 45082
rect 30472 45018 30524 45024
rect 30104 44872 30156 44878
rect 30024 44832 30104 44860
rect 30104 44814 30156 44820
rect 30012 44736 30064 44742
rect 30012 44678 30064 44684
rect 29920 43920 29972 43926
rect 29920 43862 29972 43868
rect 30024 43790 30052 44678
rect 30012 43784 30064 43790
rect 30012 43726 30064 43732
rect 30116 43382 30144 44814
rect 30196 44328 30248 44334
rect 30196 44270 30248 44276
rect 30104 43376 30156 43382
rect 30104 43318 30156 43324
rect 29000 43308 29052 43314
rect 29000 43250 29052 43256
rect 29644 43308 29696 43314
rect 29644 43250 29696 43256
rect 30116 42702 30144 43318
rect 30104 42696 30156 42702
rect 30104 42638 30156 42644
rect 29460 42628 29512 42634
rect 29460 42570 29512 42576
rect 29472 42362 29500 42570
rect 28816 42356 28868 42362
rect 28816 42298 28868 42304
rect 29460 42356 29512 42362
rect 29460 42298 29512 42304
rect 30116 42294 30144 42638
rect 30104 42288 30156 42294
rect 30104 42230 30156 42236
rect 27804 41812 27856 41818
rect 27804 41754 27856 41760
rect 30208 26234 30236 44270
rect 30576 43926 30604 46566
rect 30654 46543 30656 46552
rect 30708 46543 30710 46552
rect 30748 46572 30800 46578
rect 30656 46514 30708 46520
rect 30748 46514 30800 46520
rect 30668 45898 30696 46514
rect 30760 45966 30788 46514
rect 30748 45960 30800 45966
rect 30748 45902 30800 45908
rect 30656 45892 30708 45898
rect 30656 45834 30708 45840
rect 30760 45626 30788 45902
rect 30748 45620 30800 45626
rect 30748 45562 30800 45568
rect 30564 43920 30616 43926
rect 30564 43862 30616 43868
rect 31312 43314 31340 49286
rect 31574 49200 31630 50000
rect 31942 49200 31998 50000
rect 32310 49200 32366 50000
rect 32678 49200 32734 50000
rect 33046 49200 33102 50000
rect 33414 49200 33470 50000
rect 33782 49314 33838 50000
rect 33704 49286 33838 49314
rect 31392 45824 31444 45830
rect 31392 45766 31444 45772
rect 31404 45558 31432 45766
rect 31392 45552 31444 45558
rect 31392 45494 31444 45500
rect 31588 44418 31616 49200
rect 31956 47274 31984 49200
rect 31956 47246 32076 47274
rect 31760 47116 31812 47122
rect 31760 47058 31812 47064
rect 31944 47116 31996 47122
rect 31944 47058 31996 47064
rect 31668 46980 31720 46986
rect 31668 46922 31720 46928
rect 31680 46510 31708 46922
rect 31668 46504 31720 46510
rect 31668 46446 31720 46452
rect 31772 46102 31800 47058
rect 31852 46980 31904 46986
rect 31852 46922 31904 46928
rect 31864 46646 31892 46922
rect 31852 46640 31904 46646
rect 31852 46582 31904 46588
rect 31852 46504 31904 46510
rect 31850 46472 31852 46481
rect 31904 46472 31906 46481
rect 31850 46407 31906 46416
rect 31852 46368 31904 46374
rect 31852 46310 31904 46316
rect 31760 46096 31812 46102
rect 31760 46038 31812 46044
rect 31760 45960 31812 45966
rect 31760 45902 31812 45908
rect 31772 45286 31800 45902
rect 31864 45354 31892 46310
rect 31956 45830 31984 47058
rect 32048 46510 32076 47246
rect 32220 47048 32272 47054
rect 32220 46990 32272 46996
rect 32232 46918 32260 46990
rect 32220 46912 32272 46918
rect 32220 46854 32272 46860
rect 32036 46504 32088 46510
rect 32036 46446 32088 46452
rect 32048 46374 32076 46446
rect 32036 46368 32088 46374
rect 32036 46310 32088 46316
rect 32036 46096 32088 46102
rect 32036 46038 32088 46044
rect 31944 45824 31996 45830
rect 31944 45766 31996 45772
rect 31944 45552 31996 45558
rect 31944 45494 31996 45500
rect 31852 45348 31904 45354
rect 31852 45290 31904 45296
rect 31760 45280 31812 45286
rect 31760 45222 31812 45228
rect 31668 44872 31720 44878
rect 31772 44860 31800 45222
rect 31864 44946 31892 45290
rect 31956 45082 31984 45494
rect 31944 45076 31996 45082
rect 31944 45018 31996 45024
rect 32048 45014 32076 46038
rect 32128 46028 32180 46034
rect 32128 45970 32180 45976
rect 32036 45008 32088 45014
rect 32036 44950 32088 44956
rect 31852 44940 31904 44946
rect 31852 44882 31904 44888
rect 31720 44832 31800 44860
rect 31668 44814 31720 44820
rect 32140 44810 32168 45970
rect 32128 44804 32180 44810
rect 32128 44746 32180 44752
rect 31588 44390 31708 44418
rect 31576 44328 31628 44334
rect 31576 44270 31628 44276
rect 31588 43994 31616 44270
rect 31576 43988 31628 43994
rect 31576 43930 31628 43936
rect 31300 43308 31352 43314
rect 31300 43250 31352 43256
rect 31680 43246 31708 44390
rect 31668 43240 31720 43246
rect 31668 43182 31720 43188
rect 30656 43104 30708 43110
rect 30656 43046 30708 43052
rect 30668 42838 30696 43046
rect 30656 42832 30708 42838
rect 30656 42774 30708 42780
rect 32232 42770 32260 46854
rect 32324 45642 32352 49200
rect 32588 46504 32640 46510
rect 32588 46446 32640 46452
rect 32600 46170 32628 46446
rect 32588 46164 32640 46170
rect 32588 46106 32640 46112
rect 32324 45614 32444 45642
rect 32312 45484 32364 45490
rect 32312 45426 32364 45432
rect 32324 44538 32352 45426
rect 32312 44532 32364 44538
rect 32312 44474 32364 44480
rect 32416 43314 32444 45614
rect 32588 45484 32640 45490
rect 32588 45426 32640 45432
rect 32600 45082 32628 45426
rect 32588 45076 32640 45082
rect 32588 45018 32640 45024
rect 32496 44940 32548 44946
rect 32496 44882 32548 44888
rect 32508 44402 32536 44882
rect 32496 44396 32548 44402
rect 32496 44338 32548 44344
rect 32508 43790 32536 44338
rect 32600 43994 32628 45018
rect 32588 43988 32640 43994
rect 32588 43930 32640 43936
rect 32692 43858 32720 49200
rect 32956 46096 33008 46102
rect 32954 46064 32956 46073
rect 33008 46064 33010 46073
rect 32954 45999 33010 46008
rect 32956 45960 33008 45966
rect 32956 45902 33008 45908
rect 32968 45490 32996 45902
rect 33060 45642 33088 49200
rect 33232 47116 33284 47122
rect 33232 47058 33284 47064
rect 33244 46102 33272 47058
rect 33324 46912 33376 46918
rect 33324 46854 33376 46860
rect 33336 46102 33364 46854
rect 33232 46096 33284 46102
rect 33232 46038 33284 46044
rect 33324 46096 33376 46102
rect 33324 46038 33376 46044
rect 33060 45614 33180 45642
rect 32956 45484 33008 45490
rect 32956 45426 33008 45432
rect 32772 44872 32824 44878
rect 32772 44814 32824 44820
rect 32784 44334 32812 44814
rect 32772 44328 32824 44334
rect 32772 44270 32824 44276
rect 32680 43852 32732 43858
rect 32680 43794 32732 43800
rect 32496 43784 32548 43790
rect 32496 43726 32548 43732
rect 32784 43722 32812 44270
rect 32772 43716 32824 43722
rect 32772 43658 32824 43664
rect 33152 43314 33180 45614
rect 33244 45014 33272 46038
rect 33428 45642 33456 49200
rect 33704 46617 33732 49286
rect 33782 49200 33838 49286
rect 34150 49314 34206 50000
rect 34150 49286 34468 49314
rect 34150 49200 34206 49286
rect 33968 47116 34020 47122
rect 33968 47058 34020 47064
rect 34152 47116 34204 47122
rect 34152 47058 34204 47064
rect 33784 47048 33836 47054
rect 33784 46990 33836 46996
rect 33796 46714 33824 46990
rect 33784 46708 33836 46714
rect 33980 46696 34008 47058
rect 34060 46708 34112 46714
rect 33980 46668 34060 46696
rect 33784 46650 33836 46656
rect 34060 46650 34112 46656
rect 33506 46608 33562 46617
rect 33506 46543 33562 46552
rect 33690 46608 33746 46617
rect 34164 46578 34192 47058
rect 33690 46543 33746 46552
rect 33784 46572 33836 46578
rect 33520 46510 33548 46543
rect 33784 46514 33836 46520
rect 34152 46572 34204 46578
rect 34152 46514 34204 46520
rect 33508 46504 33560 46510
rect 33508 46446 33560 46452
rect 33796 46102 33824 46514
rect 33784 46096 33836 46102
rect 33784 46038 33836 46044
rect 34060 45960 34112 45966
rect 34164 45948 34192 46514
rect 34336 46368 34388 46374
rect 34336 46310 34388 46316
rect 34112 45920 34192 45948
rect 34060 45902 34112 45908
rect 33508 45892 33560 45898
rect 33508 45834 33560 45840
rect 33336 45614 33456 45642
rect 33232 45008 33284 45014
rect 33232 44950 33284 44956
rect 32404 43308 32456 43314
rect 32404 43250 32456 43256
rect 33140 43308 33192 43314
rect 33140 43250 33192 43256
rect 33152 42906 33180 43250
rect 33336 43246 33364 45614
rect 33416 45552 33468 45558
rect 33414 45520 33416 45529
rect 33468 45520 33470 45529
rect 33414 45455 33470 45464
rect 33520 45082 33548 45834
rect 33968 45824 34020 45830
rect 33782 45792 33838 45801
rect 33968 45766 34020 45772
rect 33782 45727 33838 45736
rect 33796 45558 33824 45727
rect 33980 45558 34008 45766
rect 33784 45552 33836 45558
rect 33704 45512 33784 45540
rect 33600 45348 33652 45354
rect 33600 45290 33652 45296
rect 33508 45076 33560 45082
rect 33508 45018 33560 45024
rect 33520 43790 33548 45018
rect 33612 44538 33640 45290
rect 33600 44532 33652 44538
rect 33600 44474 33652 44480
rect 33704 43790 33732 45512
rect 33784 45494 33836 45500
rect 33968 45552 34020 45558
rect 33968 45494 34020 45500
rect 34060 45416 34112 45422
rect 34060 45358 34112 45364
rect 33784 45076 33836 45082
rect 33784 45018 33836 45024
rect 33508 43784 33560 43790
rect 33508 43726 33560 43732
rect 33692 43784 33744 43790
rect 33692 43726 33744 43732
rect 33796 43450 33824 45018
rect 34072 43994 34100 45358
rect 34164 44810 34192 45920
rect 34348 45558 34376 46310
rect 34440 45642 34468 49286
rect 34518 49200 34574 50000
rect 34886 49200 34942 50000
rect 35254 49200 35310 50000
rect 35622 49200 35678 50000
rect 35990 49200 36046 50000
rect 36358 49200 36414 50000
rect 36726 49200 36782 50000
rect 37094 49200 37150 50000
rect 37462 49314 37518 50000
rect 37292 49286 37518 49314
rect 34532 45966 34560 49200
rect 34900 47512 34928 49200
rect 34808 47484 34928 47512
rect 34808 46714 34836 47484
rect 35268 47410 35296 49200
rect 35268 47382 35388 47410
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 35360 46918 35388 47382
rect 35440 47252 35492 47258
rect 35440 47194 35492 47200
rect 35348 46912 35400 46918
rect 35348 46854 35400 46860
rect 34796 46708 34848 46714
rect 34796 46650 34848 46656
rect 34796 46368 34848 46374
rect 34796 46310 34848 46316
rect 34520 45960 34572 45966
rect 34520 45902 34572 45908
rect 34612 45892 34664 45898
rect 34612 45834 34664 45840
rect 34440 45614 34560 45642
rect 34624 45626 34652 45834
rect 34336 45552 34388 45558
rect 34336 45494 34388 45500
rect 34152 44804 34204 44810
rect 34152 44746 34204 44752
rect 34060 43988 34112 43994
rect 34060 43930 34112 43936
rect 33784 43444 33836 43450
rect 33784 43386 33836 43392
rect 34532 43314 34560 45614
rect 34612 45620 34664 45626
rect 34612 45562 34664 45568
rect 34624 45014 34652 45562
rect 34612 45008 34664 45014
rect 34612 44950 34664 44956
rect 34624 44826 34652 44950
rect 34624 44798 34744 44826
rect 34612 44736 34664 44742
rect 34612 44678 34664 44684
rect 34624 44538 34652 44678
rect 34612 44532 34664 44538
rect 34612 44474 34664 44480
rect 34624 44334 34652 44474
rect 34612 44328 34664 44334
rect 34612 44270 34664 44276
rect 34716 43722 34744 44798
rect 34808 44470 34836 46310
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 35452 46034 35480 47194
rect 35532 46504 35584 46510
rect 35532 46446 35584 46452
rect 35544 46374 35572 46446
rect 35532 46368 35584 46374
rect 35532 46310 35584 46316
rect 35636 46322 35664 49200
rect 36004 47190 36032 49200
rect 35992 47184 36044 47190
rect 35992 47126 36044 47132
rect 36084 47048 36136 47054
rect 36084 46990 36136 46996
rect 35992 46368 36044 46374
rect 35544 46034 35572 46310
rect 35636 46294 35940 46322
rect 35992 46310 36044 46316
rect 34980 46028 35032 46034
rect 34980 45970 35032 45976
rect 35440 46028 35492 46034
rect 35440 45970 35492 45976
rect 35532 46028 35584 46034
rect 35532 45970 35584 45976
rect 35808 46028 35860 46034
rect 35808 45970 35860 45976
rect 34992 45937 35020 45970
rect 35716 45960 35768 45966
rect 34978 45928 35034 45937
rect 34978 45863 35034 45872
rect 35636 45920 35716 45948
rect 35532 45620 35584 45626
rect 35532 45562 35584 45568
rect 35440 45484 35492 45490
rect 35440 45426 35492 45432
rect 35348 45280 35400 45286
rect 35348 45222 35400 45228
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 35360 45014 35388 45222
rect 35348 45008 35400 45014
rect 35348 44950 35400 44956
rect 35072 44872 35124 44878
rect 35072 44814 35124 44820
rect 34980 44804 35032 44810
rect 34980 44746 35032 44752
rect 34992 44538 35020 44746
rect 34980 44532 35032 44538
rect 34980 44474 35032 44480
rect 34796 44464 34848 44470
rect 34796 44406 34848 44412
rect 35084 44198 35112 44814
rect 35360 44402 35388 44950
rect 35452 44538 35480 45426
rect 35440 44532 35492 44538
rect 35440 44474 35492 44480
rect 35348 44396 35400 44402
rect 35348 44338 35400 44344
rect 35072 44192 35124 44198
rect 35072 44134 35124 44140
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 35452 43994 35480 44474
rect 35440 43988 35492 43994
rect 35440 43930 35492 43936
rect 34704 43716 34756 43722
rect 34704 43658 34756 43664
rect 35440 43716 35492 43722
rect 35544 43704 35572 45562
rect 35636 44810 35664 45920
rect 35716 45902 35768 45908
rect 35716 45824 35768 45830
rect 35716 45766 35768 45772
rect 35728 45558 35756 45766
rect 35820 45665 35848 45970
rect 35806 45656 35862 45665
rect 35806 45591 35862 45600
rect 35716 45552 35768 45558
rect 35716 45494 35768 45500
rect 35808 45484 35860 45490
rect 35808 45426 35860 45432
rect 35716 45280 35768 45286
rect 35716 45222 35768 45228
rect 35624 44804 35676 44810
rect 35624 44746 35676 44752
rect 35728 44470 35756 45222
rect 35820 44742 35848 45426
rect 35808 44736 35860 44742
rect 35808 44678 35860 44684
rect 35716 44464 35768 44470
rect 35716 44406 35768 44412
rect 35716 44192 35768 44198
rect 35716 44134 35768 44140
rect 35728 43994 35756 44134
rect 35716 43988 35768 43994
rect 35716 43930 35768 43936
rect 35820 43722 35848 44678
rect 35912 43994 35940 46294
rect 36004 45966 36032 46310
rect 35992 45960 36044 45966
rect 35992 45902 36044 45908
rect 36096 45506 36124 46990
rect 36268 46572 36320 46578
rect 36268 46514 36320 46520
rect 36174 45656 36230 45665
rect 36280 45626 36308 46514
rect 36372 45626 36400 49200
rect 36636 46912 36688 46918
rect 36636 46854 36688 46860
rect 36452 46504 36504 46510
rect 36504 46464 36584 46492
rect 36452 46446 36504 46452
rect 36556 46034 36584 46464
rect 36544 46028 36596 46034
rect 36544 45970 36596 45976
rect 36452 45960 36504 45966
rect 36452 45902 36504 45908
rect 36464 45801 36492 45902
rect 36450 45792 36506 45801
rect 36450 45727 36506 45736
rect 36174 45591 36230 45600
rect 36268 45620 36320 45626
rect 36004 45490 36124 45506
rect 36188 45490 36216 45591
rect 36268 45562 36320 45568
rect 36360 45620 36412 45626
rect 36360 45562 36412 45568
rect 35992 45484 36124 45490
rect 36044 45478 36124 45484
rect 35992 45426 36044 45432
rect 36096 44266 36124 45478
rect 36176 45484 36228 45490
rect 36176 45426 36228 45432
rect 36464 45336 36492 45727
rect 36544 45348 36596 45354
rect 36464 45308 36544 45336
rect 36544 45290 36596 45296
rect 36268 44940 36320 44946
rect 36268 44882 36320 44888
rect 36280 44402 36308 44882
rect 36268 44396 36320 44402
rect 36268 44338 36320 44344
rect 36084 44260 36136 44266
rect 36084 44202 36136 44208
rect 36648 43994 36676 46854
rect 36740 45898 36768 49200
rect 36912 46912 36964 46918
rect 36912 46854 36964 46860
rect 36728 45892 36780 45898
rect 36728 45834 36780 45840
rect 36924 44810 36952 46854
rect 37108 46442 37136 49200
rect 37292 46986 37320 49286
rect 37462 49200 37518 49286
rect 37830 49200 37886 50000
rect 38198 49200 38254 50000
rect 38566 49314 38622 50000
rect 38566 49286 38700 49314
rect 38566 49200 38622 49286
rect 37844 47530 37872 49200
rect 37832 47524 37884 47530
rect 37832 47466 37884 47472
rect 37830 47288 37886 47297
rect 37830 47223 37886 47232
rect 37844 47122 37872 47223
rect 38014 47152 38070 47161
rect 37556 47116 37608 47122
rect 37556 47058 37608 47064
rect 37832 47116 37884 47122
rect 38014 47087 38070 47096
rect 37832 47058 37884 47064
rect 37280 46980 37332 46986
rect 37280 46922 37332 46928
rect 37372 46980 37424 46986
rect 37372 46922 37424 46928
rect 37292 46889 37320 46922
rect 37278 46880 37334 46889
rect 37278 46815 37334 46824
rect 37384 46646 37412 46922
rect 37464 46912 37516 46918
rect 37464 46854 37516 46860
rect 37372 46640 37424 46646
rect 37372 46582 37424 46588
rect 37096 46436 37148 46442
rect 37096 46378 37148 46384
rect 37384 45966 37412 46582
rect 37476 46578 37504 46854
rect 37464 46572 37516 46578
rect 37464 46514 37516 46520
rect 37568 46374 37596 47058
rect 37648 47048 37700 47054
rect 37648 46990 37700 46996
rect 37660 46481 37688 46990
rect 37646 46472 37702 46481
rect 37646 46407 37702 46416
rect 37556 46368 37608 46374
rect 37556 46310 37608 46316
rect 37372 45960 37424 45966
rect 37372 45902 37424 45908
rect 37568 45665 37596 46310
rect 37554 45656 37610 45665
rect 37554 45591 37610 45600
rect 37372 45484 37424 45490
rect 37372 45426 37424 45432
rect 37384 44878 37412 45426
rect 37568 45422 37596 45591
rect 37464 45416 37516 45422
rect 37462 45384 37464 45393
rect 37556 45416 37608 45422
rect 37516 45384 37518 45393
rect 37556 45358 37608 45364
rect 37462 45319 37518 45328
rect 37660 45082 37688 46407
rect 37924 46368 37976 46374
rect 37924 46310 37976 46316
rect 37936 46170 37964 46310
rect 37924 46164 37976 46170
rect 37924 46106 37976 46112
rect 38028 45966 38056 47087
rect 38108 46572 38160 46578
rect 38108 46514 38160 46520
rect 38120 46170 38148 46514
rect 38108 46164 38160 46170
rect 38108 46106 38160 46112
rect 38016 45960 38068 45966
rect 38016 45902 38068 45908
rect 37648 45076 37700 45082
rect 37648 45018 37700 45024
rect 37464 44940 37516 44946
rect 37464 44882 37516 44888
rect 37372 44872 37424 44878
rect 37372 44814 37424 44820
rect 36912 44804 36964 44810
rect 36912 44746 36964 44752
rect 36820 44736 36872 44742
rect 36820 44678 36872 44684
rect 36832 44384 36860 44678
rect 36924 44538 36952 44746
rect 37476 44538 37504 44882
rect 38028 44878 38056 45902
rect 38212 45626 38240 49200
rect 38384 47524 38436 47530
rect 38384 47466 38436 47472
rect 38396 46170 38424 47466
rect 38474 47016 38530 47025
rect 38474 46951 38530 46960
rect 38488 46510 38516 46951
rect 38672 46918 38700 49286
rect 38934 49200 38990 50000
rect 39302 49200 39358 50000
rect 39670 49314 39726 50000
rect 40038 49314 40094 50000
rect 39670 49286 39988 49314
rect 39670 49200 39726 49286
rect 38844 47048 38896 47054
rect 38842 47016 38844 47025
rect 38896 47016 38898 47025
rect 38842 46951 38898 46960
rect 38660 46912 38712 46918
rect 38660 46854 38712 46860
rect 38476 46504 38528 46510
rect 38476 46446 38528 46452
rect 38384 46164 38436 46170
rect 38384 46106 38436 46112
rect 38488 46102 38516 46446
rect 38292 46096 38344 46102
rect 38292 46038 38344 46044
rect 38476 46096 38528 46102
rect 38476 46038 38528 46044
rect 38568 46096 38620 46102
rect 38568 46038 38620 46044
rect 38108 45620 38160 45626
rect 38108 45562 38160 45568
rect 38200 45620 38252 45626
rect 38200 45562 38252 45568
rect 38120 44878 38148 45562
rect 38016 44872 38068 44878
rect 38016 44814 38068 44820
rect 38108 44872 38160 44878
rect 38108 44814 38160 44820
rect 37924 44804 37976 44810
rect 37924 44746 37976 44752
rect 36912 44532 36964 44538
rect 36912 44474 36964 44480
rect 37464 44532 37516 44538
rect 37464 44474 37516 44480
rect 36912 44396 36964 44402
rect 36832 44356 36912 44384
rect 36912 44338 36964 44344
rect 37936 44334 37964 44746
rect 38120 44538 38148 44814
rect 38304 44810 38332 46038
rect 38292 44804 38344 44810
rect 38292 44746 38344 44752
rect 38488 44742 38516 46038
rect 38580 45558 38608 46038
rect 38568 45552 38620 45558
rect 38568 45494 38620 45500
rect 38476 44736 38528 44742
rect 38476 44678 38528 44684
rect 38108 44532 38160 44538
rect 38108 44474 38160 44480
rect 37924 44328 37976 44334
rect 37924 44270 37976 44276
rect 38488 44266 38516 44678
rect 38580 44402 38608 45494
rect 38672 45082 38700 46854
rect 38844 46572 38896 46578
rect 38844 46514 38896 46520
rect 38752 46436 38804 46442
rect 38752 46378 38804 46384
rect 38660 45076 38712 45082
rect 38660 45018 38712 45024
rect 38764 44946 38792 46378
rect 38856 45966 38884 46514
rect 38948 46170 38976 49200
rect 39118 46608 39174 46617
rect 39118 46543 39120 46552
rect 39172 46543 39174 46552
rect 39120 46514 39172 46520
rect 38936 46164 38988 46170
rect 38936 46106 38988 46112
rect 38844 45960 38896 45966
rect 38844 45902 38896 45908
rect 39212 45892 39264 45898
rect 39212 45834 39264 45840
rect 39224 45422 39252 45834
rect 39316 45626 39344 49200
rect 39960 47104 39988 49286
rect 40038 49286 40356 49314
rect 40038 49200 40094 49286
rect 40222 47152 40278 47161
rect 40040 47116 40092 47122
rect 39960 47076 40040 47104
rect 40222 47087 40278 47096
rect 40040 47058 40092 47064
rect 39304 45620 39356 45626
rect 39304 45562 39356 45568
rect 39212 45416 39264 45422
rect 39212 45358 39264 45364
rect 40052 45082 40080 47058
rect 40236 47054 40264 47087
rect 40224 47048 40276 47054
rect 40224 46990 40276 46996
rect 40328 46102 40356 49286
rect 40406 49200 40462 50000
rect 40774 49314 40830 50000
rect 40774 49286 40908 49314
rect 40774 49200 40830 49286
rect 40316 46096 40368 46102
rect 40316 46038 40368 46044
rect 40420 45490 40448 49200
rect 40880 46578 40908 49286
rect 41142 49200 41198 50000
rect 41510 49200 41566 50000
rect 41878 49314 41934 50000
rect 41878 49286 42196 49314
rect 41878 49200 41934 49286
rect 40868 46572 40920 46578
rect 40868 46514 40920 46520
rect 40408 45484 40460 45490
rect 40408 45426 40460 45432
rect 40880 45082 40908 46514
rect 41156 46170 41184 49200
rect 41524 46442 41552 49200
rect 41604 47116 41656 47122
rect 41604 47058 41656 47064
rect 41512 46436 41564 46442
rect 41512 46378 41564 46384
rect 41144 46164 41196 46170
rect 41144 46106 41196 46112
rect 41616 45422 41644 47058
rect 41972 46980 42024 46986
rect 41972 46922 42024 46928
rect 41984 46889 42012 46922
rect 42168 46918 42196 49286
rect 42246 49200 42302 50000
rect 42614 49200 42670 50000
rect 42982 49200 43038 50000
rect 43350 49200 43406 50000
rect 43718 49200 43774 50000
rect 44086 49200 44142 50000
rect 44454 49200 44510 50000
rect 44822 49200 44878 50000
rect 45190 49200 45246 50000
rect 45558 49314 45614 50000
rect 45558 49286 45876 49314
rect 45558 49200 45614 49286
rect 42156 46912 42208 46918
rect 41970 46880 42026 46889
rect 42156 46854 42208 46860
rect 41970 46815 42026 46824
rect 42260 46170 42288 49200
rect 42628 46578 42656 49200
rect 42996 47054 43024 49200
rect 42984 47048 43036 47054
rect 42984 46990 43036 46996
rect 43260 46980 43312 46986
rect 43260 46922 43312 46928
rect 42616 46572 42668 46578
rect 42616 46514 42668 46520
rect 43272 46170 43300 46922
rect 43364 46578 43392 49200
rect 43444 47456 43496 47462
rect 43444 47398 43496 47404
rect 43456 47258 43484 47398
rect 43444 47252 43496 47258
rect 43444 47194 43496 47200
rect 43352 46572 43404 46578
rect 43352 46514 43404 46520
rect 43732 46510 43760 49200
rect 44100 47410 44128 49200
rect 44100 47382 44220 47410
rect 44192 47054 44220 47382
rect 44270 47288 44326 47297
rect 44270 47223 44272 47232
rect 44324 47223 44326 47232
rect 44272 47194 44324 47200
rect 43812 47048 43864 47054
rect 43812 46990 43864 46996
rect 44180 47048 44232 47054
rect 44180 46990 44232 46996
rect 43720 46504 43772 46510
rect 43720 46446 43772 46452
rect 43824 46170 43852 46990
rect 44192 46170 44220 46990
rect 44468 46578 44496 49200
rect 44836 46918 44864 49200
rect 45204 47054 45232 49200
rect 45192 47048 45244 47054
rect 45192 46990 45244 46996
rect 44824 46912 44876 46918
rect 44824 46854 44876 46860
rect 44456 46572 44508 46578
rect 44456 46514 44508 46520
rect 45204 46170 45232 46990
rect 45848 46578 45876 49286
rect 45926 49200 45982 50000
rect 45940 47258 45968 49200
rect 45928 47252 45980 47258
rect 45928 47194 45980 47200
rect 45836 46572 45888 46578
rect 45836 46514 45888 46520
rect 42248 46164 42300 46170
rect 42248 46106 42300 46112
rect 43260 46164 43312 46170
rect 43260 46106 43312 46112
rect 43812 46164 43864 46170
rect 43812 46106 43864 46112
rect 44180 46164 44232 46170
rect 44180 46106 44232 46112
rect 45192 46164 45244 46170
rect 45192 46106 45244 46112
rect 41604 45416 41656 45422
rect 41604 45358 41656 45364
rect 40040 45076 40092 45082
rect 40040 45018 40092 45024
rect 40868 45076 40920 45082
rect 40868 45018 40920 45024
rect 38752 44940 38804 44946
rect 38752 44882 38804 44888
rect 38568 44396 38620 44402
rect 38568 44338 38620 44344
rect 38476 44260 38528 44266
rect 38476 44202 38528 44208
rect 35900 43988 35952 43994
rect 35900 43930 35952 43936
rect 36636 43988 36688 43994
rect 36636 43930 36688 43936
rect 35492 43676 35572 43704
rect 35808 43716 35860 43722
rect 35440 43658 35492 43664
rect 35808 43658 35860 43664
rect 35452 43450 35480 43658
rect 35440 43444 35492 43450
rect 35440 43386 35492 43392
rect 34520 43308 34572 43314
rect 34520 43250 34572 43256
rect 33324 43240 33376 43246
rect 33324 43182 33376 43188
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 33140 42900 33192 42906
rect 33140 42842 33192 42848
rect 32220 42764 32272 42770
rect 32220 42706 32272 42712
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 30116 26206 30236 26234
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25044 7404 25096 7410
rect 25044 7346 25096 7352
rect 23112 7200 23164 7206
rect 23112 7142 23164 7148
rect 23756 7200 23808 7206
rect 23756 7142 23808 7148
rect 24584 7200 24636 7206
rect 24584 7142 24636 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 2608 800 2636 2382
rect 3160 800 3188 2382
rect 3528 800 3556 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 3896 800 3924 2382
rect 4632 1850 4660 3470
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4264 1822 4660 1850
rect 4264 800 4292 1822
rect 4724 1442 4752 2926
rect 4632 1414 4752 1442
rect 4632 800 4660 1414
rect 4908 800 4936 3470
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5184 800 5212 2790
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5460 800 5488 2450
rect 5736 800 5764 3470
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 6012 800 6040 2926
rect 6276 2848 6328 2854
rect 6276 2790 6328 2796
rect 6288 800 6316 2790
rect 6564 800 6592 3470
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 6840 800 6868 2518
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7116 800 7144 2382
rect 7392 800 7420 3470
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 7668 800 7696 2790
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 7944 800 7972 2518
rect 8220 800 8248 3470
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8496 800 8524 2790
rect 8772 800 8800 2790
rect 9048 800 9076 3470
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9312 2372 9364 2378
rect 9312 2314 9364 2320
rect 9324 800 9352 2314
rect 9600 800 9628 2790
rect 9876 800 9904 3470
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10152 800 10180 2450
rect 10428 800 10456 2790
rect 10704 800 10732 3470
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 10980 800 11008 2790
rect 11244 2576 11296 2582
rect 11244 2518 11296 2524
rect 11256 800 11284 2518
rect 11532 800 11560 3470
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11808 800 11836 2790
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 12084 800 12112 2382
rect 12268 800 12296 3878
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12544 800 12572 2450
rect 12820 800 12848 3470
rect 13096 800 13124 3878
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13360 2916 13412 2922
rect 13360 2858 13412 2864
rect 13372 800 13400 2858
rect 13648 800 13676 3470
rect 13924 800 13952 3878
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14200 800 14228 3470
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14476 800 14504 2994
rect 14740 2576 14792 2582
rect 14740 2518 14792 2524
rect 14752 800 14780 2518
rect 15028 800 15056 4558
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15304 800 15332 3878
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15488 1306 15516 2450
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15580 2038 15608 2382
rect 15568 2032 15620 2038
rect 15568 1974 15620 1980
rect 15488 1278 15608 1306
rect 15580 800 15608 1278
rect 15856 800 15884 4558
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16396 3664 16448 3670
rect 16396 3606 16448 3612
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16132 3058 16160 3470
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 16132 800 16160 2790
rect 16408 800 16436 3606
rect 16776 3534 16804 4082
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 16684 800 16712 2926
rect 16776 2514 16804 3334
rect 16764 2508 16816 2514
rect 16764 2450 16816 2456
rect 16960 800 16988 4966
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17144 2922 17172 3606
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 17236 800 17264 4014
rect 17420 2394 17448 4558
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17512 3126 17540 3878
rect 17500 3120 17552 3126
rect 17500 3062 17552 3068
rect 17420 2366 17540 2394
rect 17512 800 17540 2366
rect 17696 1986 17724 3946
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17788 3126 17816 3878
rect 17972 3738 18000 5102
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17776 3120 17828 3126
rect 17776 3062 17828 3068
rect 17972 2854 18000 3470
rect 18064 2990 18092 4558
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 17880 2514 17908 2790
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 17868 2508 17920 2514
rect 17868 2450 17920 2456
rect 17696 1958 17816 1986
rect 17788 800 17816 1958
rect 18064 800 18092 2586
rect 18340 800 18368 4966
rect 18616 800 18644 5646
rect 18984 5574 19012 6054
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 18984 5234 19012 5510
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 18800 2106 18828 2246
rect 18788 2100 18840 2106
rect 18788 2042 18840 2048
rect 18892 800 18920 2790
rect 19076 1970 19104 4626
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19064 1964 19116 1970
rect 19064 1906 19116 1912
rect 19168 800 19196 3130
rect 19260 2446 19288 3538
rect 19352 3074 19380 6054
rect 20168 5772 20220 5778
rect 20168 5714 20220 5720
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19984 5092 20036 5098
rect 19984 5034 20036 5040
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19444 4146 19472 4558
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19352 3046 19472 3074
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 19444 2122 19472 3046
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19260 2094 19472 2122
rect 19260 1714 19288 2094
rect 19708 1964 19760 1970
rect 19708 1906 19760 1912
rect 19260 1686 19472 1714
rect 19444 800 19472 1686
rect 19720 800 19748 1906
rect 19996 800 20024 5034
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 20088 4690 20116 4966
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 20180 4010 20208 5714
rect 20272 4758 20300 6054
rect 20812 5704 20864 5710
rect 20812 5646 20864 5652
rect 20260 4752 20312 4758
rect 20260 4694 20312 4700
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20272 3126 20300 3674
rect 20536 3664 20588 3670
rect 20536 3606 20588 3612
rect 20260 3120 20312 3126
rect 20260 3062 20312 3068
rect 20260 2032 20312 2038
rect 20260 1974 20312 1980
rect 20272 800 20300 1974
rect 20548 800 20576 3606
rect 20824 3602 20852 5646
rect 21192 5302 21220 6734
rect 21284 6322 21312 6734
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21284 5846 21312 6258
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22100 6180 22152 6186
rect 22100 6122 22152 6128
rect 21272 5840 21324 5846
rect 21272 5782 21324 5788
rect 21732 5568 21784 5574
rect 21732 5510 21784 5516
rect 21180 5296 21232 5302
rect 21180 5238 21232 5244
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 21088 4684 21140 4690
rect 21088 4626 21140 4632
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20640 2378 20668 3334
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 20812 2100 20864 2106
rect 20812 2042 20864 2048
rect 20824 800 20852 2042
rect 21100 800 21128 4626
rect 21376 800 21404 5102
rect 21744 3602 21772 5510
rect 22112 5234 22140 6122
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22204 5778 22232 6054
rect 22192 5772 22244 5778
rect 22192 5714 22244 5720
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22296 4758 22324 6190
rect 22388 5778 22416 6598
rect 22376 5772 22428 5778
rect 22376 5714 22428 5720
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22284 4752 22336 4758
rect 22284 4694 22336 4700
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 21732 3596 21784 3602
rect 21732 3538 21784 3544
rect 21640 2848 21692 2854
rect 21640 2790 21692 2796
rect 21652 800 21680 2790
rect 22112 2446 22140 3878
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 21928 800 21956 2246
rect 22204 800 22232 3538
rect 22296 2122 22324 4014
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 22480 3058 22508 3402
rect 22468 3052 22520 3058
rect 22468 2994 22520 3000
rect 22940 2836 22968 5714
rect 23032 5302 23060 6598
rect 23020 5296 23072 5302
rect 23020 5238 23072 5244
rect 23124 4826 23152 7142
rect 23480 5160 23532 5166
rect 23480 5102 23532 5108
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 22940 2808 23060 2836
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 22296 2094 22508 2122
rect 22480 800 22508 2094
rect 22756 800 22784 2450
rect 23032 800 23060 2808
rect 23492 2802 23520 5102
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 23308 2774 23520 2802
rect 23308 800 23336 2774
rect 23584 800 23612 4626
rect 23768 3194 23796 7142
rect 24492 6656 24544 6662
rect 24492 6598 24544 6604
rect 24504 6390 24532 6598
rect 24492 6384 24544 6390
rect 24492 6326 24544 6332
rect 24596 5302 24624 7142
rect 25056 6866 25084 7346
rect 25044 6860 25096 6866
rect 25044 6802 25096 6808
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24872 5710 24900 6598
rect 24952 6248 25004 6254
rect 24952 6190 25004 6196
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 24584 5296 24636 5302
rect 24584 5238 24636 5244
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 24044 4146 24072 5102
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24032 4140 24084 4146
rect 24032 4082 24084 4088
rect 24308 4072 24360 4078
rect 24308 4014 24360 4020
rect 24676 4072 24728 4078
rect 24676 4014 24728 4020
rect 24320 3738 24348 4014
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 23848 3392 23900 3398
rect 23848 3334 23900 3340
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23860 3126 23888 3334
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 24400 2984 24452 2990
rect 24400 2926 24452 2932
rect 23860 800 23888 2926
rect 24124 2372 24176 2378
rect 24124 2314 24176 2320
rect 24136 800 24164 2314
rect 24412 800 24440 2926
rect 24688 800 24716 4014
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 24780 3058 24808 3878
rect 24872 3534 24900 4558
rect 24860 3528 24912 3534
rect 24860 3470 24912 3476
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 24964 800 24992 6190
rect 25056 5846 25084 6802
rect 25148 6798 25176 7482
rect 25596 7200 25648 7206
rect 25596 7142 25648 7148
rect 26424 7200 26476 7206
rect 26424 7142 26476 7148
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 25044 5840 25096 5846
rect 25044 5782 25096 5788
rect 25056 4690 25084 5782
rect 25136 5636 25188 5642
rect 25136 5578 25188 5584
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 25148 3670 25176 5578
rect 25228 5160 25280 5166
rect 25228 5102 25280 5108
rect 25136 3664 25188 3670
rect 25136 3606 25188 3612
rect 25240 800 25268 5102
rect 25608 4690 25636 7142
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26252 5778 26280 6734
rect 26240 5772 26292 5778
rect 26240 5714 26292 5720
rect 25596 4684 25648 4690
rect 25596 4626 25648 4632
rect 26332 4684 26384 4690
rect 26332 4626 26384 4632
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 25516 3602 25544 3878
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 26056 3596 26108 3602
rect 26056 3538 26108 3544
rect 25504 2984 25556 2990
rect 25504 2926 25556 2932
rect 25516 800 25544 2926
rect 25780 2508 25832 2514
rect 25780 2450 25832 2456
rect 25792 800 25820 2450
rect 26068 800 26096 3538
rect 26344 800 26372 4626
rect 26436 2514 26464 7142
rect 30116 6914 30144 26206
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 29840 6886 30144 6914
rect 26700 6792 26752 6798
rect 26700 6734 26752 6740
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 27804 6792 27856 6798
rect 27804 6734 27856 6740
rect 26608 5636 26660 5642
rect 26608 5578 26660 5584
rect 26424 2508 26476 2514
rect 26424 2450 26476 2456
rect 26620 800 26648 5578
rect 26712 2514 26740 6734
rect 27540 6322 27568 6734
rect 27712 6656 27764 6662
rect 27712 6598 27764 6604
rect 27724 6390 27752 6598
rect 27712 6384 27764 6390
rect 27712 6326 27764 6332
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 27816 5574 27844 6734
rect 29184 6248 29236 6254
rect 29184 6190 29236 6196
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 27804 5568 27856 5574
rect 27804 5510 27856 5516
rect 27712 5092 27764 5098
rect 27712 5034 27764 5040
rect 27436 4072 27488 4078
rect 27436 4014 27488 4020
rect 26884 2984 26936 2990
rect 26884 2926 26936 2932
rect 26700 2508 26752 2514
rect 26700 2450 26752 2456
rect 26896 800 26924 2926
rect 27160 2372 27212 2378
rect 27160 2314 27212 2320
rect 27172 800 27200 2314
rect 27448 800 27476 4014
rect 27724 800 27752 5034
rect 27816 4622 27844 5510
rect 29012 5234 29040 5646
rect 29000 5228 29052 5234
rect 29000 5170 29052 5176
rect 27988 5160 28040 5166
rect 27988 5102 28040 5108
rect 28000 4826 28028 5102
rect 27988 4820 28040 4826
rect 27988 4762 28040 4768
rect 27804 4616 27856 4622
rect 27804 4558 27856 4564
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 27816 3534 27844 4558
rect 29012 4146 29040 4558
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 27896 4072 27948 4078
rect 27896 4014 27948 4020
rect 29092 4072 29144 4078
rect 29092 4014 29144 4020
rect 27908 3738 27936 4014
rect 27896 3732 27948 3738
rect 27896 3674 27948 3680
rect 27804 3528 27856 3534
rect 27804 3470 27856 3476
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 28264 3460 28316 3466
rect 28264 3402 28316 3408
rect 27988 3188 28040 3194
rect 27988 3130 28040 3136
rect 28000 800 28028 3130
rect 28276 800 28304 3402
rect 28816 3392 28868 3398
rect 28816 3334 28868 3340
rect 28828 3126 28856 3334
rect 28816 3120 28868 3126
rect 28816 3062 28868 3068
rect 29012 3058 29040 3470
rect 29000 3052 29052 3058
rect 29000 2994 29052 3000
rect 28540 2984 28592 2990
rect 28540 2926 28592 2932
rect 28552 800 28580 2926
rect 28816 2848 28868 2854
rect 28816 2790 28868 2796
rect 28828 800 28856 2790
rect 29104 800 29132 4014
rect 29196 3194 29224 6190
rect 29644 5568 29696 5574
rect 29644 5510 29696 5516
rect 29656 5302 29684 5510
rect 29644 5296 29696 5302
rect 29644 5238 29696 5244
rect 29736 5160 29788 5166
rect 29736 5102 29788 5108
rect 29748 4826 29776 5102
rect 29736 4820 29788 4826
rect 29736 4762 29788 4768
rect 29840 3516 29868 6886
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 30012 5160 30064 5166
rect 30012 5102 30064 5108
rect 29656 3488 29868 3516
rect 29184 3188 29236 3194
rect 29184 3130 29236 3136
rect 29368 2372 29420 2378
rect 29368 2314 29420 2320
rect 29380 800 29408 2314
rect 29656 800 29684 3488
rect 29920 3188 29972 3194
rect 29920 3130 29972 3136
rect 29932 800 29960 3130
rect 30024 2854 30052 5102
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 31300 4684 31352 4690
rect 31300 4626 31352 4632
rect 31208 4616 31260 4622
rect 31208 4558 31260 4564
rect 30748 3732 30800 3738
rect 30748 3674 30800 3680
rect 30196 3664 30248 3670
rect 30196 3606 30248 3612
rect 30012 2848 30064 2854
rect 30012 2790 30064 2796
rect 30208 800 30236 3606
rect 30472 3392 30524 3398
rect 30472 3334 30524 3340
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30392 2514 30420 2790
rect 30380 2508 30432 2514
rect 30380 2450 30432 2456
rect 30484 800 30512 3334
rect 30760 800 30788 3674
rect 31220 3602 31248 4558
rect 31312 4146 31340 4626
rect 32128 4616 32180 4622
rect 32128 4558 32180 4564
rect 32312 4616 32364 4622
rect 32312 4558 32364 4564
rect 31760 4480 31812 4486
rect 31760 4422 31812 4428
rect 31300 4140 31352 4146
rect 31300 4082 31352 4088
rect 31576 4140 31628 4146
rect 31576 4082 31628 4088
rect 31392 4072 31444 4078
rect 31392 4014 31444 4020
rect 31208 3596 31260 3602
rect 31208 3538 31260 3544
rect 31024 2916 31076 2922
rect 31024 2858 31076 2864
rect 31036 800 31064 2858
rect 31404 1986 31432 4014
rect 31312 1958 31432 1986
rect 31312 800 31340 1958
rect 31588 800 31616 4082
rect 31772 4010 31800 4422
rect 32140 4214 32168 4558
rect 32128 4208 32180 4214
rect 32128 4150 32180 4156
rect 31760 4004 31812 4010
rect 31760 3946 31812 3952
rect 31852 3936 31904 3942
rect 31852 3878 31904 3884
rect 31760 3664 31812 3670
rect 31760 3606 31812 3612
rect 31772 3398 31800 3606
rect 31760 3392 31812 3398
rect 31760 3334 31812 3340
rect 31864 2378 31892 3878
rect 32140 3534 32168 4150
rect 32324 4146 32352 4558
rect 32312 4140 32364 4146
rect 32312 4082 32364 4088
rect 34060 4004 34112 4010
rect 34060 3946 34112 3952
rect 32772 3936 32824 3942
rect 32772 3878 32824 3884
rect 33784 3936 33836 3942
rect 33784 3878 33836 3884
rect 32128 3528 32180 3534
rect 32128 3470 32180 3476
rect 32680 3528 32732 3534
rect 32680 3470 32732 3476
rect 31944 3392 31996 3398
rect 31944 3334 31996 3340
rect 31956 2582 31984 3334
rect 31944 2576 31996 2582
rect 31944 2518 31996 2524
rect 32140 2446 32168 3470
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 32220 3392 32272 3398
rect 32220 3334 32272 3340
rect 32128 2440 32180 2446
rect 32128 2382 32180 2388
rect 31852 2372 31904 2378
rect 31852 2314 31904 2320
rect 31944 2372 31996 2378
rect 31944 2314 31996 2320
rect 31956 1306 31984 2314
rect 32232 1850 32260 3334
rect 32416 2650 32444 3402
rect 32496 2848 32548 2854
rect 32496 2790 32548 2796
rect 32404 2644 32456 2650
rect 32404 2586 32456 2592
rect 31864 1278 31984 1306
rect 32140 1822 32260 1850
rect 31864 800 31892 1278
rect 32140 800 32168 1822
rect 32508 1442 32536 2790
rect 32692 2514 32720 3470
rect 32680 2508 32732 2514
rect 32680 2450 32732 2456
rect 32784 1986 32812 3878
rect 33232 3664 33284 3670
rect 33232 3606 33284 3612
rect 33048 3120 33100 3126
rect 33048 3062 33100 3068
rect 32864 3052 32916 3058
rect 32864 2994 32916 3000
rect 32876 2774 32904 2994
rect 32876 2746 32996 2774
rect 32416 1414 32536 1442
rect 32692 1958 32812 1986
rect 32416 800 32444 1414
rect 32692 800 32720 1958
rect 32968 800 32996 2746
rect 33060 2650 33088 3062
rect 33048 2644 33100 2650
rect 33048 2586 33100 2592
rect 33244 800 33272 3606
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 33508 3120 33560 3126
rect 33508 3062 33560 3068
rect 33520 800 33548 3062
rect 33612 3058 33640 3402
rect 33692 3188 33744 3194
rect 33692 3130 33744 3136
rect 33600 3052 33652 3058
rect 33600 2994 33652 3000
rect 33704 2774 33732 3130
rect 33612 2746 33732 2774
rect 33612 2650 33640 2746
rect 33600 2644 33652 2650
rect 33600 2586 33652 2592
rect 33796 800 33824 3878
rect 34072 800 34100 3946
rect 35348 3936 35400 3942
rect 35348 3878 35400 3884
rect 47308 3936 47360 3942
rect 47308 3878 47360 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34520 3596 34572 3602
rect 34520 3538 34572 3544
rect 34612 3596 34664 3602
rect 34612 3538 34664 3544
rect 34336 2916 34388 2922
rect 34336 2858 34388 2864
rect 34348 800 34376 2858
rect 34532 2650 34560 3538
rect 34520 2644 34572 2650
rect 34520 2586 34572 2592
rect 34624 800 34652 3538
rect 34796 2984 34848 2990
rect 34796 2926 34848 2932
rect 34808 1578 34836 2926
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 1986 35388 3878
rect 35440 3664 35492 3670
rect 35440 3606 35492 3612
rect 37464 3664 37516 3670
rect 37464 3606 37516 3612
rect 40684 3664 40736 3670
rect 40684 3606 40736 3612
rect 46480 3664 46532 3670
rect 46480 3606 46532 3612
rect 35176 1958 35388 1986
rect 34808 1550 34928 1578
rect 34900 800 34928 1550
rect 35176 800 35204 1958
rect 35452 800 35480 3606
rect 35992 3596 36044 3602
rect 35992 3538 36044 3544
rect 35716 3052 35768 3058
rect 35716 2994 35768 3000
rect 35728 800 35756 2994
rect 36004 800 36032 3538
rect 36544 3528 36596 3534
rect 36544 3470 36596 3476
rect 36176 3120 36228 3126
rect 36176 3062 36228 3068
rect 36188 2650 36216 3062
rect 36176 2644 36228 2650
rect 36176 2586 36228 2592
rect 36268 2440 36320 2446
rect 36268 2382 36320 2388
rect 36280 800 36308 2382
rect 36556 800 36584 3470
rect 37372 2984 37424 2990
rect 37372 2926 37424 2932
rect 36820 2916 36872 2922
rect 36820 2858 36872 2864
rect 36832 800 36860 2858
rect 37384 2650 37412 2926
rect 37372 2644 37424 2650
rect 37372 2586 37424 2592
rect 37096 2508 37148 2514
rect 37096 2450 37148 2456
rect 37108 800 37136 2450
rect 37476 1850 37504 3606
rect 37924 3528 37976 3534
rect 37924 3470 37976 3476
rect 39304 3528 39356 3534
rect 39304 3470 39356 3476
rect 40132 3528 40184 3534
rect 40132 3470 40184 3476
rect 37648 2984 37700 2990
rect 37648 2926 37700 2932
rect 37384 1822 37504 1850
rect 37384 800 37412 1822
rect 37660 800 37688 2926
rect 37936 800 37964 3470
rect 38476 2916 38528 2922
rect 38476 2858 38528 2864
rect 38200 2576 38252 2582
rect 38200 2518 38252 2524
rect 38212 800 38240 2518
rect 38488 800 38516 2858
rect 38752 2848 38804 2854
rect 38752 2790 38804 2796
rect 38764 800 38792 2790
rect 39028 2508 39080 2514
rect 39028 2450 39080 2456
rect 39040 800 39068 2450
rect 39316 800 39344 3470
rect 39856 2984 39908 2990
rect 39856 2926 39908 2932
rect 39580 2440 39632 2446
rect 39580 2382 39632 2388
rect 39592 800 39620 2382
rect 39868 800 39896 2926
rect 40144 800 40172 3470
rect 40408 2916 40460 2922
rect 40408 2858 40460 2864
rect 40420 800 40448 2858
rect 40696 800 40724 3606
rect 41236 3596 41288 3602
rect 41236 3538 41288 3544
rect 40960 2508 41012 2514
rect 40960 2450 41012 2456
rect 40972 800 41000 2450
rect 41248 800 41276 3538
rect 42616 3528 42668 3534
rect 42616 3470 42668 3476
rect 42892 3528 42944 3534
rect 42892 3470 42944 3476
rect 44548 3528 44600 3534
rect 44548 3470 44600 3476
rect 45376 3528 45428 3534
rect 45376 3470 45428 3476
rect 46204 3528 46256 3534
rect 46204 3470 46256 3476
rect 42340 2984 42392 2990
rect 42340 2926 42392 2932
rect 41788 2848 41840 2854
rect 41788 2790 41840 2796
rect 41512 2440 41564 2446
rect 41512 2382 41564 2388
rect 41524 800 41552 2382
rect 41800 800 41828 2790
rect 42064 2576 42116 2582
rect 42064 2518 42116 2524
rect 42076 800 42104 2518
rect 42352 800 42380 2926
rect 42628 800 42656 3470
rect 42904 800 42932 3470
rect 44272 2984 44324 2990
rect 44272 2926 44324 2932
rect 43168 2916 43220 2922
rect 43168 2858 43220 2864
rect 43180 800 43208 2858
rect 43720 2848 43772 2854
rect 43720 2790 43772 2796
rect 43444 2508 43496 2514
rect 43444 2450 43496 2456
rect 43456 800 43484 2450
rect 43732 800 43760 2790
rect 43996 2372 44048 2378
rect 43996 2314 44048 2320
rect 44008 800 44036 2314
rect 44284 800 44312 2926
rect 44560 800 44588 3470
rect 45100 2916 45152 2922
rect 45100 2858 45152 2864
rect 44824 2576 44876 2582
rect 44824 2518 44876 2524
rect 44836 800 44864 2518
rect 45112 800 45140 2858
rect 45388 800 45416 3470
rect 45652 2848 45704 2854
rect 45652 2790 45704 2796
rect 45664 800 45692 2790
rect 45928 2440 45980 2446
rect 45928 2382 45980 2388
rect 45940 800 45968 2382
rect 46216 800 46244 3470
rect 46492 800 46520 3606
rect 47032 3596 47084 3602
rect 47032 3538 47084 3544
rect 46756 2848 46808 2854
rect 46756 2790 46808 2796
rect 46768 800 46796 2790
rect 47044 800 47072 3538
rect 47320 800 47348 3878
rect 2410 0 2466 800
rect 2502 0 2558 800
rect 2594 0 2650 800
rect 2686 0 2742 800
rect 2778 0 2834 800
rect 2870 0 2926 800
rect 2962 0 3018 800
rect 3054 0 3110 800
rect 3146 0 3202 800
rect 3238 0 3294 800
rect 3330 0 3386 800
rect 3422 0 3478 800
rect 3514 0 3570 800
rect 3606 0 3662 800
rect 3698 0 3754 800
rect 3790 0 3846 800
rect 3882 0 3938 800
rect 3974 0 4030 800
rect 4066 0 4122 800
rect 4158 0 4214 800
rect 4250 0 4306 800
rect 4342 0 4398 800
rect 4434 0 4490 800
rect 4526 0 4582 800
rect 4618 0 4674 800
rect 4710 0 4766 800
rect 4802 0 4858 800
rect 4894 0 4950 800
rect 4986 0 5042 800
rect 5078 0 5134 800
rect 5170 0 5226 800
rect 5262 0 5318 800
rect 5354 0 5410 800
rect 5446 0 5502 800
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5722 0 5778 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6366 0 6422 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6642 0 6698 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7010 0 7066 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
<< via2 >>
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19430 46008 19486 46064
rect 19798 46008 19854 46064
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 20810 45500 20812 45520
rect 20812 45500 20864 45520
rect 20864 45500 20866 45520
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 20810 45464 20866 45500
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 21638 44940 21694 44976
rect 21638 44920 21640 44940
rect 21640 44920 21692 44940
rect 21692 44920 21694 44940
rect 22006 45328 22062 45384
rect 22374 45600 22430 45656
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 23478 45192 23534 45248
rect 24306 46452 24308 46472
rect 24308 46452 24360 46472
rect 24360 46452 24362 46472
rect 24306 46416 24362 46452
rect 24858 46588 24860 46608
rect 24860 46588 24912 46608
rect 24912 46588 24914 46608
rect 24858 46552 24914 46588
rect 26422 46552 26478 46608
rect 26054 45908 26056 45928
rect 26056 45908 26108 45928
rect 26108 45908 26110 45928
rect 26054 45872 26110 45908
rect 26790 45908 26792 45928
rect 26792 45908 26844 45928
rect 26844 45908 26846 45928
rect 26238 45620 26294 45656
rect 26238 45600 26240 45620
rect 26240 45600 26292 45620
rect 26292 45600 26294 45620
rect 26238 45192 26294 45248
rect 26422 44920 26478 44976
rect 26790 45872 26846 45908
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 27342 46552 27398 46608
rect 27526 45600 27582 45656
rect 27802 46416 27858 46472
rect 27986 45892 28042 45928
rect 27986 45872 27988 45892
rect 27988 45872 28040 45892
rect 28040 45872 28042 45892
rect 27710 42356 27766 42392
rect 27710 42336 27712 42356
rect 27712 42336 27764 42356
rect 27764 42336 27766 42356
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 29826 45872 29882 45928
rect 30654 46572 30710 46608
rect 30654 46552 30656 46572
rect 30656 46552 30708 46572
rect 30708 46552 30710 46572
rect 31850 46452 31852 46472
rect 31852 46452 31904 46472
rect 31904 46452 31906 46472
rect 31850 46416 31906 46452
rect 32954 46044 32956 46064
rect 32956 46044 33008 46064
rect 33008 46044 33010 46064
rect 32954 46008 33010 46044
rect 33506 46552 33562 46608
rect 33690 46552 33746 46608
rect 33414 45500 33416 45520
rect 33416 45500 33468 45520
rect 33468 45500 33470 45520
rect 33414 45464 33470 45500
rect 33782 45736 33838 45792
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34978 45872 35034 45928
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 35806 45600 35862 45656
rect 36174 45600 36230 45656
rect 36450 45736 36506 45792
rect 37830 47232 37886 47288
rect 38014 47096 38070 47152
rect 37278 46824 37334 46880
rect 37646 46416 37702 46472
rect 37554 45600 37610 45656
rect 37462 45364 37464 45384
rect 37464 45364 37516 45384
rect 37516 45364 37518 45384
rect 37462 45328 37518 45364
rect 38474 46960 38530 47016
rect 38842 46996 38844 47016
rect 38844 46996 38896 47016
rect 38896 46996 38898 47016
rect 38842 46960 38898 46996
rect 39118 46572 39174 46608
rect 39118 46552 39120 46572
rect 39120 46552 39172 46572
rect 39172 46552 39174 46572
rect 40222 47096 40278 47152
rect 41970 46824 42026 46880
rect 44270 47252 44326 47288
rect 44270 47232 44272 47252
rect 44272 47232 44324 47252
rect 44324 47232 44326 47252
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
<< metal3 >>
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 37825 47290 37891 47293
rect 44265 47290 44331 47293
rect 37825 47288 44331 47290
rect 37825 47232 37830 47288
rect 37886 47232 44270 47288
rect 44326 47232 44331 47288
rect 37825 47230 44331 47232
rect 37825 47227 37891 47230
rect 44265 47227 44331 47230
rect 38009 47154 38075 47157
rect 40217 47154 40283 47157
rect 38009 47152 40283 47154
rect 38009 47096 38014 47152
rect 38070 47096 40222 47152
rect 40278 47096 40283 47152
rect 38009 47094 40283 47096
rect 38009 47091 38075 47094
rect 40217 47091 40283 47094
rect 38469 47018 38535 47021
rect 38837 47018 38903 47021
rect 38469 47016 38903 47018
rect 38469 46960 38474 47016
rect 38530 46960 38842 47016
rect 38898 46960 38903 47016
rect 38469 46958 38903 46960
rect 38469 46955 38535 46958
rect 38837 46955 38903 46958
rect 37273 46882 37339 46885
rect 41965 46882 42031 46885
rect 37273 46880 42031 46882
rect 37273 46824 37278 46880
rect 37334 46824 41970 46880
rect 42026 46824 42031 46880
rect 37273 46822 42031 46824
rect 37273 46819 37339 46822
rect 41965 46819 42031 46822
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 24853 46610 24919 46613
rect 26417 46610 26483 46613
rect 27337 46610 27403 46613
rect 24853 46608 27403 46610
rect 24853 46552 24858 46608
rect 24914 46552 26422 46608
rect 26478 46552 27342 46608
rect 27398 46552 27403 46608
rect 24853 46550 27403 46552
rect 24853 46547 24919 46550
rect 26417 46547 26483 46550
rect 27337 46547 27403 46550
rect 30649 46610 30715 46613
rect 33501 46610 33567 46613
rect 30649 46608 33567 46610
rect 30649 46552 30654 46608
rect 30710 46552 33506 46608
rect 33562 46552 33567 46608
rect 30649 46550 33567 46552
rect 30649 46547 30715 46550
rect 33501 46547 33567 46550
rect 33685 46610 33751 46613
rect 39113 46610 39179 46613
rect 33685 46608 39179 46610
rect 33685 46552 33690 46608
rect 33746 46552 39118 46608
rect 39174 46552 39179 46608
rect 33685 46550 39179 46552
rect 33685 46547 33751 46550
rect 39113 46547 39179 46550
rect 24301 46474 24367 46477
rect 27797 46474 27863 46477
rect 24301 46472 27863 46474
rect 24301 46416 24306 46472
rect 24362 46416 27802 46472
rect 27858 46416 27863 46472
rect 24301 46414 27863 46416
rect 24301 46411 24367 46414
rect 27797 46411 27863 46414
rect 31845 46474 31911 46477
rect 37641 46474 37707 46477
rect 31845 46472 37707 46474
rect 31845 46416 31850 46472
rect 31906 46416 37646 46472
rect 37702 46416 37707 46472
rect 31845 46414 37707 46416
rect 31845 46411 31911 46414
rect 37641 46411 37707 46414
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 19425 46066 19491 46069
rect 19793 46066 19859 46069
rect 32949 46066 33015 46069
rect 19425 46064 33015 46066
rect 19425 46008 19430 46064
rect 19486 46008 19798 46064
rect 19854 46008 32954 46064
rect 33010 46008 33015 46064
rect 19425 46006 33015 46008
rect 19425 46003 19491 46006
rect 19793 46003 19859 46006
rect 32949 46003 33015 46006
rect 26049 45930 26115 45933
rect 26785 45930 26851 45933
rect 27981 45930 28047 45933
rect 26049 45928 28047 45930
rect 26049 45872 26054 45928
rect 26110 45872 26790 45928
rect 26846 45872 27986 45928
rect 28042 45872 28047 45928
rect 26049 45870 28047 45872
rect 26049 45867 26115 45870
rect 26785 45867 26851 45870
rect 27981 45867 28047 45870
rect 29821 45930 29887 45933
rect 34973 45930 35039 45933
rect 29821 45928 35039 45930
rect 29821 45872 29826 45928
rect 29882 45872 34978 45928
rect 35034 45872 35039 45928
rect 29821 45870 35039 45872
rect 29821 45867 29887 45870
rect 34973 45867 35039 45870
rect 33777 45794 33843 45797
rect 36445 45794 36511 45797
rect 33777 45792 36511 45794
rect 33777 45736 33782 45792
rect 33838 45736 36450 45792
rect 36506 45736 36511 45792
rect 33777 45734 36511 45736
rect 33777 45731 33843 45734
rect 36445 45731 36511 45734
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 22369 45658 22435 45661
rect 26233 45658 26299 45661
rect 22369 45656 26299 45658
rect 22369 45600 22374 45656
rect 22430 45600 26238 45656
rect 26294 45600 26299 45656
rect 22369 45598 26299 45600
rect 22369 45595 22435 45598
rect 26233 45595 26299 45598
rect 27521 45658 27587 45661
rect 27654 45658 27660 45660
rect 27521 45656 27660 45658
rect 27521 45600 27526 45656
rect 27582 45600 27660 45656
rect 27521 45598 27660 45600
rect 27521 45595 27587 45598
rect 27654 45596 27660 45598
rect 27724 45596 27730 45660
rect 35801 45658 35867 45661
rect 36169 45658 36235 45661
rect 37549 45658 37615 45661
rect 35801 45656 37615 45658
rect 35801 45600 35806 45656
rect 35862 45600 36174 45656
rect 36230 45600 37554 45656
rect 37610 45600 37615 45656
rect 35801 45598 37615 45600
rect 35801 45595 35867 45598
rect 36169 45595 36235 45598
rect 37549 45595 37615 45598
rect 20805 45522 20871 45525
rect 33409 45522 33475 45525
rect 20805 45520 33475 45522
rect 20805 45464 20810 45520
rect 20866 45464 33414 45520
rect 33470 45464 33475 45520
rect 20805 45462 33475 45464
rect 20805 45459 20871 45462
rect 33409 45459 33475 45462
rect 22001 45386 22067 45389
rect 37457 45386 37523 45389
rect 22001 45384 37523 45386
rect 22001 45328 22006 45384
rect 22062 45328 37462 45384
rect 37518 45328 37523 45384
rect 22001 45326 37523 45328
rect 22001 45323 22067 45326
rect 37457 45323 37523 45326
rect 23473 45250 23539 45253
rect 26233 45250 26299 45253
rect 23473 45248 26299 45250
rect 23473 45192 23478 45248
rect 23534 45192 26238 45248
rect 26294 45192 26299 45248
rect 23473 45190 26299 45192
rect 23473 45187 23539 45190
rect 26233 45187 26299 45190
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 21633 44978 21699 44981
rect 26417 44978 26483 44981
rect 21633 44976 26483 44978
rect 21633 44920 21638 44976
rect 21694 44920 26422 44976
rect 26478 44920 26483 44976
rect 21633 44918 26483 44920
rect 21633 44915 21699 44918
rect 26417 44915 26483 44918
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 27705 42396 27771 42397
rect 27654 42332 27660 42396
rect 27724 42394 27771 42396
rect 27724 42392 27816 42394
rect 27766 42336 27816 42392
rect 27724 42334 27816 42336
rect 27724 42332 27771 42334
rect 27705 42331 27771 42332
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 27660 45596 27724 45660
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 27660 42392 27724 42396
rect 27660 42336 27710 42392
rect 27710 42336 27724 42392
rect 27660 42332 27724 42336
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 27659 45660 27725 45661
rect 27659 45596 27660 45660
rect 27724 45596 27725 45660
rect 27659 45595 27725 45596
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 27662 42397 27722 45595
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 27659 42396 27725 42397
rect 27659 42332 27660 42396
rect 27724 42332 27725 42396
rect 27659 42331 27725 42332
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 21344 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1666199351
transform 1 0 17756 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1666199351
transform -1 0 25300 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1666199351
transform 1 0 24564 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1666199351
transform 1 0 19412 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1666199351
transform 1 0 18952 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A_N
timestamp 1666199351
transform 1 0 30360 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B
timestamp 1666199351
transform 1 0 30636 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__B1
timestamp 1666199351
transform 1 0 23368 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B1
timestamp 1666199351
transform -1 0 20424 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1666199351
transform -1 0 28520 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__B2
timestamp 1666199351
transform -1 0 23000 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A2
timestamp 1666199351
transform -1 0 22356 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1666199351
transform -1 0 18952 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1666199351
transform 1 0 19780 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A2
timestamp 1666199351
transform 1 0 29716 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A2
timestamp 1666199351
transform 1 0 34868 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A1
timestamp 1666199351
transform 1 0 26680 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1666199351
transform 1 0 21804 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1666199351
transform 1 0 19688 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A1
timestamp 1666199351
transform -1 0 27876 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A
timestamp 1666199351
transform 1 0 25300 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__B1
timestamp 1666199351
transform 1 0 26220 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A1
timestamp 1666199351
transform 1 0 29716 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A
timestamp 1666199351
transform 1 0 20332 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1666199351
transform 1 0 20976 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1666199351
transform 1 0 23920 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A2
timestamp 1666199351
transform 1 0 26128 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A2
timestamp 1666199351
transform 1 0 29440 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A1
timestamp 1666199351
transform -1 0 24840 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__C1
timestamp 1666199351
transform 1 0 23644 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666199351
transform -1 0 4048 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666199351
transform -1 0 23000 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666199351
transform -1 0 22172 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666199351
transform -1 0 27324 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666199351
transform -1 0 27876 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666199351
transform -1 0 29072 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666199351
transform -1 0 33304 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666199351
transform -1 0 32292 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1666199351
transform -1 0 34684 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1666199351
transform -1 0 33580 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1666199351
transform -1 0 35696 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1666199351
transform -1 0 36984 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1666199351
transform -1 0 38548 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1666199351
transform -1 0 42136 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1666199351
transform -1 0 39468 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1666199351
transform -1 0 40204 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1666199351
transform -1 0 40848 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1666199351
transform -1 0 43424 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1666199351
transform -1 0 43976 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1666199351
transform -1 0 44528 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1666199351
transform -1 0 45356 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 1666199351
transform 1 0 9936 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19
timestamp 1666199351
transform 1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40
timestamp 1666199351
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47
timestamp 1666199351
transform 1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1666199351
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1666199351
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1666199351
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1666199351
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1666199351
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1666199351
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1666199351
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1666199351
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1666199351
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1666199351
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124
timestamp 1666199351
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 1666199351
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1666199351
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1666199351
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152
timestamp 1666199351
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_159
timestamp 1666199351
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1666199351
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1666199351
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1666199351
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1666199351
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1666199351
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1666199351
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1666199351
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1666199351
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1666199351
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1666199351
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1666199351
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1666199351
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1666199351
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666199351
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_342
timestamp 1666199351
transform 1 0 32568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1666199351
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1666199351
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1666199351
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_370
timestamp 1666199351
transform 1 0 35144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1666199351
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1666199351
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1666199351
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_398
timestamp 1666199351
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_405
timestamp 1666199351
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1666199351
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1666199351
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_426
timestamp 1666199351
transform 1 0 40296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_433
timestamp 1666199351
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_440
timestamp 1666199351
transform 1 0 41584 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1666199351
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_454
timestamp 1666199351
transform 1 0 42872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1666199351
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_468
timestamp 1666199351
transform 1 0 44160 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1666199351
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_482
timestamp 1666199351
transform 1 0 45448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1666199351
transform 1 0 46092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_496
timestamp 1666199351
transform 1 0 46736 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1666199351
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_510
timestamp 1666199351
transform 1 0 48024 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 1666199351
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1666199351
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_33
timestamp 1666199351
transform 1 0 4140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1666199351
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_47
timestamp 1666199351
transform 1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1666199351
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1666199351
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_68
timestamp 1666199351
transform 1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1666199351
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1666199351
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_89
timestamp 1666199351
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1666199351
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1666199351
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1666199351
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1666199351
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_124
timestamp 1666199351
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_131
timestamp 1666199351
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_138
timestamp 1666199351
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1666199351
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_152
timestamp 1666199351
transform 1 0 15088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_159
timestamp 1666199351
transform 1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1666199351
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_169
timestamp 1666199351
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_175 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 17204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_197
timestamp 1666199351
transform 1 0 19228 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1666199351
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_225
timestamp 1666199351
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_231
timestamp 1666199351
transform 1 0 22356 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_253
timestamp 1666199351
transform 1 0 24380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1666199351
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1666199351
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_304
timestamp 1666199351
transform 1 0 29072 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1666199351
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1666199351
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1666199351
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_342
timestamp 1666199351
transform 1 0 32568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_349
timestamp 1666199351
transform 1 0 33212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_356
timestamp 1666199351
transform 1 0 33856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_363
timestamp 1666199351
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_370
timestamp 1666199351
transform 1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_377
timestamp 1666199351
transform 1 0 35788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_384
timestamp 1666199351
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1666199351
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_398
timestamp 1666199351
transform 1 0 37720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_405
timestamp 1666199351
transform 1 0 38364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_412
timestamp 1666199351
transform 1 0 39008 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_419
timestamp 1666199351
transform 1 0 39652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_426
timestamp 1666199351
transform 1 0 40296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_433
timestamp 1666199351
transform 1 0 40940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_440
timestamp 1666199351
transform 1 0 41584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1666199351
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_454
timestamp 1666199351
transform 1 0 42872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1666199351
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_468
timestamp 1666199351
transform 1 0 44160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_475
timestamp 1666199351
transform 1 0 44804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_482
timestamp 1666199351
transform 1 0 45448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_489
timestamp 1666199351
transform 1 0 46092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_496
timestamp 1666199351
transform 1 0 46736 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1666199351
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_510
timestamp 1666199351
transform 1 0 48024 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666199351
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666199351
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666199351
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp 1666199351
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_38
timestamp 1666199351
transform 1 0 4600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_45
timestamp 1666199351
transform 1 0 5244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_54
timestamp 1666199351
transform 1 0 6072 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_63
timestamp 1666199351
transform 1 0 6900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_72
timestamp 1666199351
transform 1 0 7728 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1666199351
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_90
timestamp 1666199351
transform 1 0 9384 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_99
timestamp 1666199351
transform 1 0 10212 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_108
timestamp 1666199351
transform 1 0 11040 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1666199351
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_124
timestamp 1666199351
transform 1 0 12512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_131
timestamp 1666199351
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1666199351
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1666199351
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_152
timestamp 1666199351
transform 1 0 15088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1666199351
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1666199351
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1666199351
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1666199351
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_187
timestamp 1666199351
transform 1 0 18308 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1666199351
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1666199351
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_204
timestamp 1666199351
transform 1 0 19872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_211
timestamp 1666199351
transform 1 0 20516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_218
timestamp 1666199351
transform 1 0 21160 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_243
timestamp 1666199351
transform 1 0 23460 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1666199351
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1666199351
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_257
timestamp 1666199351
transform 1 0 24748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_261
timestamp 1666199351
transform 1 0 25116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_286
timestamp 1666199351
transform 1 0 27416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_293
timestamp 1666199351
transform 1 0 28060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp 1666199351
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1666199351
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_332
timestamp 1666199351
transform 1 0 31648 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_339
timestamp 1666199351
transform 1 0 32292 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_346
timestamp 1666199351
transform 1 0 32936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_353
timestamp 1666199351
transform 1 0 33580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1666199351
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1666199351
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_370
timestamp 1666199351
transform 1 0 35144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_377
timestamp 1666199351
transform 1 0 35788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_384
timestamp 1666199351
transform 1 0 36432 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_391
timestamp 1666199351
transform 1 0 37076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_398
timestamp 1666199351
transform 1 0 37720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_405
timestamp 1666199351
transform 1 0 38364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_412
timestamp 1666199351
transform 1 0 39008 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1666199351
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_426
timestamp 1666199351
transform 1 0 40296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_433
timestamp 1666199351
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_440
timestamp 1666199351
transform 1 0 41584 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_447
timestamp 1666199351
transform 1 0 42228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_451
timestamp 1666199351
transform 1 0 42596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_455
timestamp 1666199351
transform 1 0 42964 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_462
timestamp 1666199351
transform 1 0 43608 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1666199351
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1666199351
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_482
timestamp 1666199351
transform 1 0 45448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_489
timestamp 1666199351
transform 1 0 46092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_496
timestamp 1666199351
transform 1 0 46736 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_503
timestamp 1666199351
transform 1 0 47380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_510
timestamp 1666199351
transform 1 0 48024 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666199351
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666199351
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666199351
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666199351
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1666199351
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666199351
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666199351
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666199351
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666199351
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666199351
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666199351
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666199351
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1666199351
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1666199351
transform 1 0 12236 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_125
timestamp 1666199351
transform 1 0 12604 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_134
timestamp 1666199351
transform 1 0 13432 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_143
timestamp 1666199351
transform 1 0 14260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_152
timestamp 1666199351
transform 1 0 15088 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_159
timestamp 1666199351
transform 1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1666199351
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1666199351
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_176
timestamp 1666199351
transform 1 0 17296 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_183
timestamp 1666199351
transform 1 0 17940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_190
timestamp 1666199351
transform 1 0 18584 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_197
timestamp 1666199351
transform 1 0 19228 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1666199351
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1666199351
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_232
timestamp 1666199351
transform 1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_239
timestamp 1666199351
transform 1 0 23092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_246
timestamp 1666199351
transform 1 0 23736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_271
timestamp 1666199351
transform 1 0 26036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1666199351
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1666199351
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_304
timestamp 1666199351
transform 1 0 29072 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1666199351
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1666199351
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1666199351
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_342
timestamp 1666199351
transform 1 0 32568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_349
timestamp 1666199351
transform 1 0 33212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_356
timestamp 1666199351
transform 1 0 33856 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_363
timestamp 1666199351
transform 1 0 34500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_370
timestamp 1666199351
transform 1 0 35144 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_377
timestamp 1666199351
transform 1 0 35788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_389
timestamp 1666199351
transform 1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1666199351
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1666199351
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1666199351
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1666199351
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1666199351
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1666199351
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1666199351
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1666199351
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1666199351
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1666199351
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1666199351
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1666199351
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_505
timestamp 1666199351
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_510
timestamp 1666199351
transform 1 0 48024 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666199351
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666199351
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666199351
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666199351
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666199351
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666199351
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666199351
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666199351
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666199351
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666199351
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666199351
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666199351
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666199351
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666199351
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666199351
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_141
timestamp 1666199351
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_149
timestamp 1666199351
transform 1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_155
timestamp 1666199351
transform 1 0 15364 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_164
timestamp 1666199351
transform 1 0 16192 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_173
timestamp 1666199351
transform 1 0 17020 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_180
timestamp 1666199351
transform 1 0 17664 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_187
timestamp 1666199351
transform 1 0 18308 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1666199351
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_197
timestamp 1666199351
transform 1 0 19228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_203
timestamp 1666199351
transform 1 0 19780 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_225
timestamp 1666199351
transform 1 0 21804 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1666199351
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_253
timestamp 1666199351
transform 1 0 24380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_262
timestamp 1666199351
transform 1 0 25208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_287
timestamp 1666199351
transform 1 0 27508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_294
timestamp 1666199351
transform 1 0 28152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1666199351
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1666199351
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1666199351
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_314
timestamp 1666199351
transform 1 0 29992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp 1666199351
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_328
timestamp 1666199351
transform 1 0 31280 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_335
timestamp 1666199351
transform 1 0 31924 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_342
timestamp 1666199351
transform 1 0 32568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_354
timestamp 1666199351
transform 1 0 33672 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1666199351
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1666199351
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1666199351
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1666199351
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1666199351
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1666199351
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1666199351
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1666199351
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1666199351
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1666199351
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1666199351
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1666199351
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1666199351
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1666199351
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1666199351
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1666199351
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_513
timestamp 1666199351
transform 1 0 48300 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666199351
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666199351
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666199351
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1666199351
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666199351
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666199351
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666199351
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666199351
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666199351
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666199351
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666199351
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666199351
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666199351
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666199351
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666199351
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666199351
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666199351
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666199351
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1666199351
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_176
timestamp 1666199351
transform 1 0 17296 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_183
timestamp 1666199351
transform 1 0 17940 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_190
timestamp 1666199351
transform 1 0 18584 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1666199351
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1666199351
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1666199351
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_249
timestamp 1666199351
transform 1 0 24012 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1666199351
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1666199351
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_304
timestamp 1666199351
transform 1 0 29072 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1666199351
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1666199351
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1666199351
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1666199351
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1666199351
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1666199351
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1666199351
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1666199351
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1666199351
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1666199351
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1666199351
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1666199351
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1666199351
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1666199351
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1666199351
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1666199351
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1666199351
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1666199351
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1666199351
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1666199351
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_505
timestamp 1666199351
transform 1 0 47564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_513
timestamp 1666199351
transform 1 0 48300 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666199351
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666199351
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666199351
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666199351
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666199351
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666199351
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666199351
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666199351
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666199351
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666199351
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666199351
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666199351
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666199351
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666199351
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666199351
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666199351
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666199351
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666199351
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666199351
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp 1666199351
transform 1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1666199351
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1666199351
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_201
timestamp 1666199351
transform 1 0 19596 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_208
timestamp 1666199351
transform 1 0 20240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1666199351
transform 1 0 20884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_225
timestamp 1666199351
transform 1 0 21804 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1666199351
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_253
timestamp 1666199351
transform 1 0 24380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_257
timestamp 1666199351
transform 1 0 24748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_264
timestamp 1666199351
transform 1 0 25392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_289
timestamp 1666199351
transform 1 0 27692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_296
timestamp 1666199351
transform 1 0 28336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1666199351
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1666199351
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1666199351
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_314
timestamp 1666199351
transform 1 0 29992 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_326
timestamp 1666199351
transform 1 0 31096 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_338
timestamp 1666199351
transform 1 0 32200 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_350
timestamp 1666199351
transform 1 0 33304 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1666199351
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1666199351
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1666199351
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1666199351
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1666199351
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1666199351
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1666199351
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1666199351
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1666199351
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1666199351
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1666199351
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1666199351
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1666199351
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1666199351
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1666199351
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1666199351
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_513
timestamp 1666199351
transform 1 0 48300 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666199351
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666199351
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666199351
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666199351
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666199351
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666199351
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666199351
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666199351
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666199351
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666199351
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666199351
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666199351
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666199351
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666199351
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666199351
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666199351
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666199351
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666199351
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666199351
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666199351
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_193
timestamp 1666199351
transform 1 0 18860 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_196
timestamp 1666199351
transform 1 0 19136 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_203
timestamp 1666199351
transform 1 0 19780 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_207
timestamp 1666199351
transform 1 0 20148 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_211
timestamp 1666199351
transform 1 0 20516 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1666199351
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_225
timestamp 1666199351
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_229
timestamp 1666199351
transform 1 0 22172 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_233
timestamp 1666199351
transform 1 0 22540 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_240
timestamp 1666199351
transform 1 0 23184 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_244
timestamp 1666199351
transform 1 0 23552 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_248
timestamp 1666199351
transform 1 0 23920 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1666199351
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1666199351
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_281
timestamp 1666199351
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_308
timestamp 1666199351
transform 1 0 29440 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_320
timestamp 1666199351
transform 1 0 30544 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1666199351
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1666199351
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1666199351
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1666199351
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1666199351
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1666199351
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1666199351
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1666199351
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1666199351
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1666199351
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1666199351
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1666199351
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1666199351
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1666199351
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1666199351
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1666199351
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1666199351
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1666199351
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1666199351
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1666199351
transform 1 0 47564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_513
timestamp 1666199351
transform 1 0 48300 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666199351
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666199351
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666199351
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666199351
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666199351
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666199351
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666199351
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666199351
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666199351
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666199351
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666199351
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666199351
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666199351
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666199351
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666199351
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666199351
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666199351
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666199351
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666199351
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666199351
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666199351
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666199351
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_209
timestamp 1666199351
transform 1 0 20332 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_217
timestamp 1666199351
transform 1 0 21068 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_221
timestamp 1666199351
transform 1 0 21436 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_229
timestamp 1666199351
transform 1 0 22172 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_233
timestamp 1666199351
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_240
timestamp 1666199351
transform 1 0 23184 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_246
timestamp 1666199351
transform 1 0 23736 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1666199351
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1666199351
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_257
timestamp 1666199351
transform 1 0 24748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_267
timestamp 1666199351
transform 1 0 25668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_274
timestamp 1666199351
transform 1 0 26312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_281
timestamp 1666199351
transform 1 0 26956 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_287
timestamp 1666199351
transform 1 0 27508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_291
timestamp 1666199351
transform 1 0 27876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_298
timestamp 1666199351
transform 1 0 28520 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1666199351
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1666199351
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1666199351
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1666199351
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1666199351
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1666199351
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1666199351
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1666199351
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1666199351
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1666199351
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1666199351
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1666199351
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1666199351
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1666199351
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1666199351
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1666199351
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1666199351
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1666199351
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1666199351
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1666199351
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1666199351
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1666199351
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_513
timestamp 1666199351
transform 1 0 48300 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666199351
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666199351
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666199351
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1666199351
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1666199351
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666199351
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666199351
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666199351
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666199351
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666199351
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666199351
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666199351
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666199351
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666199351
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666199351
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666199351
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666199351
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666199351
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666199351
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666199351
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666199351
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666199351
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666199351
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666199351
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666199351
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_237
timestamp 1666199351
transform 1 0 22908 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_242
timestamp 1666199351
transform 1 0 23368 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_249
timestamp 1666199351
transform 1 0 24012 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_253
timestamp 1666199351
transform 1 0 24380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_257
timestamp 1666199351
transform 1 0 24748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_263
timestamp 1666199351
transform 1 0 25300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_270
timestamp 1666199351
transform 1 0 25944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1666199351
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666199351
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1666199351
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1666199351
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1666199351
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1666199351
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1666199351
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1666199351
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1666199351
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1666199351
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1666199351
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1666199351
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1666199351
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1666199351
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1666199351
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1666199351
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1666199351
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1666199351
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1666199351
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1666199351
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1666199351
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1666199351
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1666199351
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1666199351
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1666199351
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_505
timestamp 1666199351
transform 1 0 47564 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_513
timestamp 1666199351
transform 1 0 48300 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666199351
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666199351
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666199351
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666199351
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666199351
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666199351
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666199351
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666199351
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666199351
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666199351
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666199351
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666199351
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666199351
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666199351
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666199351
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666199351
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666199351
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666199351
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666199351
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666199351
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666199351
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666199351
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666199351
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666199351
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1666199351
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1666199351
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666199351
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1666199351
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1666199351
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1666199351
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1666199351
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1666199351
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1666199351
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1666199351
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1666199351
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1666199351
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1666199351
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1666199351
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1666199351
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1666199351
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1666199351
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1666199351
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1666199351
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1666199351
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1666199351
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1666199351
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1666199351
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1666199351
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1666199351
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1666199351
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1666199351
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1666199351
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1666199351
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1666199351
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_513
timestamp 1666199351
transform 1 0 48300 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666199351
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666199351
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666199351
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666199351
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666199351
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666199351
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666199351
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666199351
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666199351
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666199351
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666199351
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666199351
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666199351
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666199351
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666199351
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666199351
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666199351
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666199351
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666199351
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666199351
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666199351
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666199351
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666199351
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666199351
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1666199351
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1666199351
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1666199351
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1666199351
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1666199351
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666199351
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666199351
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1666199351
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1666199351
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1666199351
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1666199351
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1666199351
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1666199351
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1666199351
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1666199351
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1666199351
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1666199351
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1666199351
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1666199351
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1666199351
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1666199351
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1666199351
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1666199351
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1666199351
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1666199351
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1666199351
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1666199351
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1666199351
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1666199351
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1666199351
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1666199351
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1666199351
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666199351
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666199351
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666199351
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666199351
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666199351
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666199351
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666199351
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666199351
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666199351
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666199351
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666199351
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666199351
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666199351
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666199351
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666199351
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666199351
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666199351
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666199351
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666199351
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666199351
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666199351
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666199351
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666199351
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1666199351
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1666199351
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1666199351
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1666199351
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1666199351
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1666199351
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1666199351
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1666199351
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1666199351
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1666199351
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1666199351
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1666199351
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1666199351
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1666199351
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1666199351
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1666199351
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1666199351
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1666199351
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1666199351
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1666199351
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1666199351
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1666199351
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1666199351
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1666199351
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1666199351
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1666199351
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1666199351
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1666199351
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1666199351
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1666199351
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1666199351
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_513
timestamp 1666199351
transform 1 0 48300 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666199351
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666199351
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1666199351
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1666199351
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1666199351
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666199351
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666199351
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666199351
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666199351
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666199351
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666199351
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666199351
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666199351
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666199351
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666199351
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666199351
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666199351
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666199351
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666199351
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666199351
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666199351
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666199351
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666199351
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666199351
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666199351
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666199351
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666199351
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666199351
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666199351
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666199351
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1666199351
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1666199351
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1666199351
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1666199351
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1666199351
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1666199351
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1666199351
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1666199351
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1666199351
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1666199351
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1666199351
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1666199351
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1666199351
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1666199351
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1666199351
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1666199351
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1666199351
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1666199351
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1666199351
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1666199351
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1666199351
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1666199351
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1666199351
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1666199351
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1666199351
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1666199351
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666199351
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1666199351
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666199351
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666199351
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666199351
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666199351
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666199351
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666199351
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666199351
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666199351
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666199351
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666199351
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666199351
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666199351
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666199351
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666199351
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666199351
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666199351
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666199351
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666199351
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666199351
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666199351
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666199351
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1666199351
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1666199351
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1666199351
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666199351
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1666199351
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1666199351
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1666199351
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1666199351
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1666199351
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1666199351
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1666199351
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1666199351
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1666199351
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1666199351
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1666199351
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1666199351
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1666199351
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1666199351
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1666199351
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1666199351
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1666199351
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1666199351
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1666199351
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1666199351
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1666199351
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1666199351
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1666199351
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1666199351
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1666199351
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1666199351
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1666199351
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_513
timestamp 1666199351
transform 1 0 48300 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666199351
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666199351
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666199351
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666199351
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1666199351
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666199351
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666199351
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666199351
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666199351
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666199351
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666199351
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666199351
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666199351
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666199351
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666199351
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666199351
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666199351
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666199351
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666199351
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666199351
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666199351
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666199351
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666199351
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666199351
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666199351
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666199351
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1666199351
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666199351
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1666199351
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666199351
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1666199351
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1666199351
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1666199351
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1666199351
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1666199351
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1666199351
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1666199351
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1666199351
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1666199351
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1666199351
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1666199351
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1666199351
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1666199351
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1666199351
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1666199351
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1666199351
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1666199351
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1666199351
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1666199351
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1666199351
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1666199351
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1666199351
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1666199351
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1666199351
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1666199351
transform 1 0 47564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_513
timestamp 1666199351
transform 1 0 48300 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666199351
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666199351
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666199351
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666199351
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666199351
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666199351
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666199351
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666199351
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666199351
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666199351
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666199351
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666199351
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666199351
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666199351
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666199351
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666199351
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666199351
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666199351
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666199351
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666199351
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666199351
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666199351
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666199351
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666199351
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1666199351
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1666199351
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666199351
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666199351
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1666199351
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1666199351
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1666199351
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1666199351
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1666199351
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1666199351
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1666199351
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1666199351
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1666199351
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1666199351
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1666199351
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1666199351
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1666199351
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1666199351
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1666199351
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1666199351
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1666199351
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1666199351
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1666199351
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1666199351
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1666199351
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1666199351
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1666199351
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1666199351
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1666199351
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1666199351
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_513
timestamp 1666199351
transform 1 0 48300 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666199351
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666199351
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1666199351
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1666199351
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1666199351
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666199351
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666199351
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666199351
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666199351
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666199351
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666199351
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666199351
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666199351
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666199351
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666199351
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666199351
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666199351
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666199351
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666199351
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666199351
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666199351
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666199351
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666199351
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666199351
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1666199351
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1666199351
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1666199351
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1666199351
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666199351
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666199351
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1666199351
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1666199351
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1666199351
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1666199351
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1666199351
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1666199351
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1666199351
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1666199351
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1666199351
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1666199351
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1666199351
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1666199351
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1666199351
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1666199351
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1666199351
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1666199351
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1666199351
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1666199351
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1666199351
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1666199351
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1666199351
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1666199351
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1666199351
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1666199351
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1666199351
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_513
timestamp 1666199351
transform 1 0 48300 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666199351
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1666199351
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666199351
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666199351
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666199351
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666199351
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666199351
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666199351
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666199351
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666199351
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666199351
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666199351
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666199351
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666199351
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666199351
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666199351
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666199351
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666199351
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666199351
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666199351
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666199351
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666199351
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666199351
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1666199351
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1666199351
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1666199351
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666199351
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1666199351
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1666199351
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1666199351
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1666199351
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1666199351
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1666199351
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1666199351
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1666199351
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1666199351
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1666199351
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1666199351
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1666199351
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1666199351
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1666199351
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1666199351
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1666199351
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1666199351
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1666199351
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1666199351
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1666199351
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1666199351
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1666199351
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1666199351
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1666199351
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1666199351
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1666199351
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1666199351
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1666199351
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666199351
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666199351
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666199351
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666199351
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666199351
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666199351
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666199351
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666199351
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666199351
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666199351
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666199351
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666199351
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666199351
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666199351
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666199351
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666199351
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666199351
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666199351
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666199351
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666199351
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666199351
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666199351
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666199351
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666199351
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666199351
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1666199351
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1666199351
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1666199351
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1666199351
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666199351
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1666199351
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1666199351
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1666199351
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1666199351
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1666199351
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1666199351
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1666199351
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1666199351
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1666199351
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1666199351
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1666199351
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1666199351
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1666199351
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1666199351
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1666199351
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1666199351
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1666199351
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1666199351
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1666199351
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1666199351
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1666199351
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1666199351
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1666199351
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1666199351
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1666199351
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1666199351
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1666199351
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1666199351
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666199351
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666199351
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666199351
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666199351
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666199351
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666199351
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666199351
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666199351
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666199351
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666199351
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666199351
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666199351
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666199351
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666199351
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666199351
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666199351
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666199351
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666199351
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666199351
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666199351
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666199351
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666199351
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1666199351
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1666199351
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1666199351
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1666199351
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1666199351
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1666199351
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1666199351
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1666199351
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1666199351
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1666199351
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1666199351
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1666199351
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1666199351
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1666199351
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1666199351
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1666199351
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1666199351
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1666199351
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1666199351
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1666199351
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1666199351
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1666199351
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1666199351
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1666199351
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1666199351
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1666199351
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1666199351
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1666199351
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1666199351
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1666199351
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_513
timestamp 1666199351
transform 1 0 48300 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666199351
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666199351
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666199351
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666199351
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666199351
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666199351
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666199351
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666199351
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666199351
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666199351
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666199351
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666199351
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666199351
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666199351
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666199351
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666199351
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666199351
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666199351
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666199351
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666199351
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666199351
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666199351
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666199351
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666199351
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1666199351
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1666199351
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1666199351
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1666199351
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1666199351
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666199351
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1666199351
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1666199351
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1666199351
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1666199351
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1666199351
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1666199351
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1666199351
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1666199351
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1666199351
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1666199351
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1666199351
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1666199351
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1666199351
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1666199351
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1666199351
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1666199351
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1666199351
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1666199351
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1666199351
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1666199351
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1666199351
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1666199351
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1666199351
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1666199351
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1666199351
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_513
timestamp 1666199351
transform 1 0 48300 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666199351
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1666199351
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666199351
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666199351
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666199351
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666199351
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666199351
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666199351
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666199351
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666199351
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666199351
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666199351
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666199351
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666199351
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666199351
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666199351
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666199351
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666199351
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666199351
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666199351
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666199351
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666199351
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666199351
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666199351
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1666199351
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1666199351
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1666199351
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1666199351
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1666199351
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1666199351
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1666199351
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1666199351
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1666199351
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1666199351
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1666199351
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1666199351
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1666199351
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1666199351
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1666199351
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1666199351
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1666199351
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1666199351
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1666199351
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1666199351
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1666199351
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1666199351
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1666199351
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1666199351
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1666199351
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1666199351
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1666199351
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1666199351
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1666199351
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1666199351
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1666199351
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666199351
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666199351
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666199351
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666199351
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666199351
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666199351
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666199351
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666199351
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666199351
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666199351
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666199351
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666199351
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666199351
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666199351
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666199351
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666199351
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666199351
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666199351
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666199351
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666199351
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666199351
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666199351
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666199351
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666199351
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1666199351
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1666199351
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1666199351
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1666199351
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1666199351
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1666199351
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1666199351
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1666199351
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1666199351
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1666199351
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1666199351
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1666199351
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1666199351
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1666199351
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1666199351
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1666199351
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1666199351
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1666199351
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1666199351
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1666199351
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1666199351
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1666199351
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1666199351
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1666199351
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1666199351
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1666199351
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1666199351
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1666199351
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1666199351
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1666199351
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1666199351
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1666199351
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666199351
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1666199351
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666199351
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666199351
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666199351
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666199351
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666199351
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666199351
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666199351
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666199351
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666199351
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666199351
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666199351
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666199351
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666199351
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666199351
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666199351
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666199351
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666199351
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666199351
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666199351
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666199351
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666199351
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1666199351
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1666199351
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1666199351
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1666199351
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1666199351
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1666199351
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1666199351
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1666199351
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1666199351
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1666199351
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1666199351
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1666199351
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1666199351
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1666199351
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1666199351
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1666199351
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1666199351
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1666199351
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1666199351
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1666199351
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1666199351
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1666199351
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1666199351
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1666199351
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1666199351
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1666199351
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1666199351
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1666199351
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1666199351
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1666199351
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1666199351
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_513
timestamp 1666199351
transform 1 0 48300 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666199351
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666199351
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666199351
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1666199351
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1666199351
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666199351
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666199351
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666199351
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666199351
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666199351
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666199351
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666199351
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666199351
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666199351
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666199351
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666199351
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666199351
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666199351
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666199351
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666199351
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666199351
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666199351
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666199351
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666199351
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1666199351
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1666199351
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1666199351
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1666199351
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1666199351
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1666199351
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1666199351
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1666199351
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1666199351
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1666199351
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1666199351
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1666199351
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1666199351
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1666199351
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1666199351
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1666199351
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1666199351
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1666199351
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1666199351
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1666199351
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1666199351
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1666199351
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1666199351
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1666199351
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1666199351
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1666199351
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1666199351
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1666199351
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1666199351
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1666199351
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_505
timestamp 1666199351
transform 1 0 47564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_513
timestamp 1666199351
transform 1 0 48300 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666199351
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666199351
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666199351
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666199351
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666199351
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666199351
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666199351
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666199351
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666199351
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666199351
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666199351
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666199351
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666199351
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666199351
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666199351
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666199351
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666199351
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666199351
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666199351
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666199351
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666199351
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666199351
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666199351
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1666199351
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1666199351
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1666199351
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1666199351
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1666199351
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1666199351
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1666199351
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1666199351
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1666199351
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1666199351
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1666199351
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1666199351
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1666199351
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1666199351
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1666199351
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1666199351
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1666199351
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1666199351
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1666199351
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1666199351
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1666199351
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1666199351
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1666199351
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1666199351
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1666199351
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1666199351
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1666199351
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1666199351
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1666199351
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1666199351
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1666199351
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_513
timestamp 1666199351
transform 1 0 48300 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666199351
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666199351
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666199351
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666199351
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666199351
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666199351
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666199351
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666199351
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666199351
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666199351
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666199351
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666199351
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666199351
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666199351
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666199351
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666199351
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666199351
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666199351
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666199351
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666199351
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666199351
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666199351
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666199351
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666199351
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1666199351
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1666199351
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1666199351
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1666199351
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1666199351
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1666199351
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1666199351
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1666199351
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1666199351
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1666199351
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1666199351
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1666199351
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1666199351
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1666199351
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1666199351
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1666199351
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1666199351
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1666199351
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1666199351
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1666199351
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1666199351
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1666199351
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1666199351
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1666199351
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1666199351
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1666199351
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1666199351
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1666199351
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1666199351
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1666199351
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1666199351
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_513
timestamp 1666199351
transform 1 0 48300 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666199351
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1666199351
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666199351
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666199351
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666199351
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666199351
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666199351
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666199351
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666199351
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666199351
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666199351
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666199351
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666199351
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666199351
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666199351
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666199351
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666199351
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666199351
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666199351
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666199351
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666199351
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666199351
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666199351
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666199351
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1666199351
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1666199351
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1666199351
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1666199351
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1666199351
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1666199351
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1666199351
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1666199351
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1666199351
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1666199351
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1666199351
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1666199351
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1666199351
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1666199351
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1666199351
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1666199351
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1666199351
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1666199351
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1666199351
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1666199351
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1666199351
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1666199351
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1666199351
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1666199351
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1666199351
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1666199351
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1666199351
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1666199351
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1666199351
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1666199351
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_513
timestamp 1666199351
transform 1 0 48300 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666199351
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1666199351
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1666199351
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1666199351
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1666199351
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1666199351
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666199351
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666199351
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666199351
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666199351
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666199351
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666199351
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666199351
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666199351
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666199351
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666199351
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666199351
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666199351
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666199351
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666199351
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666199351
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666199351
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666199351
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666199351
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1666199351
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1666199351
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1666199351
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1666199351
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1666199351
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1666199351
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1666199351
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1666199351
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1666199351
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1666199351
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1666199351
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1666199351
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1666199351
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1666199351
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1666199351
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1666199351
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1666199351
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1666199351
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1666199351
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1666199351
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1666199351
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1666199351
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1666199351
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1666199351
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1666199351
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1666199351
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1666199351
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1666199351
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1666199351
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1666199351
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1666199351
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_513
timestamp 1666199351
transform 1 0 48300 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666199351
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666199351
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666199351
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666199351
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666199351
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666199351
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666199351
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666199351
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666199351
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666199351
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666199351
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666199351
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666199351
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666199351
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666199351
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666199351
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666199351
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666199351
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666199351
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666199351
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666199351
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666199351
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666199351
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1666199351
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1666199351
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1666199351
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1666199351
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1666199351
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1666199351
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1666199351
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1666199351
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1666199351
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1666199351
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1666199351
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1666199351
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1666199351
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1666199351
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1666199351
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1666199351
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1666199351
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1666199351
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1666199351
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1666199351
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1666199351
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1666199351
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1666199351
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1666199351
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1666199351
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1666199351
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1666199351
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1666199351
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1666199351
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1666199351
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1666199351
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_513
timestamp 1666199351
transform 1 0 48300 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666199351
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666199351
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666199351
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666199351
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666199351
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666199351
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666199351
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666199351
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666199351
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666199351
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666199351
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666199351
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666199351
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666199351
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666199351
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666199351
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666199351
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666199351
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666199351
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666199351
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666199351
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666199351
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666199351
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666199351
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1666199351
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1666199351
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1666199351
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1666199351
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1666199351
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1666199351
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1666199351
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1666199351
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1666199351
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1666199351
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1666199351
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1666199351
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1666199351
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1666199351
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1666199351
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1666199351
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1666199351
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1666199351
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1666199351
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1666199351
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1666199351
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1666199351
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1666199351
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1666199351
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1666199351
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1666199351
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1666199351
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1666199351
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1666199351
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1666199351
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_505
timestamp 1666199351
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_513
timestamp 1666199351
transform 1 0 48300 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666199351
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666199351
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666199351
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666199351
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666199351
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666199351
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666199351
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666199351
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666199351
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666199351
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666199351
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666199351
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666199351
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666199351
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666199351
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666199351
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666199351
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666199351
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666199351
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666199351
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666199351
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666199351
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1666199351
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1666199351
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1666199351
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1666199351
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1666199351
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1666199351
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1666199351
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1666199351
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1666199351
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1666199351
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1666199351
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1666199351
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1666199351
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1666199351
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1666199351
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1666199351
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1666199351
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1666199351
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1666199351
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1666199351
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1666199351
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1666199351
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1666199351
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1666199351
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1666199351
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1666199351
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1666199351
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1666199351
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1666199351
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1666199351
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1666199351
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1666199351
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_513
timestamp 1666199351
transform 1 0 48300 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666199351
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666199351
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1666199351
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666199351
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666199351
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666199351
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666199351
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666199351
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666199351
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666199351
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666199351
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666199351
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666199351
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666199351
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666199351
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666199351
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666199351
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666199351
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666199351
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666199351
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666199351
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1666199351
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666199351
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666199351
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1666199351
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1666199351
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1666199351
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1666199351
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1666199351
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1666199351
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1666199351
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1666199351
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1666199351
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1666199351
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1666199351
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1666199351
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1666199351
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1666199351
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1666199351
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1666199351
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1666199351
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1666199351
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1666199351
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1666199351
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1666199351
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1666199351
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1666199351
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1666199351
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1666199351
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1666199351
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1666199351
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1666199351
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1666199351
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1666199351
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1666199351
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_513
timestamp 1666199351
transform 1 0 48300 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666199351
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666199351
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666199351
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666199351
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666199351
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666199351
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666199351
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666199351
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666199351
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666199351
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666199351
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666199351
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666199351
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666199351
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666199351
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666199351
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666199351
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666199351
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666199351
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666199351
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666199351
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666199351
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666199351
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666199351
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1666199351
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1666199351
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1666199351
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1666199351
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1666199351
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1666199351
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1666199351
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1666199351
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1666199351
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1666199351
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1666199351
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1666199351
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1666199351
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1666199351
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1666199351
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1666199351
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1666199351
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1666199351
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1666199351
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1666199351
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1666199351
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1666199351
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1666199351
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1666199351
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1666199351
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1666199351
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1666199351
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1666199351
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1666199351
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1666199351
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_513
timestamp 1666199351
transform 1 0 48300 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666199351
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666199351
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1666199351
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1666199351
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1666199351
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666199351
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666199351
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666199351
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666199351
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666199351
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666199351
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666199351
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666199351
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666199351
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666199351
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666199351
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666199351
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666199351
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666199351
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666199351
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1666199351
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1666199351
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1666199351
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1666199351
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1666199351
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1666199351
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1666199351
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1666199351
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1666199351
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1666199351
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1666199351
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1666199351
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1666199351
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1666199351
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1666199351
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1666199351
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1666199351
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1666199351
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1666199351
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1666199351
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1666199351
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1666199351
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1666199351
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1666199351
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1666199351
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1666199351
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1666199351
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1666199351
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1666199351
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1666199351
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1666199351
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1666199351
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1666199351
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1666199351
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1666199351
transform 1 0 47564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_513
timestamp 1666199351
transform 1 0 48300 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666199351
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666199351
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666199351
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666199351
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666199351
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666199351
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666199351
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666199351
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666199351
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666199351
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666199351
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666199351
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666199351
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666199351
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666199351
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666199351
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666199351
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666199351
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1666199351
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1666199351
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1666199351
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1666199351
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1666199351
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1666199351
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1666199351
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1666199351
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666199351
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1666199351
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1666199351
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1666199351
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1666199351
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1666199351
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1666199351
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1666199351
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1666199351
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1666199351
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1666199351
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1666199351
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1666199351
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1666199351
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1666199351
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1666199351
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1666199351
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1666199351
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1666199351
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1666199351
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1666199351
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1666199351
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1666199351
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1666199351
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1666199351
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1666199351
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1666199351
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1666199351
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_513
timestamp 1666199351
transform 1 0 48300 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666199351
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666199351
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1666199351
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1666199351
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1666199351
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1666199351
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666199351
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666199351
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666199351
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666199351
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666199351
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666199351
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666199351
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666199351
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666199351
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666199351
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666199351
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666199351
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1666199351
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1666199351
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1666199351
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1666199351
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1666199351
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666199351
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1666199351
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1666199351
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1666199351
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1666199351
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1666199351
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666199351
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1666199351
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1666199351
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1666199351
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1666199351
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1666199351
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1666199351
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1666199351
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1666199351
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1666199351
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1666199351
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1666199351
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1666199351
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1666199351
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1666199351
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1666199351
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1666199351
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1666199351
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1666199351
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1666199351
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1666199351
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1666199351
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1666199351
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1666199351
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1666199351
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1666199351
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_513
timestamp 1666199351
transform 1 0 48300 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666199351
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666199351
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666199351
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666199351
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666199351
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666199351
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666199351
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666199351
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666199351
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666199351
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666199351
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666199351
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666199351
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666199351
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666199351
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666199351
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1666199351
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1666199351
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1666199351
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1666199351
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666199351
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1666199351
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1666199351
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1666199351
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1666199351
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1666199351
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1666199351
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1666199351
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1666199351
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1666199351
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1666199351
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1666199351
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1666199351
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1666199351
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1666199351
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1666199351
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1666199351
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1666199351
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1666199351
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1666199351
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1666199351
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1666199351
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1666199351
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1666199351
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1666199351
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1666199351
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1666199351
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1666199351
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1666199351
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1666199351
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1666199351
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1666199351
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1666199351
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1666199351
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_513
timestamp 1666199351
transform 1 0 48300 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1666199351
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666199351
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1666199351
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1666199351
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1666199351
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1666199351
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666199351
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666199351
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666199351
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666199351
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666199351
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666199351
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666199351
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666199351
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666199351
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1666199351
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666199351
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666199351
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666199351
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1666199351
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1666199351
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1666199351
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1666199351
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666199351
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1666199351
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1666199351
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1666199351
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1666199351
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1666199351
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1666199351
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1666199351
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1666199351
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1666199351
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1666199351
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1666199351
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1666199351
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1666199351
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1666199351
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1666199351
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1666199351
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1666199351
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1666199351
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1666199351
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1666199351
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1666199351
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1666199351
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1666199351
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1666199351
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1666199351
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1666199351
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1666199351
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1666199351
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1666199351
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1666199351
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1666199351
transform 1 0 47564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_513
timestamp 1666199351
transform 1 0 48300 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666199351
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1666199351
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666199351
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666199351
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666199351
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666199351
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666199351
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666199351
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666199351
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666199351
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666199351
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666199351
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666199351
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666199351
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666199351
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666199351
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1666199351
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1666199351
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1666199351
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1666199351
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1666199351
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666199351
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1666199351
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1666199351
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1666199351
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1666199351
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1666199351
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1666199351
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1666199351
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1666199351
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1666199351
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1666199351
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1666199351
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1666199351
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1666199351
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1666199351
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1666199351
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1666199351
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1666199351
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1666199351
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1666199351
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1666199351
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1666199351
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1666199351
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1666199351
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1666199351
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1666199351
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1666199351
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1666199351
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1666199351
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1666199351
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1666199351
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1666199351
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1666199351
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_513
timestamp 1666199351
transform 1 0 48300 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666199351
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666199351
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666199351
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666199351
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666199351
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666199351
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666199351
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666199351
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666199351
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666199351
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666199351
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666199351
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666199351
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666199351
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666199351
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1666199351
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1666199351
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1666199351
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666199351
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1666199351
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1666199351
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1666199351
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1666199351
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1666199351
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1666199351
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1666199351
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1666199351
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1666199351
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1666199351
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1666199351
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666199351
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1666199351
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1666199351
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1666199351
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1666199351
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1666199351
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1666199351
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1666199351
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1666199351
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1666199351
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1666199351
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1666199351
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1666199351
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1666199351
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1666199351
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1666199351
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1666199351
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1666199351
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1666199351
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1666199351
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1666199351
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1666199351
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1666199351
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1666199351
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_505
timestamp 1666199351
transform 1 0 47564 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_513
timestamp 1666199351
transform 1 0 48300 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666199351
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1666199351
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666199351
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666199351
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666199351
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666199351
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666199351
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666199351
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666199351
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666199351
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666199351
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1666199351
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1666199351
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1666199351
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666199351
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666199351
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1666199351
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1666199351
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1666199351
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1666199351
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1666199351
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1666199351
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1666199351
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1666199351
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1666199351
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1666199351
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666199351
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1666199351
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1666199351
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1666199351
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1666199351
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1666199351
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1666199351
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1666199351
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1666199351
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1666199351
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1666199351
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1666199351
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1666199351
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1666199351
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1666199351
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1666199351
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1666199351
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1666199351
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1666199351
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1666199351
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1666199351
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1666199351
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1666199351
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1666199351
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1666199351
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1666199351
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1666199351
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1666199351
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_513
timestamp 1666199351
transform 1 0 48300 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666199351
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666199351
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1666199351
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1666199351
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1666199351
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666199351
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666199351
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666199351
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666199351
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1666199351
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666199351
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666199351
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666199351
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1666199351
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1666199351
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1666199351
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1666199351
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1666199351
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1666199351
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1666199351
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1666199351
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1666199351
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1666199351
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1666199351
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666199351
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666199351
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1666199351
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1666199351
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1666199351
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1666199351
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1666199351
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1666199351
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1666199351
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1666199351
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1666199351
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1666199351
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1666199351
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1666199351
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1666199351
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1666199351
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1666199351
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1666199351
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1666199351
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1666199351
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1666199351
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1666199351
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1666199351
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1666199351
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1666199351
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1666199351
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1666199351
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1666199351
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1666199351
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1666199351
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_505
timestamp 1666199351
transform 1 0 47564 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_513
timestamp 1666199351
transform 1 0 48300 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666199351
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1666199351
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666199351
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666199351
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666199351
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666199351
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666199351
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666199351
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666199351
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1666199351
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1666199351
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1666199351
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1666199351
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1666199351
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666199351
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666199351
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666199351
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1666199351
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1666199351
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1666199351
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1666199351
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1666199351
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1666199351
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1666199351
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1666199351
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1666199351
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666199351
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1666199351
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1666199351
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1666199351
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1666199351
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1666199351
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1666199351
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1666199351
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1666199351
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1666199351
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1666199351
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1666199351
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1666199351
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1666199351
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1666199351
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1666199351
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1666199351
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1666199351
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1666199351
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1666199351
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1666199351
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1666199351
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1666199351
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1666199351
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1666199351
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1666199351
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1666199351
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1666199351
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_513
timestamp 1666199351
transform 1 0 48300 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666199351
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666199351
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666199351
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666199351
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666199351
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666199351
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666199351
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666199351
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1666199351
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1666199351
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1666199351
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666199351
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1666199351
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1666199351
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1666199351
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1666199351
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666199351
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666199351
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666199351
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1666199351
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1666199351
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1666199351
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1666199351
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666199351
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1666199351
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1666199351
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1666199351
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1666199351
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1666199351
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1666199351
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1666199351
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1666199351
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1666199351
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1666199351
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1666199351
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1666199351
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1666199351
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1666199351
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1666199351
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1666199351
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1666199351
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1666199351
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1666199351
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1666199351
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1666199351
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1666199351
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1666199351
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1666199351
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1666199351
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1666199351
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1666199351
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1666199351
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1666199351
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1666199351
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1666199351
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1666199351
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666199351
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666199351
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666199351
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666199351
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666199351
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666199351
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666199351
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1666199351
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666199351
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1666199351
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1666199351
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1666199351
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1666199351
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1666199351
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666199351
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1666199351
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1666199351
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1666199351
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1666199351
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1666199351
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666199351
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666199351
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1666199351
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1666199351
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1666199351
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1666199351
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1666199351
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1666199351
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1666199351
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1666199351
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1666199351
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1666199351
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1666199351
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1666199351
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1666199351
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1666199351
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1666199351
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1666199351
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1666199351
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1666199351
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1666199351
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1666199351
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1666199351
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1666199351
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1666199351
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1666199351
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1666199351
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1666199351
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1666199351
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1666199351
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1666199351
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1666199351
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1666199351
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1666199351
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_513
timestamp 1666199351
transform 1 0 48300 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666199351
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666199351
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666199351
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1666199351
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1666199351
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666199351
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666199351
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1666199351
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1666199351
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1666199351
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1666199351
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666199351
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1666199351
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1666199351
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666199351
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1666199351
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1666199351
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1666199351
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1666199351
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1666199351
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1666199351
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1666199351
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1666199351
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1666199351
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1666199351
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1666199351
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1666199351
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1666199351
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1666199351
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1666199351
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1666199351
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1666199351
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1666199351
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1666199351
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1666199351
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1666199351
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1666199351
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1666199351
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1666199351
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1666199351
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1666199351
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1666199351
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1666199351
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1666199351
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1666199351
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1666199351
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1666199351
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1666199351
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1666199351
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1666199351
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1666199351
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1666199351
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1666199351
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1666199351
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_505
timestamp 1666199351
transform 1 0 47564 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_513
timestamp 1666199351
transform 1 0 48300 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666199351
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1666199351
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666199351
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666199351
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666199351
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666199351
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666199351
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666199351
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666199351
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1666199351
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1666199351
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1666199351
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1666199351
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1666199351
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666199351
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1666199351
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1666199351
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1666199351
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1666199351
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1666199351
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1666199351
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1666199351
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1666199351
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1666199351
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1666199351
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1666199351
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1666199351
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1666199351
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1666199351
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1666199351
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1666199351
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1666199351
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1666199351
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1666199351
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1666199351
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1666199351
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1666199351
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1666199351
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1666199351
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1666199351
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1666199351
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1666199351
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1666199351
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1666199351
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1666199351
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1666199351
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1666199351
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1666199351
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1666199351
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1666199351
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1666199351
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1666199351
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1666199351
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1666199351
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_513
timestamp 1666199351
transform 1 0 48300 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666199351
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666199351
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666199351
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666199351
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666199351
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666199351
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666199351
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1666199351
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1666199351
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1666199351
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1666199351
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1666199351
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1666199351
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1666199351
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1666199351
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1666199351
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1666199351
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666199351
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1666199351
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1666199351
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1666199351
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1666199351
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1666199351
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1666199351
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1666199351
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1666199351
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1666199351
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1666199351
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1666199351
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1666199351
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1666199351
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1666199351
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1666199351
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1666199351
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1666199351
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1666199351
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1666199351
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1666199351
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1666199351
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1666199351
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1666199351
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1666199351
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1666199351
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1666199351
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1666199351
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1666199351
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1666199351
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1666199351
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1666199351
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1666199351
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1666199351
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1666199351
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1666199351
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1666199351
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1666199351
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1666199351
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666199351
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666199351
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666199351
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666199351
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666199351
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666199351
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666199351
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666199351
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666199351
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1666199351
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1666199351
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1666199351
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1666199351
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1666199351
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1666199351
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1666199351
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1666199351
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1666199351
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1666199351
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1666199351
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666199351
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1666199351
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1666199351
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1666199351
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1666199351
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1666199351
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1666199351
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1666199351
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1666199351
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1666199351
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1666199351
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1666199351
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666199351
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1666199351
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1666199351
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1666199351
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1666199351
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1666199351
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1666199351
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1666199351
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1666199351
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1666199351
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1666199351
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1666199351
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1666199351
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1666199351
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1666199351
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1666199351
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1666199351
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1666199351
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1666199351
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1666199351
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1666199351
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1666199351
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_513
timestamp 1666199351
transform 1 0 48300 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666199351
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666199351
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666199351
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666199351
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666199351
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666199351
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666199351
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666199351
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666199351
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666199351
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666199351
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666199351
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666199351
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1666199351
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1666199351
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1666199351
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1666199351
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666199351
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1666199351
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1666199351
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1666199351
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1666199351
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1666199351
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666199351
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1666199351
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1666199351
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1666199351
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1666199351
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1666199351
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666199351
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1666199351
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1666199351
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1666199351
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1666199351
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1666199351
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1666199351
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1666199351
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1666199351
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1666199351
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1666199351
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1666199351
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1666199351
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1666199351
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1666199351
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1666199351
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1666199351
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1666199351
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1666199351
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1666199351
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1666199351
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1666199351
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1666199351
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1666199351
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1666199351
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1666199351
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1666199351
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666199351
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666199351
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666199351
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666199351
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666199351
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666199351
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666199351
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666199351
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666199351
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1666199351
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1666199351
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1666199351
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1666199351
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1666199351
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666199351
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1666199351
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1666199351
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1666199351
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1666199351
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1666199351
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1666199351
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1666199351
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1666199351
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1666199351
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1666199351
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1666199351
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1666199351
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1666199351
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1666199351
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1666199351
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1666199351
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1666199351
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666199351
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1666199351
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1666199351
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1666199351
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1666199351
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1666199351
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1666199351
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1666199351
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1666199351
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1666199351
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1666199351
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1666199351
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1666199351
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1666199351
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1666199351
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1666199351
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1666199351
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1666199351
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1666199351
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1666199351
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1666199351
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1666199351
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1666199351
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666199351
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666199351
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666199351
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1666199351
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1666199351
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1666199351
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666199351
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666199351
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666199351
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1666199351
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1666199351
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666199351
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666199351
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1666199351
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1666199351
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1666199351
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1666199351
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666199351
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1666199351
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1666199351
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1666199351
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1666199351
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1666199351
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1666199351
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1666199351
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1666199351
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1666199351
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1666199351
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1666199351
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1666199351
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1666199351
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1666199351
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1666199351
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1666199351
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1666199351
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1666199351
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1666199351
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1666199351
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1666199351
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1666199351
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1666199351
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1666199351
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1666199351
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1666199351
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1666199351
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1666199351
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1666199351
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1666199351
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1666199351
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1666199351
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1666199351
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1666199351
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1666199351
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1666199351
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1666199351
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1666199351
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666199351
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1666199351
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666199351
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666199351
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666199351
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666199351
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666199351
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666199351
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666199351
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666199351
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666199351
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1666199351
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1666199351
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1666199351
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666199351
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1666199351
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1666199351
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1666199351
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1666199351
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1666199351
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1666199351
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1666199351
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1666199351
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1666199351
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1666199351
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1666199351
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1666199351
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1666199351
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1666199351
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1666199351
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1666199351
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1666199351
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1666199351
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1666199351
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1666199351
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1666199351
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1666199351
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1666199351
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1666199351
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1666199351
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1666199351
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1666199351
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1666199351
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1666199351
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1666199351
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1666199351
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1666199351
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1666199351
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1666199351
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1666199351
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1666199351
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1666199351
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1666199351
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1666199351
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_513
timestamp 1666199351
transform 1 0 48300 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666199351
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666199351
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666199351
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666199351
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666199351
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666199351
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666199351
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666199351
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1666199351
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666199351
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666199351
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666199351
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1666199351
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1666199351
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666199351
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666199351
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666199351
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666199351
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1666199351
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1666199351
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1666199351
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1666199351
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1666199351
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1666199351
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1666199351
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1666199351
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1666199351
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1666199351
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1666199351
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1666199351
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1666199351
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1666199351
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1666199351
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1666199351
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1666199351
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1666199351
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1666199351
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1666199351
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1666199351
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1666199351
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1666199351
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1666199351
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1666199351
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1666199351
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1666199351
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1666199351
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1666199351
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1666199351
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1666199351
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1666199351
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1666199351
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1666199351
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1666199351
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1666199351
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1666199351
transform 1 0 47564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_513
timestamp 1666199351
transform 1 0 48300 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666199351
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666199351
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666199351
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666199351
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666199351
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666199351
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666199351
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666199351
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666199351
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666199351
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1666199351
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1666199351
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1666199351
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1666199351
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666199351
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666199351
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1666199351
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1666199351
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1666199351
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1666199351
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1666199351
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1666199351
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1666199351
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1666199351
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1666199351
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1666199351
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666199351
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1666199351
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1666199351
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1666199351
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1666199351
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1666199351
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1666199351
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1666199351
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1666199351
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1666199351
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1666199351
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1666199351
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1666199351
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1666199351
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1666199351
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1666199351
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1666199351
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1666199351
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1666199351
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1666199351
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1666199351
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1666199351
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1666199351
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1666199351
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1666199351
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1666199351
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1666199351
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1666199351
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_513
timestamp 1666199351
transform 1 0 48300 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666199351
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666199351
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1666199351
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1666199351
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1666199351
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1666199351
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666199351
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1666199351
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1666199351
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1666199351
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1666199351
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666199351
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666199351
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666199351
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1666199351
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1666199351
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1666199351
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666199351
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1666199351
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1666199351
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1666199351
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1666199351
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1666199351
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1666199351
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1666199351
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1666199351
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1666199351
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1666199351
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1666199351
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1666199351
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1666199351
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1666199351
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1666199351
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1666199351
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1666199351
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1666199351
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1666199351
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1666199351
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1666199351
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1666199351
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1666199351
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1666199351
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1666199351
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1666199351
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1666199351
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1666199351
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1666199351
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1666199351
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1666199351
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1666199351
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1666199351
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1666199351
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1666199351
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1666199351
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_505
timestamp 1666199351
transform 1 0 47564 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_513
timestamp 1666199351
transform 1 0 48300 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1666199351
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1666199351
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666199351
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1666199351
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1666199351
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1666199351
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666199351
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1666199351
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666199351
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1666199351
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1666199351
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1666199351
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1666199351
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1666199351
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666199351
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1666199351
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1666199351
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1666199351
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1666199351
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1666199351
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1666199351
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1666199351
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1666199351
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1666199351
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1666199351
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1666199351
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1666199351
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1666199351
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1666199351
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1666199351
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1666199351
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1666199351
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1666199351
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1666199351
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1666199351
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1666199351
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1666199351
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1666199351
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1666199351
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1666199351
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1666199351
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1666199351
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1666199351
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1666199351
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1666199351
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1666199351
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1666199351
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1666199351
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1666199351
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1666199351
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1666199351
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1666199351
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1666199351
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1666199351
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_513
timestamp 1666199351
transform 1 0 48300 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1666199351
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666199351
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1666199351
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1666199351
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1666199351
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1666199351
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1666199351
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1666199351
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1666199351
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1666199351
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1666199351
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666199351
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1666199351
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1666199351
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1666199351
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1666199351
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1666199351
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1666199351
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1666199351
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1666199351
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1666199351
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1666199351
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1666199351
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1666199351
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1666199351
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1666199351
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1666199351
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1666199351
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1666199351
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1666199351
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1666199351
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1666199351
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1666199351
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1666199351
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1666199351
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1666199351
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1666199351
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1666199351
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1666199351
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1666199351
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1666199351
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1666199351
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1666199351
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1666199351
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1666199351
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1666199351
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1666199351
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1666199351
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1666199351
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1666199351
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1666199351
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1666199351
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1666199351
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1666199351
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1666199351
transform 1 0 47564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_513
timestamp 1666199351
transform 1 0 48300 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1666199351
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1666199351
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1666199351
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1666199351
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1666199351
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1666199351
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1666199351
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1666199351
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666199351
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1666199351
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1666199351
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1666199351
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1666199351
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1666199351
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666199351
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1666199351
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1666199351
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1666199351
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1666199351
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1666199351
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1666199351
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1666199351
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1666199351
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1666199351
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1666199351
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1666199351
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1666199351
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1666199351
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1666199351
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1666199351
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1666199351
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1666199351
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1666199351
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1666199351
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1666199351
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1666199351
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1666199351
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1666199351
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1666199351
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1666199351
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1666199351
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1666199351
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1666199351
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1666199351
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1666199351
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1666199351
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1666199351
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1666199351
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1666199351
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1666199351
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1666199351
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1666199351
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1666199351
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1666199351
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_513
timestamp 1666199351
transform 1 0 48300 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1666199351
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1666199351
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1666199351
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1666199351
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1666199351
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1666199351
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1666199351
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1666199351
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1666199351
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1666199351
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1666199351
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666199351
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1666199351
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1666199351
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1666199351
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1666199351
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1666199351
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666199351
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1666199351
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1666199351
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1666199351
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1666199351
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1666199351
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1666199351
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1666199351
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1666199351
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1666199351
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1666199351
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1666199351
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1666199351
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1666199351
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1666199351
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1666199351
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1666199351
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1666199351
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1666199351
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1666199351
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1666199351
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1666199351
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1666199351
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1666199351
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1666199351
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1666199351
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1666199351
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1666199351
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1666199351
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1666199351
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1666199351
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1666199351
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1666199351
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1666199351
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1666199351
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1666199351
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1666199351
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1666199351
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1666199351
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1666199351
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1666199351
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1666199351
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1666199351
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1666199351
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1666199351
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1666199351
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1666199351
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1666199351
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1666199351
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1666199351
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1666199351
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1666199351
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1666199351
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1666199351
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1666199351
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1666199351
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1666199351
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1666199351
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1666199351
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1666199351
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1666199351
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1666199351
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1666199351
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1666199351
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1666199351
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1666199351
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1666199351
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1666199351
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1666199351
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1666199351
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1666199351
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1666199351
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1666199351
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1666199351
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1666199351
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1666199351
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1666199351
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1666199351
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1666199351
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1666199351
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1666199351
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1666199351
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1666199351
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1666199351
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1666199351
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1666199351
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1666199351
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1666199351
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1666199351
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1666199351
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1666199351
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1666199351
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1666199351
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1666199351
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1666199351
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1666199351
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1666199351
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1666199351
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1666199351
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1666199351
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1666199351
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1666199351
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1666199351
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1666199351
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1666199351
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666199351
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1666199351
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1666199351
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1666199351
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1666199351
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1666199351
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1666199351
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1666199351
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1666199351
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1666199351
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1666199351
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1666199351
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1666199351
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1666199351
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1666199351
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1666199351
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1666199351
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1666199351
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1666199351
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1666199351
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1666199351
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1666199351
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1666199351
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1666199351
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1666199351
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1666199351
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1666199351
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1666199351
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1666199351
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1666199351
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1666199351
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1666199351
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1666199351
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1666199351
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1666199351
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1666199351
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1666199351
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1666199351
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1666199351
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1666199351
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1666199351
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1666199351
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1666199351
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1666199351
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1666199351
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1666199351
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1666199351
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1666199351
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1666199351
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1666199351
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1666199351
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1666199351
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1666199351
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1666199351
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1666199351
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1666199351
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1666199351
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1666199351
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1666199351
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1666199351
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1666199351
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1666199351
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1666199351
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1666199351
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1666199351
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1666199351
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1666199351
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1666199351
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1666199351
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1666199351
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1666199351
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1666199351
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1666199351
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1666199351
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1666199351
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1666199351
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1666199351
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1666199351
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1666199351
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1666199351
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1666199351
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1666199351
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1666199351
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1666199351
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1666199351
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1666199351
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1666199351
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1666199351
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1666199351
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1666199351
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1666199351
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1666199351
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1666199351
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1666199351
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1666199351
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1666199351
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1666199351
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1666199351
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1666199351
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_513
timestamp 1666199351
transform 1 0 48300 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1666199351
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1666199351
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1666199351
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1666199351
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1666199351
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1666199351
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1666199351
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1666199351
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1666199351
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1666199351
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1666199351
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1666199351
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1666199351
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1666199351
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1666199351
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1666199351
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1666199351
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1666199351
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1666199351
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1666199351
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1666199351
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1666199351
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1666199351
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1666199351
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1666199351
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1666199351
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1666199351
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1666199351
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1666199351
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1666199351
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1666199351
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1666199351
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1666199351
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1666199351
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1666199351
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1666199351
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1666199351
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1666199351
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1666199351
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1666199351
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1666199351
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1666199351
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1666199351
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1666199351
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1666199351
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1666199351
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1666199351
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1666199351
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1666199351
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1666199351
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1666199351
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1666199351
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1666199351
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1666199351
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_505
timestamp 1666199351
transform 1 0 47564 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_513
timestamp 1666199351
transform 1 0 48300 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1666199351
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1666199351
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1666199351
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1666199351
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1666199351
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1666199351
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1666199351
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1666199351
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1666199351
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1666199351
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1666199351
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1666199351
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1666199351
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1666199351
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1666199351
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1666199351
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1666199351
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1666199351
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1666199351
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1666199351
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1666199351
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1666199351
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1666199351
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1666199351
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1666199351
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1666199351
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1666199351
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1666199351
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1666199351
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1666199351
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1666199351
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1666199351
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1666199351
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1666199351
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1666199351
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1666199351
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1666199351
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1666199351
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1666199351
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1666199351
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1666199351
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1666199351
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1666199351
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1666199351
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1666199351
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1666199351
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1666199351
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1666199351
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1666199351
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1666199351
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1666199351
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1666199351
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1666199351
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1666199351
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_513
timestamp 1666199351
transform 1 0 48300 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1666199351
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1666199351
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1666199351
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1666199351
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1666199351
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1666199351
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1666199351
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1666199351
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1666199351
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1666199351
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1666199351
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1666199351
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1666199351
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1666199351
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1666199351
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1666199351
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1666199351
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1666199351
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1666199351
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1666199351
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1666199351
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1666199351
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1666199351
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1666199351
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1666199351
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1666199351
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1666199351
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1666199351
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1666199351
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1666199351
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1666199351
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1666199351
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1666199351
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1666199351
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1666199351
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1666199351
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1666199351
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1666199351
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1666199351
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1666199351
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1666199351
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1666199351
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1666199351
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1666199351
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1666199351
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1666199351
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1666199351
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1666199351
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1666199351
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1666199351
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1666199351
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1666199351
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1666199351
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1666199351
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_505
timestamp 1666199351
transform 1 0 47564 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_513
timestamp 1666199351
transform 1 0 48300 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1666199351
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1666199351
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1666199351
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1666199351
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1666199351
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1666199351
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1666199351
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1666199351
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1666199351
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1666199351
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1666199351
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1666199351
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1666199351
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1666199351
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1666199351
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1666199351
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1666199351
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1666199351
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1666199351
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1666199351
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1666199351
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1666199351
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1666199351
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1666199351
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1666199351
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1666199351
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1666199351
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1666199351
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1666199351
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1666199351
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1666199351
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1666199351
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1666199351
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1666199351
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1666199351
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1666199351
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1666199351
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1666199351
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1666199351
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1666199351
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1666199351
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1666199351
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1666199351
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1666199351
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1666199351
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1666199351
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1666199351
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1666199351
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1666199351
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1666199351
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1666199351
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1666199351
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1666199351
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1666199351
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_513
timestamp 1666199351
transform 1 0 48300 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1666199351
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1666199351
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1666199351
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1666199351
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1666199351
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1666199351
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1666199351
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1666199351
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1666199351
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1666199351
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1666199351
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1666199351
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1666199351
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1666199351
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1666199351
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1666199351
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1666199351
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1666199351
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1666199351
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1666199351
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1666199351
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1666199351
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1666199351
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1666199351
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1666199351
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1666199351
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1666199351
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1666199351
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1666199351
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1666199351
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1666199351
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1666199351
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1666199351
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1666199351
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1666199351
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1666199351
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1666199351
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1666199351
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1666199351
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1666199351
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1666199351
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1666199351
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1666199351
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1666199351
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1666199351
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1666199351
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1666199351
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1666199351
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1666199351
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1666199351
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1666199351
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1666199351
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1666199351
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1666199351
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_505
timestamp 1666199351
transform 1 0 47564 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_513
timestamp 1666199351
transform 1 0 48300 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1666199351
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1666199351
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1666199351
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1666199351
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1666199351
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1666199351
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1666199351
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1666199351
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1666199351
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1666199351
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1666199351
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1666199351
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1666199351
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1666199351
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1666199351
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1666199351
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1666199351
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1666199351
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1666199351
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1666199351
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1666199351
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1666199351
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1666199351
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1666199351
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1666199351
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1666199351
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1666199351
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1666199351
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1666199351
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1666199351
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1666199351
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1666199351
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1666199351
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1666199351
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1666199351
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1666199351
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1666199351
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1666199351
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1666199351
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1666199351
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1666199351
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1666199351
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1666199351
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1666199351
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1666199351
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1666199351
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1666199351
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1666199351
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1666199351
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1666199351
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1666199351
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1666199351
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1666199351
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1666199351
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_513
timestamp 1666199351
transform 1 0 48300 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1666199351
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1666199351
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1666199351
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1666199351
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1666199351
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1666199351
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1666199351
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1666199351
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1666199351
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1666199351
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1666199351
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1666199351
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1666199351
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1666199351
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1666199351
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1666199351
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1666199351
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1666199351
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1666199351
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1666199351
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1666199351
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1666199351
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1666199351
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1666199351
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1666199351
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1666199351
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1666199351
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1666199351
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1666199351
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1666199351
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1666199351
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1666199351
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1666199351
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1666199351
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1666199351
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1666199351
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1666199351
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1666199351
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1666199351
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1666199351
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1666199351
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1666199351
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1666199351
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1666199351
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1666199351
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1666199351
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1666199351
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1666199351
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1666199351
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1666199351
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1666199351
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1666199351
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1666199351
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1666199351
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_505
timestamp 1666199351
transform 1 0 47564 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_513
timestamp 1666199351
transform 1 0 48300 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1666199351
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1666199351
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1666199351
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1666199351
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1666199351
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1666199351
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1666199351
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1666199351
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1666199351
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1666199351
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1666199351
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1666199351
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1666199351
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1666199351
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1666199351
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1666199351
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1666199351
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1666199351
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1666199351
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1666199351
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1666199351
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1666199351
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1666199351
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1666199351
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1666199351
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1666199351
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1666199351
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1666199351
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1666199351
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1666199351
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_291
timestamp 1666199351
transform 1 0 27876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_303
timestamp 1666199351
transform 1 0 28980 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1666199351
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1666199351
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1666199351
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1666199351
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1666199351
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1666199351
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1666199351
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1666199351
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1666199351
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1666199351
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1666199351
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1666199351
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1666199351
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1666199351
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1666199351
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1666199351
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1666199351
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1666199351
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1666199351
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1666199351
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1666199351
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1666199351
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_513
timestamp 1666199351
transform 1 0 48300 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1666199351
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1666199351
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1666199351
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1666199351
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1666199351
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1666199351
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1666199351
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1666199351
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1666199351
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1666199351
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1666199351
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1666199351
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1666199351
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1666199351
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1666199351
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1666199351
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1666199351
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1666199351
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1666199351
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1666199351
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1666199351
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1666199351
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1666199351
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1666199351
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1666199351
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_237
timestamp 1666199351
transform 1 0 22908 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_247
timestamp 1666199351
transform 1 0 23828 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_255
timestamp 1666199351
transform 1 0 24564 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_258
timestamp 1666199351
transform 1 0 24840 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_270
timestamp 1666199351
transform 1 0 25944 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_278
timestamp 1666199351
transform 1 0 26680 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_281
timestamp 1666199351
transform 1 0 26956 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_285
timestamp 1666199351
transform 1 0 27324 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_291
timestamp 1666199351
transform 1 0 27876 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_295
timestamp 1666199351
transform 1 0 28244 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_298
timestamp 1666199351
transform 1 0 28520 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_304
timestamp 1666199351
transform 1 0 29072 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_310
timestamp 1666199351
transform 1 0 29624 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_322
timestamp 1666199351
transform 1 0 30728 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_334
timestamp 1666199351
transform 1 0 31832 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1666199351
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1666199351
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1666199351
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1666199351
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1666199351
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1666199351
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1666199351
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1666199351
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1666199351
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1666199351
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1666199351
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1666199351
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1666199351
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1666199351
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1666199351
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1666199351
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1666199351
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1666199351
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1666199351
transform 1 0 47564 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_513
timestamp 1666199351
transform 1 0 48300 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1666199351
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1666199351
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1666199351
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1666199351
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1666199351
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1666199351
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1666199351
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1666199351
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1666199351
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1666199351
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1666199351
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1666199351
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1666199351
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1666199351
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1666199351
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1666199351
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1666199351
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1666199351
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1666199351
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1666199351
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1666199351
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1666199351
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1666199351
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_221
timestamp 1666199351
transform 1 0 21436 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_227
timestamp 1666199351
transform 1 0 21988 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_235
timestamp 1666199351
transform 1 0 22724 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_238
timestamp 1666199351
transform 1 0 23000 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_244
timestamp 1666199351
transform 1 0 23552 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1666199351
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_74_253
timestamp 1666199351
transform 1 0 24380 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_259
timestamp 1666199351
transform 1 0 24932 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_265
timestamp 1666199351
transform 1 0 25484 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_271
timestamp 1666199351
transform 1 0 26036 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_274
timestamp 1666199351
transform 1 0 26312 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_280
timestamp 1666199351
transform 1 0 26864 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_287
timestamp 1666199351
transform 1 0 27508 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_294
timestamp 1666199351
transform 1 0 28152 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1666199351
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1666199351
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_309
timestamp 1666199351
transform 1 0 29532 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_313
timestamp 1666199351
transform 1 0 29900 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_317
timestamp 1666199351
transform 1 0 30268 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_320
timestamp 1666199351
transform 1 0 30544 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_332
timestamp 1666199351
transform 1 0 31648 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_336
timestamp 1666199351
transform 1 0 32016 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_339
timestamp 1666199351
transform 1 0 32292 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_353
timestamp 1666199351
transform 1 0 33580 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_361
timestamp 1666199351
transform 1 0 34316 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1666199351
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1666199351
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1666199351
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1666199351
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1666199351
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1666199351
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1666199351
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1666199351
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1666199351
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1666199351
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1666199351
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1666199351
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1666199351
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1666199351
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1666199351
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_513
timestamp 1666199351
transform 1 0 48300 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1666199351
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1666199351
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1666199351
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1666199351
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1666199351
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1666199351
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1666199351
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1666199351
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1666199351
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1666199351
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1666199351
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1666199351
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1666199351
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1666199351
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1666199351
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1666199351
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1666199351
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1666199351
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1666199351
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1666199351
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1666199351
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1666199351
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_217
timestamp 1666199351
transform 1 0 21068 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_220
timestamp 1666199351
transform 1 0 21344 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_225
timestamp 1666199351
transform 1 0 21804 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_231
timestamp 1666199351
transform 1 0 22356 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_235
timestamp 1666199351
transform 1 0 22724 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_242
timestamp 1666199351
transform 1 0 23368 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_249
timestamp 1666199351
transform 1 0 24012 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_253
timestamp 1666199351
transform 1 0 24380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_259
timestamp 1666199351
transform 1 0 24932 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_269
timestamp 1666199351
transform 1 0 25852 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_275
timestamp 1666199351
transform 1 0 26404 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1666199351
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_281
timestamp 1666199351
transform 1 0 26956 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_289
timestamp 1666199351
transform 1 0 27692 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_296
timestamp 1666199351
transform 1 0 28336 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_303
timestamp 1666199351
transform 1 0 28980 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_310
timestamp 1666199351
transform 1 0 29624 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_317
timestamp 1666199351
transform 1 0 30268 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_323
timestamp 1666199351
transform 1 0 30820 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_327
timestamp 1666199351
transform 1 0 31188 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_331
timestamp 1666199351
transform 1 0 31556 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1666199351
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_337
timestamp 1666199351
transform 1 0 32108 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_342
timestamp 1666199351
transform 1 0 32568 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_349
timestamp 1666199351
transform 1 0 33212 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_356
timestamp 1666199351
transform 1 0 33856 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_363
timestamp 1666199351
transform 1 0 34500 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_370
timestamp 1666199351
transform 1 0 35144 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_376
timestamp 1666199351
transform 1 0 35696 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_388
timestamp 1666199351
transform 1 0 36800 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1666199351
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1666199351
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1666199351
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1666199351
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1666199351
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1666199351
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1666199351
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1666199351
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1666199351
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1666199351
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1666199351
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1666199351
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_505
timestamp 1666199351
transform 1 0 47564 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_513
timestamp 1666199351
transform 1 0 48300 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1666199351
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1666199351
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1666199351
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1666199351
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1666199351
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1666199351
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1666199351
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1666199351
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1666199351
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1666199351
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1666199351
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1666199351
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1666199351
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1666199351
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1666199351
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1666199351
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1666199351
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1666199351
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1666199351
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1666199351
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1666199351
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_197
timestamp 1666199351
transform 1 0 19228 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_205
timestamp 1666199351
transform 1 0 19964 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_211
timestamp 1666199351
transform 1 0 20516 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_215
timestamp 1666199351
transform 1 0 20884 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_218
timestamp 1666199351
transform 1 0 21160 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_225
timestamp 1666199351
transform 1 0 21804 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_232
timestamp 1666199351
transform 1 0 22448 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_238
timestamp 1666199351
transform 1 0 23000 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_242
timestamp 1666199351
transform 1 0 23368 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_250
timestamp 1666199351
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_253
timestamp 1666199351
transform 1 0 24380 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_264
timestamp 1666199351
transform 1 0 25392 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_271
timestamp 1666199351
transform 1 0 26036 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_282
timestamp 1666199351
transform 1 0 27048 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_292
timestamp 1666199351
transform 1 0 27968 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_304
timestamp 1666199351
transform 1 0 29072 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_309
timestamp 1666199351
transform 1 0 29532 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_317
timestamp 1666199351
transform 1 0 30268 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_324
timestamp 1666199351
transform 1 0 30912 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_331
timestamp 1666199351
transform 1 0 31556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_337
timestamp 1666199351
transform 1 0 32108 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_343
timestamp 1666199351
transform 1 0 32660 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_349
timestamp 1666199351
transform 1 0 33212 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_354
timestamp 1666199351
transform 1 0 33672 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_361
timestamp 1666199351
transform 1 0 34316 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_76_365
timestamp 1666199351
transform 1 0 34684 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_371
timestamp 1666199351
transform 1 0 35236 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_377
timestamp 1666199351
transform 1 0 35788 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_384
timestamp 1666199351
transform 1 0 36432 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_390
timestamp 1666199351
transform 1 0 36984 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_402
timestamp 1666199351
transform 1 0 38088 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_414
timestamp 1666199351
transform 1 0 39192 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1666199351
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1666199351
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1666199351
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1666199351
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1666199351
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1666199351
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1666199351
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1666199351
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1666199351
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_513
timestamp 1666199351
transform 1 0 48300 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1666199351
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1666199351
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1666199351
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1666199351
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1666199351
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1666199351
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1666199351
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1666199351
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1666199351
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1666199351
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1666199351
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1666199351
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1666199351
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1666199351
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1666199351
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1666199351
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1666199351
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1666199351
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1666199351
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1666199351
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_193
timestamp 1666199351
transform 1 0 18860 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_201
timestamp 1666199351
transform 1 0 19596 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_204
timestamp 1666199351
transform 1 0 19872 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_210
timestamp 1666199351
transform 1 0 20424 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1666199351
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1666199351
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_225
timestamp 1666199351
transform 1 0 21804 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_229
timestamp 1666199351
transform 1 0 22172 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_236
timestamp 1666199351
transform 1 0 22816 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_247
timestamp 1666199351
transform 1 0 23828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_253
timestamp 1666199351
transform 1 0 24380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_259
timestamp 1666199351
transform 1 0 24932 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_268
timestamp 1666199351
transform 1 0 25760 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_278
timestamp 1666199351
transform 1 0 26680 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_281
timestamp 1666199351
transform 1 0 26956 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_287
timestamp 1666199351
transform 1 0 27508 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_296
timestamp 1666199351
transform 1 0 28336 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_307
timestamp 1666199351
transform 1 0 29348 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_332
timestamp 1666199351
transform 1 0 31648 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_337
timestamp 1666199351
transform 1 0 32108 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_344
timestamp 1666199351
transform 1 0 32752 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_350
timestamp 1666199351
transform 1 0 33304 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_359
timestamp 1666199351
transform 1 0 34132 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_370
timestamp 1666199351
transform 1 0 35144 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_380
timestamp 1666199351
transform 1 0 36064 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_390
timestamp 1666199351
transform 1 0 36984 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_393
timestamp 1666199351
transform 1 0 37260 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_401
timestamp 1666199351
transform 1 0 37996 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_407
timestamp 1666199351
transform 1 0 38548 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_419
timestamp 1666199351
transform 1 0 39652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_431
timestamp 1666199351
transform 1 0 40756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_443
timestamp 1666199351
transform 1 0 41860 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1666199351
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1666199351
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1666199351
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1666199351
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1666199351
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1666199351
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1666199351
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_505
timestamp 1666199351
transform 1 0 47564 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_513
timestamp 1666199351
transform 1 0 48300 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1666199351
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1666199351
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1666199351
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1666199351
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1666199351
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1666199351
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1666199351
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1666199351
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1666199351
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1666199351
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1666199351
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1666199351
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1666199351
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1666199351
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1666199351
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1666199351
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1666199351
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1666199351
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1666199351
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_189
timestamp 1666199351
transform 1 0 18492 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_194
timestamp 1666199351
transform 1 0 18952 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_197
timestamp 1666199351
transform 1 0 19228 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_203
timestamp 1666199351
transform 1 0 19780 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_207
timestamp 1666199351
transform 1 0 20148 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_216
timestamp 1666199351
transform 1 0 20976 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_224
timestamp 1666199351
transform 1 0 21712 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_232
timestamp 1666199351
transform 1 0 22448 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_237
timestamp 1666199351
transform 1 0 22908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_247
timestamp 1666199351
transform 1 0 23828 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1666199351
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_253
timestamp 1666199351
transform 1 0 24380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_262
timestamp 1666199351
transform 1 0 25208 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_268
timestamp 1666199351
transform 1 0 25760 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_275
timestamp 1666199351
transform 1 0 26404 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_279
timestamp 1666199351
transform 1 0 26772 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_286
timestamp 1666199351
transform 1 0 27416 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_296
timestamp 1666199351
transform 1 0 28336 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_304
timestamp 1666199351
transform 1 0 29072 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_309
timestamp 1666199351
transform 1 0 29532 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_316
timestamp 1666199351
transform 1 0 30176 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_324
timestamp 1666199351
transform 1 0 30912 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_334
timestamp 1666199351
transform 1 0 31832 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_78_349
timestamp 1666199351
transform 1 0 33212 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_355
timestamp 1666199351
transform 1 0 33764 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_362
timestamp 1666199351
transform 1 0 34408 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_365
timestamp 1666199351
transform 1 0 34684 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_373
timestamp 1666199351
transform 1 0 35420 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_377
timestamp 1666199351
transform 1 0 35788 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_386
timestamp 1666199351
transform 1 0 36616 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_397
timestamp 1666199351
transform 1 0 37628 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_404
timestamp 1666199351
transform 1 0 38272 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_411
timestamp 1666199351
transform 1 0 38916 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_78_417
timestamp 1666199351
transform 1 0 39468 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_421
timestamp 1666199351
transform 1 0 39836 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_425
timestamp 1666199351
transform 1 0 40204 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_429
timestamp 1666199351
transform 1 0 40572 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_432
timestamp 1666199351
transform 1 0 40848 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_444
timestamp 1666199351
transform 1 0 41952 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_456
timestamp 1666199351
transform 1 0 43056 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_468
timestamp 1666199351
transform 1 0 44160 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1666199351
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1666199351
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1666199351
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_513
timestamp 1666199351
transform 1 0 48300 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1666199351
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1666199351
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1666199351
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1666199351
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1666199351
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1666199351
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1666199351
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1666199351
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1666199351
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1666199351
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1666199351
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1666199351
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1666199351
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1666199351
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1666199351
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1666199351
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1666199351
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1666199351
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1666199351
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_183
timestamp 1666199351
transform 1 0 17940 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_190
timestamp 1666199351
transform 1 0 18584 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_197
timestamp 1666199351
transform 1 0 19228 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_207
timestamp 1666199351
transform 1 0 20148 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_219
timestamp 1666199351
transform 1 0 21252 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1666199351
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_225
timestamp 1666199351
transform 1 0 21804 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_232
timestamp 1666199351
transform 1 0 22448 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_238
timestamp 1666199351
transform 1 0 23000 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_246
timestamp 1666199351
transform 1 0 23736 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_253
timestamp 1666199351
transform 1 0 24380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_262
timestamp 1666199351
transform 1 0 25208 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_274
timestamp 1666199351
transform 1 0 26312 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_79_281
timestamp 1666199351
transform 1 0 26956 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_289
timestamp 1666199351
transform 1 0 27692 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_300
timestamp 1666199351
transform 1 0 28704 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_311
timestamp 1666199351
transform 1 0 29716 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_315
timestamp 1666199351
transform 1 0 30084 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_323
timestamp 1666199351
transform 1 0 30820 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_327
timestamp 1666199351
transform 1 0 31188 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_334
timestamp 1666199351
transform 1 0 31832 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_337
timestamp 1666199351
transform 1 0 32108 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_346
timestamp 1666199351
transform 1 0 32936 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_350
timestamp 1666199351
transform 1 0 33304 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_359
timestamp 1666199351
transform 1 0 34132 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_365
timestamp 1666199351
transform 1 0 34684 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_375
timestamp 1666199351
transform 1 0 35604 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1666199351
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1666199351
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_393
timestamp 1666199351
transform 1 0 37260 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_401
timestamp 1666199351
transform 1 0 37996 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_410
timestamp 1666199351
transform 1 0 38824 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_417
timestamp 1666199351
transform 1 0 39468 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_424
timestamp 1666199351
transform 1 0 40112 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_431
timestamp 1666199351
transform 1 0 40756 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_438
timestamp 1666199351
transform 1 0 41400 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_446
timestamp 1666199351
transform 1 0 42136 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1666199351
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1666199351
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1666199351
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1666199351
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1666199351
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1666199351
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_505
timestamp 1666199351
transform 1 0 47564 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_513
timestamp 1666199351
transform 1 0 48300 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1666199351
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1666199351
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1666199351
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1666199351
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_41
timestamp 1666199351
transform 1 0 4876 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_49
timestamp 1666199351
transform 1 0 5612 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_55
timestamp 1666199351
transform 1 0 6164 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_67
timestamp 1666199351
transform 1 0 7268 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_79
timestamp 1666199351
transform 1 0 8372 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1666199351
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_85
timestamp 1666199351
transform 1 0 8924 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_93
timestamp 1666199351
transform 1 0 9660 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_98
timestamp 1666199351
transform 1 0 10120 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_110
timestamp 1666199351
transform 1 0 11224 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_122
timestamp 1666199351
transform 1 0 12328 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_134
timestamp 1666199351
transform 1 0 13432 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1666199351
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1666199351
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_165
timestamp 1666199351
transform 1 0 16284 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_171
timestamp 1666199351
transform 1 0 16836 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_175
timestamp 1666199351
transform 1 0 17204 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_183
timestamp 1666199351
transform 1 0 17940 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_187
timestamp 1666199351
transform 1 0 18308 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_194
timestamp 1666199351
transform 1 0 18952 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_197
timestamp 1666199351
transform 1 0 19228 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_206
timestamp 1666199351
transform 1 0 20056 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_216
timestamp 1666199351
transform 1 0 20976 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_225
timestamp 1666199351
transform 1 0 21804 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_231
timestamp 1666199351
transform 1 0 22356 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_240
timestamp 1666199351
transform 1 0 23184 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_244
timestamp 1666199351
transform 1 0 23552 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_250
timestamp 1666199351
transform 1 0 24104 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_253
timestamp 1666199351
transform 1 0 24380 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_80_266
timestamp 1666199351
transform 1 0 25576 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_280
timestamp 1666199351
transform 1 0 26864 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_291
timestamp 1666199351
transform 1 0 27876 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1666199351
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1666199351
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_309
timestamp 1666199351
transform 1 0 29532 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_313
timestamp 1666199351
transform 1 0 29900 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_323
timestamp 1666199351
transform 1 0 30820 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_80_338
timestamp 1666199351
transform 1 0 32200 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_353
timestamp 1666199351
transform 1 0 33580 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_362
timestamp 1666199351
transform 1 0 34408 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_365
timestamp 1666199351
transform 1 0 34684 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_369
timestamp 1666199351
transform 1 0 35052 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_380
timestamp 1666199351
transform 1 0 36064 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_387
timestamp 1666199351
transform 1 0 36708 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_398
timestamp 1666199351
transform 1 0 37720 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_409
timestamp 1666199351
transform 1 0 38732 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_416
timestamp 1666199351
transform 1 0 39376 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_421
timestamp 1666199351
transform 1 0 39836 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_426
timestamp 1666199351
transform 1 0 40296 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_433
timestamp 1666199351
transform 1 0 40940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_440
timestamp 1666199351
transform 1 0 41584 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_447
timestamp 1666199351
transform 1 0 42228 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_454
timestamp 1666199351
transform 1 0 42872 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_460
timestamp 1666199351
transform 1 0 43424 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_466
timestamp 1666199351
transform 1 0 43976 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_472
timestamp 1666199351
transform 1 0 44528 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_477
timestamp 1666199351
transform 1 0 44988 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_481
timestamp 1666199351
transform 1 0 45356 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_493
timestamp 1666199351
transform 1 0 46460 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_505
timestamp 1666199351
transform 1 0 47564 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_513
timestamp 1666199351
transform 1 0 48300 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1666199351
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1666199351
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_27
timestamp 1666199351
transform 1 0 3588 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_32
timestamp 1666199351
transform 1 0 4048 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_81_43
timestamp 1666199351
transform 1 0 5060 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1666199351
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_57
timestamp 1666199351
transform 1 0 6348 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_63
timestamp 1666199351
transform 1 0 6900 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_67
timestamp 1666199351
transform 1 0 7268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_79
timestamp 1666199351
transform 1 0 8372 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_87
timestamp 1666199351
transform 1 0 9108 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_91
timestamp 1666199351
transform 1 0 9476 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_99
timestamp 1666199351
transform 1 0 10212 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_103
timestamp 1666199351
transform 1 0 10580 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1666199351
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_113
timestamp 1666199351
transform 1 0 11500 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_118
timestamp 1666199351
transform 1 0 11960 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_81_127
timestamp 1666199351
transform 1 0 12788 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_135
timestamp 1666199351
transform 1 0 13524 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_139
timestamp 1666199351
transform 1 0 13892 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_147
timestamp 1666199351
transform 1 0 14628 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_151
timestamp 1666199351
transform 1 0 14996 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_159
timestamp 1666199351
transform 1 0 15732 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_163
timestamp 1666199351
transform 1 0 16100 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1666199351
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_169
timestamp 1666199351
transform 1 0 16652 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_176
timestamp 1666199351
transform 1 0 17296 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_183
timestamp 1666199351
transform 1 0 17940 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_191
timestamp 1666199351
transform 1 0 18676 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_199
timestamp 1666199351
transform 1 0 19412 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_208
timestamp 1666199351
transform 1 0 20240 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_81_222
timestamp 1666199351
transform 1 0 21528 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_225
timestamp 1666199351
transform 1 0 21804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_236
timestamp 1666199351
transform 1 0 22816 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_243
timestamp 1666199351
transform 1 0 23460 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_256
timestamp 1666199351
transform 1 0 24656 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_265
timestamp 1666199351
transform 1 0 25484 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_277
timestamp 1666199351
transform 1 0 26588 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_281
timestamp 1666199351
transform 1 0 26956 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_289
timestamp 1666199351
transform 1 0 27692 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_299
timestamp 1666199351
transform 1 0 28612 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_311
timestamp 1666199351
transform 1 0 29716 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_325
timestamp 1666199351
transform 1 0 31004 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_334
timestamp 1666199351
transform 1 0 31832 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_337
timestamp 1666199351
transform 1 0 32108 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_349
timestamp 1666199351
transform 1 0 33212 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_365
timestamp 1666199351
transform 1 0 34684 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_372
timestamp 1666199351
transform 1 0 35328 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_376
timestamp 1666199351
transform 1 0 35696 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_387
timestamp 1666199351
transform 1 0 36708 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1666199351
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_393
timestamp 1666199351
transform 1 0 37260 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_401
timestamp 1666199351
transform 1 0 37996 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_409
timestamp 1666199351
transform 1 0 38732 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_416
timestamp 1666199351
transform 1 0 39376 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_423
timestamp 1666199351
transform 1 0 40020 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_431
timestamp 1666199351
transform 1 0 40756 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_442
timestamp 1666199351
transform 1 0 41768 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_81_449
timestamp 1666199351
transform 1 0 42412 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_454
timestamp 1666199351
transform 1 0 42872 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_461
timestamp 1666199351
transform 1 0 43516 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_468
timestamp 1666199351
transform 1 0 44160 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_475
timestamp 1666199351
transform 1 0 44804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_482
timestamp 1666199351
transform 1 0 45448 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_489
timestamp 1666199351
transform 1 0 46092 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_501
timestamp 1666199351
transform 1 0 47196 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_505
timestamp 1666199351
transform 1 0 47564 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_513
timestamp 1666199351
transform 1 0 48300 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1666199351
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1666199351
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1666199351
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_29
timestamp 1666199351
transform 1 0 3772 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_42
timestamp 1666199351
transform 1 0 4968 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_50
timestamp 1666199351
transform 1 0 5704 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_82_57
timestamp 1666199351
transform 1 0 6348 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_68
timestamp 1666199351
transform 1 0 7360 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_75
timestamp 1666199351
transform 1 0 8004 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_82
timestamp 1666199351
transform 1 0 8648 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_85
timestamp 1666199351
transform 1 0 8924 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_91
timestamp 1666199351
transform 1 0 9476 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_96
timestamp 1666199351
transform 1 0 9936 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_108
timestamp 1666199351
transform 1 0 11040 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_113
timestamp 1666199351
transform 1 0 11500 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_120
timestamp 1666199351
transform 1 0 12144 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_132
timestamp 1666199351
transform 1 0 13248 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_141
timestamp 1666199351
transform 1 0 14076 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_147
timestamp 1666199351
transform 1 0 14628 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_151
timestamp 1666199351
transform 1 0 14996 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_156
timestamp 1666199351
transform 1 0 15456 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_82_166
timestamp 1666199351
transform 1 0 16376 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_169
timestamp 1666199351
transform 1 0 16652 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_173
timestamp 1666199351
transform 1 0 17020 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_178
timestamp 1666199351
transform 1 0 17480 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_186
timestamp 1666199351
transform 1 0 18216 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1666199351
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_197
timestamp 1666199351
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_207
timestamp 1666199351
transform 1 0 20148 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_214
timestamp 1666199351
transform 1 0 20792 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_222
timestamp 1666199351
transform 1 0 21528 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_225
timestamp 1666199351
transform 1 0 21804 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_232
timestamp 1666199351
transform 1 0 22448 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_238
timestamp 1666199351
transform 1 0 23000 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1666199351
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1666199351
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_259
timestamp 1666199351
transform 1 0 24932 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_271
timestamp 1666199351
transform 1 0 26036 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_278
timestamp 1666199351
transform 1 0 26680 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_281
timestamp 1666199351
transform 1 0 26956 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_293
timestamp 1666199351
transform 1 0 28060 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_306
timestamp 1666199351
transform 1 0 29256 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_82_309
timestamp 1666199351
transform 1 0 29532 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_82_322
timestamp 1666199351
transform 1 0 30728 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_328
timestamp 1666199351
transform 1 0 31280 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_334
timestamp 1666199351
transform 1 0 31832 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_337
timestamp 1666199351
transform 1 0 32108 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_349
timestamp 1666199351
transform 1 0 33212 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_359
timestamp 1666199351
transform 1 0 34132 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1666199351
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_365
timestamp 1666199351
transform 1 0 34684 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_371
timestamp 1666199351
transform 1 0 35236 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_382
timestamp 1666199351
transform 1 0 36248 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_390
timestamp 1666199351
transform 1 0 36984 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_393
timestamp 1666199351
transform 1 0 37260 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_401
timestamp 1666199351
transform 1 0 37996 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_407
timestamp 1666199351
transform 1 0 38548 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_418
timestamp 1666199351
transform 1 0 39560 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_421
timestamp 1666199351
transform 1 0 39836 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_433
timestamp 1666199351
transform 1 0 40940 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_440
timestamp 1666199351
transform 1 0 41584 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_446
timestamp 1666199351
transform 1 0 42136 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1666199351
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_455
timestamp 1666199351
transform 1 0 42964 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_463
timestamp 1666199351
transform 1 0 43700 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_467
timestamp 1666199351
transform 1 0 44068 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1666199351
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_477
timestamp 1666199351
transform 1 0 44988 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_484
timestamp 1666199351
transform 1 0 45632 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_491
timestamp 1666199351
transform 1 0 46276 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_498
timestamp 1666199351
transform 1 0 46920 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_82_505
timestamp 1666199351
transform 1 0 47564 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_513
timestamp 1666199351
transform 1 0 48300 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666199351
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666199351
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666199351
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666199351
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666199351
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666199351
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666199351
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666199351
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666199351
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666199351
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666199351
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666199351
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666199351
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666199351
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666199351
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666199351
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666199351
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666199351
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666199351
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666199351
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666199351
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666199351
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666199351
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666199351
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666199351
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666199351
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666199351
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666199351
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666199351
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666199351
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666199351
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666199351
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666199351
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666199351
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666199351
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666199351
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666199351
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666199351
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666199351
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666199351
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666199351
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666199351
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666199351
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666199351
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666199351
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666199351
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666199351
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666199351
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666199351
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666199351
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666199351
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666199351
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666199351
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666199351
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666199351
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666199351
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666199351
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666199351
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666199351
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666199351
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666199351
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666199351
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666199351
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666199351
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666199351
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666199351
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666199351
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666199351
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666199351
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666199351
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666199351
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666199351
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666199351
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666199351
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666199351
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666199351
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666199351
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666199351
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666199351
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666199351
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666199351
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666199351
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666199351
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666199351
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666199351
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666199351
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666199351
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666199351
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666199351
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666199351
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666199351
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666199351
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666199351
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666199351
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666199351
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666199351
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666199351
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666199351
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666199351
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666199351
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666199351
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666199351
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666199351
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666199351
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666199351
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666199351
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666199351
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666199351
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666199351
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666199351
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666199351
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666199351
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666199351
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666199351
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666199351
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666199351
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666199351
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666199351
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666199351
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666199351
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666199351
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666199351
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666199351
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666199351
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666199351
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666199351
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666199351
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666199351
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666199351
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666199351
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666199351
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666199351
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666199351
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666199351
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666199351
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666199351
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666199351
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666199351
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666199351
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666199351
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666199351
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666199351
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666199351
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666199351
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666199351
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666199351
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666199351
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666199351
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666199351
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666199351
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666199351
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666199351
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666199351
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666199351
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666199351
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666199351
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666199351
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666199351
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666199351
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666199351
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666199351
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666199351
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666199351
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666199351
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666199351
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666199351
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666199351
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666199351
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666199351
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666199351
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666199351
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666199351
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666199351
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666199351
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666199351
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666199351
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666199351
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666199351
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666199351
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666199351
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666199351
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666199351
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666199351
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666199351
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666199351
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666199351
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666199351
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666199351
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666199351
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666199351
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666199351
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666199351
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666199351
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666199351
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666199351
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666199351
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666199351
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666199351
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666199351
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666199351
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666199351
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666199351
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666199351
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666199351
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666199351
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666199351
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666199351
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666199351
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666199351
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666199351
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666199351
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666199351
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666199351
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666199351
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666199351
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666199351
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666199351
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666199351
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666199351
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666199351
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666199351
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666199351
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666199351
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666199351
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666199351
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666199351
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666199351
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666199351
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666199351
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666199351
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666199351
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666199351
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666199351
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666199351
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666199351
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666199351
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666199351
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666199351
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666199351
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666199351
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666199351
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666199351
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666199351
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666199351
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666199351
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666199351
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666199351
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666199351
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666199351
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666199351
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666199351
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666199351
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666199351
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666199351
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666199351
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666199351
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666199351
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666199351
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666199351
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666199351
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666199351
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666199351
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666199351
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666199351
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666199351
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666199351
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666199351
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666199351
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666199351
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666199351
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666199351
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666199351
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666199351
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666199351
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666199351
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666199351
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666199351
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666199351
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666199351
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666199351
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666199351
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666199351
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666199351
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666199351
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666199351
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666199351
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666199351
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666199351
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666199351
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666199351
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666199351
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666199351
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666199351
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666199351
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666199351
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666199351
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666199351
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666199351
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666199351
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666199351
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666199351
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666199351
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666199351
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666199351
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666199351
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666199351
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666199351
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666199351
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666199351
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666199351
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666199351
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666199351
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666199351
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666199351
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666199351
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666199351
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666199351
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666199351
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666199351
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666199351
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666199351
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666199351
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666199351
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666199351
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666199351
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666199351
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666199351
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666199351
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666199351
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666199351
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666199351
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666199351
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666199351
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666199351
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666199351
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666199351
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666199351
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666199351
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666199351
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666199351
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666199351
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666199351
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666199351
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666199351
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666199351
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666199351
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666199351
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666199351
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666199351
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666199351
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666199351
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666199351
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666199351
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666199351
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666199351
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666199351
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666199351
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666199351
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666199351
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666199351
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666199351
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666199351
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666199351
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666199351
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666199351
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666199351
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666199351
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666199351
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666199351
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666199351
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666199351
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666199351
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666199351
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666199351
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666199351
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666199351
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666199351
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666199351
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666199351
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666199351
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666199351
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666199351
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666199351
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666199351
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666199351
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666199351
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666199351
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666199351
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666199351
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666199351
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666199351
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666199351
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666199351
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666199351
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666199351
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666199351
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666199351
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666199351
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666199351
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666199351
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666199351
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666199351
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666199351
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666199351
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666199351
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666199351
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666199351
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666199351
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666199351
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666199351
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666199351
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666199351
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666199351
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666199351
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666199351
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666199351
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666199351
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666199351
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666199351
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666199351
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666199351
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666199351
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666199351
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666199351
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666199351
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666199351
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666199351
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666199351
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666199351
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666199351
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666199351
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666199351
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666199351
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666199351
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666199351
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666199351
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666199351
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666199351
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666199351
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666199351
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666199351
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666199351
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666199351
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666199351
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666199351
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666199351
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666199351
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666199351
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666199351
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666199351
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666199351
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666199351
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666199351
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666199351
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666199351
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666199351
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666199351
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666199351
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666199351
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666199351
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666199351
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666199351
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666199351
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666199351
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666199351
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666199351
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666199351
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666199351
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666199351
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666199351
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666199351
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666199351
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666199351
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666199351
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666199351
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666199351
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666199351
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666199351
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666199351
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666199351
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666199351
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666199351
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666199351
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666199351
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666199351
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666199351
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666199351
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666199351
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666199351
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666199351
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666199351
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666199351
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666199351
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666199351
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666199351
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666199351
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666199351
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666199351
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666199351
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666199351
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666199351
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666199351
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666199351
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666199351
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666199351
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666199351
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666199351
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666199351
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666199351
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666199351
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666199351
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666199351
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666199351
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666199351
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666199351
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666199351
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666199351
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666199351
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666199351
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666199351
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666199351
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666199351
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666199351
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666199351
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666199351
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666199351
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666199351
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666199351
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666199351
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666199351
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666199351
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666199351
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666199351
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666199351
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666199351
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666199351
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666199351
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666199351
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666199351
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666199351
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666199351
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666199351
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666199351
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666199351
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666199351
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666199351
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666199351
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666199351
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666199351
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666199351
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666199351
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666199351
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666199351
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666199351
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666199351
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666199351
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666199351
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666199351
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666199351
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666199351
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666199351
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666199351
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666199351
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666199351
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666199351
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666199351
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666199351
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666199351
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666199351
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666199351
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666199351
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666199351
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666199351
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666199351
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666199351
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666199351
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666199351
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666199351
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666199351
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666199351
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666199351
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666199351
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666199351
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666199351
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666199351
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666199351
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666199351
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666199351
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666199351
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666199351
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666199351
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666199351
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666199351
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666199351
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666199351
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666199351
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666199351
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666199351
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666199351
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666199351
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666199351
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666199351
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666199351
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666199351
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666199351
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666199351
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666199351
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666199351
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666199351
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666199351
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666199351
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666199351
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666199351
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666199351
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666199351
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666199351
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666199351
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666199351
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666199351
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666199351
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666199351
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666199351
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666199351
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666199351
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666199351
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666199351
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666199351
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666199351
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666199351
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666199351
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666199351
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666199351
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666199351
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666199351
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666199351
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666199351
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666199351
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666199351
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666199351
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666199351
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666199351
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666199351
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666199351
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666199351
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666199351
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666199351
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666199351
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666199351
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666199351
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666199351
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666199351
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666199351
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666199351
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666199351
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666199351
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666199351
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666199351
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666199351
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666199351
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666199351
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666199351
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666199351
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666199351
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666199351
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666199351
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666199351
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666199351
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666199351
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666199351
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666199351
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666199351
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666199351
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666199351
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666199351
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666199351
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666199351
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666199351
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666199351
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666199351
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666199351
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666199351
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666199351
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666199351
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666199351
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666199351
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666199351
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666199351
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666199351
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666199351
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666199351
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666199351
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666199351
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666199351
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666199351
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666199351
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666199351
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666199351
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666199351
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666199351
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666199351
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666199351
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666199351
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666199351
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666199351
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666199351
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666199351
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666199351
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666199351
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666199351
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666199351
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666199351
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666199351
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666199351
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666199351
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666199351
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666199351
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666199351
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666199351
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666199351
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666199351
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666199351
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666199351
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666199351
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666199351
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666199351
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666199351
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666199351
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666199351
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666199351
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666199351
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666199351
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666199351
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666199351
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666199351
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666199351
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666199351
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666199351
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666199351
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666199351
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666199351
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666199351
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666199351
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666199351
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666199351
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666199351
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666199351
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666199351
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666199351
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666199351
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666199351
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666199351
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666199351
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666199351
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666199351
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666199351
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666199351
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666199351
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666199351
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666199351
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666199351
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666199351
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666199351
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666199351
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666199351
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666199351
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666199351
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666199351
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666199351
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666199351
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666199351
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666199351
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666199351
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666199351
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666199351
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666199351
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666199351
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666199351
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666199351
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666199351
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666199351
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666199351
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666199351
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666199351
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666199351
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666199351
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666199351
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666199351
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666199351
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666199351
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666199351
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666199351
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666199351
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666199351
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666199351
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666199351
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666199351
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666199351
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666199351
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666199351
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666199351
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666199351
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666199351
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666199351
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666199351
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666199351
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666199351
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666199351
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666199351
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666199351
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666199351
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666199351
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666199351
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666199351
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666199351
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666199351
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666199351
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666199351
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666199351
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666199351
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666199351
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666199351
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666199351
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666199351
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666199351
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666199351
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666199351
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666199351
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666199351
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666199351
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666199351
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666199351
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666199351
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666199351
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666199351
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666199351
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666199351
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666199351
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666199351
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666199351
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666199351
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666199351
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666199351
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666199351
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666199351
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666199351
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666199351
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666199351
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666199351
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666199351
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666199351
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666199351
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666199351
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666199351
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666199351
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666199351
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666199351
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666199351
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666199351
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666199351
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666199351
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666199351
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666199351
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666199351
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666199351
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666199351
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666199351
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666199351
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666199351
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666199351
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666199351
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666199351
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666199351
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666199351
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666199351
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666199351
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666199351
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666199351
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666199351
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666199351
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666199351
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666199351
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666199351
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666199351
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666199351
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666199351
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666199351
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666199351
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666199351
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666199351
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666199351
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666199351
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666199351
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666199351
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666199351
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666199351
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666199351
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666199351
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666199351
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666199351
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666199351
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666199351
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666199351
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666199351
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666199351
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666199351
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666199351
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666199351
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666199351
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666199351
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666199351
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666199351
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666199351
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666199351
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666199351
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666199351
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666199351
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666199351
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666199351
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666199351
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666199351
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666199351
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666199351
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666199351
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666199351
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666199351
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666199351
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666199351
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666199351
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666199351
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666199351
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _157_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 21344 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _158_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 19596 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _159_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 24840 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _160_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 32568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1666199351
transform -1 0 31924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1666199351
transform -1 0 29992 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1666199351
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1666199351
transform -1 0 32568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1666199351
transform -1 0 28520 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1666199351
transform 1 0 27876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1666199351
transform 1 0 27784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1666199351
transform -1 0 32292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1666199351
transform -1 0 24104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _170_
timestamp 1666199351
transform 1 0 25116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1666199351
transform 1 0 28060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1666199351
transform 1 0 24932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1666199351
transform 1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1666199351
transform -1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1666199351
transform 1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1666199351
transform 1 0 24472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1666199351
transform 1 0 23828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1666199351
transform 1 0 20240 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1666199351
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1666199351
transform -1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _181_
timestamp 1666199351
transform 1 0 21252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1666199351
transform 1 0 17664 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1666199351
transform 1 0 21252 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1666199351
transform 1 0 22908 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1666199351
transform 1 0 22264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1666199351
transform 1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1666199351
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1666199351
transform 1 0 19964 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1666199351
transform 1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1666199351
transform 1 0 17020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1666199351
transform 1 0 16744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1666199351
transform 1 0 18952 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _193_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 30176 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _194_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 29072 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _195_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 28704 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _196_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 25484 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _197_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 30268 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _198_
timestamp 1666199351
transform -1 0 29348 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _199_
timestamp 1666199351
transform -1 0 24932 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _200_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 28336 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _201_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 28336 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _202_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 26864 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _203_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 25852 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _204_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 27692 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _205_
timestamp 1666199351
transform 1 0 26128 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _206_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 24104 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _207_
timestamp 1666199351
transform -1 0 24932 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _208_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 25208 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _209_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 28704 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _210_
timestamp 1666199351
transform 1 0 22540 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _211_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 23092 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _212_
timestamp 1666199351
transform -1 0 23184 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _213_
timestamp 1666199351
transform -1 0 38824 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _214_
timestamp 1666199351
transform 1 0 38088 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _215_
timestamp 1666199351
transform -1 0 37720 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _216_
timestamp 1666199351
transform -1 0 31832 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _217_
timestamp 1666199351
transform 1 0 37444 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _218_
timestamp 1666199351
transform -1 0 37628 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _219_
timestamp 1666199351
transform -1 0 32660 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _220_
timestamp 1666199351
transform -1 0 36984 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _221_
timestamp 1666199351
transform -1 0 36616 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _222_
timestamp 1666199351
transform 1 0 35052 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _223_
timestamp 1666199351
transform 1 0 33856 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _224_
timestamp 1666199351
transform 1 0 35328 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _225_
timestamp 1666199351
transform 1 0 34868 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _226_
timestamp 1666199351
transform -1 0 31832 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _227_
timestamp 1666199351
transform -1 0 32752 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _228_
timestamp 1666199351
transform -1 0 32936 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _229_
timestamp 1666199351
transform 1 0 38364 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _230_
timestamp 1666199351
transform 1 0 30544 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _231_
timestamp 1666199351
transform 1 0 31556 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _232_
timestamp 1666199351
transform -1 0 29256 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _233_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 29716 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _234_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 20976 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _235_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 22172 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1666199351
transform -1 0 28336 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _237_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 25852 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _238_
timestamp 1666199351
transform 1 0 25484 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _239_
timestamp 1666199351
transform 1 0 24932 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1666199351
transform -1 0 36708 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _241_
timestamp 1666199351
transform 1 0 33948 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _242_
timestamp 1666199351
transform 1 0 33580 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _243_
timestamp 1666199351
transform 1 0 32936 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _244_
timestamp 1666199351
transform -1 0 20056 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _245_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 18032 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _246_
timestamp 1666199351
transform 1 0 19780 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1666199351
transform 1 0 19872 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _248_
timestamp 1666199351
transform -1 0 20148 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _249_
timestamp 1666199351
transform 1 0 27416 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _250_
timestamp 1666199351
transform -1 0 27048 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _251_
timestamp 1666199351
transform 1 0 28244 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _252_
timestamp 1666199351
transform 1 0 27232 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _253_
timestamp 1666199351
transform 1 0 26312 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _254_
timestamp 1666199351
transform 1 0 35512 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _255_
timestamp 1666199351
transform 1 0 34500 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _256_
timestamp 1666199351
transform 1 0 37444 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _257_
timestamp 1666199351
transform 1 0 35420 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _258_
timestamp 1666199351
transform 1 0 37444 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _259_
timestamp 1666199351
transform -1 0 22448 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1666199351
transform 1 0 18676 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _261_
timestamp 1666199351
transform 1 0 21344 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1666199351
transform 1 0 21528 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _263_
timestamp 1666199351
transform -1 0 21528 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _264_
timestamp 1666199351
transform 1 0 27140 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _265_
timestamp 1666199351
transform 1 0 24748 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _266_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 24748 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _267_
timestamp 1666199351
transform 1 0 25300 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _268_
timestamp 1666199351
transform -1 0 25852 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _269_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 26312 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _270_
timestamp 1666199351
transform -1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _271_
timestamp 1666199351
transform -1 0 34132 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _272_
timestamp 1666199351
transform 1 0 32568 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _273_
timestamp 1666199351
transform -1 0 34408 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _274_
timestamp 1666199351
transform -1 0 33672 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _275_
timestamp 1666199351
transform 1 0 33396 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _276_
timestamp 1666199351
transform 1 0 20516 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1666199351
transform -1 0 21068 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _278_
timestamp 1666199351
transform 1 0 21988 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _279_
timestamp 1666199351
transform 1 0 22172 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _280_
timestamp 1666199351
transform 1 0 20516 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _281_
timestamp 1666199351
transform 1 0 23736 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _282_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 23828 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _283_
timestamp 1666199351
transform 1 0 23184 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _284_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 23736 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _285_
timestamp 1666199351
transform 1 0 27140 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _286_
timestamp 1666199351
transform 1 0 28060 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _287_
timestamp 1666199351
transform -1 0 23368 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _288_
timestamp 1666199351
transform 1 0 31280 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _289_
timestamp 1666199351
transform -1 0 31832 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _290_
timestamp 1666199351
transform 1 0 30176 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _291_
timestamp 1666199351
transform 1 0 37444 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _292_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 36708 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _293_
timestamp 1666199351
transform 1 0 30268 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _294_
timestamp 1666199351
transform 1 0 30084 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _295_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 24656 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _296_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 23368 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _519__194 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 20516 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _519_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 19872 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _520__195
timestamp 1666199351
transform -1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _520_
timestamp 1666199351
transform 1 0 19596 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _521__196
timestamp 1666199351
transform -1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _521_
timestamp 1666199351
transform 1 0 17296 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _522_
timestamp 1666199351
transform 1 0 17020 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _522__197
timestamp 1666199351
transform 1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _523__198
timestamp 1666199351
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _523_
timestamp 1666199351
transform 1 0 21528 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _524__199
timestamp 1666199351
transform 1 0 18676 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _524_
timestamp 1666199351
transform 1 0 19596 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _525__200
timestamp 1666199351
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _525_
timestamp 1666199351
transform 1 0 19596 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _526_
timestamp 1666199351
transform 1 0 22172 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _526__201
timestamp 1666199351
transform -1 0 22540 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _527__202
timestamp 1666199351
transform -1 0 23184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _527_
timestamp 1666199351
transform 1 0 22080 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _528__203
timestamp 1666199351
transform -1 0 23368 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _528_
timestamp 1666199351
transform 1 0 22172 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _529__204
timestamp 1666199351
transform -1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _529_
timestamp 1666199351
transform 1 0 19596 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _530__205
timestamp 1666199351
transform 1 0 18952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _530_
timestamp 1666199351
transform 1 0 22172 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _531__206
timestamp 1666199351
transform 1 0 19596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _531_
timestamp 1666199351
transform 1 0 22448 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _532_
timestamp 1666199351
transform 1 0 24104 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _532__207
timestamp 1666199351
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _533__208
timestamp 1666199351
transform 1 0 23644 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _533_
timestamp 1666199351
transform 1 0 24288 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _534_
timestamp 1666199351
transform 1 0 24380 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _534__209
timestamp 1666199351
transform 1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _535__210
timestamp 1666199351
transform 1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _535_
timestamp 1666199351
transform 1 0 24748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _536__211
timestamp 1666199351
transform -1 0 26956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _536_
timestamp 1666199351
transform -1 0 26680 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _537__212
timestamp 1666199351
transform -1 0 26680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _537_
timestamp 1666199351
transform 1 0 25484 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _538__213
timestamp 1666199351
transform -1 0 25944 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _538_
timestamp 1666199351
transform 1 0 25576 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _539__214
timestamp 1666199351
transform 1 0 26036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _539_
timestamp 1666199351
transform -1 0 27692 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _540__215
timestamp 1666199351
transform 1 0 28428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _540_
timestamp 1666199351
transform -1 0 29072 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _541__216
timestamp 1666199351
transform -1 0 32568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _541_
timestamp 1666199351
transform -1 0 29072 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _542__217
timestamp 1666199351
transform 1 0 28520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _542_
timestamp 1666199351
transform -1 0 29072 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _543__218
timestamp 1666199351
transform 1 0 28704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _543_
timestamp 1666199351
transform -1 0 29072 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _544__219
timestamp 1666199351
transform -1 0 27876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _544_
timestamp 1666199351
transform 1 0 27508 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _545__220
timestamp 1666199351
transform 1 0 31004 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _545_
timestamp 1666199351
transform -1 0 31648 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _546__221
timestamp 1666199351
transform -1 0 33212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _546_
timestamp 1666199351
transform -1 0 31372 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _547_
timestamp 1666199351
transform 1 0 29440 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _547__222
timestamp 1666199351
transform -1 0 29992 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _548__223
timestamp 1666199351
transform 1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _548_
timestamp 1666199351
transform -1 0 31372 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _549__224
timestamp 1666199351
transform -1 0 32936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _549_
timestamp 1666199351
transform -1 0 31648 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _550_
timestamp 1666199351
transform -1 0 31648 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _550__225
timestamp 1666199351
transform 1 0 30636 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 4048 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666199351
transform -1 0 22816 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666199351
transform -1 0 24380 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1666199351
transform 1 0 27140 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1666199351
transform 1 0 27876 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 28704 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1666199351
transform 1 0 29808 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1666199351
transform 1 0 32292 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1666199351
transform 1 0 32292 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1666199351
transform -1 0 33856 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1666199351
transform -1 0 35144 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1666199351
transform -1 0 36248 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1666199351
transform 1 0 37996 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1666199351
transform -1 0 36984 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1666199351
transform 1 0 38640 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1666199351
transform 1 0 40020 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1666199351
transform 1 0 40848 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input18 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 42964 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1666199351
transform -1 0 43700 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1666199351
transform -1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1666199351
transform -1 0 45632 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  macro_golden_37
timestamp 1666199351
transform -1 0 42228 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_38
timestamp 1666199351
transform -1 0 42872 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_39
timestamp 1666199351
transform -1 0 44160 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_40
timestamp 1666199351
transform -1 0 45448 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_41
timestamp 1666199351
transform -1 0 46092 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_42
timestamp 1666199351
transform 1 0 5796 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_43
timestamp 1666199351
transform 1 0 7084 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_44
timestamp 1666199351
transform -1 0 8648 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_45
timestamp 1666199351
transform -1 0 26036 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_46
timestamp 1666199351
transform -1 0 26680 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_47
timestamp 1666199351
transform -1 0 27508 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_48
timestamp 1666199351
transform -1 0 28796 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_49
timestamp 1666199351
transform -1 0 30268 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_50
timestamp 1666199351
transform -1 0 31556 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_51
timestamp 1666199351
transform -1 0 32568 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_52
timestamp 1666199351
transform -1 0 34316 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_53
timestamp 1666199351
transform -1 0 39376 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_54
timestamp 1666199351
transform -1 0 40020 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_55
timestamp 1666199351
transform -1 0 41584 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_56
timestamp 1666199351
transform -1 0 38916 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_57
timestamp 1666199351
transform -1 0 40112 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_58
timestamp 1666199351
transform -1 0 40756 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_59
timestamp 1666199351
transform -1 0 41400 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_60
timestamp 1666199351
transform -1 0 42872 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_61
timestamp 1666199351
transform -1 0 43516 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_62
timestamp 1666199351
transform -1 0 44804 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_63
timestamp 1666199351
transform -1 0 46276 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_64
timestamp 1666199351
transform -1 0 46920 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_65
timestamp 1666199351
transform -1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_66
timestamp 1666199351
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_67
timestamp 1666199351
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_68
timestamp 1666199351
transform -1 0 13432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_69
timestamp 1666199351
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_70
timestamp 1666199351
transform 1 0 12880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_71
timestamp 1666199351
transform -1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_72
timestamp 1666199351
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_73
timestamp 1666199351
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_74
timestamp 1666199351
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_75
timestamp 1666199351
transform -1 0 15364 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_76
timestamp 1666199351
transform 1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_77
timestamp 1666199351
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_78
timestamp 1666199351
transform -1 0 16192 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_79
timestamp 1666199351
transform 1 0 13524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_80
timestamp 1666199351
transform 1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_81
timestamp 1666199351
transform 1 0 14168 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_82
timestamp 1666199351
transform -1 0 17296 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_83
timestamp 1666199351
transform 1 0 15456 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_84
timestamp 1666199351
transform 1 0 16744 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_85
timestamp 1666199351
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_86
timestamp 1666199351
transform 1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_87
timestamp 1666199351
transform 1 0 17664 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_88
timestamp 1666199351
transform -1 0 18952 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_89
timestamp 1666199351
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_90
timestamp 1666199351
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_91
timestamp 1666199351
transform -1 0 19780 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_92
timestamp 1666199351
transform 1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_93
timestamp 1666199351
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_94
timestamp 1666199351
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_95
timestamp 1666199351
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_96
timestamp 1666199351
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_97
timestamp 1666199351
transform -1 0 33856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_98
timestamp 1666199351
transform -1 0 33856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_99
timestamp 1666199351
transform -1 0 35144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_100
timestamp 1666199351
transform -1 0 33580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_101
timestamp 1666199351
transform -1 0 34500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_102
timestamp 1666199351
transform -1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_103
timestamp 1666199351
transform -1 0 32568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_104
timestamp 1666199351
transform -1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_105
timestamp 1666199351
transform -1 0 34224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_106
timestamp 1666199351
transform -1 0 35144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_107
timestamp 1666199351
transform -1 0 33856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_108
timestamp 1666199351
transform -1 0 35788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_109
timestamp 1666199351
transform -1 0 35144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_110
timestamp 1666199351
transform -1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_111
timestamp 1666199351
transform -1 0 34500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_112
timestamp 1666199351
transform -1 0 35144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_113
timestamp 1666199351
transform -1 0 36432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_114
timestamp 1666199351
transform -1 0 35788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_115
timestamp 1666199351
transform -1 0 37720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_116
timestamp 1666199351
transform -1 0 35788 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_117
timestamp 1666199351
transform -1 0 36432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_118
timestamp 1666199351
transform -1 0 37720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_119
timestamp 1666199351
transform -1 0 37076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_120
timestamp 1666199351
transform -1 0 38364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_121
timestamp 1666199351
transform -1 0 37720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_122
timestamp 1666199351
transform -1 0 38364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_123
timestamp 1666199351
transform -1 0 39008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_124
timestamp 1666199351
transform -1 0 38364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_125
timestamp 1666199351
transform -1 0 39008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_126
timestamp 1666199351
transform -1 0 39008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_127
timestamp 1666199351
transform -1 0 40296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_128
timestamp 1666199351
transform -1 0 39652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_129
timestamp 1666199351
transform -1 0 40296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_130
timestamp 1666199351
transform -1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_131
timestamp 1666199351
transform -1 0 40296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_132
timestamp 1666199351
transform -1 0 41584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_133
timestamp 1666199351
transform -1 0 40940 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_134
timestamp 1666199351
transform -1 0 40940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_135
timestamp 1666199351
transform -1 0 41584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_136
timestamp 1666199351
transform -1 0 41584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_137
timestamp 1666199351
transform -1 0 42872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_138
timestamp 1666199351
transform -1 0 42228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_139
timestamp 1666199351
transform -1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_140
timestamp 1666199351
transform -1 0 42872 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_141
timestamp 1666199351
transform -1 0 44160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_142
timestamp 1666199351
transform -1 0 43516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_143
timestamp 1666199351
transform -1 0 42964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_144
timestamp 1666199351
transform -1 0 43608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_145
timestamp 1666199351
transform -1 0 44160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_146
timestamp 1666199351
transform -1 0 45448 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_147
timestamp 1666199351
transform -1 0 44804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_148
timestamp 1666199351
transform -1 0 46092 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_149
timestamp 1666199351
transform -1 0 45448 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_150
timestamp 1666199351
transform -1 0 45448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_151
timestamp 1666199351
transform -1 0 46736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_152
timestamp 1666199351
transform -1 0 46092 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_153
timestamp 1666199351
transform -1 0 46092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_154
timestamp 1666199351
transform -1 0 46736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_155
timestamp 1666199351
transform -1 0 48024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_156
timestamp 1666199351
transform -1 0 46736 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_157
timestamp 1666199351
transform -1 0 47380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_158
timestamp 1666199351
transform -1 0 48024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_159
timestamp 1666199351
transform -1 0 48024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_160
timestamp 1666199351
transform -1 0 48024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_161
timestamp 1666199351
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_162
timestamp 1666199351
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_163
timestamp 1666199351
transform 1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_164
timestamp 1666199351
transform 1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_165
timestamp 1666199351
transform -1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_166
timestamp 1666199351
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_167
timestamp 1666199351
transform -1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_168
timestamp 1666199351
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_169
timestamp 1666199351
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_170
timestamp 1666199351
transform -1 0 6072 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_171
timestamp 1666199351
transform 1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_172
timestamp 1666199351
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_173
timestamp 1666199351
transform -1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_174
timestamp 1666199351
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_175
timestamp 1666199351
transform 1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_176
timestamp 1666199351
transform -1 0 7728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_177
timestamp 1666199351
transform 1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_178
timestamp 1666199351
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_179
timestamp 1666199351
transform -1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_180
timestamp 1666199351
transform 1 0 7728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_181
timestamp 1666199351
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_182
timestamp 1666199351
transform -1 0 9384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_183
timestamp 1666199351
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_184
timestamp 1666199351
transform 1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_185
timestamp 1666199351
transform -1 0 10212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_186
timestamp 1666199351
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_187
timestamp 1666199351
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_188
timestamp 1666199351
transform -1 0 11040 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_189
timestamp 1666199351
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_190
timestamp 1666199351
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_191
timestamp 1666199351
transform -1 0 11868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_192
timestamp 1666199351
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_193
timestamp 1666199351
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_226
timestamp 1666199351
transform -1 0 5060 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_227
timestamp 1666199351
transform -1 0 6164 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_228
timestamp 1666199351
transform -1 0 7268 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_229
timestamp 1666199351
transform 1 0 7728 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_230
timestamp 1666199351
transform -1 0 9476 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_231
timestamp 1666199351
transform -1 0 10580 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_232
timestamp 1666199351
transform -1 0 11960 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_233
timestamp 1666199351
transform -1 0 12788 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_234
timestamp 1666199351
transform -1 0 13892 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_235
timestamp 1666199351
transform -1 0 14996 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_236
timestamp 1666199351
transform -1 0 16100 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_237
timestamp 1666199351
transform -1 0 17204 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_238
timestamp 1666199351
transform 1 0 17020 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_239
timestamp 1666199351
transform 1 0 18308 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_240
timestamp 1666199351
transform 1 0 18952 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_241
timestamp 1666199351
transform 1 0 17664 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_242
timestamp 1666199351
transform -1 0 22724 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_243
timestamp 1666199351
transform 1 0 23092 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_244
timestamp 1666199351
transform -1 0 24932 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_245
timestamp 1666199351
transform 1 0 23184 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_246
timestamp 1666199351
transform 1 0 20516 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_247
timestamp 1666199351
transform -1 0 28980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_248
timestamp 1666199351
transform -1 0 29624 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_249
timestamp 1666199351
transform -1 0 35328 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_250
timestamp 1666199351
transform -1 0 31556 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_251
timestamp 1666199351
transform -1 0 33212 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_252
timestamp 1666199351
transform -1 0 34500 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_253
timestamp 1666199351
transform -1 0 39376 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_254
timestamp 1666199351
transform -1 0 36432 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_255
timestamp 1666199351
transform -1 0 39468 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_256
timestamp 1666199351
transform -1 0 40296 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_257
timestamp 1666199351
transform -1 0 40940 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_golden_258
timestamp 1666199351
transform -1 0 41584 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1666199351
transform -1 0 5704 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1666199351
transform -1 0 16376 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1666199351
transform -1 0 17480 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1666199351
transform -1 0 18676 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1666199351
transform -1 0 18216 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1666199351
transform -1 0 19412 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1666199351
transform -1 0 18952 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1666199351
transform 1 0 21160 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1666199351
transform 1 0 24564 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1666199351
transform -1 0 9936 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1666199351
transform -1 0 11040 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1666199351
transform -1 0 12144 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1666199351
transform -1 0 13248 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1666199351
transform -1 0 14628 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1666199351
transform -1 0 15456 0 1 46784
box -38 -48 406 592
<< labels >>
flabel metal2 s 3974 49200 4030 50000 0 FreeSans 224 90 0 0 io_active
port 0 nsew signal input
flabel metal2 s 4342 49200 4398 50000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 15382 49200 15438 50000 0 FreeSans 224 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s 16486 49200 16542 50000 0 FreeSans 224 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal2 s 17590 49200 17646 50000 0 FreeSans 224 90 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 18694 49200 18750 50000 0 FreeSans 224 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 19798 49200 19854 50000 0 FreeSans 224 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal2 s 20902 49200 20958 50000 0 FreeSans 224 90 0 0 io_in[15]
port 7 nsew signal input
flabel metal2 s 22006 49200 22062 50000 0 FreeSans 224 90 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 23110 49200 23166 50000 0 FreeSans 224 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 24214 49200 24270 50000 0 FreeSans 224 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 25318 49200 25374 50000 0 FreeSans 224 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal2 s 5446 49200 5502 50000 0 FreeSans 224 90 0 0 io_in[1]
port 12 nsew signal input
flabel metal2 s 26422 49200 26478 50000 0 FreeSans 224 90 0 0 io_in[20]
port 13 nsew signal input
flabel metal2 s 27526 49200 27582 50000 0 FreeSans 224 90 0 0 io_in[21]
port 14 nsew signal input
flabel metal2 s 28630 49200 28686 50000 0 FreeSans 224 90 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 29734 49200 29790 50000 0 FreeSans 224 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 30838 49200 30894 50000 0 FreeSans 224 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 31942 49200 31998 50000 0 FreeSans 224 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 33046 49200 33102 50000 0 FreeSans 224 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal2 s 34150 49200 34206 50000 0 FreeSans 224 90 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 35254 49200 35310 50000 0 FreeSans 224 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 36358 49200 36414 50000 0 FreeSans 224 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 6550 49200 6606 50000 0 FreeSans 224 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal2 s 37462 49200 37518 50000 0 FreeSans 224 90 0 0 io_in[30]
port 24 nsew signal input
flabel metal2 s 38566 49200 38622 50000 0 FreeSans 224 90 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 39670 49200 39726 50000 0 FreeSans 224 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal2 s 40774 49200 40830 50000 0 FreeSans 224 90 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 41878 49200 41934 50000 0 FreeSans 224 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 42982 49200 43038 50000 0 FreeSans 224 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal2 s 44086 49200 44142 50000 0 FreeSans 224 90 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 45190 49200 45246 50000 0 FreeSans 224 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 7654 49200 7710 50000 0 FreeSans 224 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal2 s 8758 49200 8814 50000 0 FreeSans 224 90 0 0 io_in[4]
port 33 nsew signal input
flabel metal2 s 9862 49200 9918 50000 0 FreeSans 224 90 0 0 io_in[5]
port 34 nsew signal input
flabel metal2 s 10966 49200 11022 50000 0 FreeSans 224 90 0 0 io_in[6]
port 35 nsew signal input
flabel metal2 s 12070 49200 12126 50000 0 FreeSans 224 90 0 0 io_in[7]
port 36 nsew signal input
flabel metal2 s 13174 49200 13230 50000 0 FreeSans 224 90 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 14278 49200 14334 50000 0 FreeSans 224 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 4710 49200 4766 50000 0 FreeSans 224 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal2 s 15750 49200 15806 50000 0 FreeSans 224 90 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal2 s 16854 49200 16910 50000 0 FreeSans 224 90 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal2 s 17958 49200 18014 50000 0 FreeSans 224 90 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal2 s 19062 49200 19118 50000 0 FreeSans 224 90 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal2 s 20166 49200 20222 50000 0 FreeSans 224 90 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 21270 49200 21326 50000 0 FreeSans 224 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal2 s 22374 49200 22430 50000 0 FreeSans 224 90 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 23478 49200 23534 50000 0 FreeSans 224 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 24582 49200 24638 50000 0 FreeSans 224 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 25686 49200 25742 50000 0 FreeSans 224 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal2 s 5814 49200 5870 50000 0 FreeSans 224 90 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal2 s 26790 49200 26846 50000 0 FreeSans 224 90 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal2 s 27894 49200 27950 50000 0 FreeSans 224 90 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 28998 49200 29054 50000 0 FreeSans 224 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 30102 49200 30158 50000 0 FreeSans 224 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 31206 49200 31262 50000 0 FreeSans 224 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal2 s 32310 49200 32366 50000 0 FreeSans 224 90 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal2 s 33414 49200 33470 50000 0 FreeSans 224 90 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 34518 49200 34574 50000 0 FreeSans 224 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal2 s 35622 49200 35678 50000 0 FreeSans 224 90 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal2 s 36726 49200 36782 50000 0 FreeSans 224 90 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 6918 49200 6974 50000 0 FreeSans 224 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal2 s 37830 49200 37886 50000 0 FreeSans 224 90 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal2 s 38934 49200 38990 50000 0 FreeSans 224 90 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal2 s 40038 49200 40094 50000 0 FreeSans 224 90 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal2 s 41142 49200 41198 50000 0 FreeSans 224 90 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal2 s 42246 49200 42302 50000 0 FreeSans 224 90 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal2 s 43350 49200 43406 50000 0 FreeSans 224 90 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal2 s 44454 49200 44510 50000 0 FreeSans 224 90 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal2 s 45558 49200 45614 50000 0 FreeSans 224 90 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 8022 49200 8078 50000 0 FreeSans 224 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal2 s 9126 49200 9182 50000 0 FreeSans 224 90 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal2 s 10230 49200 10286 50000 0 FreeSans 224 90 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal2 s 11334 49200 11390 50000 0 FreeSans 224 90 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 12438 49200 12494 50000 0 FreeSans 224 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 13542 49200 13598 50000 0 FreeSans 224 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 14646 49200 14702 50000 0 FreeSans 224 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal2 s 5078 49200 5134 50000 0 FreeSans 224 90 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal2 s 16118 49200 16174 50000 0 FreeSans 224 90 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal2 s 17222 49200 17278 50000 0 FreeSans 224 90 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal2 s 18326 49200 18382 50000 0 FreeSans 224 90 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal2 s 19430 49200 19486 50000 0 FreeSans 224 90 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal2 s 20534 49200 20590 50000 0 FreeSans 224 90 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal2 s 21638 49200 21694 50000 0 FreeSans 224 90 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal2 s 22742 49200 22798 50000 0 FreeSans 224 90 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 23846 49200 23902 50000 0 FreeSans 224 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal2 s 24950 49200 25006 50000 0 FreeSans 224 90 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal2 s 26054 49200 26110 50000 0 FreeSans 224 90 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 6182 49200 6238 50000 0 FreeSans 224 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 27158 49200 27214 50000 0 FreeSans 224 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal2 s 28262 49200 28318 50000 0 FreeSans 224 90 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 29366 49200 29422 50000 0 FreeSans 224 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal2 s 30470 49200 30526 50000 0 FreeSans 224 90 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 31574 49200 31630 50000 0 FreeSans 224 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 32678 49200 32734 50000 0 FreeSans 224 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal2 s 33782 49200 33838 50000 0 FreeSans 224 90 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 34886 49200 34942 50000 0 FreeSans 224 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 35990 49200 36046 50000 0 FreeSans 224 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal2 s 37094 49200 37150 50000 0 FreeSans 224 90 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 7286 49200 7342 50000 0 FreeSans 224 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal2 s 38198 49200 38254 50000 0 FreeSans 224 90 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal2 s 39302 49200 39358 50000 0 FreeSans 224 90 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal2 s 40406 49200 40462 50000 0 FreeSans 224 90 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal2 s 41510 49200 41566 50000 0 FreeSans 224 90 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal2 s 42614 49200 42670 50000 0 FreeSans 224 90 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal2 s 43718 49200 43774 50000 0 FreeSans 224 90 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 44822 49200 44878 50000 0 FreeSans 224 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal2 s 45926 49200 45982 50000 0 FreeSans 224 90 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal2 s 8390 49200 8446 50000 0 FreeSans 224 90 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal2 s 9494 49200 9550 50000 0 FreeSans 224 90 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 10598 49200 10654 50000 0 FreeSans 224 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 11702 49200 11758 50000 0 FreeSans 224 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal2 s 12806 49200 12862 50000 0 FreeSans 224 90 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 13910 49200 13966 50000 0 FreeSans 224 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal2 s 15014 49200 15070 50000 0 FreeSans 224 90 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 115 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 116 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 117 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 118 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 119 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 120 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 121 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 122 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 123 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 124 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 125 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 126 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 127 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 128 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 129 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 130 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 131 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 132 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 133 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 134 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 135 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 136 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 137 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 138 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 139 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 140 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 141 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 142 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 143 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 144 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 145 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 146 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 147 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 148 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 149 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 150 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 151 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 152 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 153 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 154 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 155 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 156 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 157 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 158 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 159 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 160 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 161 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 162 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 163 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 164 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 165 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 166 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 167 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 168 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 169 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 170 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 171 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 172 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 173 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 174 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 175 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 176 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 177 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 178 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 179 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 180 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 181 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 182 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 183 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 184 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 185 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 186 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 187 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 188 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 189 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 190 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 191 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 192 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 193 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 194 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 195 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 196 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 197 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 198 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 199 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 200 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 201 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 202 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 203 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 204 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 205 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 206 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 207 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 208 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 209 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 210 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 211 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 212 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 213 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 214 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 215 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 216 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 217 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 218 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 219 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 220 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 221 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 222 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 223 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 224 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 225 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 226 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 227 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 228 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 229 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 230 nsew signal input
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 231 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 232 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 233 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 234 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 235 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 236 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 237 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 238 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 239 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 240 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 241 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 242 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 243 nsew signal tristate
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 244 nsew signal tristate
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 245 nsew signal tristate
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 246 nsew signal tristate
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 247 nsew signal tristate
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 248 nsew signal tristate
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 249 nsew signal tristate
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 250 nsew signal tristate
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 251 nsew signal tristate
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 252 nsew signal tristate
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 253 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 254 nsew signal tristate
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 255 nsew signal tristate
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 256 nsew signal tristate
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 257 nsew signal tristate
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 258 nsew signal tristate
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 259 nsew signal tristate
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 260 nsew signal tristate
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 261 nsew signal tristate
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 262 nsew signal tristate
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 263 nsew signal tristate
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 264 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 265 nsew signal tristate
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 266 nsew signal tristate
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 267 nsew signal tristate
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 268 nsew signal tristate
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 269 nsew signal tristate
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 270 nsew signal tristate
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 271 nsew signal tristate
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 272 nsew signal tristate
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 273 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 274 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 275 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 276 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 277 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 278 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 279 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 280 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 281 nsew signal tristate
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 282 nsew signal tristate
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 283 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 284 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 285 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 286 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 287 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 288 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 289 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 290 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 291 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 292 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 293 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 294 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 295 nsew signal tristate
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 296 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 297 nsew signal tristate
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 298 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 299 nsew signal tristate
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 300 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 301 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 302 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 303 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 304 nsew signal tristate
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 305 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 306 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 307 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 308 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 309 nsew signal tristate
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 310 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 311 nsew signal tristate
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 312 nsew signal tristate
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 313 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 314 nsew signal tristate
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 315 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 316 nsew signal tristate
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 317 nsew signal tristate
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 318 nsew signal tristate
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 319 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 320 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 321 nsew signal tristate
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 322 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 323 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 324 nsew signal tristate
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 325 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 326 nsew signal tristate
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 327 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 328 nsew signal tristate
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 329 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 330 nsew signal tristate
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 331 nsew signal tristate
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 332 nsew signal tristate
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 333 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 334 nsew signal tristate
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 335 nsew signal tristate
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 336 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 337 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 338 nsew signal tristate
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 339 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 340 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 341 nsew signal tristate
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 342 nsew signal tristate
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 343 nsew signal tristate
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 344 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 345 nsew signal tristate
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 346 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 347 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 348 nsew signal tristate
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 349 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 350 nsew signal tristate
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 351 nsew signal tristate
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 352 nsew signal tristate
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 353 nsew signal tristate
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 354 nsew signal tristate
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 355 nsew signal tristate
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 356 nsew signal tristate
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 357 nsew signal tristate
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 358 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 359 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 360 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 361 nsew signal tristate
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 362 nsew signal tristate
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 363 nsew signal tristate
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 364 nsew signal tristate
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 365 nsew signal tristate
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 366 nsew signal tristate
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 367 nsew signal tristate
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 368 nsew signal tristate
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 369 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 370 nsew signal tristate
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 371 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 372 nsew signal input
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 373 nsew signal input
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 374 nsew signal input
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 375 nsew signal input
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 376 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 377 nsew signal input
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 378 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 379 nsew signal input
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 380 nsew signal input
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 381 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 382 nsew signal input
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 383 nsew signal input
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 384 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 385 nsew signal input
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 386 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 387 nsew signal input
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 388 nsew signal input
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 389 nsew signal input
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 390 nsew signal input
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 391 nsew signal input
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 392 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 393 nsew signal input
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 394 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 395 nsew signal input
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 396 nsew signal input
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 397 nsew signal input
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 398 nsew signal input
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 399 nsew signal input
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 400 nsew signal input
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 401 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 402 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 403 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 404 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 405 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 406 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 407 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 408 nsew signal input
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 409 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 410 nsew signal input
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 411 nsew signal input
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 412 nsew signal input
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 413 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 414 nsew signal input
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 415 nsew signal input
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 416 nsew signal input
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 417 nsew signal input
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 418 nsew signal input
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 419 nsew signal input
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 420 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 421 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 422 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 423 nsew signal input
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 424 nsew signal input
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 425 nsew signal input
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 426 nsew signal input
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 427 nsew signal input
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 428 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 429 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 430 nsew signal input
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 431 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 432 nsew signal input
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 433 nsew signal input
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 434 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 435 nsew signal input
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 436 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 437 nsew signal input
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 438 nsew signal input
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 439 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 440 nsew signal input
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 441 nsew signal input
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 442 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 443 nsew signal input
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 444 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 445 nsew signal input
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 446 nsew signal input
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 447 nsew signal input
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 448 nsew signal input
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 449 nsew signal input
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 450 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 451 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 452 nsew signal input
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 453 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 454 nsew signal input
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 455 nsew signal input
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 456 nsew signal input
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 457 nsew signal input
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 458 nsew signal input
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 459 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 460 nsew signal input
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 461 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 462 nsew signal input
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 463 nsew signal input
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 464 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 465 nsew signal input
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 466 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 467 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 468 nsew signal input
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 469 nsew signal input
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 470 nsew signal input
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 471 nsew signal input
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 472 nsew signal input
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 473 nsew signal input
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 474 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 475 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 476 nsew signal input
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 477 nsew signal input
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 478 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 479 nsew signal input
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 480 nsew signal input
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 481 nsew signal input
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 482 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 483 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 484 nsew signal input
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 485 nsew signal input
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 486 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 487 nsew signal input
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 488 nsew signal input
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 489 nsew signal input
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 490 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 491 nsew signal input
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 492 nsew signal input
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 493 nsew signal input
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 494 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 495 nsew signal input
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 496 nsew signal input
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 497 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 498 nsew signal input
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 34928 2128 35248 47376 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 19568 2128 19888 47376 0 FreeSans 1920 90 0 0 vssd1
port 500 nsew ground bidirectional
flabel metal2 s 2410 0 2466 800 0 FreeSans 224 90 0 0 wb_clk_i
port 501 nsew signal input
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 wb_rst_i
port 502 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 503 nsew signal tristate
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 504 nsew signal input
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 505 nsew signal input
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 506 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 507 nsew signal input
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 508 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 509 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 510 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 511 nsew signal input
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 512 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 513 nsew signal input
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 514 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 515 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 516 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 517 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 518 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 519 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 520 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 521 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 522 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 523 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 524 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 525 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 526 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 527 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 528 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 529 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 530 nsew signal input
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 531 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 532 nsew signal input
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 533 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 534 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 535 nsew signal input
flabel metal2 s 2686 0 2742 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 536 nsew signal input
flabel metal2 s 3054 0 3110 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 537 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 538 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 539 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 540 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 541 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 542 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 543 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 544 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 545 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 546 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 547 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 548 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 549 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 550 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 551 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 552 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 553 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 554 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 555 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 556 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 557 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 558 nsew signal input
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 559 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 560 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 561 nsew signal input
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 562 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 563 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 564 nsew signal input
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 565 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 566 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 567 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 568 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 569 nsew signal tristate
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 570 nsew signal tristate
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 571 nsew signal tristate
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 572 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 573 nsew signal tristate
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 574 nsew signal tristate
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 575 nsew signal tristate
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 576 nsew signal tristate
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 577 nsew signal tristate
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 578 nsew signal tristate
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 579 nsew signal tristate
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 580 nsew signal tristate
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 581 nsew signal tristate
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 582 nsew signal tristate
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 583 nsew signal tristate
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 584 nsew signal tristate
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 585 nsew signal tristate
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 586 nsew signal tristate
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 587 nsew signal tristate
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 588 nsew signal tristate
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 589 nsew signal tristate
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 590 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 591 nsew signal tristate
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 592 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 593 nsew signal tristate
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 594 nsew signal tristate
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 595 nsew signal tristate
flabel metal2 s 4894 0 4950 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 596 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 597 nsew signal tristate
flabel metal2 s 5446 0 5502 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 598 nsew signal tristate
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 599 nsew signal tristate
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 600 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 601 nsew signal input
flabel metal2 s 3606 0 3662 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 602 nsew signal input
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 603 nsew signal input
flabel metal2 s 4342 0 4398 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 604 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 605 nsew signal input
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 wbs_we_i
port 606 nsew signal input
rlabel metal1 24978 47328 24978 47328 0 vccd1
rlabel metal1 24978 46784 24978 46784 0 vssd1
rlabel metal1 29900 44710 29900 44710 0 _000_
rlabel metal1 28842 45390 28842 45390 0 _001_
rlabel metal1 25622 46546 25622 46546 0 _002_
rlabel metal1 23598 45458 23598 45458 0 _003_
rlabel metal1 29716 43962 29716 43962 0 _004_
rlabel metal1 25116 43826 25116 43826 0 _005_
rlabel metal1 24702 43418 24702 43418 0 _006_
rlabel metal1 27554 44710 27554 44710 0 _007_
rlabel metal1 27600 44166 27600 44166 0 _008_
rlabel metal2 26910 44234 26910 44234 0 _009_
rlabel metal2 26634 44540 26634 44540 0 _010_
rlabel metal1 27462 43962 27462 43962 0 _011_
rlabel metal2 25346 44030 25346 44030 0 _012_
rlabel metal1 23736 44914 23736 44914 0 _013_
rlabel metal1 24242 44166 24242 44166 0 _014_
rlabel metal1 22862 44812 22862 44812 0 _015_
rlabel metal2 23506 45305 23506 45305 0 _016_
rlabel metal1 20838 45900 20838 45900 0 _017_
rlabel metal1 20930 45968 20930 45968 0 _018_
rlabel metal2 22770 46342 22770 46342 0 _019_
rlabel metal2 38870 46240 38870 46240 0 _020_
rlabel metal2 38134 46342 38134 46342 0 _021_
rlabel metal1 31602 46580 31602 46580 0 _022_
rlabel metal1 31832 46002 31832 46002 0 _023_
rlabel metal2 37490 44710 37490 44710 0 _024_
rlabel metal1 33488 44914 33488 44914 0 _025_
rlabel metal2 32614 44710 32614 44710 0 _026_
rlabel metal1 35512 43962 35512 43962 0 _027_
rlabel metal1 35880 44710 35880 44710 0 _028_
rlabel metal1 35282 44880 35282 44880 0 _029_
rlabel via1 34638 44506 34638 44506 0 _030_
rlabel metal1 35374 44166 35374 44166 0 _031_
rlabel metal1 32706 45492 32706 45492 0 _032_
rlabel metal1 31832 44914 31832 44914 0 _033_
rlabel metal2 32338 44982 32338 44982 0 _034_
rlabel metal2 31786 45390 31786 45390 0 _035_
rlabel metal1 32522 46002 32522 46002 0 _036_
rlabel metal2 29394 45764 29394 45764 0 _037_
rlabel metal2 29210 46308 29210 46308 0 _038_
rlabel metal1 22816 46478 22816 46478 0 _039_
rlabel metal1 28244 46546 28244 46546 0 _040_
rlabel metal1 25806 46682 25806 46682 0 _041_
rlabel metal1 25484 46002 25484 46002 0 _042_
rlabel metal1 20148 46546 20148 46546 0 _043_
rlabel metal2 30682 46206 30682 46206 0 _044_
rlabel metal1 33902 46682 33902 46682 0 _045_
rlabel metal1 33396 46002 33396 46002 0 _046_
rlabel metal2 19826 45985 19826 45985 0 _047_
rlabel metal1 18262 45968 18262 45968 0 _048_
rlabel metal2 20102 45594 20102 45594 0 _049_
rlabel metal1 26818 43792 26818 43792 0 _050_
rlabel metal1 26634 43962 26634 43962 0 _051_
rlabel metal1 27881 45944 27881 45944 0 _052_
rlabel metal1 26542 45900 26542 45900 0 _053_
rlabel metal2 21574 46240 21574 46240 0 _054_
rlabel metal1 34730 44336 34730 44336 0 _055_
rlabel metal1 35098 44472 35098 44472 0 _056_
rlabel metal2 36018 46138 36018 46138 0 _057_
rlabel metal1 37674 45492 37674 45492 0 _058_
rlabel metal2 22034 45448 22034 45448 0 _059_
rlabel metal1 19320 45934 19320 45934 0 _060_
rlabel metal2 21758 44778 21758 44778 0 _061_
rlabel metal1 26588 45526 26588 45526 0 _062_
rlabel metal1 26082 45390 26082 45390 0 _063_
rlabel metal1 25484 43826 25484 43826 0 _064_
rlabel metal1 25760 44506 25760 44506 0 _065_
rlabel metal1 25668 43146 25668 43146 0 _066_
rlabel metal1 22310 45458 22310 45458 0 _067_
rlabel metal1 33718 45390 33718 45390 0 _068_
rlabel metal1 33672 44506 33672 44506 0 _069_
rlabel metal1 33350 45050 33350 45050 0 _070_
rlabel via1 33971 45526 33971 45526 0 _071_
rlabel metal2 34086 44676 34086 44676 0 _072_
rlabel metal1 20746 45560 20746 45560 0 _073_
rlabel metal2 20838 44540 20838 44540 0 _074_
rlabel metal2 22402 44506 22402 44506 0 _075_
rlabel metal1 23598 44370 23598 44370 0 _076_
rlabel metal2 23322 44506 23322 44506 0 _077_
rlabel metal1 24012 44506 24012 44506 0 _078_
rlabel metal1 23736 43418 23736 43418 0 _079_
rlabel viali 24426 46545 24426 46545 0 _080_
rlabel via2 24334 46461 24334 46461 0 _081_
rlabel metal1 23276 43962 23276 43962 0 _082_
rlabel metal1 30866 45458 30866 45458 0 _083_
rlabel metal1 30912 45050 30912 45050 0 _084_
rlabel metal2 30774 46240 30774 46240 0 _085_
rlabel metal1 37076 46546 37076 46546 0 _086_
rlabel metal1 30314 46444 30314 46444 0 _087_
rlabel metal2 30314 46784 30314 46784 0 _088_
rlabel metal1 19228 5542 19228 5542 0 _089_
rlabel metal1 24058 3570 24058 3570 0 _090_
rlabel metal1 18492 3502 18492 3502 0 _091_
rlabel metal1 22632 6766 22632 6766 0 _092_
rlabel metal2 20102 4828 20102 4828 0 _093_
rlabel metal1 17434 3706 17434 3706 0 _094_
rlabel metal2 17526 3502 17526 3502 0 _095_
rlabel metal2 16790 2924 16790 2924 0 _096_
rlabel metal2 21758 4556 21758 4556 0 _097_
rlabel metal1 19136 4046 19136 4046 0 _098_
rlabel metal2 17894 2652 17894 2652 0 _099_
rlabel metal2 22402 6188 22402 6188 0 _100_
rlabel metal1 22678 5270 22678 5270 0 _101_
rlabel metal1 22402 4692 22402 4692 0 _102_
rlabel metal1 19642 2958 19642 2958 0 _103_
rlabel metal1 21528 2346 21528 2346 0 _104_
rlabel metal1 21482 3094 21482 3094 0 _105_
rlabel metal1 22356 3706 22356 3706 0 _106_
rlabel metal2 24518 6494 24518 6494 0 _107_
rlabel metal2 24610 6222 24610 6222 0 _108_
rlabel metal1 24426 3094 24426 3094 0 _109_
rlabel metal2 26450 4828 26450 4828 0 _110_
rlabel metal1 25346 3434 25346 3434 0 _111_
rlabel metal1 25438 4522 25438 4522 0 _112_
rlabel metal1 27830 5610 27830 5610 0 _113_
rlabel metal2 28842 3230 28842 3230 0 _114_
rlabel metal1 28842 2516 28842 2516 0 _115_
rlabel metal2 27922 3876 27922 3876 0 _116_
rlabel metal2 28014 4964 28014 4964 0 _117_
rlabel metal2 27738 6494 27738 6494 0 _118_
rlabel metal1 31924 3434 31924 3434 0 _119_
rlabel metal1 32108 3094 32108 3094 0 _120_
rlabel metal2 29670 5406 29670 5406 0 _121_
rlabel metal1 31142 4012 31142 4012 0 _122_
rlabel metal1 31648 2346 31648 2346 0 _123_
rlabel metal1 29578 46580 29578 46580 0 _124_
rlabel metal2 4094 48195 4094 48195 0 io_active
rlabel metal1 22632 44370 22632 44370 0 io_in[18]
rlabel metal1 24150 45492 24150 45492 0 io_in[19]
rlabel metal2 27186 44676 27186 44676 0 io_in[20]
rlabel via2 27738 42347 27738 42347 0 io_in[21]
rlabel metal2 28842 46529 28842 46529 0 io_in[22]
rlabel metal1 29808 47022 29808 47022 0 io_in[23]
rlabel metal1 32292 47022 32292 47022 0 io_in[24]
rlabel metal1 32200 46478 32200 46478 0 io_in[25]
rlabel metal1 33396 43282 33396 43282 0 io_in[26]
rlabel metal1 34730 43282 34730 43282 0 io_in[27]
rlabel metal1 36202 46954 36202 46954 0 io_in[28]
rlabel metal1 38180 44846 38180 44846 0 io_in[29]
rlabel metal2 41998 46903 41998 46903 0 io_in[30]
rlabel metal1 39008 45050 39008 45050 0 io_in[31]
rlabel metal2 40020 47090 40020 47090 0 io_in[32]
rlabel metal2 40894 47923 40894 47923 0 io_in[33]
rlabel metal1 42918 46988 42918 46988 0 io_in[34]
rlabel metal1 43332 47022 43332 47022 0 io_in[35]
rlabel metal1 44344 47022 44344 47022 0 io_in[36]
rlabel metal2 45218 47712 45218 47712 0 io_in[37]
rlabel metal1 5290 47226 5290 47226 0 io_out[0]
rlabel metal2 16146 48256 16146 48256 0 io_out[10]
rlabel metal2 17250 48256 17250 48256 0 io_out[11]
rlabel metal2 18446 47991 18446 47991 0 io_out[12]
rlabel metal1 18722 47226 18722 47226 0 io_out[13]
rlabel metal1 19872 46682 19872 46682 0 io_out[14]
rlabel metal1 19458 47158 19458 47158 0 io_out[15]
rlabel metal2 22770 48256 22770 48256 0 io_out[16]
rlabel metal1 24334 47226 24334 47226 0 io_out[17]
rlabel metal2 9706 47651 9706 47651 0 io_out[4]
rlabel metal2 10810 48263 10810 48263 0 io_out[5]
rlabel metal2 11914 48263 11914 48263 0 io_out[6]
rlabel metal2 13018 48263 13018 48263 0 io_out[7]
rlabel metal1 14168 47226 14168 47226 0 io_out[8]
rlabel metal2 15226 47651 15226 47651 0 io_out[9]
rlabel metal2 21114 2710 21114 2710 0 la_data_out[32]
rlabel metal2 21390 2948 21390 2948 0 la_data_out[33]
rlabel metal2 21666 1792 21666 1792 0 la_data_out[34]
rlabel metal2 21942 1520 21942 1520 0 la_data_out[35]
rlabel metal2 22218 2166 22218 2166 0 la_data_out[36]
rlabel metal2 22494 1435 22494 1435 0 la_data_out[37]
rlabel metal2 22770 1622 22770 1622 0 la_data_out[38]
rlabel metal2 23046 1792 23046 1792 0 la_data_out[39]
rlabel metal2 23322 1775 23322 1775 0 la_data_out[40]
rlabel metal2 23598 2710 23598 2710 0 la_data_out[41]
rlabel metal2 23874 1860 23874 1860 0 la_data_out[42]
rlabel metal2 24150 1554 24150 1554 0 la_data_out[43]
rlabel metal2 24426 1860 24426 1860 0 la_data_out[44]
rlabel metal2 24702 2404 24702 2404 0 la_data_out[45]
rlabel metal2 24978 3492 24978 3492 0 la_data_out[46]
rlabel metal2 25254 2948 25254 2948 0 la_data_out[47]
rlabel metal2 25530 1860 25530 1860 0 la_data_out[48]
rlabel metal2 25806 1622 25806 1622 0 la_data_out[49]
rlabel metal2 26082 2166 26082 2166 0 la_data_out[50]
rlabel metal2 26358 2710 26358 2710 0 la_data_out[51]
rlabel metal2 26634 3186 26634 3186 0 la_data_out[52]
rlabel metal2 26910 1860 26910 1860 0 la_data_out[53]
rlabel metal2 27186 1554 27186 1554 0 la_data_out[54]
rlabel metal2 27462 2404 27462 2404 0 la_data_out[55]
rlabel metal2 27738 2914 27738 2914 0 la_data_out[56]
rlabel metal2 28014 1962 28014 1962 0 la_data_out[57]
rlabel metal2 28290 2098 28290 2098 0 la_data_out[58]
rlabel metal2 28566 1860 28566 1860 0 la_data_out[59]
rlabel metal2 28842 1792 28842 1792 0 la_data_out[60]
rlabel metal2 29118 2404 29118 2404 0 la_data_out[61]
rlabel metal2 29394 1554 29394 1554 0 la_data_out[62]
rlabel metal2 29670 2132 29670 2132 0 la_data_out[63]
rlabel metal2 11730 47260 11730 47260 0 net1
rlabel metal1 33902 45050 33902 45050 0 net10
rlabel metal2 30774 2234 30774 2234 0 net100
rlabel metal2 31050 1826 31050 1826 0 net101
rlabel metal2 31326 1367 31326 1367 0 net102
rlabel metal2 31602 2438 31602 2438 0 net103
rlabel metal2 31878 1027 31878 1027 0 net104
rlabel metal2 32154 1299 32154 1299 0 net105
rlabel metal2 32430 1095 32430 1095 0 net106
rlabel metal2 32706 1367 32706 1367 0 net107
rlabel metal2 32982 1761 32982 1761 0 net108
rlabel metal1 34086 3638 34086 3638 0 net109
rlabel metal1 35282 45526 35282 45526 0 net11
rlabel metal1 34868 3094 34868 3094 0 net110
rlabel metal1 34040 3910 34040 3910 0 net111
rlabel metal1 34500 3978 34500 3978 0 net112
rlabel metal1 35282 2890 35282 2890 0 net113
rlabel metal1 35098 3570 35098 3570 0 net114
rlabel metal1 37444 2618 37444 2618 0 net115
rlabel metal2 35190 1367 35190 1367 0 net116
rlabel metal1 35834 3638 35834 3638 0 net117
rlabel metal1 36616 3026 36616 3026 0 net118
rlabel metal1 36432 3570 36432 3570 0 net119
rlabel via1 36018 45475 36018 45475 0 net12
rlabel metal2 36294 1588 36294 1588 0 net120
rlabel metal1 37030 3502 37030 3502 0 net121
rlabel metal1 37490 2890 37490 2890 0 net122
rlabel metal2 37122 1622 37122 1622 0 net123
rlabel metal2 37398 1299 37398 1299 0 net124
rlabel metal1 38226 2958 38226 2958 0 net125
rlabel metal1 38364 3502 38364 3502 0 net126
rlabel metal2 38226 1656 38226 1656 0 net127
rlabel metal1 38962 2890 38962 2890 0 net128
rlabel metal1 39422 2822 39422 2822 0 net129
rlabel metal2 37674 46036 37674 46036 0 net13
rlabel metal2 39054 1622 39054 1622 0 net130
rlabel metal1 39698 3502 39698 3502 0 net131
rlabel metal2 39606 1588 39606 1588 0 net132
rlabel metal1 40296 2958 40296 2958 0 net133
rlabel metal1 40434 3502 40434 3502 0 net134
rlabel metal1 40894 2890 40894 2890 0 net135
rlabel metal1 41032 3638 41032 3638 0 net136
rlabel metal2 40986 1622 40986 1622 0 net137
rlabel metal2 41262 2166 41262 2166 0 net138
rlabel metal2 41538 1588 41538 1588 0 net139
rlabel metal1 36432 44846 36432 44846 0 net14
rlabel metal2 41814 1792 41814 1792 0 net140
rlabel metal2 42090 1656 42090 1656 0 net141
rlabel metal2 42366 1860 42366 1860 0 net142
rlabel metal2 42642 2132 42642 2132 0 net143
rlabel metal2 42918 2132 42918 2132 0 net144
rlabel metal2 43194 1826 43194 1826 0 net145
rlabel metal2 43470 1622 43470 1622 0 net146
rlabel metal2 43746 1792 43746 1792 0 net147
rlabel metal2 44022 1554 44022 1554 0 net148
rlabel metal2 44298 1860 44298 1860 0 net149
rlabel metal1 38226 46478 38226 46478 0 net15
rlabel metal2 44574 2132 44574 2132 0 net150
rlabel metal2 44850 1656 44850 1656 0 net151
rlabel metal2 45126 1826 45126 1826 0 net152
rlabel metal2 45402 2132 45402 2132 0 net153
rlabel metal2 45678 1792 45678 1792 0 net154
rlabel metal2 45954 1588 45954 1588 0 net155
rlabel metal2 46230 2132 46230 2132 0 net156
rlabel metal2 46506 2200 46506 2200 0 net157
rlabel metal2 46782 1792 46782 1792 0 net158
rlabel metal2 47058 2166 47058 2166 0 net159
rlabel metal1 38186 45934 38186 45934 0 net16
rlabel metal2 47334 2336 47334 2336 0 net160
rlabel metal2 2622 1588 2622 1588 0 net161
rlabel metal2 3174 1588 3174 1588 0 net162
rlabel metal2 3542 1792 3542 1792 0 net163
rlabel metal2 3910 1588 3910 1588 0 net164
rlabel metal2 4278 1299 4278 1299 0 net165
rlabel metal2 4646 1095 4646 1095 0 net166
rlabel metal2 4922 2132 4922 2132 0 net167
rlabel metal2 5198 1792 5198 1792 0 net168
rlabel metal2 5474 1622 5474 1622 0 net169
rlabel metal1 37444 45934 37444 45934 0 net17
rlabel metal2 5750 2132 5750 2132 0 net170
rlabel metal2 6026 1860 6026 1860 0 net171
rlabel metal2 6302 1792 6302 1792 0 net172
rlabel metal2 6578 2132 6578 2132 0 net173
rlabel metal2 6854 1656 6854 1656 0 net174
rlabel metal2 7130 1588 7130 1588 0 net175
rlabel metal2 7406 2132 7406 2132 0 net176
rlabel metal2 7682 1792 7682 1792 0 net177
rlabel metal2 7958 1656 7958 1656 0 net178
rlabel metal2 8234 2132 8234 2132 0 net179
rlabel metal1 35236 46002 35236 46002 0 net18
rlabel metal2 8510 1792 8510 1792 0 net180
rlabel metal2 8786 1792 8786 1792 0 net181
rlabel metal2 9062 2132 9062 2132 0 net182
rlabel metal2 9338 1554 9338 1554 0 net183
rlabel metal2 9614 1792 9614 1792 0 net184
rlabel metal2 9890 2132 9890 2132 0 net185
rlabel metal2 10166 1622 10166 1622 0 net186
rlabel metal2 10442 1792 10442 1792 0 net187
rlabel metal2 10718 2132 10718 2132 0 net188
rlabel metal2 10994 1792 10994 1792 0 net189
rlabel metal2 43470 47328 43470 47328 0 net19
rlabel metal2 11270 1656 11270 1656 0 net190
rlabel metal2 11546 2132 11546 2132 0 net191
rlabel metal2 11822 1792 11822 1792 0 net192
rlabel metal2 12098 1588 12098 1588 0 net193
rlabel metal1 19918 4692 19918 4692 0 net194
rlabel metal1 19642 5236 19642 5236 0 net195
rlabel metal1 17710 2958 17710 2958 0 net196
rlabel metal1 16698 2414 16698 2414 0 net197
rlabel metal1 21206 3570 21206 3570 0 net198
rlabel metal1 19550 4114 19550 4114 0 net199
rlabel metal2 25990 44744 25990 44744 0 net2
rlabel metal1 37720 46342 37720 46342 0 net20
rlabel metal1 19458 2414 19458 2414 0 net200
rlabel metal2 22218 5916 22218 5916 0 net201
rlabel metal2 22126 5678 22126 5678 0 net202
rlabel metal1 22678 4794 22678 4794 0 net203
rlabel metal1 21712 3162 21712 3162 0 net204
rlabel metal1 22172 2414 22172 2414 0 net205
rlabel metal2 22494 3230 22494 3230 0 net206
rlabel metal1 23276 4046 23276 4046 0 net207
rlabel metal1 24104 6222 24104 6222 0 net208
rlabel metal1 23874 4114 23874 4114 0 net209
rlabel metal1 43470 47090 43470 47090 0 net21
rlabel metal2 24794 3468 24794 3468 0 net210
rlabel metal1 26680 2482 26680 2482 0 net211
rlabel metal2 25530 3740 25530 3740 0 net212
rlabel metal1 25668 7174 25668 7174 0 net213
rlabel metal1 26956 5746 26956 5746 0 net214
rlabel metal2 29026 3264 29026 3264 0 net215
rlabel metal1 29716 2482 29716 2482 0 net216
rlabel metal2 29026 4352 29026 4352 0 net217
rlabel metal2 29026 5440 29026 5440 0 net218
rlabel metal2 27554 6528 27554 6528 0 net219
rlabel metal2 5658 46750 5658 46750 0 net22
rlabel metal1 31418 3570 31418 3570 0 net220
rlabel metal1 32154 2958 32154 2958 0 net221
rlabel metal2 29762 4964 29762 4964 0 net222
rlabel metal2 31326 4386 31326 4386 0 net223
rlabel metal1 32154 2482 32154 2482 0 net224
rlabel metal1 31234 43962 31234 43962 0 net225
rlabel metal2 4830 47923 4830 47923 0 net226
rlabel metal2 5934 47719 5934 47719 0 net227
rlabel metal2 7038 47923 7038 47923 0 net228
rlabel metal2 7958 48263 7958 48263 0 net229
rlabel metal2 18078 46614 18078 46614 0 net23
rlabel metal2 9246 47923 9246 47923 0 net230
rlabel metal2 10350 47923 10350 47923 0 net231
rlabel metal1 11546 46546 11546 46546 0 net232
rlabel metal2 12558 47923 12558 47923 0 net233
rlabel metal2 13662 47923 13662 47923 0 net234
rlabel metal2 14766 47923 14766 47923 0 net235
rlabel metal2 15870 47923 15870 47923 0 net236
rlabel metal2 16974 47719 16974 47719 0 net237
rlabel metal1 17618 46546 17618 46546 0 net238
rlabel metal1 18814 45458 18814 45458 0 net239
rlabel metal2 18722 46512 18722 46512 0 net24
rlabel metal1 19688 45390 19688 45390 0 net240
rlabel metal1 18354 46342 18354 46342 0 net241
rlabel metal2 22494 44727 22494 44727 0 net242
rlabel metal1 23368 43282 23368 43282 0 net243
rlabel metal2 24702 44336 24702 44336 0 net244
rlabel metal1 23552 46546 23552 46546 0 net245
rlabel metal2 26818 48222 26818 48222 0 net246
rlabel metal1 28336 43214 28336 43214 0 net247
rlabel metal1 29210 43282 29210 43282 0 net248
rlabel metal1 35098 46580 35098 46580 0 net249
rlabel metal1 21022 44472 21022 44472 0 net25
rlabel metal2 31326 46291 31326 46291 0 net250
rlabel metal1 32706 43282 32706 43282 0 net251
rlabel metal1 33810 43214 33810 43214 0 net252
rlabel metal1 39238 45934 39238 45934 0 net253
rlabel metal1 36064 43962 36064 43962 0 net254
rlabel metal2 39238 45628 39238 45628 0 net255
rlabel metal1 39468 46002 39468 46002 0 net256
rlabel metal1 39836 46138 39836 46138 0 net257
rlabel metal1 40848 46070 40848 46070 0 net258
rlabel metal2 18170 47226 18170 47226 0 net26
rlabel metal2 19366 45798 19366 45798 0 net27
rlabel metal2 20930 45118 20930 45118 0 net28
rlabel metal2 21114 44608 21114 44608 0 net29
rlabel metal1 26680 44846 26680 44846 0 net3
rlabel metal1 24150 47090 24150 47090 0 net30
rlabel metal2 9890 46410 9890 46410 0 net31
rlabel metal2 10994 47430 10994 47430 0 net32
rlabel metal1 12098 46988 12098 46988 0 net33
rlabel metal2 21482 46920 21482 46920 0 net34
rlabel metal1 20470 45254 20470 45254 0 net35
rlabel metal2 15410 47396 15410 47396 0 net36
rlabel metal2 41170 47712 41170 47712 0 net37
rlabel metal1 42458 46138 42458 46138 0 net38
rlabel metal1 43654 46546 43654 46546 0 net39
rlabel metal2 27646 46240 27646 46240 0 net4
rlabel metal1 44850 46546 44850 46546 0 net40
rlabel metal2 45862 47923 45862 47923 0 net41
rlabel metal2 6026 47923 6026 47923 0 net42
rlabel metal2 7314 48256 7314 48256 0 net43
rlabel metal2 8418 48256 8418 48256 0 net44
rlabel metal1 25438 43962 25438 43962 0 net45
rlabel metal1 26266 47226 26266 47226 0 net46
rlabel metal2 27278 46019 27278 46019 0 net47
rlabel metal1 28428 42738 28428 42738 0 net48
rlabel metal1 29854 43282 29854 43282 0 net49
rlabel metal1 27232 46546 27232 46546 0 net5
rlabel metal1 30958 43894 30958 43894 0 net50
rlabel metal2 31694 43809 31694 43809 0 net51
rlabel metal1 33396 43826 33396 43826 0 net52
rlabel via2 39146 46563 39146 46563 0 net53
rlabel metal1 39790 46614 39790 46614 0 net54
rlabel metal1 38686 47158 38686 47158 0 net55
rlabel metal1 38732 44914 38732 44914 0 net56
rlabel metal1 39468 45458 39468 45458 0 net57
rlabel metal1 40296 45390 40296 45390 0 net58
rlabel metal1 40802 45458 40802 45458 0 net59
rlabel metal1 29394 43826 29394 43826 0 net6
rlabel metal1 42090 46410 42090 46410 0 net60
rlabel metal1 42964 46546 42964 46546 0 net61
rlabel metal1 44160 46478 44160 46478 0 net62
rlabel metal1 45494 46920 45494 46920 0 net63
rlabel metal1 46322 47226 46322 47226 0 net64
rlabel metal2 12282 2336 12282 2336 0 net65
rlabel metal2 12558 1622 12558 1622 0 net66
rlabel metal2 12834 2132 12834 2132 0 net67
rlabel metal2 13110 2336 13110 2336 0 net68
rlabel metal2 13386 1826 13386 1826 0 net69
rlabel metal1 29716 45390 29716 45390 0 net7
rlabel metal2 13662 2132 13662 2132 0 net70
rlabel metal2 13938 2336 13938 2336 0 net71
rlabel metal2 14214 2132 14214 2132 0 net72
rlabel metal2 14490 1894 14490 1894 0 net73
rlabel metal2 14766 1656 14766 1656 0 net74
rlabel metal2 15042 2676 15042 2676 0 net75
rlabel metal2 15318 2336 15318 2336 0 net76
rlabel metal2 15594 1027 15594 1027 0 net77
rlabel metal2 15870 2676 15870 2676 0 net78
rlabel metal2 16146 1792 16146 1792 0 net79
rlabel metal2 31970 46444 31970 46444 0 net8
rlabel metal2 16422 2200 16422 2200 0 net80
rlabel metal2 16698 1860 16698 1860 0 net81
rlabel metal2 16974 2880 16974 2880 0 net82
rlabel metal2 17250 2404 17250 2404 0 net83
rlabel metal2 17526 1571 17526 1571 0 net84
rlabel metal2 17802 1367 17802 1367 0 net85
rlabel metal2 18078 1690 18078 1690 0 net86
rlabel metal2 18354 2880 18354 2880 0 net87
rlabel metal2 18630 3220 18630 3220 0 net88
rlabel metal2 18906 1792 18906 1792 0 net89
rlabel metal2 32614 46308 32614 46308 0 net9
rlabel metal2 19182 1962 19182 1962 0 net90
rlabel metal2 19458 1231 19458 1231 0 net91
rlabel metal2 19734 1350 19734 1350 0 net92
rlabel metal2 20010 2914 20010 2914 0 net93
rlabel metal2 20286 1384 20286 1384 0 net94
rlabel metal2 20562 2200 20562 2200 0 net95
rlabel metal2 20838 1418 20838 1418 0 net96
rlabel metal2 29946 1962 29946 1962 0 net97
rlabel metal2 30222 2200 30222 2200 0 net98
rlabel metal2 30498 2064 30498 2064 0 net99
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
