magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -36 538 512 1177
<< locali >>
rect 0 1103 476 1137
rect 64 501 98 567
rect 183 517 217 551
rect 0 -17 476 17
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0
timestamp 1666199351
transform 1 0 0 0 1 0
box -36 -17 512 1177
<< labels >>
rlabel locali s 200 534 200 534 4 Z
port 1 nsew
rlabel locali s 81 534 81 534 4 A
port 2 nsew
rlabel locali s 238 0 238 0 4 gnd
port 3 nsew
rlabel locali s 238 1120 238 1120 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 476 1120
string GDS_END 62650
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 61822
<< end >>
