magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 98 157 459 203
rect 1 21 459 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 174 47 204 177
rect 349 47 379 177
<< scpmoshvt >>
rect 79 413 109 497
rect 246 297 276 497
rect 349 297 379 497
<< ndiff >>
rect 124 131 174 177
rect 27 106 79 131
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 89 174 131
rect 109 55 119 89
rect 153 55 174 89
rect 109 47 174 55
rect 204 47 349 177
rect 379 161 433 177
rect 379 127 389 161
rect 423 127 433 161
rect 379 93 433 127
rect 379 59 389 93
rect 423 59 433 93
rect 379 47 433 59
<< pdiff >>
rect 27 472 79 497
rect 27 438 35 472
rect 69 438 79 472
rect 27 413 79 438
rect 109 488 246 497
rect 109 454 121 488
rect 155 454 189 488
rect 223 454 246 488
rect 109 413 246 454
rect 124 297 246 413
rect 276 297 349 497
rect 379 477 433 497
rect 379 443 391 477
rect 425 443 433 477
rect 379 297 433 443
<< ndiffc >>
rect 35 72 69 106
rect 119 55 153 89
rect 389 127 423 161
rect 389 59 423 93
<< pdiffc >>
rect 35 438 69 472
rect 121 454 155 488
rect 189 454 223 488
rect 391 443 425 477
<< poly >>
rect 79 497 109 523
rect 246 497 276 523
rect 349 497 379 523
rect 79 261 109 413
rect 22 249 109 261
rect 22 215 38 249
rect 72 222 109 249
rect 246 265 276 297
rect 349 265 379 297
rect 246 249 300 265
rect 72 215 204 222
rect 22 203 204 215
rect 79 192 204 203
rect 246 215 256 249
rect 290 215 300 249
rect 246 199 300 215
rect 349 249 439 265
rect 349 215 395 249
rect 429 215 439 249
rect 349 199 439 215
rect 79 131 109 192
rect 174 177 204 192
rect 349 177 379 199
rect 79 21 109 47
rect 174 21 204 47
rect 349 21 379 47
<< polycont >>
rect 38 215 72 249
rect 256 215 290 249
rect 395 215 429 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 17 472 69 493
rect 17 438 35 472
rect 103 488 290 527
rect 103 454 121 488
rect 155 454 189 488
rect 223 454 290 488
rect 103 447 290 454
rect 324 477 443 493
rect 17 413 69 438
rect 324 443 391 477
rect 425 443 443 477
rect 324 425 443 443
rect 17 379 290 413
rect 17 249 109 345
rect 17 215 38 249
rect 72 215 109 249
rect 17 199 109 215
rect 143 249 290 379
rect 143 215 256 249
rect 143 165 290 215
rect 17 131 290 165
rect 324 161 359 425
rect 395 249 443 391
rect 429 215 443 249
rect 395 195 443 215
rect 17 106 69 131
rect 17 72 35 106
rect 324 127 389 161
rect 423 127 443 161
rect 17 51 69 72
rect 103 89 290 97
rect 103 55 119 89
rect 153 55 290 89
rect 103 17 290 55
rect 324 93 443 127
rect 324 59 389 93
rect 423 59 443 93
rect 324 51 443 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 TE
port 2 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 TE
port 2 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 398 357 432 391 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 398 289 432 323 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 398 425 432 459 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 398 85 432 119 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 einvp_1
rlabel metal1 s 0 -48 460 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 2024636
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2020124
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 11.500 0.000 
<< end >>
