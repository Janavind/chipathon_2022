magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1169 203
rect 30 -17 64 21
<< locali >>
rect 98 153 156 335
rect 190 153 256 285
rect 379 289 1179 345
rect 1135 171 1179 289
rect 829 123 1179 171
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 353 69 493
rect 103 369 186 527
rect 220 353 271 493
rect 313 421 362 493
rect 396 455 462 527
rect 496 421 530 493
rect 564 455 630 527
rect 664 421 1179 493
rect 313 387 1179 421
rect 379 379 1179 387
rect 17 133 64 353
rect 220 319 345 353
rect 290 255 345 319
rect 290 205 762 255
rect 796 205 1101 255
rect 17 56 69 133
rect 290 119 345 205
rect 103 17 186 119
rect 220 51 345 119
rect 379 131 795 171
rect 379 51 435 131
rect 469 17 535 97
rect 569 55 603 131
rect 637 17 703 97
rect 737 89 795 131
rect 737 51 1147 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< obsm1 >>
rect 17 252 76 261
rect 850 252 908 261
rect 17 224 908 252
rect 17 215 76 224
rect 850 215 908 224
<< labels >>
rlabel locali s 98 153 156 335 6 A
port 1 nsew signal input
rlabel locali s 190 153 256 285 6 TE_B
port 2 nsew signal input
rlabel metal1 s 0 -48 1196 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 1169 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 829 123 1179 171 6 Z
port 7 nsew signal output
rlabel locali s 1135 171 1179 289 6 Z
port 7 nsew signal output
rlabel locali s 379 289 1179 345 6 Z
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1196 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2956310
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2946864
<< end >>
