magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< dnwell >>
rect -2476 -1400 2776 7401
<< nwell >>
rect -2076 6801 2376 7001
rect -2076 -799 -1876 6801
rect -10 0 310 6000
rect 2176 -799 2376 6801
rect -2076 -999 2376 -799
<< pwell >>
rect -3084 7875 3384 8009
rect -3084 -1874 -2950 7875
rect -1102 -26 -374 6026
rect 674 -26 1402 6026
rect 3250 -1874 3384 7875
rect -3084 -2008 3384 -1874
<< obsactive >>
rect -3158 -2082 3458 8083
<< locali >>
rect -3058 7959 3358 7983
rect -3058 7925 -2927 7959
rect -2893 7925 -2855 7959
rect -2821 7925 -2783 7959
rect -2749 7925 -2711 7959
rect -2677 7925 -2639 7959
rect -2605 7925 -2567 7959
rect -2533 7925 -2495 7959
rect -2461 7925 -2423 7959
rect -2389 7925 -2351 7959
rect -2317 7925 -2279 7959
rect -2245 7925 -2207 7959
rect -2173 7925 -2135 7959
rect -2101 7925 -2063 7959
rect -2029 7925 -1991 7959
rect -1957 7925 -1919 7959
rect -1885 7925 -1847 7959
rect -1813 7925 -1775 7959
rect -1741 7925 -1703 7959
rect -1669 7925 -1631 7959
rect -1597 7925 -1559 7959
rect -1525 7925 -1487 7959
rect -1453 7925 -1415 7959
rect -1381 7925 -1343 7959
rect -1309 7925 -1271 7959
rect -1237 7925 -1199 7959
rect -1165 7925 -1127 7959
rect -1093 7925 -1055 7959
rect -1021 7925 -983 7959
rect -949 7925 -911 7959
rect -877 7925 -839 7959
rect -805 7925 -767 7959
rect -733 7925 -695 7959
rect -661 7925 -623 7959
rect -589 7925 -551 7959
rect -517 7925 -479 7959
rect -445 7925 -407 7959
rect -373 7925 -335 7959
rect -301 7925 -263 7959
rect -229 7925 -191 7959
rect -157 7925 -119 7959
rect -85 7925 -47 7959
rect -13 7925 25 7959
rect 59 7925 97 7959
rect 131 7925 169 7959
rect 203 7925 241 7959
rect 275 7925 313 7959
rect 347 7925 385 7959
rect 419 7925 457 7959
rect 491 7925 529 7959
rect 563 7925 601 7959
rect 635 7925 673 7959
rect 707 7925 745 7959
rect 779 7925 817 7959
rect 851 7925 889 7959
rect 923 7925 961 7959
rect 995 7925 1033 7959
rect 1067 7925 1105 7959
rect 1139 7925 1177 7959
rect 1211 7925 1249 7959
rect 1283 7925 1321 7959
rect 1355 7925 1393 7959
rect 1427 7925 1465 7959
rect 1499 7925 1537 7959
rect 1571 7925 1609 7959
rect 1643 7925 1681 7959
rect 1715 7925 1753 7959
rect 1787 7925 1825 7959
rect 1859 7925 1897 7959
rect 1931 7925 1969 7959
rect 2003 7925 2041 7959
rect 2075 7925 2113 7959
rect 2147 7925 2185 7959
rect 2219 7925 2257 7959
rect 2291 7925 2329 7959
rect 2363 7925 2401 7959
rect 2435 7925 2473 7959
rect 2507 7925 2545 7959
rect 2579 7925 2617 7959
rect 2651 7925 2689 7959
rect 2723 7925 2761 7959
rect 2795 7925 2833 7959
rect 2867 7925 2905 7959
rect 2939 7925 2977 7959
rect 3011 7925 3049 7959
rect 3083 7925 3121 7959
rect 3155 7925 3193 7959
rect 3227 7925 3358 7959
rect -3058 7901 3358 7925
rect -3058 7877 -2976 7901
rect -3058 7843 -3034 7877
rect -3000 7843 -2976 7877
rect -3058 7805 -2976 7843
rect -3058 7771 -3034 7805
rect -3000 7771 -2976 7805
rect -3058 7733 -2976 7771
rect -3058 7699 -3034 7733
rect -3000 7699 -2976 7733
rect -3058 7661 -2976 7699
rect -3058 7627 -3034 7661
rect -3000 7627 -2976 7661
rect -3058 7589 -2976 7627
rect -3058 7555 -3034 7589
rect -3000 7555 -2976 7589
rect -3058 7517 -2976 7555
rect -3058 7483 -3034 7517
rect -3000 7483 -2976 7517
rect -3058 7445 -2976 7483
rect -3058 7411 -3034 7445
rect -3000 7411 -2976 7445
rect -3058 7373 -2976 7411
rect -3058 7339 -3034 7373
rect -3000 7339 -2976 7373
rect -3058 7301 -2976 7339
rect -3058 7267 -3034 7301
rect -3000 7267 -2976 7301
rect -3058 7229 -2976 7267
rect -3058 7195 -3034 7229
rect -3000 7195 -2976 7229
rect -3058 7157 -2976 7195
rect -3058 7123 -3034 7157
rect -3000 7123 -2976 7157
rect -3058 7085 -2976 7123
rect -3058 7051 -3034 7085
rect -3000 7051 -2976 7085
rect -3058 7013 -2976 7051
rect -3058 6979 -3034 7013
rect -3000 6979 -2976 7013
rect -3058 6941 -2976 6979
rect -3058 6907 -3034 6941
rect -3000 6907 -2976 6941
rect -3058 6869 -2976 6907
rect -3058 6835 -3034 6869
rect -3000 6835 -2976 6869
rect -3058 6797 -2976 6835
rect -3058 6763 -3034 6797
rect -3000 6763 -2976 6797
rect -3058 6725 -2976 6763
rect -3058 6691 -3034 6725
rect -3000 6691 -2976 6725
rect -3058 6653 -2976 6691
rect -3058 6619 -3034 6653
rect -3000 6619 -2976 6653
rect -3058 6581 -2976 6619
rect -3058 6547 -3034 6581
rect -3000 6547 -2976 6581
rect -3058 6509 -2976 6547
rect -3058 6475 -3034 6509
rect -3000 6475 -2976 6509
rect -3058 6437 -2976 6475
rect -3058 6403 -3034 6437
rect -3000 6403 -2976 6437
rect -3058 6365 -2976 6403
rect -3058 6331 -3034 6365
rect -3000 6331 -2976 6365
rect -3058 6293 -2976 6331
rect -3058 6259 -3034 6293
rect -3000 6259 -2976 6293
rect -3058 6221 -2976 6259
rect -3058 6187 -3034 6221
rect -3000 6187 -2976 6221
rect -3058 6149 -2976 6187
rect -3058 6115 -3034 6149
rect -3000 6115 -2976 6149
rect -3058 6077 -2976 6115
rect -3058 6043 -3034 6077
rect -3000 6043 -2976 6077
rect -3058 6005 -2976 6043
rect -3058 5971 -3034 6005
rect -3000 5971 -2976 6005
rect 3276 7877 3358 7901
rect 3276 7843 3300 7877
rect 3334 7843 3358 7877
rect 3276 7805 3358 7843
rect 3276 7771 3300 7805
rect 3334 7771 3358 7805
rect 3276 7733 3358 7771
rect 3276 7699 3300 7733
rect 3334 7699 3358 7733
rect 3276 7661 3358 7699
rect 3276 7627 3300 7661
rect 3334 7627 3358 7661
rect 3276 7589 3358 7627
rect 3276 7555 3300 7589
rect 3334 7555 3358 7589
rect 3276 7517 3358 7555
rect 3276 7483 3300 7517
rect 3334 7483 3358 7517
rect 3276 7445 3358 7483
rect 3276 7411 3300 7445
rect 3334 7411 3358 7445
rect 3276 7373 3358 7411
rect 3276 7339 3300 7373
rect 3334 7339 3358 7373
rect 3276 7301 3358 7339
rect 3276 7267 3300 7301
rect 3334 7267 3358 7301
rect 3276 7229 3358 7267
rect 3276 7195 3300 7229
rect 3334 7195 3358 7229
rect 3276 7157 3358 7195
rect 3276 7123 3300 7157
rect 3334 7123 3358 7157
rect 3276 7085 3358 7123
rect 3276 7051 3300 7085
rect 3334 7051 3358 7085
rect 3276 7013 3358 7051
rect 3276 6979 3300 7013
rect 3334 6979 3358 7013
rect 3276 6941 3358 6979
rect 3276 6907 3300 6941
rect 3334 6907 3358 6941
rect 3276 6869 3358 6907
rect 3276 6835 3300 6869
rect 3334 6835 3358 6869
rect 3276 6797 3358 6835
rect 3276 6763 3300 6797
rect 3334 6763 3358 6797
rect 3276 6725 3358 6763
rect 3276 6691 3300 6725
rect 3334 6691 3358 6725
rect 3276 6653 3358 6691
rect 3276 6619 3300 6653
rect 3334 6619 3358 6653
rect 3276 6581 3358 6619
rect 3276 6547 3300 6581
rect 3334 6547 3358 6581
rect 3276 6509 3358 6547
rect 3276 6475 3300 6509
rect 3334 6475 3358 6509
rect 3276 6437 3358 6475
rect 3276 6403 3300 6437
rect 3334 6403 3358 6437
rect 3276 6365 3358 6403
rect 3276 6331 3300 6365
rect 3334 6331 3358 6365
rect 3276 6293 3358 6331
rect 3276 6259 3300 6293
rect 3334 6259 3358 6293
rect 3276 6221 3358 6259
rect 3276 6187 3300 6221
rect 3334 6187 3358 6221
rect 3276 6149 3358 6187
rect 3276 6115 3300 6149
rect 3334 6115 3358 6149
rect 3276 6077 3358 6115
rect 3276 6043 3300 6077
rect 3334 6043 3358 6077
rect 3276 6005 3358 6043
rect -3058 5933 -2976 5971
rect -3058 5899 -3034 5933
rect -3000 5899 -2976 5933
rect -3058 5861 -2976 5899
rect -3058 5827 -3034 5861
rect -3000 5827 -2976 5861
rect -3058 5789 -2976 5827
rect -3058 5755 -3034 5789
rect -3000 5755 -2976 5789
rect -3058 5717 -2976 5755
rect -3058 5683 -3034 5717
rect -3000 5683 -2976 5717
rect -3058 5645 -2976 5683
rect -3058 5611 -3034 5645
rect -3000 5611 -2976 5645
rect -3058 5573 -2976 5611
rect -3058 5539 -3034 5573
rect -3000 5539 -2976 5573
rect -3058 5501 -2976 5539
rect -3058 5467 -3034 5501
rect -3000 5467 -2976 5501
rect -3058 5429 -2976 5467
rect -3058 5395 -3034 5429
rect -3000 5395 -2976 5429
rect -3058 5357 -2976 5395
rect -3058 5323 -3034 5357
rect -3000 5323 -2976 5357
rect -3058 5285 -2976 5323
rect -3058 5251 -3034 5285
rect -3000 5251 -2976 5285
rect -3058 5213 -2976 5251
rect -3058 5179 -3034 5213
rect -3000 5179 -2976 5213
rect -3058 5141 -2976 5179
rect -3058 5107 -3034 5141
rect -3000 5107 -2976 5141
rect -3058 5069 -2976 5107
rect -3058 5035 -3034 5069
rect -3000 5035 -2976 5069
rect -3058 4997 -2976 5035
rect -3058 4963 -3034 4997
rect -3000 4963 -2976 4997
rect -3058 4925 -2976 4963
rect -3058 4891 -3034 4925
rect -3000 4891 -2976 4925
rect -3058 4853 -2976 4891
rect -3058 4819 -3034 4853
rect -3000 4819 -2976 4853
rect -3058 4781 -2976 4819
rect -3058 4747 -3034 4781
rect -3000 4747 -2976 4781
rect -3058 4709 -2976 4747
rect -3058 4675 -3034 4709
rect -3000 4675 -2976 4709
rect -3058 4637 -2976 4675
rect -3058 4603 -3034 4637
rect -3000 4603 -2976 4637
rect -3058 4565 -2976 4603
rect -3058 4531 -3034 4565
rect -3000 4531 -2976 4565
rect -3058 4493 -2976 4531
rect -3058 4459 -3034 4493
rect -3000 4459 -2976 4493
rect -3058 4421 -2976 4459
rect -3058 4387 -3034 4421
rect -3000 4387 -2976 4421
rect -3058 4349 -2976 4387
rect -3058 4315 -3034 4349
rect -3000 4315 -2976 4349
rect -3058 4277 -2976 4315
rect -3058 4243 -3034 4277
rect -3000 4243 -2976 4277
rect -3058 4205 -2976 4243
rect -3058 4171 -3034 4205
rect -3000 4171 -2976 4205
rect -3058 4133 -2976 4171
rect -3058 4099 -3034 4133
rect -3000 4099 -2976 4133
rect -3058 4061 -2976 4099
rect -3058 4027 -3034 4061
rect -3000 4027 -2976 4061
rect -3058 3989 -2976 4027
rect -3058 3955 -3034 3989
rect -3000 3955 -2976 3989
rect -3058 3917 -2976 3955
rect -3058 3883 -3034 3917
rect -3000 3883 -2976 3917
rect -3058 3845 -2976 3883
rect -3058 3811 -3034 3845
rect -3000 3811 -2976 3845
rect -3058 3773 -2976 3811
rect -3058 3739 -3034 3773
rect -3000 3739 -2976 3773
rect -3058 3701 -2976 3739
rect -3058 3667 -3034 3701
rect -3000 3667 -2976 3701
rect -3058 3629 -2976 3667
rect -3058 3595 -3034 3629
rect -3000 3595 -2976 3629
rect -3058 3557 -2976 3595
rect -3058 3523 -3034 3557
rect -3000 3523 -2976 3557
rect -3058 3485 -2976 3523
rect -3058 3451 -3034 3485
rect -3000 3451 -2976 3485
rect -3058 3413 -2976 3451
rect -3058 3379 -3034 3413
rect -3000 3379 -2976 3413
rect -3058 3341 -2976 3379
rect -3058 3307 -3034 3341
rect -3000 3307 -2976 3341
rect -3058 3269 -2976 3307
rect -3058 3235 -3034 3269
rect -3000 3235 -2976 3269
rect -3058 3197 -2976 3235
rect -3058 3163 -3034 3197
rect -3000 3163 -2976 3197
rect -3058 3125 -2976 3163
rect -3058 3091 -3034 3125
rect -3000 3091 -2976 3125
rect -3058 3053 -2976 3091
rect -3058 3019 -3034 3053
rect -3000 3019 -2976 3053
rect -3058 2981 -2976 3019
rect -3058 2947 -3034 2981
rect -3000 2947 -2976 2981
rect -3058 2909 -2976 2947
rect -3058 2875 -3034 2909
rect -3000 2875 -2976 2909
rect -3058 2837 -2976 2875
rect -3058 2803 -3034 2837
rect -3000 2803 -2976 2837
rect -3058 2765 -2976 2803
rect -3058 2731 -3034 2765
rect -3000 2731 -2976 2765
rect -3058 2693 -2976 2731
rect -3058 2659 -3034 2693
rect -3000 2659 -2976 2693
rect -3058 2621 -2976 2659
rect -3058 2587 -3034 2621
rect -3000 2587 -2976 2621
rect -3058 2549 -2976 2587
rect -3058 2515 -3034 2549
rect -3000 2515 -2976 2549
rect -3058 2477 -2976 2515
rect -3058 2443 -3034 2477
rect -3000 2443 -2976 2477
rect -3058 2405 -2976 2443
rect -3058 2371 -3034 2405
rect -3000 2371 -2976 2405
rect -3058 2333 -2976 2371
rect -3058 2299 -3034 2333
rect -3000 2299 -2976 2333
rect -3058 2261 -2976 2299
rect -3058 2227 -3034 2261
rect -3000 2227 -2976 2261
rect -3058 2189 -2976 2227
rect -3058 2155 -3034 2189
rect -3000 2155 -2976 2189
rect -3058 2117 -2976 2155
rect -3058 2083 -3034 2117
rect -3000 2083 -2976 2117
rect -3058 2045 -2976 2083
rect -3058 2011 -3034 2045
rect -3000 2011 -2976 2045
rect -3058 1973 -2976 2011
rect -3058 1939 -3034 1973
rect -3000 1939 -2976 1973
rect -3058 1901 -2976 1939
rect -3058 1867 -3034 1901
rect -3000 1867 -2976 1901
rect -3058 1829 -2976 1867
rect -3058 1795 -3034 1829
rect -3000 1795 -2976 1829
rect -3058 1757 -2976 1795
rect -3058 1723 -3034 1757
rect -3000 1723 -2976 1757
rect -3058 1685 -2976 1723
rect -3058 1651 -3034 1685
rect -3000 1651 -2976 1685
rect -3058 1613 -2976 1651
rect -3058 1579 -3034 1613
rect -3000 1579 -2976 1613
rect -3058 1541 -2976 1579
rect -3058 1507 -3034 1541
rect -3000 1507 -2976 1541
rect -3058 1469 -2976 1507
rect -3058 1435 -3034 1469
rect -3000 1435 -2976 1469
rect -3058 1397 -2976 1435
rect -3058 1363 -3034 1397
rect -3000 1363 -2976 1397
rect -3058 1325 -2976 1363
rect -3058 1291 -3034 1325
rect -3000 1291 -2976 1325
rect -3058 1253 -2976 1291
rect -3058 1219 -3034 1253
rect -3000 1219 -2976 1253
rect -3058 1181 -2976 1219
rect -3058 1147 -3034 1181
rect -3000 1147 -2976 1181
rect -3058 1109 -2976 1147
rect -3058 1075 -3034 1109
rect -3000 1075 -2976 1109
rect -3058 1037 -2976 1075
rect -3058 1003 -3034 1037
rect -3000 1003 -2976 1037
rect -3058 965 -2976 1003
rect -3058 931 -3034 965
rect -3000 931 -2976 965
rect -3058 893 -2976 931
rect -3058 859 -3034 893
rect -3000 859 -2976 893
rect -3058 821 -2976 859
rect -3058 787 -3034 821
rect -3000 787 -2976 821
rect -3058 749 -2976 787
rect -3058 715 -3034 749
rect -3000 715 -2976 749
rect -3058 677 -2976 715
rect -3058 643 -3034 677
rect -3000 643 -2976 677
rect -3058 605 -2976 643
rect -3058 571 -3034 605
rect -3000 571 -2976 605
rect -3058 533 -2976 571
rect -3058 499 -3034 533
rect -3000 499 -2976 533
rect -3058 461 -2976 499
rect -3058 427 -3034 461
rect -3000 427 -2976 461
rect -3058 389 -2976 427
rect -3058 355 -3034 389
rect -3000 355 -2976 389
rect -3058 317 -2976 355
rect -3058 283 -3034 317
rect -3000 283 -2976 317
rect -3058 245 -2976 283
rect -3058 211 -3034 245
rect -3000 211 -2976 245
rect -3058 173 -2976 211
rect -3058 139 -3034 173
rect -3000 139 -2976 173
rect -3058 101 -2976 139
rect -3058 67 -3034 101
rect -3000 67 -2976 101
rect -3058 29 -2976 67
rect -3058 -5 -3034 29
rect -3000 -5 -2976 29
rect -1068 5969 -934 5991
rect -1068 31 -1054 5969
rect -948 31 -934 5969
rect -1068 9 -934 31
rect -830 5969 -696 5991
rect -830 31 -816 5969
rect -710 31 -696 5969
rect 996 5969 1130 5991
rect 15 5933 285 5957
rect 15 67 25 5933
rect 275 67 285 5933
rect 15 43 285 67
rect -830 9 -696 31
rect 996 31 1010 5969
rect 1116 31 1130 5969
rect 996 9 1130 31
rect 1234 5969 1368 5991
rect 1234 31 1248 5969
rect 1354 31 1368 5969
rect 1234 9 1368 31
rect 3276 5971 3300 6005
rect 3334 5971 3358 6005
rect 3276 5933 3358 5971
rect 3276 5899 3300 5933
rect 3334 5899 3358 5933
rect 3276 5861 3358 5899
rect 3276 5827 3300 5861
rect 3334 5827 3358 5861
rect 3276 5789 3358 5827
rect 3276 5755 3300 5789
rect 3334 5755 3358 5789
rect 3276 5717 3358 5755
rect 3276 5683 3300 5717
rect 3334 5683 3358 5717
rect 3276 5645 3358 5683
rect 3276 5611 3300 5645
rect 3334 5611 3358 5645
rect 3276 5573 3358 5611
rect 3276 5539 3300 5573
rect 3334 5539 3358 5573
rect 3276 5501 3358 5539
rect 3276 5467 3300 5501
rect 3334 5467 3358 5501
rect 3276 5429 3358 5467
rect 3276 5395 3300 5429
rect 3334 5395 3358 5429
rect 3276 5357 3358 5395
rect 3276 5323 3300 5357
rect 3334 5323 3358 5357
rect 3276 5285 3358 5323
rect 3276 5251 3300 5285
rect 3334 5251 3358 5285
rect 3276 5213 3358 5251
rect 3276 5179 3300 5213
rect 3334 5179 3358 5213
rect 3276 5141 3358 5179
rect 3276 5107 3300 5141
rect 3334 5107 3358 5141
rect 3276 5069 3358 5107
rect 3276 5035 3300 5069
rect 3334 5035 3358 5069
rect 3276 4997 3358 5035
rect 3276 4963 3300 4997
rect 3334 4963 3358 4997
rect 3276 4925 3358 4963
rect 3276 4891 3300 4925
rect 3334 4891 3358 4925
rect 3276 4853 3358 4891
rect 3276 4819 3300 4853
rect 3334 4819 3358 4853
rect 3276 4781 3358 4819
rect 3276 4747 3300 4781
rect 3334 4747 3358 4781
rect 3276 4709 3358 4747
rect 3276 4675 3300 4709
rect 3334 4675 3358 4709
rect 3276 4637 3358 4675
rect 3276 4603 3300 4637
rect 3334 4603 3358 4637
rect 3276 4565 3358 4603
rect 3276 4531 3300 4565
rect 3334 4531 3358 4565
rect 3276 4493 3358 4531
rect 3276 4459 3300 4493
rect 3334 4459 3358 4493
rect 3276 4421 3358 4459
rect 3276 4387 3300 4421
rect 3334 4387 3358 4421
rect 3276 4349 3358 4387
rect 3276 4315 3300 4349
rect 3334 4315 3358 4349
rect 3276 4277 3358 4315
rect 3276 4243 3300 4277
rect 3334 4243 3358 4277
rect 3276 4205 3358 4243
rect 3276 4171 3300 4205
rect 3334 4171 3358 4205
rect 3276 4133 3358 4171
rect 3276 4099 3300 4133
rect 3334 4099 3358 4133
rect 3276 4061 3358 4099
rect 3276 4027 3300 4061
rect 3334 4027 3358 4061
rect 3276 3989 3358 4027
rect 3276 3955 3300 3989
rect 3334 3955 3358 3989
rect 3276 3917 3358 3955
rect 3276 3883 3300 3917
rect 3334 3883 3358 3917
rect 3276 3845 3358 3883
rect 3276 3811 3300 3845
rect 3334 3811 3358 3845
rect 3276 3773 3358 3811
rect 3276 3739 3300 3773
rect 3334 3739 3358 3773
rect 3276 3701 3358 3739
rect 3276 3667 3300 3701
rect 3334 3667 3358 3701
rect 3276 3629 3358 3667
rect 3276 3595 3300 3629
rect 3334 3595 3358 3629
rect 3276 3557 3358 3595
rect 3276 3523 3300 3557
rect 3334 3523 3358 3557
rect 3276 3485 3358 3523
rect 3276 3451 3300 3485
rect 3334 3451 3358 3485
rect 3276 3413 3358 3451
rect 3276 3379 3300 3413
rect 3334 3379 3358 3413
rect 3276 3341 3358 3379
rect 3276 3307 3300 3341
rect 3334 3307 3358 3341
rect 3276 3269 3358 3307
rect 3276 3235 3300 3269
rect 3334 3235 3358 3269
rect 3276 3197 3358 3235
rect 3276 3163 3300 3197
rect 3334 3163 3358 3197
rect 3276 3125 3358 3163
rect 3276 3091 3300 3125
rect 3334 3091 3358 3125
rect 3276 3053 3358 3091
rect 3276 3019 3300 3053
rect 3334 3019 3358 3053
rect 3276 2981 3358 3019
rect 3276 2947 3300 2981
rect 3334 2947 3358 2981
rect 3276 2909 3358 2947
rect 3276 2875 3300 2909
rect 3334 2875 3358 2909
rect 3276 2837 3358 2875
rect 3276 2803 3300 2837
rect 3334 2803 3358 2837
rect 3276 2765 3358 2803
rect 3276 2731 3300 2765
rect 3334 2731 3358 2765
rect 3276 2693 3358 2731
rect 3276 2659 3300 2693
rect 3334 2659 3358 2693
rect 3276 2621 3358 2659
rect 3276 2587 3300 2621
rect 3334 2587 3358 2621
rect 3276 2549 3358 2587
rect 3276 2515 3300 2549
rect 3334 2515 3358 2549
rect 3276 2477 3358 2515
rect 3276 2443 3300 2477
rect 3334 2443 3358 2477
rect 3276 2405 3358 2443
rect 3276 2371 3300 2405
rect 3334 2371 3358 2405
rect 3276 2333 3358 2371
rect 3276 2299 3300 2333
rect 3334 2299 3358 2333
rect 3276 2261 3358 2299
rect 3276 2227 3300 2261
rect 3334 2227 3358 2261
rect 3276 2189 3358 2227
rect 3276 2155 3300 2189
rect 3334 2155 3358 2189
rect 3276 2117 3358 2155
rect 3276 2083 3300 2117
rect 3334 2083 3358 2117
rect 3276 2045 3358 2083
rect 3276 2011 3300 2045
rect 3334 2011 3358 2045
rect 3276 1973 3358 2011
rect 3276 1939 3300 1973
rect 3334 1939 3358 1973
rect 3276 1901 3358 1939
rect 3276 1867 3300 1901
rect 3334 1867 3358 1901
rect 3276 1829 3358 1867
rect 3276 1795 3300 1829
rect 3334 1795 3358 1829
rect 3276 1757 3358 1795
rect 3276 1723 3300 1757
rect 3334 1723 3358 1757
rect 3276 1685 3358 1723
rect 3276 1651 3300 1685
rect 3334 1651 3358 1685
rect 3276 1613 3358 1651
rect 3276 1579 3300 1613
rect 3334 1579 3358 1613
rect 3276 1541 3358 1579
rect 3276 1507 3300 1541
rect 3334 1507 3358 1541
rect 3276 1469 3358 1507
rect 3276 1435 3300 1469
rect 3334 1435 3358 1469
rect 3276 1397 3358 1435
rect 3276 1363 3300 1397
rect 3334 1363 3358 1397
rect 3276 1325 3358 1363
rect 3276 1291 3300 1325
rect 3334 1291 3358 1325
rect 3276 1253 3358 1291
rect 3276 1219 3300 1253
rect 3334 1219 3358 1253
rect 3276 1181 3358 1219
rect 3276 1147 3300 1181
rect 3334 1147 3358 1181
rect 3276 1109 3358 1147
rect 3276 1075 3300 1109
rect 3334 1075 3358 1109
rect 3276 1037 3358 1075
rect 3276 1003 3300 1037
rect 3334 1003 3358 1037
rect 3276 965 3358 1003
rect 3276 931 3300 965
rect 3334 931 3358 965
rect 3276 893 3358 931
rect 3276 859 3300 893
rect 3334 859 3358 893
rect 3276 821 3358 859
rect 3276 787 3300 821
rect 3334 787 3358 821
rect 3276 749 3358 787
rect 3276 715 3300 749
rect 3334 715 3358 749
rect 3276 677 3358 715
rect 3276 643 3300 677
rect 3334 643 3358 677
rect 3276 605 3358 643
rect 3276 571 3300 605
rect 3334 571 3358 605
rect 3276 533 3358 571
rect 3276 499 3300 533
rect 3334 499 3358 533
rect 3276 461 3358 499
rect 3276 427 3300 461
rect 3334 427 3358 461
rect 3276 389 3358 427
rect 3276 355 3300 389
rect 3334 355 3358 389
rect 3276 317 3358 355
rect 3276 283 3300 317
rect 3334 283 3358 317
rect 3276 245 3358 283
rect 3276 211 3300 245
rect 3334 211 3358 245
rect 3276 173 3358 211
rect 3276 139 3300 173
rect 3334 139 3358 173
rect 3276 101 3358 139
rect 3276 67 3300 101
rect 3334 67 3358 101
rect 3276 29 3358 67
rect -3058 -43 -2976 -5
rect -3058 -77 -3034 -43
rect -3000 -77 -2976 -43
rect -3058 -115 -2976 -77
rect -3058 -149 -3034 -115
rect -3000 -149 -2976 -115
rect -3058 -187 -2976 -149
rect -3058 -221 -3034 -187
rect -3000 -221 -2976 -187
rect -3058 -259 -2976 -221
rect -3058 -293 -3034 -259
rect -3000 -293 -2976 -259
rect -3058 -331 -2976 -293
rect -3058 -365 -3034 -331
rect -3000 -365 -2976 -331
rect -3058 -403 -2976 -365
rect -3058 -437 -3034 -403
rect -3000 -437 -2976 -403
rect -3058 -475 -2976 -437
rect 3276 -5 3300 29
rect 3334 -5 3358 29
rect 3276 -43 3358 -5
rect 3276 -77 3300 -43
rect 3334 -77 3358 -43
rect 3276 -115 3358 -77
rect 3276 -149 3300 -115
rect 3334 -149 3358 -115
rect 3276 -187 3358 -149
rect 3276 -221 3300 -187
rect 3334 -221 3358 -187
rect 3276 -259 3358 -221
rect 3276 -293 3300 -259
rect 3334 -293 3358 -259
rect 3276 -331 3358 -293
rect 3276 -365 3300 -331
rect 3334 -365 3358 -331
rect 3276 -403 3358 -365
rect 3276 -437 3300 -403
rect 3334 -437 3358 -403
rect -3058 -509 -3034 -475
rect -3000 -509 -2976 -475
rect -3058 -547 -2976 -509
rect -3058 -581 -3034 -547
rect -3000 -581 -2976 -547
rect -3058 -619 -2976 -581
rect -3058 -653 -3034 -619
rect -3000 -653 -2976 -619
rect -3058 -691 -2976 -653
rect -209 -459 555 -443
rect -209 -493 -180 -459
rect -146 -493 -106 -459
rect -72 -493 -32 -459
rect 2 -493 42 -459
rect 76 -493 116 -459
rect 150 -493 190 -459
rect 224 -493 264 -459
rect 298 -493 338 -459
rect 372 -493 412 -459
rect 446 -493 486 -459
rect 520 -493 555 -459
rect -209 -533 555 -493
rect -209 -567 -180 -533
rect -146 -567 -106 -533
rect -72 -567 -32 -533
rect 2 -567 42 -533
rect 76 -567 116 -533
rect 150 -567 190 -533
rect 224 -567 264 -533
rect 298 -567 338 -533
rect 372 -567 412 -533
rect 446 -567 486 -533
rect 520 -567 555 -533
rect -209 -607 555 -567
rect -209 -641 -180 -607
rect -146 -641 -106 -607
rect -72 -641 -32 -607
rect 2 -641 42 -607
rect 76 -641 116 -607
rect 150 -641 190 -607
rect 224 -641 264 -607
rect 298 -641 338 -607
rect 372 -641 412 -607
rect 446 -641 486 -607
rect 520 -641 555 -607
rect -209 -657 555 -641
rect 3276 -475 3358 -437
rect 3276 -509 3300 -475
rect 3334 -509 3358 -475
rect 3276 -547 3358 -509
rect 3276 -581 3300 -547
rect 3334 -581 3358 -547
rect 3276 -619 3358 -581
rect 3276 -653 3300 -619
rect 3334 -653 3358 -619
rect -3058 -725 -3034 -691
rect -3000 -725 -2976 -691
rect -3058 -763 -2976 -725
rect -3058 -797 -3034 -763
rect -3000 -797 -2976 -763
rect -3058 -835 -2976 -797
rect -3058 -869 -3034 -835
rect -3000 -869 -2976 -835
rect -3058 -907 -2976 -869
rect -3058 -941 -3034 -907
rect -3000 -941 -2976 -907
rect -3058 -979 -2976 -941
rect -3058 -1013 -3034 -979
rect -3000 -1013 -2976 -979
rect -3058 -1051 -2976 -1013
rect -3058 -1085 -3034 -1051
rect -3000 -1085 -2976 -1051
rect -3058 -1123 -2976 -1085
rect -3058 -1157 -3034 -1123
rect -3000 -1157 -2976 -1123
rect -3058 -1195 -2976 -1157
rect -3058 -1229 -3034 -1195
rect -3000 -1229 -2976 -1195
rect -3058 -1267 -2976 -1229
rect -3058 -1301 -3034 -1267
rect -3000 -1301 -2976 -1267
rect -3058 -1339 -2976 -1301
rect -3058 -1373 -3034 -1339
rect -3000 -1373 -2976 -1339
rect -3058 -1411 -2976 -1373
rect -3058 -1445 -3034 -1411
rect -3000 -1445 -2976 -1411
rect -3058 -1483 -2976 -1445
rect -3058 -1517 -3034 -1483
rect -3000 -1517 -2976 -1483
rect -3058 -1555 -2976 -1517
rect -3058 -1589 -3034 -1555
rect -3000 -1589 -2976 -1555
rect -3058 -1627 -2976 -1589
rect -3058 -1661 -3034 -1627
rect -3000 -1661 -2976 -1627
rect -3058 -1699 -2976 -1661
rect -3058 -1733 -3034 -1699
rect -3000 -1733 -2976 -1699
rect -3058 -1771 -2976 -1733
rect -3058 -1805 -3034 -1771
rect -3000 -1805 -2976 -1771
rect -3058 -1843 -2976 -1805
rect -3058 -1877 -3034 -1843
rect -3000 -1877 -2976 -1843
rect -3058 -1900 -2976 -1877
rect 3276 -691 3358 -653
rect 3276 -725 3300 -691
rect 3334 -725 3358 -691
rect 3276 -763 3358 -725
rect 3276 -797 3300 -763
rect 3334 -797 3358 -763
rect 3276 -835 3358 -797
rect 3276 -869 3300 -835
rect 3334 -869 3358 -835
rect 3276 -907 3358 -869
rect 3276 -941 3300 -907
rect 3334 -941 3358 -907
rect 3276 -979 3358 -941
rect 3276 -1013 3300 -979
rect 3334 -1013 3358 -979
rect 3276 -1051 3358 -1013
rect 3276 -1085 3300 -1051
rect 3334 -1085 3358 -1051
rect 3276 -1123 3358 -1085
rect 3276 -1157 3300 -1123
rect 3334 -1157 3358 -1123
rect 3276 -1195 3358 -1157
rect 3276 -1229 3300 -1195
rect 3334 -1229 3358 -1195
rect 3276 -1267 3358 -1229
rect 3276 -1301 3300 -1267
rect 3334 -1301 3358 -1267
rect 3276 -1339 3358 -1301
rect 3276 -1373 3300 -1339
rect 3334 -1373 3358 -1339
rect 3276 -1411 3358 -1373
rect 3276 -1445 3300 -1411
rect 3334 -1445 3358 -1411
rect 3276 -1483 3358 -1445
rect 3276 -1517 3300 -1483
rect 3334 -1517 3358 -1483
rect 3276 -1555 3358 -1517
rect 3276 -1589 3300 -1555
rect 3334 -1589 3358 -1555
rect 3276 -1627 3358 -1589
rect 3276 -1661 3300 -1627
rect 3334 -1661 3358 -1627
rect 3276 -1699 3358 -1661
rect 3276 -1733 3300 -1699
rect 3334 -1733 3358 -1699
rect 3276 -1771 3358 -1733
rect 3276 -1805 3300 -1771
rect 3334 -1805 3358 -1771
rect 3276 -1843 3358 -1805
rect 3276 -1877 3300 -1843
rect 3334 -1877 3358 -1843
rect 3276 -1900 3358 -1877
rect -3058 -1924 3358 -1900
rect -3058 -1958 -2927 -1924
rect -2893 -1958 -2855 -1924
rect -2821 -1958 -2783 -1924
rect -2749 -1958 -2711 -1924
rect -2677 -1958 -2639 -1924
rect -2605 -1958 -2567 -1924
rect -2533 -1958 -2495 -1924
rect -2461 -1958 -2423 -1924
rect -2389 -1958 -2351 -1924
rect -2317 -1958 -2279 -1924
rect -2245 -1958 -2207 -1924
rect -2173 -1958 -2135 -1924
rect -2101 -1958 -2063 -1924
rect -2029 -1958 -1991 -1924
rect -1957 -1958 -1919 -1924
rect -1885 -1958 -1847 -1924
rect -1813 -1958 -1775 -1924
rect -1741 -1958 -1703 -1924
rect -1669 -1958 -1631 -1924
rect -1597 -1958 -1559 -1924
rect -1525 -1958 -1487 -1924
rect -1453 -1958 -1415 -1924
rect -1381 -1958 -1343 -1924
rect -1309 -1958 -1271 -1924
rect -1237 -1958 -1199 -1924
rect -1165 -1958 -1127 -1924
rect -1093 -1958 -1055 -1924
rect -1021 -1958 -983 -1924
rect -949 -1958 -911 -1924
rect -877 -1958 -839 -1924
rect -805 -1958 -767 -1924
rect -733 -1958 -695 -1924
rect -661 -1958 -623 -1924
rect -589 -1958 -551 -1924
rect -517 -1958 -479 -1924
rect -445 -1958 -407 -1924
rect -373 -1958 -335 -1924
rect -301 -1958 -263 -1924
rect -229 -1958 -191 -1924
rect -157 -1958 -119 -1924
rect -85 -1958 -47 -1924
rect -13 -1958 25 -1924
rect 59 -1958 97 -1924
rect 131 -1958 169 -1924
rect 203 -1958 241 -1924
rect 275 -1958 313 -1924
rect 347 -1958 385 -1924
rect 419 -1958 457 -1924
rect 491 -1958 529 -1924
rect 563 -1958 601 -1924
rect 635 -1958 673 -1924
rect 707 -1958 745 -1924
rect 779 -1958 817 -1924
rect 851 -1958 889 -1924
rect 923 -1958 961 -1924
rect 995 -1958 1033 -1924
rect 1067 -1958 1105 -1924
rect 1139 -1958 1177 -1924
rect 1211 -1958 1249 -1924
rect 1283 -1958 1321 -1924
rect 1355 -1958 1393 -1924
rect 1427 -1958 1465 -1924
rect 1499 -1958 1537 -1924
rect 1571 -1958 1609 -1924
rect 1643 -1958 1681 -1924
rect 1715 -1958 1753 -1924
rect 1787 -1958 1825 -1924
rect 1859 -1958 1897 -1924
rect 1931 -1958 1969 -1924
rect 2003 -1958 2041 -1924
rect 2075 -1958 2113 -1924
rect 2147 -1958 2185 -1924
rect 2219 -1958 2257 -1924
rect 2291 -1958 2329 -1924
rect 2363 -1958 2401 -1924
rect 2435 -1958 2473 -1924
rect 2507 -1958 2545 -1924
rect 2579 -1958 2617 -1924
rect 2651 -1958 2689 -1924
rect 2723 -1958 2761 -1924
rect 2795 -1958 2833 -1924
rect 2867 -1958 2905 -1924
rect 2939 -1958 2977 -1924
rect 3011 -1958 3049 -1924
rect 3083 -1958 3121 -1924
rect 3155 -1958 3193 -1924
rect 3227 -1958 3358 -1924
rect -3058 -1982 3358 -1958
<< viali >>
rect -2927 7925 -2893 7959
rect -2855 7925 -2821 7959
rect -2783 7925 -2749 7959
rect -2711 7925 -2677 7959
rect -2639 7925 -2605 7959
rect -2567 7925 -2533 7959
rect -2495 7925 -2461 7959
rect -2423 7925 -2389 7959
rect -2351 7925 -2317 7959
rect -2279 7925 -2245 7959
rect -2207 7925 -2173 7959
rect -2135 7925 -2101 7959
rect -2063 7925 -2029 7959
rect -1991 7925 -1957 7959
rect -1919 7925 -1885 7959
rect -1847 7925 -1813 7959
rect -1775 7925 -1741 7959
rect -1703 7925 -1669 7959
rect -1631 7925 -1597 7959
rect -1559 7925 -1525 7959
rect -1487 7925 -1453 7959
rect -1415 7925 -1381 7959
rect -1343 7925 -1309 7959
rect -1271 7925 -1237 7959
rect -1199 7925 -1165 7959
rect -1127 7925 -1093 7959
rect -1055 7925 -1021 7959
rect -983 7925 -949 7959
rect -911 7925 -877 7959
rect -839 7925 -805 7959
rect -767 7925 -733 7959
rect -695 7925 -661 7959
rect -623 7925 -589 7959
rect -551 7925 -517 7959
rect -479 7925 -445 7959
rect -407 7925 -373 7959
rect -335 7925 -301 7959
rect -263 7925 -229 7959
rect -191 7925 -157 7959
rect -119 7925 -85 7959
rect -47 7925 -13 7959
rect 25 7925 59 7959
rect 97 7925 131 7959
rect 169 7925 203 7959
rect 241 7925 275 7959
rect 313 7925 347 7959
rect 385 7925 419 7959
rect 457 7925 491 7959
rect 529 7925 563 7959
rect 601 7925 635 7959
rect 673 7925 707 7959
rect 745 7925 779 7959
rect 817 7925 851 7959
rect 889 7925 923 7959
rect 961 7925 995 7959
rect 1033 7925 1067 7959
rect 1105 7925 1139 7959
rect 1177 7925 1211 7959
rect 1249 7925 1283 7959
rect 1321 7925 1355 7959
rect 1393 7925 1427 7959
rect 1465 7925 1499 7959
rect 1537 7925 1571 7959
rect 1609 7925 1643 7959
rect 1681 7925 1715 7959
rect 1753 7925 1787 7959
rect 1825 7925 1859 7959
rect 1897 7925 1931 7959
rect 1969 7925 2003 7959
rect 2041 7925 2075 7959
rect 2113 7925 2147 7959
rect 2185 7925 2219 7959
rect 2257 7925 2291 7959
rect 2329 7925 2363 7959
rect 2401 7925 2435 7959
rect 2473 7925 2507 7959
rect 2545 7925 2579 7959
rect 2617 7925 2651 7959
rect 2689 7925 2723 7959
rect 2761 7925 2795 7959
rect 2833 7925 2867 7959
rect 2905 7925 2939 7959
rect 2977 7925 3011 7959
rect 3049 7925 3083 7959
rect 3121 7925 3155 7959
rect 3193 7925 3227 7959
rect -3034 7843 -3000 7877
rect -3034 7771 -3000 7805
rect -3034 7699 -3000 7733
rect -3034 7627 -3000 7661
rect -3034 7555 -3000 7589
rect -3034 7483 -3000 7517
rect -3034 7411 -3000 7445
rect -3034 7339 -3000 7373
rect -3034 7267 -3000 7301
rect -3034 7195 -3000 7229
rect -3034 7123 -3000 7157
rect -3034 7051 -3000 7085
rect -3034 6979 -3000 7013
rect -3034 6907 -3000 6941
rect -3034 6835 -3000 6869
rect -3034 6763 -3000 6797
rect -3034 6691 -3000 6725
rect -3034 6619 -3000 6653
rect -3034 6547 -3000 6581
rect -3034 6475 -3000 6509
rect -3034 6403 -3000 6437
rect -3034 6331 -3000 6365
rect -3034 6259 -3000 6293
rect -3034 6187 -3000 6221
rect -3034 6115 -3000 6149
rect -3034 6043 -3000 6077
rect -3034 5971 -3000 6005
rect 3300 7843 3334 7877
rect 3300 7771 3334 7805
rect 3300 7699 3334 7733
rect 3300 7627 3334 7661
rect 3300 7555 3334 7589
rect 3300 7483 3334 7517
rect 3300 7411 3334 7445
rect 3300 7339 3334 7373
rect 3300 7267 3334 7301
rect 3300 7195 3334 7229
rect 3300 7123 3334 7157
rect 3300 7051 3334 7085
rect 3300 6979 3334 7013
rect 3300 6907 3334 6941
rect 3300 6835 3334 6869
rect 3300 6763 3334 6797
rect 3300 6691 3334 6725
rect 3300 6619 3334 6653
rect 3300 6547 3334 6581
rect 3300 6475 3334 6509
rect 3300 6403 3334 6437
rect 3300 6331 3334 6365
rect 3300 6259 3334 6293
rect 3300 6187 3334 6221
rect 3300 6115 3334 6149
rect 3300 6043 3334 6077
rect -3034 5899 -3000 5933
rect -3034 5827 -3000 5861
rect -3034 5755 -3000 5789
rect -3034 5683 -3000 5717
rect -3034 5611 -3000 5645
rect -3034 5539 -3000 5573
rect -3034 5467 -3000 5501
rect -3034 5395 -3000 5429
rect -3034 5323 -3000 5357
rect -3034 5251 -3000 5285
rect -3034 5179 -3000 5213
rect -3034 5107 -3000 5141
rect -3034 5035 -3000 5069
rect -3034 4963 -3000 4997
rect -3034 4891 -3000 4925
rect -3034 4819 -3000 4853
rect -3034 4747 -3000 4781
rect -3034 4675 -3000 4709
rect -3034 4603 -3000 4637
rect -3034 4531 -3000 4565
rect -3034 4459 -3000 4493
rect -3034 4387 -3000 4421
rect -3034 4315 -3000 4349
rect -3034 4243 -3000 4277
rect -3034 4171 -3000 4205
rect -3034 4099 -3000 4133
rect -3034 4027 -3000 4061
rect -3034 3955 -3000 3989
rect -3034 3883 -3000 3917
rect -3034 3811 -3000 3845
rect -3034 3739 -3000 3773
rect -3034 3667 -3000 3701
rect -3034 3595 -3000 3629
rect -3034 3523 -3000 3557
rect -3034 3451 -3000 3485
rect -3034 3379 -3000 3413
rect -3034 3307 -3000 3341
rect -3034 3235 -3000 3269
rect -3034 3163 -3000 3197
rect -3034 3091 -3000 3125
rect -3034 3019 -3000 3053
rect -3034 2947 -3000 2981
rect -3034 2875 -3000 2909
rect -3034 2803 -3000 2837
rect -3034 2731 -3000 2765
rect -3034 2659 -3000 2693
rect -3034 2587 -3000 2621
rect -3034 2515 -3000 2549
rect -3034 2443 -3000 2477
rect -3034 2371 -3000 2405
rect -3034 2299 -3000 2333
rect -3034 2227 -3000 2261
rect -3034 2155 -3000 2189
rect -3034 2083 -3000 2117
rect -3034 2011 -3000 2045
rect -3034 1939 -3000 1973
rect -3034 1867 -3000 1901
rect -3034 1795 -3000 1829
rect -3034 1723 -3000 1757
rect -3034 1651 -3000 1685
rect -3034 1579 -3000 1613
rect -3034 1507 -3000 1541
rect -3034 1435 -3000 1469
rect -3034 1363 -3000 1397
rect -3034 1291 -3000 1325
rect -3034 1219 -3000 1253
rect -3034 1147 -3000 1181
rect -3034 1075 -3000 1109
rect -3034 1003 -3000 1037
rect -3034 931 -3000 965
rect -3034 859 -3000 893
rect -3034 787 -3000 821
rect -3034 715 -3000 749
rect -3034 643 -3000 677
rect -3034 571 -3000 605
rect -3034 499 -3000 533
rect -3034 427 -3000 461
rect -3034 355 -3000 389
rect -3034 283 -3000 317
rect -3034 211 -3000 245
rect -3034 139 -3000 173
rect -3034 67 -3000 101
rect -3034 -5 -3000 29
rect -1054 31 -948 5969
rect -816 31 -710 5969
rect 25 67 275 5933
rect 1010 31 1116 5969
rect 1248 31 1354 5969
rect 3300 5971 3334 6005
rect 3300 5899 3334 5933
rect 3300 5827 3334 5861
rect 3300 5755 3334 5789
rect 3300 5683 3334 5717
rect 3300 5611 3334 5645
rect 3300 5539 3334 5573
rect 3300 5467 3334 5501
rect 3300 5395 3334 5429
rect 3300 5323 3334 5357
rect 3300 5251 3334 5285
rect 3300 5179 3334 5213
rect 3300 5107 3334 5141
rect 3300 5035 3334 5069
rect 3300 4963 3334 4997
rect 3300 4891 3334 4925
rect 3300 4819 3334 4853
rect 3300 4747 3334 4781
rect 3300 4675 3334 4709
rect 3300 4603 3334 4637
rect 3300 4531 3334 4565
rect 3300 4459 3334 4493
rect 3300 4387 3334 4421
rect 3300 4315 3334 4349
rect 3300 4243 3334 4277
rect 3300 4171 3334 4205
rect 3300 4099 3334 4133
rect 3300 4027 3334 4061
rect 3300 3955 3334 3989
rect 3300 3883 3334 3917
rect 3300 3811 3334 3845
rect 3300 3739 3334 3773
rect 3300 3667 3334 3701
rect 3300 3595 3334 3629
rect 3300 3523 3334 3557
rect 3300 3451 3334 3485
rect 3300 3379 3334 3413
rect 3300 3307 3334 3341
rect 3300 3235 3334 3269
rect 3300 3163 3334 3197
rect 3300 3091 3334 3125
rect 3300 3019 3334 3053
rect 3300 2947 3334 2981
rect 3300 2875 3334 2909
rect 3300 2803 3334 2837
rect 3300 2731 3334 2765
rect 3300 2659 3334 2693
rect 3300 2587 3334 2621
rect 3300 2515 3334 2549
rect 3300 2443 3334 2477
rect 3300 2371 3334 2405
rect 3300 2299 3334 2333
rect 3300 2227 3334 2261
rect 3300 2155 3334 2189
rect 3300 2083 3334 2117
rect 3300 2011 3334 2045
rect 3300 1939 3334 1973
rect 3300 1867 3334 1901
rect 3300 1795 3334 1829
rect 3300 1723 3334 1757
rect 3300 1651 3334 1685
rect 3300 1579 3334 1613
rect 3300 1507 3334 1541
rect 3300 1435 3334 1469
rect 3300 1363 3334 1397
rect 3300 1291 3334 1325
rect 3300 1219 3334 1253
rect 3300 1147 3334 1181
rect 3300 1075 3334 1109
rect 3300 1003 3334 1037
rect 3300 931 3334 965
rect 3300 859 3334 893
rect 3300 787 3334 821
rect 3300 715 3334 749
rect 3300 643 3334 677
rect 3300 571 3334 605
rect 3300 499 3334 533
rect 3300 427 3334 461
rect 3300 355 3334 389
rect 3300 283 3334 317
rect 3300 211 3334 245
rect 3300 139 3334 173
rect 3300 67 3334 101
rect -3034 -77 -3000 -43
rect -3034 -149 -3000 -115
rect -3034 -221 -3000 -187
rect -3034 -293 -3000 -259
rect -3034 -365 -3000 -331
rect -3034 -437 -3000 -403
rect 3300 -5 3334 29
rect 3300 -77 3334 -43
rect 3300 -149 3334 -115
rect 3300 -221 3334 -187
rect 3300 -293 3334 -259
rect 3300 -365 3334 -331
rect 3300 -437 3334 -403
rect -3034 -509 -3000 -475
rect -3034 -581 -3000 -547
rect -3034 -653 -3000 -619
rect -180 -493 -146 -459
rect -106 -493 -72 -459
rect -32 -493 2 -459
rect 42 -493 76 -459
rect 116 -493 150 -459
rect 190 -493 224 -459
rect 264 -493 298 -459
rect 338 -493 372 -459
rect 412 -493 446 -459
rect 486 -493 520 -459
rect -180 -567 -146 -533
rect -106 -567 -72 -533
rect -32 -567 2 -533
rect 42 -567 76 -533
rect 116 -567 150 -533
rect 190 -567 224 -533
rect 264 -567 298 -533
rect 338 -567 372 -533
rect 412 -567 446 -533
rect 486 -567 520 -533
rect -180 -641 -146 -607
rect -106 -641 -72 -607
rect -32 -641 2 -607
rect 42 -641 76 -607
rect 116 -641 150 -607
rect 190 -641 224 -607
rect 264 -641 298 -607
rect 338 -641 372 -607
rect 412 -641 446 -607
rect 486 -641 520 -607
rect 3300 -509 3334 -475
rect 3300 -581 3334 -547
rect 3300 -653 3334 -619
rect -3034 -725 -3000 -691
rect -3034 -797 -3000 -763
rect -3034 -869 -3000 -835
rect -3034 -941 -3000 -907
rect -3034 -1013 -3000 -979
rect -3034 -1085 -3000 -1051
rect -3034 -1157 -3000 -1123
rect -3034 -1229 -3000 -1195
rect -3034 -1301 -3000 -1267
rect -3034 -1373 -3000 -1339
rect -3034 -1445 -3000 -1411
rect -3034 -1517 -3000 -1483
rect -3034 -1589 -3000 -1555
rect -3034 -1661 -3000 -1627
rect -3034 -1733 -3000 -1699
rect -3034 -1805 -3000 -1771
rect -3034 -1877 -3000 -1843
rect 3300 -725 3334 -691
rect 3300 -797 3334 -763
rect 3300 -869 3334 -835
rect 3300 -941 3334 -907
rect 3300 -1013 3334 -979
rect 3300 -1085 3334 -1051
rect 3300 -1157 3334 -1123
rect 3300 -1229 3334 -1195
rect 3300 -1301 3334 -1267
rect 3300 -1373 3334 -1339
rect 3300 -1445 3334 -1411
rect 3300 -1517 3334 -1483
rect 3300 -1589 3334 -1555
rect 3300 -1661 3334 -1627
rect 3300 -1733 3334 -1699
rect 3300 -1805 3334 -1771
rect 3300 -1877 3334 -1843
rect -2927 -1958 -2893 -1924
rect -2855 -1958 -2821 -1924
rect -2783 -1958 -2749 -1924
rect -2711 -1958 -2677 -1924
rect -2639 -1958 -2605 -1924
rect -2567 -1958 -2533 -1924
rect -2495 -1958 -2461 -1924
rect -2423 -1958 -2389 -1924
rect -2351 -1958 -2317 -1924
rect -2279 -1958 -2245 -1924
rect -2207 -1958 -2173 -1924
rect -2135 -1958 -2101 -1924
rect -2063 -1958 -2029 -1924
rect -1991 -1958 -1957 -1924
rect -1919 -1958 -1885 -1924
rect -1847 -1958 -1813 -1924
rect -1775 -1958 -1741 -1924
rect -1703 -1958 -1669 -1924
rect -1631 -1958 -1597 -1924
rect -1559 -1958 -1525 -1924
rect -1487 -1958 -1453 -1924
rect -1415 -1958 -1381 -1924
rect -1343 -1958 -1309 -1924
rect -1271 -1958 -1237 -1924
rect -1199 -1958 -1165 -1924
rect -1127 -1958 -1093 -1924
rect -1055 -1958 -1021 -1924
rect -983 -1958 -949 -1924
rect -911 -1958 -877 -1924
rect -839 -1958 -805 -1924
rect -767 -1958 -733 -1924
rect -695 -1958 -661 -1924
rect -623 -1958 -589 -1924
rect -551 -1958 -517 -1924
rect -479 -1958 -445 -1924
rect -407 -1958 -373 -1924
rect -335 -1958 -301 -1924
rect -263 -1958 -229 -1924
rect -191 -1958 -157 -1924
rect -119 -1958 -85 -1924
rect -47 -1958 -13 -1924
rect 25 -1958 59 -1924
rect 97 -1958 131 -1924
rect 169 -1958 203 -1924
rect 241 -1958 275 -1924
rect 313 -1958 347 -1924
rect 385 -1958 419 -1924
rect 457 -1958 491 -1924
rect 529 -1958 563 -1924
rect 601 -1958 635 -1924
rect 673 -1958 707 -1924
rect 745 -1958 779 -1924
rect 817 -1958 851 -1924
rect 889 -1958 923 -1924
rect 961 -1958 995 -1924
rect 1033 -1958 1067 -1924
rect 1105 -1958 1139 -1924
rect 1177 -1958 1211 -1924
rect 1249 -1958 1283 -1924
rect 1321 -1958 1355 -1924
rect 1393 -1958 1427 -1924
rect 1465 -1958 1499 -1924
rect 1537 -1958 1571 -1924
rect 1609 -1958 1643 -1924
rect 1681 -1958 1715 -1924
rect 1753 -1958 1787 -1924
rect 1825 -1958 1859 -1924
rect 1897 -1958 1931 -1924
rect 1969 -1958 2003 -1924
rect 2041 -1958 2075 -1924
rect 2113 -1958 2147 -1924
rect 2185 -1958 2219 -1924
rect 2257 -1958 2291 -1924
rect 2329 -1958 2363 -1924
rect 2401 -1958 2435 -1924
rect 2473 -1958 2507 -1924
rect 2545 -1958 2579 -1924
rect 2617 -1958 2651 -1924
rect 2689 -1958 2723 -1924
rect 2761 -1958 2795 -1924
rect 2833 -1958 2867 -1924
rect 2905 -1958 2939 -1924
rect 2977 -1958 3011 -1924
rect 3049 -1958 3083 -1924
rect 3121 -1958 3155 -1924
rect 3193 -1958 3227 -1924
<< metal1 >>
rect -3058 7959 3358 7983
rect -3058 7925 -2927 7959
rect -2893 7925 -2855 7959
rect -2821 7925 -2783 7959
rect -2749 7925 -2711 7959
rect -2677 7925 -2639 7959
rect -2605 7925 -2567 7959
rect -2533 7925 -2495 7959
rect -2461 7925 -2423 7959
rect -2389 7925 -2351 7959
rect -2317 7925 -2279 7959
rect -2245 7925 -2207 7959
rect -2173 7925 -2135 7959
rect -2101 7925 -2063 7959
rect -2029 7925 -1991 7959
rect -1957 7925 -1919 7959
rect -1885 7925 -1847 7959
rect -1813 7925 -1775 7959
rect -1741 7925 -1703 7959
rect -1669 7925 -1631 7959
rect -1597 7925 -1559 7959
rect -1525 7925 -1487 7959
rect -1453 7925 -1415 7959
rect -1381 7925 -1343 7959
rect -1309 7925 -1271 7959
rect -1237 7925 -1199 7959
rect -1165 7925 -1127 7959
rect -1093 7925 -1055 7959
rect -1021 7925 -983 7959
rect -949 7925 -911 7959
rect -877 7925 -839 7959
rect -805 7925 -767 7959
rect -733 7925 -695 7959
rect -661 7925 -623 7959
rect -589 7925 -551 7959
rect -517 7925 -479 7959
rect -445 7925 -407 7959
rect -373 7925 -335 7959
rect -301 7925 -263 7959
rect -229 7925 -191 7959
rect -157 7925 -119 7959
rect -85 7925 -47 7959
rect -13 7925 25 7959
rect 59 7925 97 7959
rect 131 7925 169 7959
rect 203 7925 241 7959
rect 275 7925 313 7959
rect 347 7925 385 7959
rect 419 7925 457 7959
rect 491 7925 529 7959
rect 563 7925 601 7959
rect 635 7925 673 7959
rect 707 7925 745 7959
rect 779 7925 817 7959
rect 851 7925 889 7959
rect 923 7925 961 7959
rect 995 7925 1033 7959
rect 1067 7925 1105 7959
rect 1139 7925 1177 7959
rect 1211 7925 1249 7959
rect 1283 7925 1321 7959
rect 1355 7925 1393 7959
rect 1427 7925 1465 7959
rect 1499 7925 1537 7959
rect 1571 7925 1609 7959
rect 1643 7925 1681 7959
rect 1715 7925 1753 7959
rect 1787 7925 1825 7959
rect 1859 7925 1897 7959
rect 1931 7925 1969 7959
rect 2003 7925 2041 7959
rect 2075 7925 2113 7959
rect 2147 7925 2185 7959
rect 2219 7925 2257 7959
rect 2291 7925 2329 7959
rect 2363 7925 2401 7959
rect 2435 7925 2473 7959
rect 2507 7925 2545 7959
rect 2579 7925 2617 7959
rect 2651 7925 2689 7959
rect 2723 7925 2761 7959
rect 2795 7925 2833 7959
rect 2867 7925 2905 7959
rect 2939 7925 2977 7959
rect 3011 7925 3049 7959
rect 3083 7925 3121 7959
rect 3155 7925 3193 7959
rect 3227 7925 3358 7959
rect -3058 7901 3358 7925
rect -3058 7877 -2976 7901
rect -3058 7843 -3034 7877
rect -3000 7843 -2976 7877
rect -3058 7805 -2976 7843
rect -3058 7771 -3034 7805
rect -3000 7771 -2976 7805
rect -3058 7733 -2976 7771
rect -3058 7699 -3034 7733
rect -3000 7699 -2976 7733
rect -3058 7661 -2976 7699
rect -3058 7627 -3034 7661
rect -3000 7627 -2976 7661
rect -3058 7589 -2976 7627
rect -3058 7555 -3034 7589
rect -3000 7555 -2976 7589
rect -3058 7517 -2976 7555
rect -3058 7483 -3034 7517
rect -3000 7483 -2976 7517
rect -3058 7445 -2976 7483
rect -3058 7411 -3034 7445
rect -3000 7411 -2976 7445
rect -3058 7373 -2976 7411
rect -3058 7339 -3034 7373
rect -3000 7339 -2976 7373
rect -3058 7301 -2976 7339
rect -3058 7267 -3034 7301
rect -3000 7267 -2976 7301
rect -3058 7229 -2976 7267
rect -3058 7195 -3034 7229
rect -3000 7195 -2976 7229
rect -3058 7157 -2976 7195
rect -3058 7123 -3034 7157
rect -3000 7123 -2976 7157
rect -3058 7085 -2976 7123
rect -3058 7051 -3034 7085
rect -3000 7051 -2976 7085
rect -3058 7013 -2976 7051
rect -3058 6979 -3034 7013
rect -3000 6979 -2976 7013
rect -3058 6941 -2976 6979
rect -3058 6907 -3034 6941
rect -3000 6907 -2976 6941
rect -3058 6869 -2976 6907
rect -3058 6835 -3034 6869
rect -3000 6835 -2976 6869
rect -3058 6797 -2976 6835
rect -3058 6763 -3034 6797
rect -3000 6763 -2976 6797
rect -3058 6725 -2976 6763
rect -3058 6691 -3034 6725
rect -3000 6691 -2976 6725
rect -3058 6653 -2976 6691
rect -3058 6619 -3034 6653
rect -3000 6619 -2976 6653
rect -3058 6581 -2976 6619
rect -3058 6547 -3034 6581
rect -3000 6547 -2976 6581
rect -3058 6509 -2976 6547
rect -3058 6475 -3034 6509
rect -3000 6475 -2976 6509
rect -3058 6437 -2976 6475
rect -3058 6403 -3034 6437
rect -3000 6403 -2976 6437
rect -3058 6365 -2976 6403
rect -3058 6331 -3034 6365
rect -3000 6331 -2976 6365
rect -3058 6293 -2976 6331
rect -3058 6259 -3034 6293
rect -3000 6259 -2976 6293
rect -3058 6221 -2976 6259
rect -3058 6187 -3034 6221
rect -3000 6187 -2976 6221
rect -3058 6149 -2976 6187
rect -3058 6115 -3034 6149
rect -3000 6115 -2976 6149
rect -3058 6077 -2976 6115
rect -3058 6043 -3034 6077
rect -3000 6043 -2976 6077
rect -3058 6005 -2976 6043
rect -3058 5971 -3034 6005
rect -3000 5971 -2976 6005
rect 3276 7877 3358 7901
rect 3276 7843 3300 7877
rect 3334 7843 3358 7877
rect 3276 7805 3358 7843
rect 3276 7771 3300 7805
rect 3334 7771 3358 7805
rect 3276 7733 3358 7771
rect 3276 7699 3300 7733
rect 3334 7699 3358 7733
rect 3276 7661 3358 7699
rect 3276 7627 3300 7661
rect 3334 7627 3358 7661
rect 3276 7589 3358 7627
rect 3276 7555 3300 7589
rect 3334 7555 3358 7589
rect 3276 7517 3358 7555
rect 3276 7483 3300 7517
rect 3334 7483 3358 7517
rect 3276 7445 3358 7483
rect 3276 7411 3300 7445
rect 3334 7411 3358 7445
rect 3276 7373 3358 7411
rect 3276 7339 3300 7373
rect 3334 7339 3358 7373
rect 3276 7301 3358 7339
rect 3276 7267 3300 7301
rect 3334 7267 3358 7301
rect 3276 7229 3358 7267
rect 3276 7195 3300 7229
rect 3334 7195 3358 7229
rect 3276 7157 3358 7195
rect 3276 7123 3300 7157
rect 3334 7123 3358 7157
rect 3276 7085 3358 7123
rect 3276 7051 3300 7085
rect 3334 7051 3358 7085
rect 3276 7013 3358 7051
rect 3276 6979 3300 7013
rect 3334 6979 3358 7013
rect 3276 6941 3358 6979
rect 3276 6907 3300 6941
rect 3334 6907 3358 6941
rect 3276 6869 3358 6907
rect 3276 6835 3300 6869
rect 3334 6835 3358 6869
rect 3276 6797 3358 6835
rect 3276 6763 3300 6797
rect 3334 6763 3358 6797
rect 3276 6725 3358 6763
rect 3276 6691 3300 6725
rect 3334 6691 3358 6725
rect 3276 6653 3358 6691
rect 3276 6619 3300 6653
rect 3334 6619 3358 6653
rect 3276 6581 3358 6619
rect 3276 6547 3300 6581
rect 3334 6547 3358 6581
rect 3276 6509 3358 6547
rect 3276 6475 3300 6509
rect 3334 6475 3358 6509
rect 3276 6437 3358 6475
rect 3276 6403 3300 6437
rect 3334 6403 3358 6437
rect 3276 6365 3358 6403
rect 3276 6331 3300 6365
rect 3334 6331 3358 6365
rect 3276 6293 3358 6331
rect 3276 6259 3300 6293
rect 3334 6259 3358 6293
rect 3276 6221 3358 6259
rect 3276 6187 3300 6221
rect 3334 6187 3358 6221
rect 3276 6149 3358 6187
rect 3276 6115 3300 6149
rect 3334 6115 3358 6149
rect 3276 6077 3358 6115
rect 3276 6043 3300 6077
rect 3334 6043 3358 6077
rect 3276 6005 3358 6043
rect -3058 5933 -2976 5971
rect -3058 5899 -3034 5933
rect -3000 5899 -2976 5933
rect -3058 5861 -2976 5899
rect -3058 5827 -3034 5861
rect -3000 5827 -2976 5861
rect -3058 5789 -2976 5827
rect -3058 5755 -3034 5789
rect -3000 5755 -2976 5789
rect -3058 5717 -2976 5755
rect -3058 5683 -3034 5717
rect -3000 5683 -2976 5717
rect -3058 5645 -2976 5683
rect -3058 5611 -3034 5645
rect -3000 5611 -2976 5645
rect -3058 5573 -2976 5611
rect -3058 5539 -3034 5573
rect -3000 5539 -2976 5573
rect -3058 5501 -2976 5539
rect -3058 5467 -3034 5501
rect -3000 5467 -2976 5501
rect -3058 5429 -2976 5467
rect -3058 5395 -3034 5429
rect -3000 5395 -2976 5429
rect -3058 5357 -2976 5395
rect -3058 5323 -3034 5357
rect -3000 5323 -2976 5357
rect -3058 5285 -2976 5323
rect -3058 5251 -3034 5285
rect -3000 5251 -2976 5285
rect -3058 5213 -2976 5251
rect -3058 5179 -3034 5213
rect -3000 5179 -2976 5213
rect -3058 5141 -2976 5179
rect -3058 5107 -3034 5141
rect -3000 5107 -2976 5141
rect -3058 5069 -2976 5107
rect -3058 5035 -3034 5069
rect -3000 5035 -2976 5069
rect -3058 4997 -2976 5035
rect -3058 4963 -3034 4997
rect -3000 4963 -2976 4997
rect -3058 4925 -2976 4963
rect -3058 4891 -3034 4925
rect -3000 4891 -2976 4925
rect -3058 4853 -2976 4891
rect -3058 4819 -3034 4853
rect -3000 4819 -2976 4853
rect -3058 4781 -2976 4819
rect -3058 4747 -3034 4781
rect -3000 4747 -2976 4781
rect -3058 4709 -2976 4747
rect -3058 4675 -3034 4709
rect -3000 4675 -2976 4709
rect -3058 4637 -2976 4675
rect -3058 4603 -3034 4637
rect -3000 4603 -2976 4637
rect -3058 4565 -2976 4603
rect -3058 4531 -3034 4565
rect -3000 4531 -2976 4565
rect -3058 4493 -2976 4531
rect -3058 4459 -3034 4493
rect -3000 4459 -2976 4493
rect -3058 4421 -2976 4459
rect -3058 4387 -3034 4421
rect -3000 4387 -2976 4421
rect -3058 4349 -2976 4387
rect -3058 4315 -3034 4349
rect -3000 4315 -2976 4349
rect -3058 4277 -2976 4315
rect -3058 4243 -3034 4277
rect -3000 4243 -2976 4277
rect -3058 4205 -2976 4243
rect -3058 4171 -3034 4205
rect -3000 4171 -2976 4205
rect -3058 4133 -2976 4171
rect -3058 4099 -3034 4133
rect -3000 4099 -2976 4133
rect -3058 4061 -2976 4099
rect -3058 4027 -3034 4061
rect -3000 4027 -2976 4061
rect -3058 3989 -2976 4027
rect -3058 3955 -3034 3989
rect -3000 3955 -2976 3989
rect -3058 3917 -2976 3955
rect -3058 3883 -3034 3917
rect -3000 3883 -2976 3917
rect -3058 3845 -2976 3883
rect -3058 3811 -3034 3845
rect -3000 3811 -2976 3845
rect -3058 3773 -2976 3811
rect -3058 3739 -3034 3773
rect -3000 3739 -2976 3773
rect -3058 3701 -2976 3739
rect -3058 3667 -3034 3701
rect -3000 3667 -2976 3701
rect -3058 3629 -2976 3667
rect -3058 3595 -3034 3629
rect -3000 3595 -2976 3629
rect -3058 3557 -2976 3595
rect -3058 3523 -3034 3557
rect -3000 3523 -2976 3557
rect -3058 3485 -2976 3523
rect -3058 3451 -3034 3485
rect -3000 3451 -2976 3485
rect -3058 3413 -2976 3451
rect -3058 3379 -3034 3413
rect -3000 3379 -2976 3413
rect -3058 3341 -2976 3379
rect -3058 3307 -3034 3341
rect -3000 3307 -2976 3341
rect -3058 3269 -2976 3307
rect -3058 3235 -3034 3269
rect -3000 3235 -2976 3269
rect -3058 3197 -2976 3235
rect -3058 3163 -3034 3197
rect -3000 3163 -2976 3197
rect -3058 3125 -2976 3163
rect -3058 3091 -3034 3125
rect -3000 3091 -2976 3125
rect -3058 3053 -2976 3091
rect -3058 3019 -3034 3053
rect -3000 3019 -2976 3053
rect -3058 2981 -2976 3019
rect -3058 2947 -3034 2981
rect -3000 2947 -2976 2981
rect -3058 2909 -2976 2947
rect -3058 2875 -3034 2909
rect -3000 2875 -2976 2909
rect -3058 2837 -2976 2875
rect -3058 2803 -3034 2837
rect -3000 2803 -2976 2837
rect -3058 2765 -2976 2803
rect -3058 2731 -3034 2765
rect -3000 2731 -2976 2765
rect -3058 2693 -2976 2731
rect -3058 2659 -3034 2693
rect -3000 2659 -2976 2693
rect -3058 2621 -2976 2659
rect -3058 2587 -3034 2621
rect -3000 2587 -2976 2621
rect -3058 2549 -2976 2587
rect -3058 2515 -3034 2549
rect -3000 2515 -2976 2549
rect -3058 2477 -2976 2515
rect -3058 2443 -3034 2477
rect -3000 2443 -2976 2477
rect -3058 2405 -2976 2443
rect -3058 2371 -3034 2405
rect -3000 2371 -2976 2405
rect -3058 2333 -2976 2371
rect -3058 2299 -3034 2333
rect -3000 2299 -2976 2333
rect -3058 2261 -2976 2299
rect -3058 2227 -3034 2261
rect -3000 2227 -2976 2261
rect -3058 2189 -2976 2227
rect -3058 2155 -3034 2189
rect -3000 2155 -2976 2189
rect -3058 2117 -2976 2155
rect -3058 2083 -3034 2117
rect -3000 2083 -2976 2117
rect -3058 2045 -2976 2083
rect -3058 2011 -3034 2045
rect -3000 2011 -2976 2045
rect -3058 1973 -2976 2011
rect -3058 1939 -3034 1973
rect -3000 1939 -2976 1973
rect -3058 1901 -2976 1939
rect -3058 1867 -3034 1901
rect -3000 1867 -2976 1901
rect -3058 1829 -2976 1867
rect -3058 1795 -3034 1829
rect -3000 1795 -2976 1829
rect -3058 1757 -2976 1795
rect -3058 1723 -3034 1757
rect -3000 1723 -2976 1757
rect -3058 1685 -2976 1723
rect -3058 1651 -3034 1685
rect -3000 1651 -2976 1685
rect -3058 1613 -2976 1651
rect -3058 1579 -3034 1613
rect -3000 1579 -2976 1613
rect -3058 1541 -2976 1579
rect -3058 1507 -3034 1541
rect -3000 1507 -2976 1541
rect -3058 1469 -2976 1507
rect -3058 1435 -3034 1469
rect -3000 1435 -2976 1469
rect -3058 1397 -2976 1435
rect -3058 1363 -3034 1397
rect -3000 1363 -2976 1397
rect -3058 1325 -2976 1363
rect -3058 1291 -3034 1325
rect -3000 1291 -2976 1325
rect -3058 1253 -2976 1291
rect -3058 1219 -3034 1253
rect -3000 1219 -2976 1253
rect -3058 1181 -2976 1219
rect -3058 1147 -3034 1181
rect -3000 1147 -2976 1181
rect -3058 1109 -2976 1147
rect -3058 1075 -3034 1109
rect -3000 1075 -2976 1109
rect -3058 1037 -2976 1075
rect -3058 1003 -3034 1037
rect -3000 1003 -2976 1037
rect -3058 965 -2976 1003
rect -3058 931 -3034 965
rect -3000 931 -2976 965
rect -3058 893 -2976 931
rect -3058 859 -3034 893
rect -3000 859 -2976 893
rect -3058 821 -2976 859
rect -3058 787 -3034 821
rect -3000 787 -2976 821
rect -3058 749 -2976 787
rect -3058 715 -3034 749
rect -3000 715 -2976 749
rect -3058 677 -2976 715
rect -3058 643 -3034 677
rect -3000 643 -2976 677
rect -3058 605 -2976 643
rect -3058 571 -3034 605
rect -3000 571 -2976 605
rect -3058 533 -2976 571
rect -3058 499 -3034 533
rect -3000 499 -2976 533
rect -3058 461 -2976 499
rect -3058 427 -3034 461
rect -3000 427 -2976 461
rect -3058 389 -2976 427
rect -3058 355 -3034 389
rect -3000 355 -2976 389
rect -3058 317 -2976 355
rect -3058 283 -3034 317
rect -3000 283 -2976 317
rect -3058 245 -2976 283
rect -3058 211 -3034 245
rect -3000 211 -2976 245
rect -3058 173 -2976 211
rect -3058 139 -3034 173
rect -3000 139 -2976 173
rect -3058 101 -2976 139
rect -3058 67 -3034 101
rect -3000 67 -2976 101
rect -3058 29 -2976 67
rect -3058 -5 -3034 29
rect -3000 -5 -2976 29
rect -1066 5969 -936 5981
rect -1066 31 -1054 5969
rect -948 31 -936 5969
rect -1066 19 -936 31
rect -828 5969 -698 5981
rect -828 31 -816 5969
rect -710 31 -698 5969
rect 998 5969 1128 5981
rect 13 5939 287 5945
rect 13 5933 28 5939
rect 272 5933 287 5939
rect 13 67 25 5933
rect 275 67 287 5933
rect 13 63 28 67
rect 272 63 287 67
rect 13 55 287 63
rect -828 19 -698 31
rect 998 31 1010 5969
rect 1116 31 1128 5969
rect 998 19 1128 31
rect 1236 5969 1366 5981
rect 1236 31 1248 5969
rect 1354 31 1366 5969
rect 1236 19 1366 31
rect 3276 5971 3300 6005
rect 3334 5971 3358 6005
rect 3276 5933 3358 5971
rect 3276 5899 3300 5933
rect 3334 5899 3358 5933
rect 3276 5861 3358 5899
rect 3276 5827 3300 5861
rect 3334 5827 3358 5861
rect 3276 5789 3358 5827
rect 3276 5755 3300 5789
rect 3334 5755 3358 5789
rect 3276 5717 3358 5755
rect 3276 5683 3300 5717
rect 3334 5683 3358 5717
rect 3276 5645 3358 5683
rect 3276 5611 3300 5645
rect 3334 5611 3358 5645
rect 3276 5573 3358 5611
rect 3276 5539 3300 5573
rect 3334 5539 3358 5573
rect 3276 5501 3358 5539
rect 3276 5467 3300 5501
rect 3334 5467 3358 5501
rect 3276 5429 3358 5467
rect 3276 5395 3300 5429
rect 3334 5395 3358 5429
rect 3276 5357 3358 5395
rect 3276 5323 3300 5357
rect 3334 5323 3358 5357
rect 3276 5285 3358 5323
rect 3276 5251 3300 5285
rect 3334 5251 3358 5285
rect 3276 5213 3358 5251
rect 3276 5179 3300 5213
rect 3334 5179 3358 5213
rect 3276 5141 3358 5179
rect 3276 5107 3300 5141
rect 3334 5107 3358 5141
rect 3276 5069 3358 5107
rect 3276 5035 3300 5069
rect 3334 5035 3358 5069
rect 3276 4997 3358 5035
rect 3276 4963 3300 4997
rect 3334 4963 3358 4997
rect 3276 4925 3358 4963
rect 3276 4891 3300 4925
rect 3334 4891 3358 4925
rect 3276 4853 3358 4891
rect 3276 4819 3300 4853
rect 3334 4819 3358 4853
rect 3276 4781 3358 4819
rect 3276 4747 3300 4781
rect 3334 4747 3358 4781
rect 3276 4709 3358 4747
rect 3276 4675 3300 4709
rect 3334 4675 3358 4709
rect 3276 4637 3358 4675
rect 3276 4603 3300 4637
rect 3334 4603 3358 4637
rect 3276 4565 3358 4603
rect 3276 4531 3300 4565
rect 3334 4531 3358 4565
rect 3276 4493 3358 4531
rect 3276 4459 3300 4493
rect 3334 4459 3358 4493
rect 3276 4421 3358 4459
rect 3276 4387 3300 4421
rect 3334 4387 3358 4421
rect 3276 4349 3358 4387
rect 3276 4315 3300 4349
rect 3334 4315 3358 4349
rect 3276 4277 3358 4315
rect 3276 4243 3300 4277
rect 3334 4243 3358 4277
rect 3276 4205 3358 4243
rect 3276 4171 3300 4205
rect 3334 4171 3358 4205
rect 3276 4133 3358 4171
rect 3276 4099 3300 4133
rect 3334 4099 3358 4133
rect 3276 4061 3358 4099
rect 3276 4027 3300 4061
rect 3334 4027 3358 4061
rect 3276 3989 3358 4027
rect 3276 3955 3300 3989
rect 3334 3955 3358 3989
rect 3276 3917 3358 3955
rect 3276 3883 3300 3917
rect 3334 3883 3358 3917
rect 3276 3845 3358 3883
rect 3276 3811 3300 3845
rect 3334 3811 3358 3845
rect 3276 3773 3358 3811
rect 3276 3739 3300 3773
rect 3334 3739 3358 3773
rect 3276 3701 3358 3739
rect 3276 3667 3300 3701
rect 3334 3667 3358 3701
rect 3276 3629 3358 3667
rect 3276 3595 3300 3629
rect 3334 3595 3358 3629
rect 3276 3557 3358 3595
rect 3276 3523 3300 3557
rect 3334 3523 3358 3557
rect 3276 3485 3358 3523
rect 3276 3451 3300 3485
rect 3334 3451 3358 3485
rect 3276 3413 3358 3451
rect 3276 3379 3300 3413
rect 3334 3379 3358 3413
rect 3276 3341 3358 3379
rect 3276 3307 3300 3341
rect 3334 3307 3358 3341
rect 3276 3269 3358 3307
rect 3276 3235 3300 3269
rect 3334 3235 3358 3269
rect 3276 3197 3358 3235
rect 3276 3163 3300 3197
rect 3334 3163 3358 3197
rect 3276 3125 3358 3163
rect 3276 3091 3300 3125
rect 3334 3091 3358 3125
rect 3276 3053 3358 3091
rect 3276 3019 3300 3053
rect 3334 3019 3358 3053
rect 3276 2981 3358 3019
rect 3276 2947 3300 2981
rect 3334 2947 3358 2981
rect 3276 2909 3358 2947
rect 3276 2875 3300 2909
rect 3334 2875 3358 2909
rect 3276 2837 3358 2875
rect 3276 2803 3300 2837
rect 3334 2803 3358 2837
rect 3276 2765 3358 2803
rect 3276 2731 3300 2765
rect 3334 2731 3358 2765
rect 3276 2693 3358 2731
rect 3276 2659 3300 2693
rect 3334 2659 3358 2693
rect 3276 2621 3358 2659
rect 3276 2587 3300 2621
rect 3334 2587 3358 2621
rect 3276 2549 3358 2587
rect 3276 2515 3300 2549
rect 3334 2515 3358 2549
rect 3276 2477 3358 2515
rect 3276 2443 3300 2477
rect 3334 2443 3358 2477
rect 3276 2405 3358 2443
rect 3276 2371 3300 2405
rect 3334 2371 3358 2405
rect 3276 2333 3358 2371
rect 3276 2299 3300 2333
rect 3334 2299 3358 2333
rect 3276 2261 3358 2299
rect 3276 2227 3300 2261
rect 3334 2227 3358 2261
rect 3276 2189 3358 2227
rect 3276 2155 3300 2189
rect 3334 2155 3358 2189
rect 3276 2117 3358 2155
rect 3276 2083 3300 2117
rect 3334 2083 3358 2117
rect 3276 2045 3358 2083
rect 3276 2011 3300 2045
rect 3334 2011 3358 2045
rect 3276 1973 3358 2011
rect 3276 1939 3300 1973
rect 3334 1939 3358 1973
rect 3276 1901 3358 1939
rect 3276 1867 3300 1901
rect 3334 1867 3358 1901
rect 3276 1829 3358 1867
rect 3276 1795 3300 1829
rect 3334 1795 3358 1829
rect 3276 1757 3358 1795
rect 3276 1723 3300 1757
rect 3334 1723 3358 1757
rect 3276 1685 3358 1723
rect 3276 1651 3300 1685
rect 3334 1651 3358 1685
rect 3276 1613 3358 1651
rect 3276 1579 3300 1613
rect 3334 1579 3358 1613
rect 3276 1541 3358 1579
rect 3276 1507 3300 1541
rect 3334 1507 3358 1541
rect 3276 1469 3358 1507
rect 3276 1435 3300 1469
rect 3334 1435 3358 1469
rect 3276 1397 3358 1435
rect 3276 1363 3300 1397
rect 3334 1363 3358 1397
rect 3276 1325 3358 1363
rect 3276 1291 3300 1325
rect 3334 1291 3358 1325
rect 3276 1253 3358 1291
rect 3276 1219 3300 1253
rect 3334 1219 3358 1253
rect 3276 1181 3358 1219
rect 3276 1147 3300 1181
rect 3334 1147 3358 1181
rect 3276 1109 3358 1147
rect 3276 1075 3300 1109
rect 3334 1075 3358 1109
rect 3276 1037 3358 1075
rect 3276 1003 3300 1037
rect 3334 1003 3358 1037
rect 3276 965 3358 1003
rect 3276 931 3300 965
rect 3334 931 3358 965
rect 3276 893 3358 931
rect 3276 859 3300 893
rect 3334 859 3358 893
rect 3276 821 3358 859
rect 3276 787 3300 821
rect 3334 787 3358 821
rect 3276 749 3358 787
rect 3276 715 3300 749
rect 3334 715 3358 749
rect 3276 677 3358 715
rect 3276 643 3300 677
rect 3334 643 3358 677
rect 3276 605 3358 643
rect 3276 571 3300 605
rect 3334 571 3358 605
rect 3276 533 3358 571
rect 3276 499 3300 533
rect 3334 499 3358 533
rect 3276 461 3358 499
rect 3276 427 3300 461
rect 3334 427 3358 461
rect 3276 389 3358 427
rect 3276 355 3300 389
rect 3334 355 3358 389
rect 3276 317 3358 355
rect 3276 283 3300 317
rect 3334 283 3358 317
rect 3276 245 3358 283
rect 3276 211 3300 245
rect 3334 211 3358 245
rect 3276 173 3358 211
rect 3276 139 3300 173
rect 3334 139 3358 173
rect 3276 101 3358 139
rect 3276 67 3300 101
rect 3334 67 3358 101
rect 3276 29 3358 67
rect -3058 -43 -2976 -5
rect -3058 -77 -3034 -43
rect -3000 -77 -2976 -43
rect -3058 -115 -2976 -77
rect -3058 -149 -3034 -115
rect -3000 -149 -2976 -115
rect -3058 -187 -2976 -149
rect -3058 -221 -3034 -187
rect -3000 -221 -2976 -187
rect -3058 -259 -2976 -221
rect -3058 -293 -3034 -259
rect -3000 -293 -2976 -259
rect -3058 -331 -2976 -293
rect -3058 -365 -3034 -331
rect -3000 -365 -2976 -331
rect -3058 -403 -2976 -365
rect -3058 -437 -3034 -403
rect -3000 -437 -2976 -403
rect -3058 -475 -2976 -437
rect 3276 -5 3300 29
rect 3334 -5 3358 29
rect 3276 -43 3358 -5
rect 3276 -77 3300 -43
rect 3334 -77 3358 -43
rect 3276 -115 3358 -77
rect 3276 -149 3300 -115
rect 3334 -149 3358 -115
rect 3276 -187 3358 -149
rect 3276 -221 3300 -187
rect 3334 -221 3358 -187
rect 3276 -259 3358 -221
rect 3276 -293 3300 -259
rect 3334 -293 3358 -259
rect 3276 -331 3358 -293
rect 3276 -365 3300 -331
rect 3334 -365 3358 -331
rect 3276 -403 3358 -365
rect 3276 -437 3300 -403
rect 3334 -437 3358 -403
rect -3058 -509 -3034 -475
rect -3000 -509 -2976 -475
rect -3058 -547 -2976 -509
rect -3058 -581 -3034 -547
rect -3000 -581 -2976 -547
rect -3058 -619 -2976 -581
rect -3058 -653 -3034 -619
rect -3000 -653 -2976 -619
rect -3058 -691 -2976 -653
rect -209 -450 555 -443
rect -209 -502 -189 -450
rect -137 -502 -115 -450
rect -63 -502 -41 -450
rect 11 -502 33 -450
rect 85 -502 107 -450
rect 159 -502 181 -450
rect 233 -502 255 -450
rect 307 -502 329 -450
rect 381 -502 403 -450
rect 455 -502 477 -450
rect 529 -502 555 -450
rect -209 -524 555 -502
rect -209 -576 -189 -524
rect -137 -576 -115 -524
rect -63 -576 -41 -524
rect 11 -576 33 -524
rect 85 -576 107 -524
rect 159 -576 181 -524
rect 233 -576 255 -524
rect 307 -576 329 -524
rect 381 -576 403 -524
rect 455 -576 477 -524
rect 529 -576 555 -524
rect -209 -598 555 -576
rect -209 -650 -189 -598
rect -137 -650 -115 -598
rect -63 -650 -41 -598
rect 11 -650 33 -598
rect 85 -650 107 -598
rect 159 -650 181 -598
rect 233 -650 255 -598
rect 307 -650 329 -598
rect 381 -650 403 -598
rect 455 -650 477 -598
rect 529 -650 555 -598
rect -209 -657 555 -650
rect 3276 -475 3358 -437
rect 3276 -509 3300 -475
rect 3334 -509 3358 -475
rect 3276 -547 3358 -509
rect 3276 -581 3300 -547
rect 3334 -581 3358 -547
rect 3276 -619 3358 -581
rect 3276 -653 3300 -619
rect 3334 -653 3358 -619
rect -3058 -725 -3034 -691
rect -3000 -725 -2976 -691
rect -3058 -763 -2976 -725
rect -3058 -797 -3034 -763
rect -3000 -797 -2976 -763
rect -3058 -835 -2976 -797
rect -3058 -869 -3034 -835
rect -3000 -869 -2976 -835
rect -3058 -907 -2976 -869
rect -3058 -941 -3034 -907
rect -3000 -941 -2976 -907
rect -3058 -979 -2976 -941
rect -3058 -1013 -3034 -979
rect -3000 -1013 -2976 -979
rect -3058 -1051 -2976 -1013
rect -3058 -1085 -3034 -1051
rect -3000 -1085 -2976 -1051
rect -3058 -1123 -2976 -1085
rect -3058 -1157 -3034 -1123
rect -3000 -1157 -2976 -1123
rect -3058 -1195 -2976 -1157
rect -3058 -1229 -3034 -1195
rect -3000 -1229 -2976 -1195
rect -3058 -1267 -2976 -1229
rect -3058 -1301 -3034 -1267
rect -3000 -1301 -2976 -1267
rect -3058 -1339 -2976 -1301
rect -3058 -1373 -3034 -1339
rect -3000 -1373 -2976 -1339
rect -3058 -1411 -2976 -1373
rect -3058 -1445 -3034 -1411
rect -3000 -1445 -2976 -1411
rect -3058 -1483 -2976 -1445
rect -3058 -1517 -3034 -1483
rect -3000 -1517 -2976 -1483
rect -3058 -1555 -2976 -1517
rect -3058 -1589 -3034 -1555
rect -3000 -1589 -2976 -1555
rect -3058 -1627 -2976 -1589
rect -3058 -1661 -3034 -1627
rect -3000 -1661 -2976 -1627
rect -3058 -1699 -2976 -1661
rect -3058 -1733 -3034 -1699
rect -3000 -1733 -2976 -1699
rect -3058 -1771 -2976 -1733
rect -3058 -1805 -3034 -1771
rect -3000 -1805 -2976 -1771
rect -3058 -1843 -2976 -1805
rect -3058 -1877 -3034 -1843
rect -3000 -1877 -2976 -1843
rect -3058 -1900 -2976 -1877
rect 3276 -691 3358 -653
rect 3276 -725 3300 -691
rect 3334 -725 3358 -691
rect 3276 -763 3358 -725
rect 3276 -797 3300 -763
rect 3334 -797 3358 -763
rect 3276 -835 3358 -797
rect 3276 -869 3300 -835
rect 3334 -869 3358 -835
rect 3276 -907 3358 -869
rect 3276 -941 3300 -907
rect 3334 -941 3358 -907
rect 3276 -979 3358 -941
rect 3276 -1013 3300 -979
rect 3334 -1013 3358 -979
rect 3276 -1051 3358 -1013
rect 3276 -1085 3300 -1051
rect 3334 -1085 3358 -1051
rect 3276 -1123 3358 -1085
rect 3276 -1157 3300 -1123
rect 3334 -1157 3358 -1123
rect 3276 -1195 3358 -1157
rect 3276 -1229 3300 -1195
rect 3334 -1229 3358 -1195
rect 3276 -1267 3358 -1229
rect 3276 -1301 3300 -1267
rect 3334 -1301 3358 -1267
rect 3276 -1339 3358 -1301
rect 3276 -1373 3300 -1339
rect 3334 -1373 3358 -1339
rect 3276 -1411 3358 -1373
rect 3276 -1445 3300 -1411
rect 3334 -1445 3358 -1411
rect 3276 -1483 3358 -1445
rect 3276 -1517 3300 -1483
rect 3334 -1517 3358 -1483
rect 3276 -1555 3358 -1517
rect 3276 -1589 3300 -1555
rect 3334 -1589 3358 -1555
rect 3276 -1627 3358 -1589
rect 3276 -1661 3300 -1627
rect 3334 -1661 3358 -1627
rect 3276 -1699 3358 -1661
rect 3276 -1733 3300 -1699
rect 3334 -1733 3358 -1699
rect 3276 -1771 3358 -1733
rect 3276 -1805 3300 -1771
rect 3334 -1805 3358 -1771
rect 3276 -1843 3358 -1805
rect 3276 -1877 3300 -1843
rect 3334 -1877 3358 -1843
rect 3276 -1900 3358 -1877
rect -3058 -1924 3358 -1900
rect -3058 -1958 -2927 -1924
rect -2893 -1958 -2855 -1924
rect -2821 -1958 -2783 -1924
rect -2749 -1958 -2711 -1924
rect -2677 -1958 -2639 -1924
rect -2605 -1958 -2567 -1924
rect -2533 -1958 -2495 -1924
rect -2461 -1958 -2423 -1924
rect -2389 -1958 -2351 -1924
rect -2317 -1958 -2279 -1924
rect -2245 -1958 -2207 -1924
rect -2173 -1958 -2135 -1924
rect -2101 -1958 -2063 -1924
rect -2029 -1958 -1991 -1924
rect -1957 -1958 -1919 -1924
rect -1885 -1958 -1847 -1924
rect -1813 -1958 -1775 -1924
rect -1741 -1958 -1703 -1924
rect -1669 -1958 -1631 -1924
rect -1597 -1958 -1559 -1924
rect -1525 -1958 -1487 -1924
rect -1453 -1958 -1415 -1924
rect -1381 -1958 -1343 -1924
rect -1309 -1958 -1271 -1924
rect -1237 -1958 -1199 -1924
rect -1165 -1958 -1127 -1924
rect -1093 -1958 -1055 -1924
rect -1021 -1958 -983 -1924
rect -949 -1958 -911 -1924
rect -877 -1958 -839 -1924
rect -805 -1958 -767 -1924
rect -733 -1958 -695 -1924
rect -661 -1958 -623 -1924
rect -589 -1958 -551 -1924
rect -517 -1958 -479 -1924
rect -445 -1958 -407 -1924
rect -373 -1958 -335 -1924
rect -301 -1958 -263 -1924
rect -229 -1958 -191 -1924
rect -157 -1958 -119 -1924
rect -85 -1958 -47 -1924
rect -13 -1958 25 -1924
rect 59 -1958 97 -1924
rect 131 -1958 169 -1924
rect 203 -1958 241 -1924
rect 275 -1958 313 -1924
rect 347 -1958 385 -1924
rect 419 -1958 457 -1924
rect 491 -1958 529 -1924
rect 563 -1958 601 -1924
rect 635 -1958 673 -1924
rect 707 -1958 745 -1924
rect 779 -1958 817 -1924
rect 851 -1958 889 -1924
rect 923 -1958 961 -1924
rect 995 -1958 1033 -1924
rect 1067 -1958 1105 -1924
rect 1139 -1958 1177 -1924
rect 1211 -1958 1249 -1924
rect 1283 -1958 1321 -1924
rect 1355 -1958 1393 -1924
rect 1427 -1958 1465 -1924
rect 1499 -1958 1537 -1924
rect 1571 -1958 1609 -1924
rect 1643 -1958 1681 -1924
rect 1715 -1958 1753 -1924
rect 1787 -1958 1825 -1924
rect 1859 -1958 1897 -1924
rect 1931 -1958 1969 -1924
rect 2003 -1958 2041 -1924
rect 2075 -1958 2113 -1924
rect 2147 -1958 2185 -1924
rect 2219 -1958 2257 -1924
rect 2291 -1958 2329 -1924
rect 2363 -1958 2401 -1924
rect 2435 -1958 2473 -1924
rect 2507 -1958 2545 -1924
rect 2579 -1958 2617 -1924
rect 2651 -1958 2689 -1924
rect 2723 -1958 2761 -1924
rect 2795 -1958 2833 -1924
rect 2867 -1958 2905 -1924
rect 2939 -1958 2977 -1924
rect 3011 -1958 3049 -1924
rect 3083 -1958 3121 -1924
rect 3155 -1958 3193 -1924
rect 3227 -1958 3358 -1924
rect -3058 -1982 3358 -1958
<< via1 >>
rect 28 5933 272 5939
rect 28 67 272 5933
rect 28 63 272 67
rect -189 -459 -137 -450
rect -189 -493 -180 -459
rect -180 -493 -146 -459
rect -146 -493 -137 -459
rect -189 -502 -137 -493
rect -115 -459 -63 -450
rect -115 -493 -106 -459
rect -106 -493 -72 -459
rect -72 -493 -63 -459
rect -115 -502 -63 -493
rect -41 -459 11 -450
rect -41 -493 -32 -459
rect -32 -493 2 -459
rect 2 -493 11 -459
rect -41 -502 11 -493
rect 33 -459 85 -450
rect 33 -493 42 -459
rect 42 -493 76 -459
rect 76 -493 85 -459
rect 33 -502 85 -493
rect 107 -459 159 -450
rect 107 -493 116 -459
rect 116 -493 150 -459
rect 150 -493 159 -459
rect 107 -502 159 -493
rect 181 -459 233 -450
rect 181 -493 190 -459
rect 190 -493 224 -459
rect 224 -493 233 -459
rect 181 -502 233 -493
rect 255 -459 307 -450
rect 255 -493 264 -459
rect 264 -493 298 -459
rect 298 -493 307 -459
rect 255 -502 307 -493
rect 329 -459 381 -450
rect 329 -493 338 -459
rect 338 -493 372 -459
rect 372 -493 381 -459
rect 329 -502 381 -493
rect 403 -459 455 -450
rect 403 -493 412 -459
rect 412 -493 446 -459
rect 446 -493 455 -459
rect 403 -502 455 -493
rect 477 -459 529 -450
rect 477 -493 486 -459
rect 486 -493 520 -459
rect 520 -493 529 -459
rect 477 -502 529 -493
rect -189 -533 -137 -524
rect -189 -567 -180 -533
rect -180 -567 -146 -533
rect -146 -567 -137 -533
rect -189 -576 -137 -567
rect -115 -533 -63 -524
rect -115 -567 -106 -533
rect -106 -567 -72 -533
rect -72 -567 -63 -533
rect -115 -576 -63 -567
rect -41 -533 11 -524
rect -41 -567 -32 -533
rect -32 -567 2 -533
rect 2 -567 11 -533
rect -41 -576 11 -567
rect 33 -533 85 -524
rect 33 -567 42 -533
rect 42 -567 76 -533
rect 76 -567 85 -533
rect 33 -576 85 -567
rect 107 -533 159 -524
rect 107 -567 116 -533
rect 116 -567 150 -533
rect 150 -567 159 -533
rect 107 -576 159 -567
rect 181 -533 233 -524
rect 181 -567 190 -533
rect 190 -567 224 -533
rect 224 -567 233 -533
rect 181 -576 233 -567
rect 255 -533 307 -524
rect 255 -567 264 -533
rect 264 -567 298 -533
rect 298 -567 307 -533
rect 255 -576 307 -567
rect 329 -533 381 -524
rect 329 -567 338 -533
rect 338 -567 372 -533
rect 372 -567 381 -533
rect 329 -576 381 -567
rect 403 -533 455 -524
rect 403 -567 412 -533
rect 412 -567 446 -533
rect 446 -567 455 -533
rect 403 -576 455 -567
rect 477 -533 529 -524
rect 477 -567 486 -533
rect 486 -567 520 -533
rect 520 -567 529 -533
rect 477 -576 529 -567
rect -189 -607 -137 -598
rect -189 -641 -180 -607
rect -180 -641 -146 -607
rect -146 -641 -137 -607
rect -189 -650 -137 -641
rect -115 -607 -63 -598
rect -115 -641 -106 -607
rect -106 -641 -72 -607
rect -72 -641 -63 -607
rect -115 -650 -63 -641
rect -41 -607 11 -598
rect -41 -641 -32 -607
rect -32 -641 2 -607
rect 2 -641 11 -607
rect -41 -650 11 -641
rect 33 -607 85 -598
rect 33 -641 42 -607
rect 42 -641 76 -607
rect 76 -641 85 -607
rect 33 -650 85 -641
rect 107 -607 159 -598
rect 107 -641 116 -607
rect 116 -641 150 -607
rect 150 -641 159 -607
rect 107 -650 159 -641
rect 181 -607 233 -598
rect 181 -641 190 -607
rect 190 -641 224 -607
rect 224 -641 233 -607
rect 181 -650 233 -641
rect 255 -607 307 -598
rect 255 -641 264 -607
rect 264 -641 298 -607
rect 298 -641 307 -607
rect 255 -650 307 -641
rect 329 -607 381 -598
rect 329 -641 338 -607
rect 338 -641 372 -607
rect 372 -641 381 -607
rect 329 -650 381 -641
rect 403 -607 455 -598
rect 403 -641 412 -607
rect 412 -641 446 -607
rect 446 -641 455 -607
rect 403 -650 455 -641
rect 477 -607 529 -598
rect 477 -641 486 -607
rect 486 -641 520 -607
rect 520 -641 529 -607
rect 477 -650 529 -641
<< metal2 >>
rect 22 5939 278 5945
rect 22 63 28 5939
rect 272 63 278 5939
rect 22 57 278 63
rect -209 -450 555 -443
rect -209 -502 -189 -450
rect -137 -502 -115 -450
rect -63 -502 -41 -450
rect 11 -502 33 -450
rect 85 -502 107 -450
rect 159 -502 181 -450
rect 233 -502 255 -450
rect 307 -502 329 -450
rect 381 -502 403 -450
rect 455 -502 477 -450
rect 529 -502 555 -450
rect -209 -524 555 -502
rect -209 -576 -189 -524
rect -137 -576 -115 -524
rect -63 -576 -41 -524
rect 11 -576 33 -524
rect 85 -576 107 -524
rect 159 -576 181 -524
rect 233 -576 255 -524
rect 307 -576 329 -524
rect 381 -576 403 -524
rect 455 -576 477 -524
rect 529 -576 555 -524
rect -209 -598 555 -576
rect -209 -650 -189 -598
rect -137 -650 -115 -598
rect -63 -650 -41 -598
rect 11 -650 33 -598
rect 85 -650 107 -598
rect 159 -650 181 -598
rect 233 -650 255 -598
rect 307 -650 329 -598
rect 381 -650 403 -598
rect 455 -650 477 -598
rect 529 -650 555 -598
rect -209 -657 555 -650
<< labels >>
flabel comment s -763 206 -763 206 0 FreeSans 2000 0 0 0 S
flabel comment s 1062 206 1062 206 0 FreeSans 2000 0 0 0 S
flabel comment s 158 206 158 206 0 FreeSans 2000 0 0 0 D
<< properties >>
string GDS_END 5099456
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 4857928
<< end >>
