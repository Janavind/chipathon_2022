magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< pwell >>
rect -40 -8 1998 1322
<< mvnmos >>
rect 179 126 1779 1126
<< mvndiff >>
rect 126 1056 179 1126
rect 126 1022 134 1056
rect 168 1022 179 1056
rect 126 988 179 1022
rect 126 954 134 988
rect 168 954 179 988
rect 126 920 179 954
rect 126 886 134 920
rect 168 886 179 920
rect 126 852 179 886
rect 126 818 134 852
rect 168 818 179 852
rect 126 784 179 818
rect 126 750 134 784
rect 168 750 179 784
rect 126 716 179 750
rect 126 682 134 716
rect 168 682 179 716
rect 126 648 179 682
rect 126 614 134 648
rect 168 614 179 648
rect 126 580 179 614
rect 126 546 134 580
rect 168 546 179 580
rect 126 512 179 546
rect 126 478 134 512
rect 168 478 179 512
rect 126 444 179 478
rect 126 410 134 444
rect 168 410 179 444
rect 126 376 179 410
rect 126 342 134 376
rect 168 342 179 376
rect 126 308 179 342
rect 126 274 134 308
rect 168 274 179 308
rect 126 240 179 274
rect 126 206 134 240
rect 168 206 179 240
rect 126 172 179 206
rect 126 138 134 172
rect 168 138 179 172
rect 126 126 179 138
rect 1779 1056 1832 1126
rect 1779 1022 1790 1056
rect 1824 1022 1832 1056
rect 1779 988 1832 1022
rect 1779 954 1790 988
rect 1824 954 1832 988
rect 1779 920 1832 954
rect 1779 886 1790 920
rect 1824 886 1832 920
rect 1779 852 1832 886
rect 1779 818 1790 852
rect 1824 818 1832 852
rect 1779 784 1832 818
rect 1779 750 1790 784
rect 1824 750 1832 784
rect 1779 716 1832 750
rect 1779 682 1790 716
rect 1824 682 1832 716
rect 1779 648 1832 682
rect 1779 614 1790 648
rect 1824 614 1832 648
rect 1779 580 1832 614
rect 1779 546 1790 580
rect 1824 546 1832 580
rect 1779 512 1832 546
rect 1779 478 1790 512
rect 1824 478 1832 512
rect 1779 444 1832 478
rect 1779 410 1790 444
rect 1824 410 1832 444
rect 1779 376 1832 410
rect 1779 342 1790 376
rect 1824 342 1832 376
rect 1779 308 1832 342
rect 1779 274 1790 308
rect 1824 274 1832 308
rect 1779 240 1832 274
rect 1779 206 1790 240
rect 1824 206 1832 240
rect 1779 172 1832 206
rect 1779 138 1790 172
rect 1824 138 1832 172
rect 1779 126 1832 138
<< mvndiffc >>
rect 134 1022 168 1056
rect 134 954 168 988
rect 134 886 168 920
rect 134 818 168 852
rect 134 750 168 784
rect 134 682 168 716
rect 134 614 168 648
rect 134 546 168 580
rect 134 478 168 512
rect 134 410 168 444
rect 134 342 168 376
rect 134 274 168 308
rect 134 206 168 240
rect 134 138 168 172
rect 1790 1022 1824 1056
rect 1790 954 1824 988
rect 1790 886 1824 920
rect 1790 818 1824 852
rect 1790 750 1824 784
rect 1790 682 1824 716
rect 1790 614 1824 648
rect 1790 546 1824 580
rect 1790 478 1824 512
rect 1790 410 1824 444
rect 1790 342 1824 376
rect 1790 274 1824 308
rect 1790 206 1824 240
rect 1790 138 1824 172
<< mvpsubdiff >>
rect -14 1228 20 1296
rect 54 1262 88 1296
rect 122 1262 156 1296
rect 190 1262 224 1296
rect 258 1262 292 1296
rect 326 1262 360 1296
rect 394 1262 428 1296
rect 462 1262 496 1296
rect 530 1262 564 1296
rect 598 1262 632 1296
rect 666 1262 700 1296
rect 734 1262 768 1296
rect 802 1262 836 1296
rect 870 1262 904 1296
rect 938 1262 972 1296
rect 1006 1262 1040 1296
rect 1074 1262 1108 1296
rect 1142 1262 1176 1296
rect 1210 1262 1244 1296
rect 1278 1262 1312 1296
rect 1346 1262 1380 1296
rect 1414 1262 1448 1296
rect 1482 1262 1516 1296
rect 1550 1262 1584 1296
rect 1618 1262 1652 1296
rect 1686 1262 1720 1296
rect 1754 1262 1788 1296
rect 1822 1262 1856 1296
rect 1890 1262 1972 1296
rect 1938 1228 1972 1262
rect -14 1160 20 1194
rect 1938 1160 1972 1194
rect -14 1092 20 1126
rect -14 1024 20 1058
rect -14 956 20 990
rect -14 888 20 922
rect -14 820 20 854
rect -14 752 20 786
rect -14 684 20 718
rect -14 616 20 650
rect -14 548 20 582
rect -14 480 20 514
rect -14 412 20 446
rect -14 344 20 378
rect -14 276 20 310
rect -14 208 20 242
rect -14 140 20 174
rect 1938 1092 1972 1126
rect 1938 1024 1972 1058
rect 1938 956 1972 990
rect 1938 888 1972 922
rect 1938 820 1972 854
rect 1938 752 1972 786
rect 1938 684 1972 718
rect 1938 616 1972 650
rect 1938 548 1972 582
rect 1938 480 1972 514
rect 1938 412 1972 446
rect 1938 344 1972 378
rect 1938 276 1972 310
rect 1938 208 1972 242
rect 1938 140 1972 174
rect -14 18 20 106
rect 1938 52 1972 106
rect 54 18 88 52
rect 122 18 156 52
rect 190 18 224 52
rect 258 18 292 52
rect 326 18 360 52
rect 394 18 428 52
rect 462 18 496 52
rect 530 18 564 52
rect 598 18 632 52
rect 666 18 700 52
rect 734 18 768 52
rect 802 18 836 52
rect 870 18 904 52
rect 938 18 972 52
rect 1006 18 1040 52
rect 1074 18 1108 52
rect 1142 18 1176 52
rect 1210 18 1244 52
rect 1278 18 1312 52
rect 1346 18 1380 52
rect 1414 18 1448 52
rect 1482 18 1516 52
rect 1550 18 1584 52
rect 1618 18 1652 52
rect 1686 18 1720 52
rect 1754 18 1788 52
rect 1822 18 1856 52
rect 1890 18 1972 52
<< mvpsubdiffcont >>
rect 20 1262 54 1296
rect 88 1262 122 1296
rect 156 1262 190 1296
rect 224 1262 258 1296
rect 292 1262 326 1296
rect 360 1262 394 1296
rect 428 1262 462 1296
rect 496 1262 530 1296
rect 564 1262 598 1296
rect 632 1262 666 1296
rect 700 1262 734 1296
rect 768 1262 802 1296
rect 836 1262 870 1296
rect 904 1262 938 1296
rect 972 1262 1006 1296
rect 1040 1262 1074 1296
rect 1108 1262 1142 1296
rect 1176 1262 1210 1296
rect 1244 1262 1278 1296
rect 1312 1262 1346 1296
rect 1380 1262 1414 1296
rect 1448 1262 1482 1296
rect 1516 1262 1550 1296
rect 1584 1262 1618 1296
rect 1652 1262 1686 1296
rect 1720 1262 1754 1296
rect 1788 1262 1822 1296
rect 1856 1262 1890 1296
rect -14 1194 20 1228
rect -14 1126 20 1160
rect 1938 1194 1972 1228
rect 1938 1126 1972 1160
rect -14 1058 20 1092
rect -14 990 20 1024
rect -14 922 20 956
rect -14 854 20 888
rect -14 786 20 820
rect -14 718 20 752
rect -14 650 20 684
rect -14 582 20 616
rect -14 514 20 548
rect -14 446 20 480
rect -14 378 20 412
rect -14 310 20 344
rect -14 242 20 276
rect -14 174 20 208
rect -14 106 20 140
rect 1938 1058 1972 1092
rect 1938 990 1972 1024
rect 1938 922 1972 956
rect 1938 854 1972 888
rect 1938 786 1972 820
rect 1938 718 1972 752
rect 1938 650 1972 684
rect 1938 582 1972 616
rect 1938 514 1972 548
rect 1938 446 1972 480
rect 1938 378 1972 412
rect 1938 310 1972 344
rect 1938 242 1972 276
rect 1938 174 1972 208
rect 1938 106 1972 140
rect 20 18 54 52
rect 88 18 122 52
rect 156 18 190 52
rect 224 18 258 52
rect 292 18 326 52
rect 360 18 394 52
rect 428 18 462 52
rect 496 18 530 52
rect 564 18 598 52
rect 632 18 666 52
rect 700 18 734 52
rect 768 18 802 52
rect 836 18 870 52
rect 904 18 938 52
rect 972 18 1006 52
rect 1040 18 1074 52
rect 1108 18 1142 52
rect 1176 18 1210 52
rect 1244 18 1278 52
rect 1312 18 1346 52
rect 1380 18 1414 52
rect 1448 18 1482 52
rect 1516 18 1550 52
rect 1584 18 1618 52
rect 1652 18 1686 52
rect 1720 18 1754 52
rect 1788 18 1822 52
rect 1856 18 1890 52
<< poly >>
rect 179 1202 1779 1218
rect 179 1168 199 1202
rect 233 1168 267 1202
rect 301 1168 335 1202
rect 369 1168 403 1202
rect 437 1168 471 1202
rect 505 1168 539 1202
rect 573 1168 607 1202
rect 641 1168 675 1202
rect 709 1168 743 1202
rect 777 1168 811 1202
rect 845 1168 879 1202
rect 913 1168 947 1202
rect 981 1168 1015 1202
rect 1049 1168 1083 1202
rect 1117 1168 1151 1202
rect 1185 1168 1219 1202
rect 1253 1168 1287 1202
rect 1321 1168 1355 1202
rect 1389 1168 1423 1202
rect 1457 1168 1491 1202
rect 1525 1168 1559 1202
rect 1593 1168 1627 1202
rect 1661 1168 1695 1202
rect 1729 1168 1779 1202
rect 179 1126 1779 1168
rect 179 100 1779 126
<< polycont >>
rect 199 1168 233 1202
rect 267 1168 301 1202
rect 335 1168 369 1202
rect 403 1168 437 1202
rect 471 1168 505 1202
rect 539 1168 573 1202
rect 607 1168 641 1202
rect 675 1168 709 1202
rect 743 1168 777 1202
rect 811 1168 845 1202
rect 879 1168 913 1202
rect 947 1168 981 1202
rect 1015 1168 1049 1202
rect 1083 1168 1117 1202
rect 1151 1168 1185 1202
rect 1219 1168 1253 1202
rect 1287 1168 1321 1202
rect 1355 1168 1389 1202
rect 1423 1168 1457 1202
rect 1491 1168 1525 1202
rect 1559 1168 1593 1202
rect 1627 1168 1661 1202
rect 1695 1168 1729 1202
<< locali >>
rect 20 1296 1938 1302
rect -14 1262 20 1296
rect 66 1262 88 1296
rect 138 1262 156 1296
rect 210 1262 224 1296
rect 282 1262 292 1296
rect 354 1262 360 1296
rect 426 1262 428 1296
rect 462 1262 464 1296
rect 530 1262 536 1296
rect 598 1262 608 1296
rect 666 1262 680 1296
rect 734 1262 752 1296
rect 802 1262 824 1296
rect 870 1262 896 1296
rect 938 1262 968 1296
rect 1006 1262 1040 1296
rect 1074 1262 1108 1296
rect 1146 1262 1176 1296
rect 1218 1262 1244 1296
rect 1290 1262 1312 1296
rect 1362 1262 1380 1296
rect 1434 1262 1448 1296
rect 1506 1262 1516 1296
rect 1578 1262 1584 1296
rect 1650 1262 1652 1296
rect 1686 1262 1688 1296
rect 1754 1262 1760 1296
rect 1822 1262 1832 1296
rect 1890 1262 1972 1296
rect -14 1256 1972 1262
rect -14 1228 20 1256
rect 1938 1228 1972 1256
rect -14 1160 20 1194
rect 179 1202 1779 1208
rect 179 1168 191 1202
rect 233 1168 263 1202
rect 301 1168 335 1202
rect 369 1168 403 1202
rect 441 1168 471 1202
rect 513 1168 539 1202
rect 585 1168 607 1202
rect 657 1168 675 1202
rect 729 1168 743 1202
rect 801 1168 811 1202
rect 873 1168 879 1202
rect 945 1168 947 1202
rect 981 1168 983 1202
rect 1049 1168 1055 1202
rect 1117 1168 1127 1202
rect 1185 1168 1199 1202
rect 1253 1168 1271 1202
rect 1321 1168 1343 1202
rect 1389 1168 1415 1202
rect 1457 1168 1487 1202
rect 1525 1168 1559 1202
rect 1593 1168 1627 1202
rect 1665 1168 1695 1202
rect 1737 1168 1779 1202
rect 179 1162 1779 1168
rect -14 1092 20 1126
rect 1938 1160 1972 1194
rect 1938 1092 1972 1126
rect -14 1024 20 1058
rect -14 956 20 990
rect -14 888 20 922
rect -20 854 -14 859
rect 134 1056 168 1072
rect 134 988 168 1022
rect 134 920 168 954
rect 134 859 168 886
rect 1790 1056 1824 1072
rect 1790 988 1824 1022
rect 1790 920 1824 954
rect 1790 859 1824 886
rect 1938 1024 1972 1058
rect 1938 956 1972 990
rect 1938 888 1972 922
rect 20 854 26 859
rect -20 847 26 854
rect -20 786 -14 847
rect 20 786 26 847
rect -20 775 26 786
rect -20 718 -14 775
rect 20 718 26 775
rect -20 703 26 718
rect -20 650 -14 703
rect 20 650 26 703
rect -20 631 26 650
rect -20 582 -14 631
rect 20 582 26 631
rect -20 559 26 582
rect -20 514 -14 559
rect 20 514 26 559
rect -20 487 26 514
rect -20 446 -14 487
rect 20 446 26 487
rect -20 415 26 446
rect -20 378 -14 415
rect 20 378 26 415
rect -20 344 26 378
rect -20 309 -14 344
rect 20 309 26 344
rect -20 276 26 309
rect -20 237 -14 276
rect 20 237 26 276
rect 126 852 172 859
rect 126 847 134 852
rect 126 813 132 847
rect 168 818 172 852
rect 166 813 172 818
rect 126 784 172 813
rect 126 775 134 784
rect 126 741 132 775
rect 168 750 172 784
rect 166 741 172 750
rect 126 716 172 741
rect 126 703 134 716
rect 126 669 132 703
rect 168 682 172 716
rect 166 669 172 682
rect 126 648 172 669
rect 126 631 134 648
rect 126 597 132 631
rect 168 614 172 648
rect 166 597 172 614
rect 126 580 172 597
rect 126 559 134 580
rect 126 525 132 559
rect 168 546 172 580
rect 166 525 172 546
rect 126 512 172 525
rect 126 487 134 512
rect 126 453 132 487
rect 168 478 172 512
rect 166 453 172 478
rect 126 444 172 453
rect 126 415 134 444
rect 126 381 132 415
rect 168 410 172 444
rect 166 381 172 410
rect 126 376 172 381
rect 126 343 134 376
rect 126 309 132 343
rect 168 342 172 376
rect 166 309 172 342
rect 126 308 172 309
rect 126 274 134 308
rect 168 274 172 308
rect 126 269 172 274
rect 1785 852 1831 859
rect 1785 818 1790 852
rect 1824 847 1831 852
rect 1785 813 1791 818
rect 1825 813 1831 847
rect 1785 784 1831 813
rect 1785 750 1790 784
rect 1824 775 1831 784
rect 1785 741 1791 750
rect 1825 741 1831 775
rect 1785 716 1831 741
rect 1785 682 1790 716
rect 1824 703 1831 716
rect 1785 669 1791 682
rect 1825 669 1831 703
rect 1785 648 1831 669
rect 1785 614 1790 648
rect 1824 631 1831 648
rect 1785 597 1791 614
rect 1825 597 1831 631
rect 1785 580 1831 597
rect 1785 546 1790 580
rect 1824 559 1831 580
rect 1785 525 1791 546
rect 1825 525 1831 559
rect 1785 512 1831 525
rect 1785 478 1790 512
rect 1824 487 1831 512
rect 1785 453 1791 478
rect 1825 453 1831 487
rect 1785 444 1831 453
rect 1785 410 1790 444
rect 1824 415 1831 444
rect 1785 381 1791 410
rect 1825 381 1831 415
rect 1785 376 1831 381
rect 1785 342 1790 376
rect 1824 343 1831 376
rect 1785 309 1791 342
rect 1825 309 1831 343
rect 1785 308 1831 309
rect 1785 274 1790 308
rect 1824 274 1831 308
rect 1785 269 1831 274
rect 1932 854 1938 859
rect 1972 854 1978 859
rect 1932 847 1978 854
rect 1932 786 1938 847
rect 1972 786 1978 847
rect 1932 775 1978 786
rect 1932 718 1938 775
rect 1972 718 1978 775
rect 1932 703 1978 718
rect 1932 650 1938 703
rect 1972 650 1978 703
rect 1932 631 1978 650
rect 1932 582 1938 631
rect 1972 582 1978 631
rect 1932 559 1978 582
rect 1932 514 1938 559
rect 1972 514 1978 559
rect 1932 487 1978 514
rect 1932 446 1938 487
rect 1972 446 1978 487
rect 1932 415 1978 446
rect 1932 378 1938 415
rect 1972 378 1978 415
rect 1932 344 1978 378
rect 1932 309 1938 344
rect 1972 309 1978 344
rect 1932 276 1978 309
rect -20 208 26 237
rect -20 165 -14 208
rect 20 165 26 208
rect -20 140 26 165
rect -20 93 -14 140
rect 20 93 26 140
rect 134 240 168 269
rect 134 172 168 206
rect 134 122 168 138
rect 1790 240 1824 269
rect 1790 172 1824 206
rect 1790 122 1824 138
rect 1932 237 1938 276
rect 1972 237 1978 276
rect 1932 208 1978 237
rect 1932 165 1938 208
rect 1972 165 1978 208
rect 1932 140 1978 165
rect -20 58 26 93
rect 1932 93 1938 140
rect 1972 93 1978 140
rect 1932 58 1978 93
rect -20 52 1978 58
rect -20 18 20 52
rect 66 18 88 52
rect 138 18 156 52
rect 210 18 224 52
rect 282 18 292 52
rect 354 18 360 52
rect 426 18 428 52
rect 462 18 464 52
rect 530 18 536 52
rect 598 18 608 52
rect 666 18 680 52
rect 734 18 752 52
rect 802 18 824 52
rect 870 18 896 52
rect 938 18 968 52
rect 1006 18 1040 52
rect 1074 18 1108 52
rect 1146 18 1176 52
rect 1218 18 1244 52
rect 1290 18 1312 52
rect 1362 18 1380 52
rect 1434 18 1448 52
rect 1506 18 1516 52
rect 1578 18 1584 52
rect 1650 18 1652 52
rect 1686 18 1688 52
rect 1754 18 1760 52
rect 1822 18 1832 52
rect 1890 18 1978 52
rect -20 12 1978 18
<< viali >>
rect 32 1262 54 1296
rect 54 1262 66 1296
rect 104 1262 122 1296
rect 122 1262 138 1296
rect 176 1262 190 1296
rect 190 1262 210 1296
rect 248 1262 258 1296
rect 258 1262 282 1296
rect 320 1262 326 1296
rect 326 1262 354 1296
rect 392 1262 394 1296
rect 394 1262 426 1296
rect 464 1262 496 1296
rect 496 1262 498 1296
rect 536 1262 564 1296
rect 564 1262 570 1296
rect 608 1262 632 1296
rect 632 1262 642 1296
rect 680 1262 700 1296
rect 700 1262 714 1296
rect 752 1262 768 1296
rect 768 1262 786 1296
rect 824 1262 836 1296
rect 836 1262 858 1296
rect 896 1262 904 1296
rect 904 1262 930 1296
rect 968 1262 972 1296
rect 972 1262 1002 1296
rect 1040 1262 1074 1296
rect 1112 1262 1142 1296
rect 1142 1262 1146 1296
rect 1184 1262 1210 1296
rect 1210 1262 1218 1296
rect 1256 1262 1278 1296
rect 1278 1262 1290 1296
rect 1328 1262 1346 1296
rect 1346 1262 1362 1296
rect 1400 1262 1414 1296
rect 1414 1262 1434 1296
rect 1472 1262 1482 1296
rect 1482 1262 1506 1296
rect 1544 1262 1550 1296
rect 1550 1262 1578 1296
rect 1616 1262 1618 1296
rect 1618 1262 1650 1296
rect 1688 1262 1720 1296
rect 1720 1262 1722 1296
rect 1760 1262 1788 1296
rect 1788 1262 1794 1296
rect 1832 1262 1856 1296
rect 1856 1262 1866 1296
rect 191 1168 199 1202
rect 199 1168 225 1202
rect 263 1168 267 1202
rect 267 1168 297 1202
rect 335 1168 369 1202
rect 407 1168 437 1202
rect 437 1168 441 1202
rect 479 1168 505 1202
rect 505 1168 513 1202
rect 551 1168 573 1202
rect 573 1168 585 1202
rect 623 1168 641 1202
rect 641 1168 657 1202
rect 695 1168 709 1202
rect 709 1168 729 1202
rect 767 1168 777 1202
rect 777 1168 801 1202
rect 839 1168 845 1202
rect 845 1168 873 1202
rect 911 1168 913 1202
rect 913 1168 945 1202
rect 983 1168 1015 1202
rect 1015 1168 1017 1202
rect 1055 1168 1083 1202
rect 1083 1168 1089 1202
rect 1127 1168 1151 1202
rect 1151 1168 1161 1202
rect 1199 1168 1219 1202
rect 1219 1168 1233 1202
rect 1271 1168 1287 1202
rect 1287 1168 1305 1202
rect 1343 1168 1355 1202
rect 1355 1168 1377 1202
rect 1415 1168 1423 1202
rect 1423 1168 1449 1202
rect 1487 1168 1491 1202
rect 1491 1168 1521 1202
rect 1559 1168 1593 1202
rect 1631 1168 1661 1202
rect 1661 1168 1665 1202
rect 1703 1168 1729 1202
rect 1729 1168 1737 1202
rect -14 820 20 847
rect -14 813 20 820
rect -14 752 20 775
rect -14 741 20 752
rect -14 684 20 703
rect -14 669 20 684
rect -14 616 20 631
rect -14 597 20 616
rect -14 548 20 559
rect -14 525 20 548
rect -14 480 20 487
rect -14 453 20 480
rect -14 412 20 415
rect -14 381 20 412
rect -14 310 20 343
rect -14 309 20 310
rect -14 242 20 271
rect -14 237 20 242
rect 132 818 134 847
rect 134 818 166 847
rect 132 813 166 818
rect 132 750 134 775
rect 134 750 166 775
rect 132 741 166 750
rect 132 682 134 703
rect 134 682 166 703
rect 132 669 166 682
rect 132 614 134 631
rect 134 614 166 631
rect 132 597 166 614
rect 132 546 134 559
rect 134 546 166 559
rect 132 525 166 546
rect 132 478 134 487
rect 134 478 166 487
rect 132 453 166 478
rect 132 410 134 415
rect 134 410 166 415
rect 132 381 166 410
rect 132 342 134 343
rect 134 342 166 343
rect 132 309 166 342
rect 1791 818 1824 847
rect 1824 818 1825 847
rect 1791 813 1825 818
rect 1791 750 1824 775
rect 1824 750 1825 775
rect 1791 741 1825 750
rect 1791 682 1824 703
rect 1824 682 1825 703
rect 1791 669 1825 682
rect 1791 614 1824 631
rect 1824 614 1825 631
rect 1791 597 1825 614
rect 1791 546 1824 559
rect 1824 546 1825 559
rect 1791 525 1825 546
rect 1791 478 1824 487
rect 1824 478 1825 487
rect 1791 453 1825 478
rect 1791 410 1824 415
rect 1824 410 1825 415
rect 1791 381 1825 410
rect 1791 342 1824 343
rect 1824 342 1825 343
rect 1791 309 1825 342
rect 1938 820 1972 847
rect 1938 813 1972 820
rect 1938 752 1972 775
rect 1938 741 1972 752
rect 1938 684 1972 703
rect 1938 669 1972 684
rect 1938 616 1972 631
rect 1938 597 1972 616
rect 1938 548 1972 559
rect 1938 525 1972 548
rect 1938 480 1972 487
rect 1938 453 1972 480
rect 1938 412 1972 415
rect 1938 381 1972 412
rect 1938 310 1972 343
rect 1938 309 1972 310
rect -14 174 20 199
rect -14 165 20 174
rect -14 106 20 127
rect -14 93 20 106
rect 1938 242 1972 271
rect 1938 237 1972 242
rect 1938 174 1972 199
rect 1938 165 1972 174
rect 1938 106 1972 127
rect 1938 93 1972 106
rect 32 18 54 52
rect 54 18 66 52
rect 104 18 122 52
rect 122 18 138 52
rect 176 18 190 52
rect 190 18 210 52
rect 248 18 258 52
rect 258 18 282 52
rect 320 18 326 52
rect 326 18 354 52
rect 392 18 394 52
rect 394 18 426 52
rect 464 18 496 52
rect 496 18 498 52
rect 536 18 564 52
rect 564 18 570 52
rect 608 18 632 52
rect 632 18 642 52
rect 680 18 700 52
rect 700 18 714 52
rect 752 18 768 52
rect 768 18 786 52
rect 824 18 836 52
rect 836 18 858 52
rect 896 18 904 52
rect 904 18 930 52
rect 968 18 972 52
rect 972 18 1002 52
rect 1040 18 1074 52
rect 1112 18 1142 52
rect 1142 18 1146 52
rect 1184 18 1210 52
rect 1210 18 1218 52
rect 1256 18 1278 52
rect 1278 18 1290 52
rect 1328 18 1346 52
rect 1346 18 1362 52
rect 1400 18 1414 52
rect 1414 18 1434 52
rect 1472 18 1482 52
rect 1482 18 1506 52
rect 1544 18 1550 52
rect 1550 18 1578 52
rect 1616 18 1618 52
rect 1618 18 1650 52
rect 1688 18 1720 52
rect 1720 18 1722 52
rect 1760 18 1788 52
rect 1788 18 1794 52
rect 1832 18 1856 52
rect 1856 18 1866 52
<< metal1 >>
rect -14 1296 1972 1302
rect -14 1262 32 1296
rect 66 1262 104 1296
rect 138 1262 176 1296
rect 210 1262 248 1296
rect 282 1262 320 1296
rect 354 1262 392 1296
rect 426 1262 464 1296
rect 498 1262 536 1296
rect 570 1262 608 1296
rect 642 1262 680 1296
rect 714 1262 752 1296
rect 786 1262 824 1296
rect 858 1262 896 1296
rect 930 1262 968 1296
rect 1002 1262 1040 1296
rect 1074 1262 1112 1296
rect 1146 1262 1184 1296
rect 1218 1262 1256 1296
rect 1290 1262 1328 1296
rect 1362 1262 1400 1296
rect 1434 1262 1472 1296
rect 1506 1262 1544 1296
rect 1578 1262 1616 1296
rect 1650 1262 1688 1296
rect 1722 1262 1760 1296
rect 1794 1262 1832 1296
rect 1866 1262 1972 1296
rect -14 1256 1972 1262
rect -22 1202 1980 1211
rect -22 1168 191 1202
rect 225 1168 263 1202
rect 297 1168 335 1202
rect 369 1168 407 1202
rect 441 1168 479 1202
rect 513 1168 551 1202
rect 585 1168 623 1202
rect 657 1168 695 1202
rect 729 1168 767 1202
rect 801 1168 839 1202
rect 873 1168 911 1202
rect 945 1168 983 1202
rect 1017 1168 1055 1202
rect 1089 1168 1127 1202
rect 1161 1168 1199 1202
rect 1233 1168 1271 1202
rect 1305 1168 1343 1202
rect 1377 1168 1415 1202
rect 1449 1168 1487 1202
rect 1521 1168 1559 1202
rect 1593 1168 1631 1202
rect 1665 1168 1703 1202
rect 1737 1168 1980 1202
rect -22 1159 1980 1168
rect -20 847 1978 859
rect -20 813 -14 847
rect 20 813 132 847
rect 166 813 1791 847
rect 1825 813 1938 847
rect 1972 813 1978 847
rect -20 775 1978 813
rect -20 741 -14 775
rect 20 741 132 775
rect 166 741 1791 775
rect 1825 741 1938 775
rect 1972 741 1978 775
rect -20 703 1978 741
rect -20 669 -14 703
rect 20 669 132 703
rect 166 669 1791 703
rect 1825 669 1938 703
rect 1972 669 1978 703
rect -20 631 1978 669
rect -20 597 -14 631
rect 20 597 132 631
rect 166 597 1791 631
rect 1825 597 1938 631
rect 1972 597 1978 631
rect -20 559 1978 597
rect -20 525 -14 559
rect 20 525 132 559
rect 166 525 1791 559
rect 1825 525 1938 559
rect 1972 525 1978 559
rect -20 487 1978 525
rect -20 453 -14 487
rect 20 453 132 487
rect 166 453 1791 487
rect 1825 453 1938 487
rect 1972 453 1978 487
rect -20 415 1978 453
rect -20 381 -14 415
rect 20 381 132 415
rect 166 381 1791 415
rect 1825 381 1938 415
rect 1972 381 1978 415
rect -20 343 1978 381
rect -20 309 -14 343
rect 20 309 132 343
rect 166 309 1791 343
rect 1825 309 1938 343
rect 1972 309 1978 343
rect -20 271 1978 309
rect -20 237 -14 271
rect 20 269 1938 271
rect 20 237 28 269
tri 28 237 60 269 nw
tri 1898 237 1930 269 ne
rect 1930 237 1938 269
rect 1972 237 1978 271
rect -20 199 26 237
tri 26 235 28 237 nw
tri 1930 235 1932 237 ne
rect -20 165 -14 199
rect 20 165 26 199
rect -20 127 26 165
rect -20 93 -14 127
rect 20 93 26 127
rect -20 58 26 93
rect 1932 199 1978 237
rect 1932 165 1938 199
rect 1972 165 1978 199
rect 1932 127 1978 165
rect 1932 93 1938 127
rect 1972 93 1978 127
tri 26 58 60 92 sw
tri 1898 58 1932 92 se
rect 1932 58 1978 93
rect -20 52 1978 58
rect -20 18 32 52
rect 66 18 104 52
rect 138 18 176 52
rect 210 18 248 52
rect 282 18 320 52
rect 354 18 392 52
rect 426 18 464 52
rect 498 18 536 52
rect 570 18 608 52
rect 642 18 680 52
rect 714 18 752 52
rect 786 18 824 52
rect 858 18 896 52
rect 930 18 968 52
rect 1002 18 1040 52
rect 1074 18 1112 52
rect 1146 18 1184 52
rect 1218 18 1256 52
rect 1290 18 1328 52
rect 1362 18 1400 52
rect 1434 18 1472 52
rect 1506 18 1544 52
rect 1578 18 1616 52
rect 1650 18 1688 52
rect 1722 18 1760 52
rect 1794 18 1832 52
rect 1866 18 1978 52
rect -20 12 1978 18
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808680  sky130_fd_pr__model__nfet_highvoltage__example_55959141808680_0
timestamp 1666199351
transform 1 0 179 0 1 126
box -1 0 1601 1
<< properties >>
string GDS_END 11822256
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 11804982
<< end >>
