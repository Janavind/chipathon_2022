magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< obsli1 >>
rect 34 3292 1958 3358
rect 34 100 100 3292
rect 260 3066 1732 3132
rect 260 326 326 3066
rect 662 2664 1330 2730
rect 662 728 728 2664
rect 895 895 1097 2497
rect 1264 728 1330 2664
rect 662 662 1330 728
rect 1666 326 1732 3066
rect 260 260 1732 326
rect 1892 100 1958 3292
rect 34 34 1958 100
<< obsm1 >>
rect 38 3296 1954 3354
rect 38 96 96 3296
rect 264 3070 1728 3128
rect 264 322 322 3070
rect 666 2668 1326 2726
rect 666 724 724 2668
rect 895 911 1097 2481
rect 1268 724 1326 2668
rect 666 666 1326 724
rect 1670 322 1728 3070
rect 264 264 1728 322
rect 1896 96 1954 3296
rect 38 38 1954 96
<< properties >>
string FIXED_BBOX 26 26 1966 3366
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8872010
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8811326
<< end >>
