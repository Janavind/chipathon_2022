magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -66 377 1122 897
<< pwell >>
rect 4 43 1047 283
rect -26 -43 1082 43
<< mvnmos >>
rect 83 107 183 257
rect 419 107 519 257
rect 561 107 661 257
rect 722 107 822 257
rect 864 107 964 257
<< mvpmos >>
rect 87 443 187 743
rect 405 443 505 743
rect 561 443 661 743
rect 717 443 817 743
rect 873 443 973 743
<< mvndiff >>
rect 30 245 83 257
rect 30 211 38 245
rect 72 211 83 245
rect 30 153 83 211
rect 30 119 38 153
rect 72 119 83 153
rect 30 107 83 119
rect 183 249 419 257
rect 183 215 194 249
rect 228 215 286 249
rect 320 215 374 249
rect 408 215 419 249
rect 183 149 419 215
rect 183 115 194 149
rect 228 115 286 149
rect 320 115 374 149
rect 408 115 419 149
rect 183 107 419 115
rect 519 107 561 257
rect 661 249 722 257
rect 661 215 677 249
rect 711 215 722 249
rect 661 149 722 215
rect 661 115 677 149
rect 711 115 722 149
rect 661 107 722 115
rect 822 107 864 257
rect 964 249 1021 257
rect 964 215 975 249
rect 1009 215 1021 249
rect 964 149 1021 215
rect 964 115 975 149
rect 1009 115 1021 149
rect 964 107 1021 115
<< mvpdiff >>
rect 30 735 87 743
rect 30 701 42 735
rect 76 701 87 735
rect 30 652 87 701
rect 30 618 42 652
rect 76 618 87 652
rect 30 568 87 618
rect 30 534 42 568
rect 76 534 87 568
rect 30 485 87 534
rect 30 451 42 485
rect 76 451 87 485
rect 30 443 87 451
rect 187 735 244 743
rect 187 701 198 735
rect 232 701 244 735
rect 187 652 244 701
rect 187 618 198 652
rect 232 618 244 652
rect 187 568 244 618
rect 187 534 198 568
rect 232 534 244 568
rect 187 485 244 534
rect 187 451 198 485
rect 232 451 244 485
rect 187 443 244 451
rect 316 735 405 743
rect 316 701 328 735
rect 362 701 405 735
rect 316 652 405 701
rect 316 618 328 652
rect 362 618 405 652
rect 316 568 405 618
rect 316 534 328 568
rect 362 534 405 568
rect 316 485 405 534
rect 316 451 328 485
rect 362 451 405 485
rect 316 443 405 451
rect 505 691 561 743
rect 505 657 516 691
rect 550 657 561 691
rect 505 623 561 657
rect 505 589 516 623
rect 550 589 561 623
rect 505 553 561 589
rect 505 519 516 553
rect 550 519 561 553
rect 505 485 561 519
rect 505 451 516 485
rect 550 451 561 485
rect 505 443 561 451
rect 661 735 717 743
rect 661 701 672 735
rect 706 701 717 735
rect 661 652 717 701
rect 661 618 672 652
rect 706 618 717 652
rect 661 568 717 618
rect 661 534 672 568
rect 706 534 717 568
rect 661 485 717 534
rect 661 451 672 485
rect 706 451 717 485
rect 661 443 717 451
rect 817 735 873 743
rect 817 701 828 735
rect 862 701 873 735
rect 817 654 873 701
rect 817 620 828 654
rect 862 620 873 654
rect 817 571 873 620
rect 817 537 828 571
rect 862 537 873 571
rect 817 490 873 537
rect 817 456 828 490
rect 862 456 873 490
rect 817 443 873 456
rect 973 731 1026 743
rect 973 697 984 731
rect 1018 697 1026 731
rect 973 651 1026 697
rect 973 617 984 651
rect 1018 617 1026 651
rect 973 569 1026 617
rect 973 535 984 569
rect 1018 535 1026 569
rect 973 489 1026 535
rect 973 455 984 489
rect 1018 455 1026 489
rect 973 443 1026 455
<< mvndiffc >>
rect 38 211 72 245
rect 38 119 72 153
rect 194 215 228 249
rect 286 215 320 249
rect 374 215 408 249
rect 194 115 228 149
rect 286 115 320 149
rect 374 115 408 149
rect 677 215 711 249
rect 677 115 711 149
rect 975 215 1009 249
rect 975 115 1009 149
<< mvpdiffc >>
rect 42 701 76 735
rect 42 618 76 652
rect 42 534 76 568
rect 42 451 76 485
rect 198 701 232 735
rect 198 618 232 652
rect 198 534 232 568
rect 198 451 232 485
rect 328 701 362 735
rect 328 618 362 652
rect 328 534 362 568
rect 328 451 362 485
rect 516 657 550 691
rect 516 589 550 623
rect 516 519 550 553
rect 516 451 550 485
rect 672 701 706 735
rect 672 618 706 652
rect 672 534 706 568
rect 672 451 706 485
rect 828 701 862 735
rect 828 620 862 654
rect 828 537 862 571
rect 828 456 862 490
rect 984 697 1018 731
rect 984 617 1018 651
rect 984 535 1018 569
rect 984 455 1018 489
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
<< poly >>
rect 87 743 187 769
rect 405 743 505 769
rect 561 743 661 769
rect 717 743 817 769
rect 873 743 973 769
rect 87 421 187 443
rect 83 335 187 421
rect 405 417 505 443
rect 83 301 133 335
rect 167 301 187 335
rect 83 279 187 301
rect 394 395 519 417
rect 394 361 414 395
rect 448 361 519 395
rect 394 283 519 361
rect 83 257 183 279
rect 419 257 519 283
rect 561 334 661 443
rect 561 300 607 334
rect 641 300 661 334
rect 561 257 661 300
rect 717 417 817 443
rect 873 417 973 443
rect 717 343 822 417
rect 717 309 737 343
rect 771 309 822 343
rect 717 283 822 309
rect 722 257 822 283
rect 864 343 1035 417
rect 864 309 981 343
rect 1015 309 1035 343
rect 864 283 1035 309
rect 864 257 964 283
rect 83 81 183 107
rect 419 81 519 107
rect 561 81 661 107
rect 722 81 822 107
rect 864 81 964 107
<< polycont >>
rect 133 301 167 335
rect 414 361 448 395
rect 607 300 641 334
rect 737 309 771 343
rect 981 309 1015 343
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 21 735 76 751
rect 21 701 42 735
rect 21 652 76 701
rect 21 618 42 652
rect 21 568 76 618
rect 21 534 42 568
rect 21 485 76 534
rect 21 451 42 485
rect 21 245 76 451
rect 112 735 292 751
rect 112 701 113 735
rect 147 701 185 735
rect 232 701 257 735
rect 291 701 292 735
rect 112 652 292 701
rect 112 618 198 652
rect 232 618 292 652
rect 112 568 292 618
rect 112 534 198 568
rect 232 534 292 568
rect 112 485 292 534
rect 112 451 198 485
rect 232 451 292 485
rect 112 435 292 451
rect 328 735 706 761
rect 362 727 672 735
rect 328 652 362 701
rect 656 701 672 727
rect 500 657 516 691
rect 550 657 566 691
rect 328 568 362 618
rect 328 485 362 534
rect 328 435 362 451
rect 398 395 464 652
rect 398 361 414 395
rect 448 361 464 395
rect 398 355 464 361
rect 500 623 566 657
rect 500 589 516 623
rect 550 589 566 623
rect 500 553 566 589
rect 500 519 516 553
rect 550 519 566 553
rect 500 485 566 519
rect 500 451 516 485
rect 550 451 566 485
rect 117 335 183 351
rect 117 301 133 335
rect 167 319 183 335
rect 500 319 566 451
rect 656 652 706 701
rect 656 618 672 652
rect 656 568 706 618
rect 656 534 672 568
rect 656 485 706 534
rect 656 451 672 485
rect 742 735 932 751
rect 742 701 748 735
rect 782 701 820 735
rect 862 701 892 735
rect 926 701 932 735
rect 742 654 932 701
rect 742 620 828 654
rect 862 620 932 654
rect 742 571 932 620
rect 742 537 828 571
rect 862 537 932 571
rect 742 490 932 537
rect 742 456 828 490
rect 862 456 932 490
rect 968 731 1034 747
rect 968 697 984 731
rect 1018 697 1034 731
rect 968 651 1034 697
rect 968 617 984 651
rect 1018 617 1034 651
rect 968 569 1034 617
rect 968 535 984 569
rect 1018 535 1034 569
rect 968 489 1034 535
rect 656 420 706 451
rect 968 455 984 489
rect 1018 455 1034 489
rect 968 420 1034 455
rect 656 386 1034 420
rect 607 334 641 350
rect 167 301 571 319
rect 117 285 571 301
rect 21 211 38 245
rect 72 211 76 245
rect 21 153 76 211
rect 21 119 38 153
rect 72 119 76 153
rect 21 99 76 119
rect 110 215 194 249
rect 228 215 286 249
rect 320 215 374 249
rect 408 215 452 249
rect 110 149 452 215
rect 110 115 194 149
rect 228 115 286 149
rect 320 115 374 149
rect 408 115 452 149
rect 110 113 452 115
rect 110 79 120 113
rect 154 79 192 113
rect 226 79 264 113
rect 298 79 336 113
rect 370 79 408 113
rect 442 79 452 113
rect 537 126 571 285
rect 697 343 929 350
rect 697 309 737 343
rect 771 309 929 343
rect 697 301 929 309
rect 965 343 1031 350
rect 965 309 981 343
rect 1015 309 1031 343
rect 965 301 1031 309
rect 607 162 641 300
rect 677 249 727 265
rect 711 215 727 249
rect 677 149 727 215
rect 537 115 677 126
rect 711 115 727 149
rect 537 92 727 115
rect 763 249 1025 265
rect 763 215 975 249
rect 1009 215 1025 249
rect 763 149 1025 215
rect 763 115 975 149
rect 1009 115 1025 149
rect 763 113 1025 115
rect 110 73 452 79
rect 763 79 769 113
rect 803 79 841 113
rect 875 79 913 113
rect 947 79 985 113
rect 1019 79 1025 113
rect 763 73 1025 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 113 701 147 735
rect 185 701 198 735
rect 198 701 219 735
rect 257 701 291 735
rect 748 701 782 735
rect 820 701 828 735
rect 828 701 854 735
rect 892 701 926 735
rect 120 79 154 113
rect 192 79 226 113
rect 264 79 298 113
rect 336 79 370 113
rect 408 79 442 113
rect 769 79 803 113
rect 841 79 875 113
rect 913 79 947 113
rect 985 79 1019 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 831 1056 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 0 791 1056 797
rect 0 735 1056 763
rect 0 701 113 735
rect 147 701 185 735
rect 219 701 257 735
rect 291 701 748 735
rect 782 701 820 735
rect 854 701 892 735
rect 926 701 1056 735
rect 0 689 1056 701
rect 0 113 1056 125
rect 0 79 120 113
rect 154 79 192 113
rect 226 79 264 113
rect 298 79 336 113
rect 370 79 408 113
rect 442 79 769 113
rect 803 79 841 113
rect 875 79 913 113
rect 947 79 985 113
rect 1019 79 1056 113
rect 0 51 1056 79
rect 0 17 1056 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -23 1056 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a22o_1
flabel metal1 s 0 51 1056 125 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 0 0 1056 23 0 FreeSans 340 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 0 689 1056 763 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 791 1056 814 0 FreeSans 340 0 0 0 VPB
port 7 nsew power bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 415 612 449 646 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 612 65 646 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1056 814
string GDS_END 783842
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 769994
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
