magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect 0 0 466 672
<< pmos >>
rect 89 36 119 636
rect 175 36 205 636
rect 261 36 291 636
rect 347 36 377 636
<< pdiff >>
rect 36 605 89 636
rect 36 571 44 605
rect 78 571 89 605
rect 36 533 89 571
rect 36 499 44 533
rect 78 499 89 533
rect 36 461 89 499
rect 36 427 44 461
rect 78 427 89 461
rect 36 389 89 427
rect 36 355 44 389
rect 78 355 89 389
rect 36 317 89 355
rect 36 283 44 317
rect 78 283 89 317
rect 36 245 89 283
rect 36 211 44 245
rect 78 211 89 245
rect 36 173 89 211
rect 36 139 44 173
rect 78 139 89 173
rect 36 101 89 139
rect 36 67 44 101
rect 78 67 89 101
rect 36 36 89 67
rect 119 605 175 636
rect 119 571 130 605
rect 164 571 175 605
rect 119 533 175 571
rect 119 499 130 533
rect 164 499 175 533
rect 119 461 175 499
rect 119 427 130 461
rect 164 427 175 461
rect 119 389 175 427
rect 119 355 130 389
rect 164 355 175 389
rect 119 317 175 355
rect 119 283 130 317
rect 164 283 175 317
rect 119 245 175 283
rect 119 211 130 245
rect 164 211 175 245
rect 119 173 175 211
rect 119 139 130 173
rect 164 139 175 173
rect 119 101 175 139
rect 119 67 130 101
rect 164 67 175 101
rect 119 36 175 67
rect 205 605 261 636
rect 205 571 216 605
rect 250 571 261 605
rect 205 533 261 571
rect 205 499 216 533
rect 250 499 261 533
rect 205 461 261 499
rect 205 427 216 461
rect 250 427 261 461
rect 205 389 261 427
rect 205 355 216 389
rect 250 355 261 389
rect 205 317 261 355
rect 205 283 216 317
rect 250 283 261 317
rect 205 245 261 283
rect 205 211 216 245
rect 250 211 261 245
rect 205 173 261 211
rect 205 139 216 173
rect 250 139 261 173
rect 205 101 261 139
rect 205 67 216 101
rect 250 67 261 101
rect 205 36 261 67
rect 291 605 347 636
rect 291 571 302 605
rect 336 571 347 605
rect 291 533 347 571
rect 291 499 302 533
rect 336 499 347 533
rect 291 461 347 499
rect 291 427 302 461
rect 336 427 347 461
rect 291 389 347 427
rect 291 355 302 389
rect 336 355 347 389
rect 291 317 347 355
rect 291 283 302 317
rect 336 283 347 317
rect 291 245 347 283
rect 291 211 302 245
rect 336 211 347 245
rect 291 173 347 211
rect 291 139 302 173
rect 336 139 347 173
rect 291 101 347 139
rect 291 67 302 101
rect 336 67 347 101
rect 291 36 347 67
rect 377 605 430 636
rect 377 571 388 605
rect 422 571 430 605
rect 377 533 430 571
rect 377 499 388 533
rect 422 499 430 533
rect 377 461 430 499
rect 377 427 388 461
rect 422 427 430 461
rect 377 389 430 427
rect 377 355 388 389
rect 422 355 430 389
rect 377 317 430 355
rect 377 283 388 317
rect 422 283 430 317
rect 377 245 430 283
rect 377 211 388 245
rect 422 211 430 245
rect 377 173 430 211
rect 377 139 388 173
rect 422 139 430 173
rect 377 101 430 139
rect 377 67 388 101
rect 422 67 430 101
rect 377 36 430 67
<< pdiffc >>
rect 44 571 78 605
rect 44 499 78 533
rect 44 427 78 461
rect 44 355 78 389
rect 44 283 78 317
rect 44 211 78 245
rect 44 139 78 173
rect 44 67 78 101
rect 130 571 164 605
rect 130 499 164 533
rect 130 427 164 461
rect 130 355 164 389
rect 130 283 164 317
rect 130 211 164 245
rect 130 139 164 173
rect 130 67 164 101
rect 216 571 250 605
rect 216 499 250 533
rect 216 427 250 461
rect 216 355 250 389
rect 216 283 250 317
rect 216 211 250 245
rect 216 139 250 173
rect 216 67 250 101
rect 302 571 336 605
rect 302 499 336 533
rect 302 427 336 461
rect 302 355 336 389
rect 302 283 336 317
rect 302 211 336 245
rect 302 139 336 173
rect 302 67 336 101
rect 388 571 422 605
rect 388 499 422 533
rect 388 427 422 461
rect 388 355 422 389
rect 388 283 422 317
rect 388 211 422 245
rect 388 139 422 173
rect 388 67 422 101
<< poly >>
rect 89 719 377 735
rect 89 685 114 719
rect 148 685 182 719
rect 216 685 250 719
rect 284 685 318 719
rect 352 685 377 719
rect 89 662 377 685
rect 89 636 119 662
rect 175 636 205 662
rect 261 636 291 662
rect 347 636 377 662
rect 89 10 119 36
rect 175 10 205 36
rect 261 10 291 36
rect 347 10 377 36
<< polycont >>
rect 114 685 148 719
rect 182 685 216 719
rect 250 685 284 719
rect 318 685 352 719
<< locali >>
rect 98 719 368 735
rect 98 685 108 719
rect 148 685 180 719
rect 216 685 250 719
rect 286 685 318 719
rect 358 685 368 719
rect 98 667 368 685
rect 44 605 78 621
rect 44 533 78 571
rect 44 461 78 499
rect 44 389 78 427
rect 44 317 78 355
rect 44 245 78 283
rect 44 173 78 211
rect 44 101 78 139
rect 44 51 78 67
rect 130 605 164 621
rect 130 533 164 571
rect 130 461 164 499
rect 130 389 164 427
rect 130 317 164 355
rect 130 245 164 283
rect 130 173 164 211
rect 130 101 164 139
rect 130 51 164 67
rect 216 605 250 621
rect 216 533 250 571
rect 216 461 250 499
rect 216 389 250 427
rect 216 317 250 355
rect 216 245 250 283
rect 216 173 250 211
rect 216 101 250 139
rect 216 51 250 67
rect 302 605 336 621
rect 302 533 336 571
rect 302 461 336 499
rect 302 389 336 427
rect 302 317 336 355
rect 302 245 336 283
rect 302 173 336 211
rect 302 101 336 139
rect 302 51 336 67
rect 388 605 422 621
rect 388 533 422 571
rect 388 461 422 499
rect 388 389 422 427
rect 388 317 422 355
rect 388 245 422 283
rect 388 173 422 211
rect 388 101 422 139
rect 388 51 422 67
<< viali >>
rect 108 685 114 719
rect 114 685 142 719
rect 180 685 182 719
rect 182 685 214 719
rect 252 685 284 719
rect 284 685 286 719
rect 324 685 352 719
rect 352 685 358 719
rect 44 571 78 605
rect 44 499 78 533
rect 44 427 78 461
rect 44 355 78 389
rect 44 283 78 317
rect 44 211 78 245
rect 44 139 78 173
rect 44 67 78 101
rect 130 571 164 605
rect 130 499 164 533
rect 130 427 164 461
rect 130 355 164 389
rect 130 283 164 317
rect 130 211 164 245
rect 130 139 164 173
rect 130 67 164 101
rect 216 571 250 605
rect 216 499 250 533
rect 216 427 250 461
rect 216 355 250 389
rect 216 283 250 317
rect 216 211 250 245
rect 216 139 250 173
rect 216 67 250 101
rect 302 571 336 605
rect 302 499 336 533
rect 302 427 336 461
rect 302 355 336 389
rect 302 283 336 317
rect 302 211 336 245
rect 302 139 336 173
rect 302 67 336 101
rect 388 571 422 605
rect 388 499 422 533
rect 388 427 422 461
rect 388 355 422 389
rect 388 283 422 317
rect 388 211 422 245
rect 388 139 422 173
rect 388 67 422 101
<< metal1 >>
rect 96 719 370 731
rect 96 685 108 719
rect 142 685 180 719
rect 214 685 252 719
rect 286 685 324 719
rect 358 685 370 719
rect 96 673 370 685
rect 38 605 84 621
rect 38 571 44 605
rect 78 571 84 605
rect 38 533 84 571
rect 38 499 44 533
rect 78 499 84 533
rect 38 461 84 499
rect 38 427 44 461
rect 78 427 84 461
rect 38 389 84 427
rect 38 355 44 389
rect 78 355 84 389
rect 38 317 84 355
rect 38 283 44 317
rect 78 283 84 317
rect 38 245 84 283
rect 38 211 44 245
rect 78 211 84 245
rect 38 173 84 211
rect 38 139 44 173
rect 78 139 84 173
rect 38 101 84 139
rect 38 67 44 101
rect 78 67 84 101
rect 38 -29 84 67
rect 121 610 173 621
rect 121 546 173 558
rect 121 461 173 494
rect 121 427 130 461
rect 164 427 173 461
rect 121 389 173 427
rect 121 355 130 389
rect 164 355 173 389
rect 121 317 173 355
rect 121 283 130 317
rect 164 283 173 317
rect 121 245 173 283
rect 121 211 130 245
rect 164 211 173 245
rect 121 173 173 211
rect 121 139 130 173
rect 164 139 173 173
rect 121 101 173 139
rect 121 67 130 101
rect 164 67 173 101
rect 121 51 173 67
rect 210 605 256 621
rect 210 571 216 605
rect 250 571 256 605
rect 210 533 256 571
rect 210 499 216 533
rect 250 499 256 533
rect 210 461 256 499
rect 210 427 216 461
rect 250 427 256 461
rect 210 389 256 427
rect 210 355 216 389
rect 250 355 256 389
rect 210 317 256 355
rect 210 283 216 317
rect 250 283 256 317
rect 210 245 256 283
rect 210 211 216 245
rect 250 211 256 245
rect 210 173 256 211
rect 210 139 216 173
rect 250 139 256 173
rect 210 101 256 139
rect 210 67 216 101
rect 250 67 256 101
rect 210 -29 256 67
rect 293 610 345 621
rect 293 546 345 558
rect 293 461 345 494
rect 293 427 302 461
rect 336 427 345 461
rect 293 389 345 427
rect 293 355 302 389
rect 336 355 345 389
rect 293 317 345 355
rect 293 283 302 317
rect 336 283 345 317
rect 293 245 345 283
rect 293 211 302 245
rect 336 211 345 245
rect 293 173 345 211
rect 293 139 302 173
rect 336 139 345 173
rect 293 101 345 139
rect 293 67 302 101
rect 336 67 345 101
rect 293 51 345 67
rect 382 605 428 621
rect 382 571 388 605
rect 422 571 428 605
rect 382 533 428 571
rect 382 499 388 533
rect 422 499 428 533
rect 382 461 428 499
rect 382 427 388 461
rect 422 427 428 461
rect 382 389 428 427
rect 382 355 388 389
rect 422 355 428 389
rect 382 317 428 355
rect 382 283 388 317
rect 422 283 428 317
rect 382 245 428 283
rect 382 211 388 245
rect 422 211 428 245
rect 382 173 428 211
rect 382 139 388 173
rect 422 139 428 173
rect 382 101 428 139
rect 382 67 388 101
rect 422 67 428 101
rect 382 -29 428 67
rect 38 -89 428 -29
<< via1 >>
rect 121 605 173 610
rect 121 571 130 605
rect 130 571 164 605
rect 164 571 173 605
rect 121 558 173 571
rect 121 533 173 546
rect 121 499 130 533
rect 130 499 164 533
rect 164 499 173 533
rect 121 494 173 499
rect 293 605 345 610
rect 293 571 302 605
rect 302 571 336 605
rect 336 571 345 605
rect 293 558 345 571
rect 293 533 345 546
rect 293 499 302 533
rect 302 499 336 533
rect 336 499 345 533
rect 293 494 345 499
<< metal2 >>
rect 114 620 180 629
rect 114 564 119 620
rect 175 564 180 620
rect 114 558 121 564
rect 173 558 180 564
rect 114 546 180 558
rect 114 540 121 546
rect 173 540 180 546
rect 114 484 119 540
rect 175 484 180 540
rect 114 475 180 484
rect 286 620 352 629
rect 286 564 291 620
rect 347 564 352 620
rect 286 558 293 564
rect 345 558 352 564
rect 286 546 352 558
rect 286 540 293 546
rect 345 540 352 546
rect 286 484 291 540
rect 347 484 352 540
rect 286 475 352 484
<< via2 >>
rect 119 610 175 620
rect 119 564 121 610
rect 121 564 173 610
rect 173 564 175 610
rect 119 494 121 540
rect 121 494 173 540
rect 173 494 175 540
rect 119 484 175 494
rect 291 610 347 620
rect 291 564 293 610
rect 293 564 345 610
rect 345 564 347 610
rect 291 494 293 540
rect 293 494 345 540
rect 345 494 347 540
rect 291 484 347 494
<< metal3 >>
rect 114 620 352 629
rect 114 564 119 620
rect 175 564 291 620
rect 347 564 352 620
rect 114 563 352 564
rect 114 540 180 563
rect 114 484 119 540
rect 175 484 180 540
rect 114 475 180 484
rect 286 540 352 563
rect 286 484 291 540
rect 347 484 352 540
rect 286 475 352 484
<< labels >>
flabel metal3 s 114 563 352 629 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 96 673 370 731 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel metal1 s 38 -89 428 -29 0 FreeSans 400 0 0 0 SOURCE
port 3 nsew
flabel nwell s 84 663 88 671 0 FreeSans 400 0 0 0 BULK
port 4 nsew
<< properties >>
string GDS_END 9148738
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9138218
string path 0.950 -1.475 10.700 -1.475 
<< end >>
