magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< metal4 >>
rect -3360 39427 -2720 39451
rect 24000 39427 24640 39451
rect -3360 39416 24640 39427
rect -3360 39180 -3087 39416
rect -2851 39180 -2765 39416
rect -2529 39180 -2443 39416
rect -2207 39180 -2121 39416
rect -1885 39180 -1799 39416
rect -1563 39180 -1477 39416
rect -1241 39180 -1155 39416
rect -919 39180 -833 39416
rect -597 39180 -511 39416
rect -275 39180 -189 39416
rect 47 39180 133 39416
rect 369 39180 455 39416
rect 691 39180 777 39416
rect 1013 39180 1099 39416
rect 1335 39180 1421 39416
rect 1657 39180 1743 39416
rect 1979 39180 2065 39416
rect 2301 39180 2387 39416
rect 2623 39180 2709 39416
rect 2945 39180 3031 39416
rect 3267 39180 3353 39416
rect 3589 39180 3675 39416
rect 3911 39180 3997 39416
rect 4233 39180 4318 39416
rect 4554 39180 4639 39416
rect 4875 39180 4960 39416
rect 5196 39180 5281 39416
rect 5517 39180 5602 39416
rect 5838 39180 5923 39416
rect 6159 39180 6244 39416
rect 6480 39180 6565 39416
rect 6801 39180 6886 39416
rect 7122 39180 7207 39416
rect 7443 39180 7528 39416
rect 7764 39180 7849 39416
rect 8085 39180 8170 39416
rect 8406 39180 8491 39416
rect 8727 39180 8812 39416
rect 9048 39180 9133 39416
rect 9369 39180 9454 39416
rect 9690 39180 9775 39416
rect 10011 39180 10096 39416
rect 10332 39180 10417 39416
rect 10653 39180 10738 39416
rect 10974 39180 11059 39416
rect 11295 39180 11380 39416
rect 11616 39180 11701 39416
rect 11937 39180 12022 39416
rect 12258 39180 12343 39416
rect 12579 39180 12664 39416
rect 12900 39180 12985 39416
rect 13221 39180 13306 39416
rect 13542 39180 13627 39416
rect 13863 39180 13948 39416
rect 14184 39180 14269 39416
rect 14505 39180 14590 39416
rect 14826 39180 14911 39416
rect 15147 39180 15232 39416
rect 15468 39180 15553 39416
rect 15789 39180 15874 39416
rect 16110 39180 16195 39416
rect 16431 39180 16516 39416
rect 16752 39180 16837 39416
rect 17073 39180 17158 39416
rect 17394 39180 17479 39416
rect 17715 39180 17800 39416
rect 18036 39180 18121 39416
rect 18357 39180 18442 39416
rect 18678 39180 18763 39416
rect 18999 39180 19084 39416
rect 19320 39180 19405 39416
rect 19641 39180 19726 39416
rect 19962 39180 20047 39416
rect 20283 39180 20368 39416
rect 20604 39180 20689 39416
rect 20925 39180 21010 39416
rect 21246 39180 21331 39416
rect 21567 39180 21652 39416
rect 21888 39180 21973 39416
rect 22209 39180 22294 39416
rect 22530 39180 22615 39416
rect 22851 39180 22936 39416
rect 23172 39180 23257 39416
rect 23493 39180 23578 39416
rect 23814 39180 23899 39416
rect 24135 39180 24220 39416
rect 24456 39180 24640 39416
rect -3360 39092 24640 39180
rect -3360 38856 -3087 39092
rect -2851 38856 -2765 39092
rect -2529 38856 -2443 39092
rect -2207 38856 -2121 39092
rect -1885 38856 -1799 39092
rect -1563 38856 -1477 39092
rect -1241 38856 -1155 39092
rect -919 38856 -833 39092
rect -597 38856 -511 39092
rect -275 38856 -189 39092
rect 47 38856 133 39092
rect 369 38856 455 39092
rect 691 38856 777 39092
rect 1013 38856 1099 39092
rect 1335 38856 1421 39092
rect 1657 38856 1743 39092
rect 1979 38856 2065 39092
rect 2301 38856 2387 39092
rect 2623 38856 2709 39092
rect 2945 38856 3031 39092
rect 3267 38856 3353 39092
rect 3589 38856 3675 39092
rect 3911 38856 3997 39092
rect 4233 38856 4318 39092
rect 4554 38856 4639 39092
rect 4875 38856 4960 39092
rect 5196 38856 5281 39092
rect 5517 38856 5602 39092
rect 5838 38856 5923 39092
rect 6159 38856 6244 39092
rect 6480 38856 6565 39092
rect 6801 38856 6886 39092
rect 7122 38856 7207 39092
rect 7443 38856 7528 39092
rect 7764 38856 7849 39092
rect 8085 38856 8170 39092
rect 8406 38856 8491 39092
rect 8727 38856 8812 39092
rect 9048 38856 9133 39092
rect 9369 38856 9454 39092
rect 9690 38856 9775 39092
rect 10011 38856 10096 39092
rect 10332 38856 10417 39092
rect 10653 38856 10738 39092
rect 10974 38856 11059 39092
rect 11295 38856 11380 39092
rect 11616 38856 11701 39092
rect 11937 38856 12022 39092
rect 12258 38856 12343 39092
rect 12579 38856 12664 39092
rect 12900 38856 12985 39092
rect 13221 38856 13306 39092
rect 13542 38856 13627 39092
rect 13863 38856 13948 39092
rect 14184 38856 14269 39092
rect 14505 38856 14590 39092
rect 14826 38856 14911 39092
rect 15147 38856 15232 39092
rect 15468 38856 15553 39092
rect 15789 38856 15874 39092
rect 16110 38856 16195 39092
rect 16431 38856 16516 39092
rect 16752 38856 16837 39092
rect 17073 38856 17158 39092
rect 17394 38856 17479 39092
rect 17715 38856 17800 39092
rect 18036 38856 18121 39092
rect 18357 38856 18442 39092
rect 18678 38856 18763 39092
rect 18999 38856 19084 39092
rect 19320 38856 19405 39092
rect 19641 38856 19726 39092
rect 19962 38856 20047 39092
rect 20283 38856 20368 39092
rect 20604 38856 20689 39092
rect 20925 38856 21010 39092
rect 21246 38856 21331 39092
rect 21567 38856 21652 39092
rect 21888 38856 21973 39092
rect 22209 38856 22294 39092
rect 22530 38856 22615 39092
rect 22851 38856 22936 39092
rect 23172 38856 23257 39092
rect 23493 38856 23578 39092
rect 23814 38856 23899 39092
rect 24135 38856 24220 39092
rect 24456 38856 24640 39092
rect -3360 38768 24640 38856
rect -3360 38532 -3087 38768
rect -2851 38532 -2765 38768
rect -2529 38532 -2443 38768
rect -2207 38532 -2121 38768
rect -1885 38532 -1799 38768
rect -1563 38532 -1477 38768
rect -1241 38532 -1155 38768
rect -919 38532 -833 38768
rect -597 38532 -511 38768
rect -275 38532 -189 38768
rect 47 38532 133 38768
rect 369 38532 455 38768
rect 691 38532 777 38768
rect 1013 38532 1099 38768
rect 1335 38532 1421 38768
rect 1657 38532 1743 38768
rect 1979 38532 2065 38768
rect 2301 38532 2387 38768
rect 2623 38532 2709 38768
rect 2945 38532 3031 38768
rect 3267 38532 3353 38768
rect 3589 38532 3675 38768
rect 3911 38532 3997 38768
rect 4233 38532 4318 38768
rect 4554 38532 4639 38768
rect 4875 38532 4960 38768
rect 5196 38532 5281 38768
rect 5517 38532 5602 38768
rect 5838 38532 5923 38768
rect 6159 38532 6244 38768
rect 6480 38532 6565 38768
rect 6801 38532 6886 38768
rect 7122 38532 7207 38768
rect 7443 38532 7528 38768
rect 7764 38532 7849 38768
rect 8085 38532 8170 38768
rect 8406 38532 8491 38768
rect 8727 38532 8812 38768
rect 9048 38532 9133 38768
rect 9369 38532 9454 38768
rect 9690 38532 9775 38768
rect 10011 38532 10096 38768
rect 10332 38532 10417 38768
rect 10653 38532 10738 38768
rect 10974 38532 11059 38768
rect 11295 38532 11380 38768
rect 11616 38532 11701 38768
rect 11937 38532 12022 38768
rect 12258 38532 12343 38768
rect 12579 38532 12664 38768
rect 12900 38532 12985 38768
rect 13221 38532 13306 38768
rect 13542 38532 13627 38768
rect 13863 38532 13948 38768
rect 14184 38532 14269 38768
rect 14505 38532 14590 38768
rect 14826 38532 14911 38768
rect 15147 38532 15232 38768
rect 15468 38532 15553 38768
rect 15789 38532 15874 38768
rect 16110 38532 16195 38768
rect 16431 38532 16516 38768
rect 16752 38532 16837 38768
rect 17073 38532 17158 38768
rect 17394 38532 17479 38768
rect 17715 38532 17800 38768
rect 18036 38532 18121 38768
rect 18357 38532 18442 38768
rect 18678 38532 18763 38768
rect 18999 38532 19084 38768
rect 19320 38532 19405 38768
rect 19641 38532 19726 38768
rect 19962 38532 20047 38768
rect 20283 38532 20368 38768
rect 20604 38532 20689 38768
rect 20925 38532 21010 38768
rect 21246 38532 21331 38768
rect 21567 38532 21652 38768
rect 21888 38532 21973 38768
rect 22209 38532 22294 38768
rect 22530 38532 22615 38768
rect 22851 38532 22936 38768
rect 23172 38532 23257 38768
rect 23493 38532 23578 38768
rect 23814 38532 23899 38768
rect 24135 38532 24220 38768
rect 24456 38532 24640 38768
rect -3360 38444 24640 38532
rect -3360 38208 -3087 38444
rect -2851 38208 -2765 38444
rect -2529 38208 -2443 38444
rect -2207 38208 -2121 38444
rect -1885 38208 -1799 38444
rect -1563 38208 -1477 38444
rect -1241 38208 -1155 38444
rect -919 38208 -833 38444
rect -597 38208 -511 38444
rect -275 38208 -189 38444
rect 47 38208 133 38444
rect 369 38208 455 38444
rect 691 38208 777 38444
rect 1013 38208 1099 38444
rect 1335 38208 1421 38444
rect 1657 38208 1743 38444
rect 1979 38208 2065 38444
rect 2301 38208 2387 38444
rect 2623 38208 2709 38444
rect 2945 38208 3031 38444
rect 3267 38208 3353 38444
rect 3589 38208 3675 38444
rect 3911 38208 3997 38444
rect 4233 38208 4318 38444
rect 4554 38208 4639 38444
rect 4875 38208 4960 38444
rect 5196 38208 5281 38444
rect 5517 38208 5602 38444
rect 5838 38208 5923 38444
rect 6159 38208 6244 38444
rect 6480 38208 6565 38444
rect 6801 38208 6886 38444
rect 7122 38208 7207 38444
rect 7443 38208 7528 38444
rect 7764 38208 7849 38444
rect 8085 38208 8170 38444
rect 8406 38208 8491 38444
rect 8727 38208 8812 38444
rect 9048 38208 9133 38444
rect 9369 38208 9454 38444
rect 9690 38208 9775 38444
rect 10011 38208 10096 38444
rect 10332 38208 10417 38444
rect 10653 38208 10738 38444
rect 10974 38208 11059 38444
rect 11295 38208 11380 38444
rect 11616 38208 11701 38444
rect 11937 38208 12022 38444
rect 12258 38208 12343 38444
rect 12579 38208 12664 38444
rect 12900 38208 12985 38444
rect 13221 38208 13306 38444
rect 13542 38208 13627 38444
rect 13863 38208 13948 38444
rect 14184 38208 14269 38444
rect 14505 38208 14590 38444
rect 14826 38208 14911 38444
rect 15147 38208 15232 38444
rect 15468 38208 15553 38444
rect 15789 38208 15874 38444
rect 16110 38208 16195 38444
rect 16431 38208 16516 38444
rect 16752 38208 16837 38444
rect 17073 38208 17158 38444
rect 17394 38208 17479 38444
rect 17715 38208 17800 38444
rect 18036 38208 18121 38444
rect 18357 38208 18442 38444
rect 18678 38208 18763 38444
rect 18999 38208 19084 38444
rect 19320 38208 19405 38444
rect 19641 38208 19726 38444
rect 19962 38208 20047 38444
rect 20283 38208 20368 38444
rect 20604 38208 20689 38444
rect 20925 38208 21010 38444
rect 21246 38208 21331 38444
rect 21567 38208 21652 38444
rect 21888 38208 21973 38444
rect 22209 38208 22294 38444
rect 22530 38208 22615 38444
rect 22851 38208 22936 38444
rect 23172 38208 23257 38444
rect 23493 38208 23578 38444
rect 23814 38208 23899 38444
rect 24135 38208 24220 38444
rect 24456 38208 24640 38444
rect -3360 38120 24640 38208
rect -3360 37884 -3087 38120
rect -2851 37884 -2765 38120
rect -2529 37884 -2443 38120
rect -2207 37884 -2121 38120
rect -1885 37884 -1799 38120
rect -1563 37884 -1477 38120
rect -1241 37884 -1155 38120
rect -919 37884 -833 38120
rect -597 37884 -511 38120
rect -275 37884 -189 38120
rect 47 37884 133 38120
rect 369 37884 455 38120
rect 691 37884 777 38120
rect 1013 37884 1099 38120
rect 1335 37884 1421 38120
rect 1657 37884 1743 38120
rect 1979 37884 2065 38120
rect 2301 37884 2387 38120
rect 2623 37884 2709 38120
rect 2945 37884 3031 38120
rect 3267 37884 3353 38120
rect 3589 37884 3675 38120
rect 3911 37884 3997 38120
rect 4233 37884 4318 38120
rect 4554 37884 4639 38120
rect 4875 37884 4960 38120
rect 5196 37884 5281 38120
rect 5517 37884 5602 38120
rect 5838 37884 5923 38120
rect 6159 37884 6244 38120
rect 6480 37884 6565 38120
rect 6801 37884 6886 38120
rect 7122 37884 7207 38120
rect 7443 37884 7528 38120
rect 7764 37884 7849 38120
rect 8085 37884 8170 38120
rect 8406 37884 8491 38120
rect 8727 37884 8812 38120
rect 9048 37884 9133 38120
rect 9369 37884 9454 38120
rect 9690 37884 9775 38120
rect 10011 37884 10096 38120
rect 10332 37884 10417 38120
rect 10653 37884 10738 38120
rect 10974 37884 11059 38120
rect 11295 37884 11380 38120
rect 11616 37884 11701 38120
rect 11937 37884 12022 38120
rect 12258 37884 12343 38120
rect 12579 37884 12664 38120
rect 12900 37884 12985 38120
rect 13221 37884 13306 38120
rect 13542 37884 13627 38120
rect 13863 37884 13948 38120
rect 14184 37884 14269 38120
rect 14505 37884 14590 38120
rect 14826 37884 14911 38120
rect 15147 37884 15232 38120
rect 15468 37884 15553 38120
rect 15789 37884 15874 38120
rect 16110 37884 16195 38120
rect 16431 37884 16516 38120
rect 16752 37884 16837 38120
rect 17073 37884 17158 38120
rect 17394 37884 17479 38120
rect 17715 37884 17800 38120
rect 18036 37884 18121 38120
rect 18357 37884 18442 38120
rect 18678 37884 18763 38120
rect 18999 37884 19084 38120
rect 19320 37884 19405 38120
rect 19641 37884 19726 38120
rect 19962 37884 20047 38120
rect 20283 37884 20368 38120
rect 20604 37884 20689 38120
rect 20925 37884 21010 38120
rect 21246 37884 21331 38120
rect 21567 37884 21652 38120
rect 21888 37884 21973 38120
rect 22209 37884 22294 38120
rect 22530 37884 22615 38120
rect 22851 37884 22936 38120
rect 23172 37884 23257 38120
rect 23493 37884 23578 38120
rect 23814 37884 23899 38120
rect 24135 37884 24220 38120
rect 24456 37884 24640 38120
rect -3360 37796 24640 37884
rect -3360 37560 -3087 37796
rect -2851 37560 -2765 37796
rect -2529 37560 -2443 37796
rect -2207 37560 -2121 37796
rect -1885 37560 -1799 37796
rect -1563 37560 -1477 37796
rect -1241 37560 -1155 37796
rect -919 37560 -833 37796
rect -597 37560 -511 37796
rect -275 37560 -189 37796
rect 47 37560 133 37796
rect 369 37560 455 37796
rect 691 37560 777 37796
rect 1013 37560 1099 37796
rect 1335 37560 1421 37796
rect 1657 37560 1743 37796
rect 1979 37560 2065 37796
rect 2301 37560 2387 37796
rect 2623 37560 2709 37796
rect 2945 37560 3031 37796
rect 3267 37560 3353 37796
rect 3589 37560 3675 37796
rect 3911 37560 3997 37796
rect 4233 37560 4318 37796
rect 4554 37560 4639 37796
rect 4875 37560 4960 37796
rect 5196 37560 5281 37796
rect 5517 37560 5602 37796
rect 5838 37560 5923 37796
rect 6159 37560 6244 37796
rect 6480 37560 6565 37796
rect 6801 37560 6886 37796
rect 7122 37560 7207 37796
rect 7443 37560 7528 37796
rect 7764 37560 7849 37796
rect 8085 37560 8170 37796
rect 8406 37560 8491 37796
rect 8727 37560 8812 37796
rect 9048 37560 9133 37796
rect 9369 37560 9454 37796
rect 9690 37560 9775 37796
rect 10011 37560 10096 37796
rect 10332 37560 10417 37796
rect 10653 37560 10738 37796
rect 10974 37560 11059 37796
rect 11295 37560 11380 37796
rect 11616 37560 11701 37796
rect 11937 37560 12022 37796
rect 12258 37560 12343 37796
rect 12579 37560 12664 37796
rect 12900 37560 12985 37796
rect 13221 37560 13306 37796
rect 13542 37560 13627 37796
rect 13863 37560 13948 37796
rect 14184 37560 14269 37796
rect 14505 37560 14590 37796
rect 14826 37560 14911 37796
rect 15147 37560 15232 37796
rect 15468 37560 15553 37796
rect 15789 37560 15874 37796
rect 16110 37560 16195 37796
rect 16431 37560 16516 37796
rect 16752 37560 16837 37796
rect 17073 37560 17158 37796
rect 17394 37560 17479 37796
rect 17715 37560 17800 37796
rect 18036 37560 18121 37796
rect 18357 37560 18442 37796
rect 18678 37560 18763 37796
rect 18999 37560 19084 37796
rect 19320 37560 19405 37796
rect 19641 37560 19726 37796
rect 19962 37560 20047 37796
rect 20283 37560 20368 37796
rect 20604 37560 20689 37796
rect 20925 37560 21010 37796
rect 21246 37560 21331 37796
rect 21567 37560 21652 37796
rect 21888 37560 21973 37796
rect 22209 37560 22294 37796
rect 22530 37560 22615 37796
rect 22851 37560 22936 37796
rect 23172 37560 23257 37796
rect 23493 37560 23578 37796
rect 23814 37560 23899 37796
rect 24135 37560 24220 37796
rect 24456 37560 24640 37796
rect -3360 37472 24640 37560
rect -3360 37236 -3087 37472
rect -2851 37236 -2765 37472
rect -2529 37236 -2443 37472
rect -2207 37236 -2121 37472
rect -1885 37236 -1799 37472
rect -1563 37236 -1477 37472
rect -1241 37236 -1155 37472
rect -919 37236 -833 37472
rect -597 37236 -511 37472
rect -275 37236 -189 37472
rect 47 37236 133 37472
rect 369 37236 455 37472
rect 691 37236 777 37472
rect 1013 37236 1099 37472
rect 1335 37236 1421 37472
rect 1657 37236 1743 37472
rect 1979 37236 2065 37472
rect 2301 37236 2387 37472
rect 2623 37236 2709 37472
rect 2945 37236 3031 37472
rect 3267 37236 3353 37472
rect 3589 37236 3675 37472
rect 3911 37236 3997 37472
rect 4233 37236 4318 37472
rect 4554 37236 4639 37472
rect 4875 37236 4960 37472
rect 5196 37236 5281 37472
rect 5517 37236 5602 37472
rect 5838 37236 5923 37472
rect 6159 37236 6244 37472
rect 6480 37236 6565 37472
rect 6801 37236 6886 37472
rect 7122 37236 7207 37472
rect 7443 37236 7528 37472
rect 7764 37236 7849 37472
rect 8085 37236 8170 37472
rect 8406 37236 8491 37472
rect 8727 37236 8812 37472
rect 9048 37236 9133 37472
rect 9369 37236 9454 37472
rect 9690 37236 9775 37472
rect 10011 37236 10096 37472
rect 10332 37236 10417 37472
rect 10653 37236 10738 37472
rect 10974 37236 11059 37472
rect 11295 37236 11380 37472
rect 11616 37236 11701 37472
rect 11937 37236 12022 37472
rect 12258 37236 12343 37472
rect 12579 37236 12664 37472
rect 12900 37236 12985 37472
rect 13221 37236 13306 37472
rect 13542 37236 13627 37472
rect 13863 37236 13948 37472
rect 14184 37236 14269 37472
rect 14505 37236 14590 37472
rect 14826 37236 14911 37472
rect 15147 37236 15232 37472
rect 15468 37236 15553 37472
rect 15789 37236 15874 37472
rect 16110 37236 16195 37472
rect 16431 37236 16516 37472
rect 16752 37236 16837 37472
rect 17073 37236 17158 37472
rect 17394 37236 17479 37472
rect 17715 37236 17800 37472
rect 18036 37236 18121 37472
rect 18357 37236 18442 37472
rect 18678 37236 18763 37472
rect 18999 37236 19084 37472
rect 19320 37236 19405 37472
rect 19641 37236 19726 37472
rect 19962 37236 20047 37472
rect 20283 37236 20368 37472
rect 20604 37236 20689 37472
rect 20925 37236 21010 37472
rect 21246 37236 21331 37472
rect 21567 37236 21652 37472
rect 21888 37236 21973 37472
rect 22209 37236 22294 37472
rect 22530 37236 22615 37472
rect 22851 37236 22936 37472
rect 23172 37236 23257 37472
rect 23493 37236 23578 37472
rect 23814 37236 23899 37472
rect 24135 37236 24220 37472
rect 24456 37236 24640 37472
rect -3360 37148 24640 37236
rect -3360 36912 -3087 37148
rect -2851 36912 -2765 37148
rect -2529 36912 -2443 37148
rect -2207 36912 -2121 37148
rect -1885 36912 -1799 37148
rect -1563 36912 -1477 37148
rect -1241 36912 -1155 37148
rect -919 36912 -833 37148
rect -597 36912 -511 37148
rect -275 36912 -189 37148
rect 47 36912 133 37148
rect 369 36912 455 37148
rect 691 36912 777 37148
rect 1013 36912 1099 37148
rect 1335 36912 1421 37148
rect 1657 36912 1743 37148
rect 1979 36912 2065 37148
rect 2301 36912 2387 37148
rect 2623 36912 2709 37148
rect 2945 36912 3031 37148
rect 3267 36912 3353 37148
rect 3589 36912 3675 37148
rect 3911 36912 3997 37148
rect 4233 36912 4318 37148
rect 4554 36912 4639 37148
rect 4875 36912 4960 37148
rect 5196 36912 5281 37148
rect 5517 36912 5602 37148
rect 5838 36912 5923 37148
rect 6159 36912 6244 37148
rect 6480 36912 6565 37148
rect 6801 36912 6886 37148
rect 7122 36912 7207 37148
rect 7443 36912 7528 37148
rect 7764 36912 7849 37148
rect 8085 36912 8170 37148
rect 8406 36912 8491 37148
rect 8727 36912 8812 37148
rect 9048 36912 9133 37148
rect 9369 36912 9454 37148
rect 9690 36912 9775 37148
rect 10011 36912 10096 37148
rect 10332 36912 10417 37148
rect 10653 36912 10738 37148
rect 10974 36912 11059 37148
rect 11295 36912 11380 37148
rect 11616 36912 11701 37148
rect 11937 36912 12022 37148
rect 12258 36912 12343 37148
rect 12579 36912 12664 37148
rect 12900 36912 12985 37148
rect 13221 36912 13306 37148
rect 13542 36912 13627 37148
rect 13863 36912 13948 37148
rect 14184 36912 14269 37148
rect 14505 36912 14590 37148
rect 14826 36912 14911 37148
rect 15147 36912 15232 37148
rect 15468 36912 15553 37148
rect 15789 36912 15874 37148
rect 16110 36912 16195 37148
rect 16431 36912 16516 37148
rect 16752 36912 16837 37148
rect 17073 36912 17158 37148
rect 17394 36912 17479 37148
rect 17715 36912 17800 37148
rect 18036 36912 18121 37148
rect 18357 36912 18442 37148
rect 18678 36912 18763 37148
rect 18999 36912 19084 37148
rect 19320 36912 19405 37148
rect 19641 36912 19726 37148
rect 19962 36912 20047 37148
rect 20283 36912 20368 37148
rect 20604 36912 20689 37148
rect 20925 36912 21010 37148
rect 21246 36912 21331 37148
rect 21567 36912 21652 37148
rect 21888 36912 21973 37148
rect 22209 36912 22294 37148
rect 22530 36912 22615 37148
rect 22851 36912 22936 37148
rect 23172 36912 23257 37148
rect 23493 36912 23578 37148
rect 23814 36912 23899 37148
rect 24135 36912 24220 37148
rect 24456 36912 24640 37148
rect -3360 36824 24640 36912
rect -3360 36588 -3087 36824
rect -2851 36588 -2765 36824
rect -2529 36588 -2443 36824
rect -2207 36588 -2121 36824
rect -1885 36588 -1799 36824
rect -1563 36588 -1477 36824
rect -1241 36588 -1155 36824
rect -919 36588 -833 36824
rect -597 36588 -511 36824
rect -275 36588 -189 36824
rect 47 36588 133 36824
rect 369 36588 455 36824
rect 691 36588 777 36824
rect 1013 36588 1099 36824
rect 1335 36588 1421 36824
rect 1657 36588 1743 36824
rect 1979 36588 2065 36824
rect 2301 36588 2387 36824
rect 2623 36588 2709 36824
rect 2945 36588 3031 36824
rect 3267 36588 3353 36824
rect 3589 36588 3675 36824
rect 3911 36588 3997 36824
rect 4233 36588 4318 36824
rect 4554 36588 4639 36824
rect 4875 36588 4960 36824
rect 5196 36588 5281 36824
rect 5517 36588 5602 36824
rect 5838 36588 5923 36824
rect 6159 36588 6244 36824
rect 6480 36588 6565 36824
rect 6801 36588 6886 36824
rect 7122 36588 7207 36824
rect 7443 36588 7528 36824
rect 7764 36588 7849 36824
rect 8085 36588 8170 36824
rect 8406 36588 8491 36824
rect 8727 36588 8812 36824
rect 9048 36588 9133 36824
rect 9369 36588 9454 36824
rect 9690 36588 9775 36824
rect 10011 36588 10096 36824
rect 10332 36588 10417 36824
rect 10653 36588 10738 36824
rect 10974 36588 11059 36824
rect 11295 36588 11380 36824
rect 11616 36588 11701 36824
rect 11937 36588 12022 36824
rect 12258 36588 12343 36824
rect 12579 36588 12664 36824
rect 12900 36588 12985 36824
rect 13221 36588 13306 36824
rect 13542 36588 13627 36824
rect 13863 36588 13948 36824
rect 14184 36588 14269 36824
rect 14505 36588 14590 36824
rect 14826 36588 14911 36824
rect 15147 36588 15232 36824
rect 15468 36588 15553 36824
rect 15789 36588 15874 36824
rect 16110 36588 16195 36824
rect 16431 36588 16516 36824
rect 16752 36588 16837 36824
rect 17073 36588 17158 36824
rect 17394 36588 17479 36824
rect 17715 36588 17800 36824
rect 18036 36588 18121 36824
rect 18357 36588 18442 36824
rect 18678 36588 18763 36824
rect 18999 36588 19084 36824
rect 19320 36588 19405 36824
rect 19641 36588 19726 36824
rect 19962 36588 20047 36824
rect 20283 36588 20368 36824
rect 20604 36588 20689 36824
rect 20925 36588 21010 36824
rect 21246 36588 21331 36824
rect 21567 36588 21652 36824
rect 21888 36588 21973 36824
rect 22209 36588 22294 36824
rect 22530 36588 22615 36824
rect 22851 36588 22936 36824
rect 23172 36588 23257 36824
rect 23493 36588 23578 36824
rect 23814 36588 23899 36824
rect 24135 36588 24220 36824
rect 24456 36588 24640 36824
rect -3360 36500 24640 36588
rect -3360 36264 -3087 36500
rect -2851 36264 -2765 36500
rect -2529 36264 -2443 36500
rect -2207 36264 -2121 36500
rect -1885 36264 -1799 36500
rect -1563 36264 -1477 36500
rect -1241 36264 -1155 36500
rect -919 36264 -833 36500
rect -597 36264 -511 36500
rect -275 36264 -189 36500
rect 47 36264 133 36500
rect 369 36264 455 36500
rect 691 36264 777 36500
rect 1013 36264 1099 36500
rect 1335 36264 1421 36500
rect 1657 36264 1743 36500
rect 1979 36264 2065 36500
rect 2301 36264 2387 36500
rect 2623 36264 2709 36500
rect 2945 36264 3031 36500
rect 3267 36264 3353 36500
rect 3589 36264 3675 36500
rect 3911 36264 3997 36500
rect 4233 36264 4318 36500
rect 4554 36264 4639 36500
rect 4875 36264 4960 36500
rect 5196 36264 5281 36500
rect 5517 36264 5602 36500
rect 5838 36264 5923 36500
rect 6159 36264 6244 36500
rect 6480 36264 6565 36500
rect 6801 36264 6886 36500
rect 7122 36264 7207 36500
rect 7443 36264 7528 36500
rect 7764 36264 7849 36500
rect 8085 36264 8170 36500
rect 8406 36264 8491 36500
rect 8727 36264 8812 36500
rect 9048 36264 9133 36500
rect 9369 36264 9454 36500
rect 9690 36264 9775 36500
rect 10011 36264 10096 36500
rect 10332 36264 10417 36500
rect 10653 36264 10738 36500
rect 10974 36264 11059 36500
rect 11295 36264 11380 36500
rect 11616 36264 11701 36500
rect 11937 36264 12022 36500
rect 12258 36264 12343 36500
rect 12579 36264 12664 36500
rect 12900 36264 12985 36500
rect 13221 36264 13306 36500
rect 13542 36264 13627 36500
rect 13863 36264 13948 36500
rect 14184 36264 14269 36500
rect 14505 36264 14590 36500
rect 14826 36264 14911 36500
rect 15147 36264 15232 36500
rect 15468 36264 15553 36500
rect 15789 36264 15874 36500
rect 16110 36264 16195 36500
rect 16431 36264 16516 36500
rect 16752 36264 16837 36500
rect 17073 36264 17158 36500
rect 17394 36264 17479 36500
rect 17715 36264 17800 36500
rect 18036 36264 18121 36500
rect 18357 36264 18442 36500
rect 18678 36264 18763 36500
rect 18999 36264 19084 36500
rect 19320 36264 19405 36500
rect 19641 36264 19726 36500
rect 19962 36264 20047 36500
rect 20283 36264 20368 36500
rect 20604 36264 20689 36500
rect 20925 36264 21010 36500
rect 21246 36264 21331 36500
rect 21567 36264 21652 36500
rect 21888 36264 21973 36500
rect 22209 36264 22294 36500
rect 22530 36264 22615 36500
rect 22851 36264 22936 36500
rect 23172 36264 23257 36500
rect 23493 36264 23578 36500
rect 23814 36264 23899 36500
rect 24135 36264 24220 36500
rect 24456 36264 24640 36500
rect -3360 36176 24640 36264
rect -3360 35940 -3087 36176
rect -2851 35940 -2765 36176
rect -2529 35940 -2443 36176
rect -2207 35940 -2121 36176
rect -1885 35940 -1799 36176
rect -1563 35940 -1477 36176
rect -1241 35940 -1155 36176
rect -919 35940 -833 36176
rect -597 35940 -511 36176
rect -275 35940 -189 36176
rect 47 35940 133 36176
rect 369 35940 455 36176
rect 691 35940 777 36176
rect 1013 35940 1099 36176
rect 1335 35940 1421 36176
rect 1657 35940 1743 36176
rect 1979 35940 2065 36176
rect 2301 35940 2387 36176
rect 2623 35940 2709 36176
rect 2945 35940 3031 36176
rect 3267 35940 3353 36176
rect 3589 35940 3675 36176
rect 3911 35940 3997 36176
rect 4233 35940 4318 36176
rect 4554 35940 4639 36176
rect 4875 35940 4960 36176
rect 5196 35940 5281 36176
rect 5517 35940 5602 36176
rect 5838 35940 5923 36176
rect 6159 35940 6244 36176
rect 6480 35940 6565 36176
rect 6801 35940 6886 36176
rect 7122 35940 7207 36176
rect 7443 35940 7528 36176
rect 7764 35940 7849 36176
rect 8085 35940 8170 36176
rect 8406 35940 8491 36176
rect 8727 35940 8812 36176
rect 9048 35940 9133 36176
rect 9369 35940 9454 36176
rect 9690 35940 9775 36176
rect 10011 35940 10096 36176
rect 10332 35940 10417 36176
rect 10653 35940 10738 36176
rect 10974 35940 11059 36176
rect 11295 35940 11380 36176
rect 11616 35940 11701 36176
rect 11937 35940 12022 36176
rect 12258 35940 12343 36176
rect 12579 35940 12664 36176
rect 12900 35940 12985 36176
rect 13221 35940 13306 36176
rect 13542 35940 13627 36176
rect 13863 35940 13948 36176
rect 14184 35940 14269 36176
rect 14505 35940 14590 36176
rect 14826 35940 14911 36176
rect 15147 35940 15232 36176
rect 15468 35940 15553 36176
rect 15789 35940 15874 36176
rect 16110 35940 16195 36176
rect 16431 35940 16516 36176
rect 16752 35940 16837 36176
rect 17073 35940 17158 36176
rect 17394 35940 17479 36176
rect 17715 35940 17800 36176
rect 18036 35940 18121 36176
rect 18357 35940 18442 36176
rect 18678 35940 18763 36176
rect 18999 35940 19084 36176
rect 19320 35940 19405 36176
rect 19641 35940 19726 36176
rect 19962 35940 20047 36176
rect 20283 35940 20368 36176
rect 20604 35940 20689 36176
rect 20925 35940 21010 36176
rect 21246 35940 21331 36176
rect 21567 35940 21652 36176
rect 21888 35940 21973 36176
rect 22209 35940 22294 36176
rect 22530 35940 22615 36176
rect 22851 35940 22936 36176
rect 23172 35940 23257 36176
rect 23493 35940 23578 36176
rect 23814 35940 23899 36176
rect 24135 35940 24220 36176
rect 24456 35940 24640 36176
rect -3360 35852 24640 35940
rect -3360 35616 -3087 35852
rect -2851 35616 -2765 35852
rect -2529 35616 -2443 35852
rect -2207 35616 -2121 35852
rect -1885 35616 -1799 35852
rect -1563 35616 -1477 35852
rect -1241 35616 -1155 35852
rect -919 35616 -833 35852
rect -597 35616 -511 35852
rect -275 35616 -189 35852
rect 47 35616 133 35852
rect 369 35616 455 35852
rect 691 35616 777 35852
rect 1013 35616 1099 35852
rect 1335 35616 1421 35852
rect 1657 35616 1743 35852
rect 1979 35616 2065 35852
rect 2301 35616 2387 35852
rect 2623 35616 2709 35852
rect 2945 35616 3031 35852
rect 3267 35616 3353 35852
rect 3589 35616 3675 35852
rect 3911 35616 3997 35852
rect 4233 35616 4318 35852
rect 4554 35616 4639 35852
rect 4875 35616 4960 35852
rect 5196 35616 5281 35852
rect 5517 35616 5602 35852
rect 5838 35616 5923 35852
rect 6159 35616 6244 35852
rect 6480 35616 6565 35852
rect 6801 35616 6886 35852
rect 7122 35616 7207 35852
rect 7443 35616 7528 35852
rect 7764 35616 7849 35852
rect 8085 35616 8170 35852
rect 8406 35616 8491 35852
rect 8727 35616 8812 35852
rect 9048 35616 9133 35852
rect 9369 35616 9454 35852
rect 9690 35616 9775 35852
rect 10011 35616 10096 35852
rect 10332 35616 10417 35852
rect 10653 35616 10738 35852
rect 10974 35616 11059 35852
rect 11295 35616 11380 35852
rect 11616 35616 11701 35852
rect 11937 35616 12022 35852
rect 12258 35616 12343 35852
rect 12579 35616 12664 35852
rect 12900 35616 12985 35852
rect 13221 35616 13306 35852
rect 13542 35616 13627 35852
rect 13863 35616 13948 35852
rect 14184 35616 14269 35852
rect 14505 35616 14590 35852
rect 14826 35616 14911 35852
rect 15147 35616 15232 35852
rect 15468 35616 15553 35852
rect 15789 35616 15874 35852
rect 16110 35616 16195 35852
rect 16431 35616 16516 35852
rect 16752 35616 16837 35852
rect 17073 35616 17158 35852
rect 17394 35616 17479 35852
rect 17715 35616 17800 35852
rect 18036 35616 18121 35852
rect 18357 35616 18442 35852
rect 18678 35616 18763 35852
rect 18999 35616 19084 35852
rect 19320 35616 19405 35852
rect 19641 35616 19726 35852
rect 19962 35616 20047 35852
rect 20283 35616 20368 35852
rect 20604 35616 20689 35852
rect 20925 35616 21010 35852
rect 21246 35616 21331 35852
rect 21567 35616 21652 35852
rect 21888 35616 21973 35852
rect 22209 35616 22294 35852
rect 22530 35616 22615 35852
rect 22851 35616 22936 35852
rect 23172 35616 23257 35852
rect 23493 35616 23578 35852
rect 23814 35616 23899 35852
rect 24135 35616 24220 35852
rect 24456 35616 24640 35852
rect -3360 35528 24640 35616
rect -3360 35292 -3087 35528
rect -2851 35292 -2765 35528
rect -2529 35292 -2443 35528
rect -2207 35292 -2121 35528
rect -1885 35292 -1799 35528
rect -1563 35292 -1477 35528
rect -1241 35292 -1155 35528
rect -919 35292 -833 35528
rect -597 35292 -511 35528
rect -275 35292 -189 35528
rect 47 35292 133 35528
rect 369 35292 455 35528
rect 691 35292 777 35528
rect 1013 35292 1099 35528
rect 1335 35292 1421 35528
rect 1657 35292 1743 35528
rect 1979 35292 2065 35528
rect 2301 35292 2387 35528
rect 2623 35292 2709 35528
rect 2945 35292 3031 35528
rect 3267 35292 3353 35528
rect 3589 35292 3675 35528
rect 3911 35292 3997 35528
rect 4233 35292 4318 35528
rect 4554 35292 4639 35528
rect 4875 35292 4960 35528
rect 5196 35292 5281 35528
rect 5517 35292 5602 35528
rect 5838 35292 5923 35528
rect 6159 35292 6244 35528
rect 6480 35292 6565 35528
rect 6801 35292 6886 35528
rect 7122 35292 7207 35528
rect 7443 35292 7528 35528
rect 7764 35292 7849 35528
rect 8085 35292 8170 35528
rect 8406 35292 8491 35528
rect 8727 35292 8812 35528
rect 9048 35292 9133 35528
rect 9369 35292 9454 35528
rect 9690 35292 9775 35528
rect 10011 35292 10096 35528
rect 10332 35292 10417 35528
rect 10653 35292 10738 35528
rect 10974 35292 11059 35528
rect 11295 35292 11380 35528
rect 11616 35292 11701 35528
rect 11937 35292 12022 35528
rect 12258 35292 12343 35528
rect 12579 35292 12664 35528
rect 12900 35292 12985 35528
rect 13221 35292 13306 35528
rect 13542 35292 13627 35528
rect 13863 35292 13948 35528
rect 14184 35292 14269 35528
rect 14505 35292 14590 35528
rect 14826 35292 14911 35528
rect 15147 35292 15232 35528
rect 15468 35292 15553 35528
rect 15789 35292 15874 35528
rect 16110 35292 16195 35528
rect 16431 35292 16516 35528
rect 16752 35292 16837 35528
rect 17073 35292 17158 35528
rect 17394 35292 17479 35528
rect 17715 35292 17800 35528
rect 18036 35292 18121 35528
rect 18357 35292 18442 35528
rect 18678 35292 18763 35528
rect 18999 35292 19084 35528
rect 19320 35292 19405 35528
rect 19641 35292 19726 35528
rect 19962 35292 20047 35528
rect 20283 35292 20368 35528
rect 20604 35292 20689 35528
rect 20925 35292 21010 35528
rect 21246 35292 21331 35528
rect 21567 35292 21652 35528
rect 21888 35292 21973 35528
rect 22209 35292 22294 35528
rect 22530 35292 22615 35528
rect 22851 35292 22936 35528
rect 23172 35292 23257 35528
rect 23493 35292 23578 35528
rect 23814 35292 23899 35528
rect 24135 35292 24220 35528
rect 24456 35292 24640 35528
rect -3360 35204 24640 35292
rect -3360 34968 -3087 35204
rect -2851 34968 -2765 35204
rect -2529 34968 -2443 35204
rect -2207 34968 -2121 35204
rect -1885 34968 -1799 35204
rect -1563 34968 -1477 35204
rect -1241 34968 -1155 35204
rect -919 34968 -833 35204
rect -597 34968 -511 35204
rect -275 34968 -189 35204
rect 47 34968 133 35204
rect 369 34968 455 35204
rect 691 34968 777 35204
rect 1013 34968 1099 35204
rect 1335 34968 1421 35204
rect 1657 34968 1743 35204
rect 1979 34968 2065 35204
rect 2301 34968 2387 35204
rect 2623 34968 2709 35204
rect 2945 34968 3031 35204
rect 3267 34968 3353 35204
rect 3589 34968 3675 35204
rect 3911 34968 3997 35204
rect 4233 34968 4318 35204
rect 4554 34968 4639 35204
rect 4875 34968 4960 35204
rect 5196 34968 5281 35204
rect 5517 34968 5602 35204
rect 5838 34968 5923 35204
rect 6159 34968 6244 35204
rect 6480 34968 6565 35204
rect 6801 34968 6886 35204
rect 7122 34968 7207 35204
rect 7443 34968 7528 35204
rect 7764 34968 7849 35204
rect 8085 34968 8170 35204
rect 8406 34968 8491 35204
rect 8727 34968 8812 35204
rect 9048 34968 9133 35204
rect 9369 34968 9454 35204
rect 9690 34968 9775 35204
rect 10011 34968 10096 35204
rect 10332 34968 10417 35204
rect 10653 34968 10738 35204
rect 10974 34968 11059 35204
rect 11295 34968 11380 35204
rect 11616 34968 11701 35204
rect 11937 34968 12022 35204
rect 12258 34968 12343 35204
rect 12579 34968 12664 35204
rect 12900 34968 12985 35204
rect 13221 34968 13306 35204
rect 13542 34968 13627 35204
rect 13863 34968 13948 35204
rect 14184 34968 14269 35204
rect 14505 34968 14590 35204
rect 14826 34968 14911 35204
rect 15147 34968 15232 35204
rect 15468 34968 15553 35204
rect 15789 34968 15874 35204
rect 16110 34968 16195 35204
rect 16431 34968 16516 35204
rect 16752 34968 16837 35204
rect 17073 34968 17158 35204
rect 17394 34968 17479 35204
rect 17715 34968 17800 35204
rect 18036 34968 18121 35204
rect 18357 34968 18442 35204
rect 18678 34968 18763 35204
rect 18999 34968 19084 35204
rect 19320 34968 19405 35204
rect 19641 34968 19726 35204
rect 19962 34968 20047 35204
rect 20283 34968 20368 35204
rect 20604 34968 20689 35204
rect 20925 34968 21010 35204
rect 21246 34968 21331 35204
rect 21567 34968 21652 35204
rect 21888 34968 21973 35204
rect 22209 34968 22294 35204
rect 22530 34968 22615 35204
rect 22851 34968 22936 35204
rect 23172 34968 23257 35204
rect 23493 34968 23578 35204
rect 23814 34968 23899 35204
rect 24135 34968 24220 35204
rect 24456 34968 24640 35204
rect -3360 34880 24640 34968
rect -3360 34644 -3087 34880
rect -2851 34644 -2765 34880
rect -2529 34644 -2443 34880
rect -2207 34644 -2121 34880
rect -1885 34644 -1799 34880
rect -1563 34644 -1477 34880
rect -1241 34644 -1155 34880
rect -919 34644 -833 34880
rect -597 34644 -511 34880
rect -275 34644 -189 34880
rect 47 34644 133 34880
rect 369 34644 455 34880
rect 691 34644 777 34880
rect 1013 34644 1099 34880
rect 1335 34644 1421 34880
rect 1657 34644 1743 34880
rect 1979 34644 2065 34880
rect 2301 34644 2387 34880
rect 2623 34644 2709 34880
rect 2945 34644 3031 34880
rect 3267 34644 3353 34880
rect 3589 34644 3675 34880
rect 3911 34644 3997 34880
rect 4233 34644 4318 34880
rect 4554 34644 4639 34880
rect 4875 34644 4960 34880
rect 5196 34644 5281 34880
rect 5517 34644 5602 34880
rect 5838 34644 5923 34880
rect 6159 34644 6244 34880
rect 6480 34644 6565 34880
rect 6801 34644 6886 34880
rect 7122 34644 7207 34880
rect 7443 34644 7528 34880
rect 7764 34644 7849 34880
rect 8085 34644 8170 34880
rect 8406 34644 8491 34880
rect 8727 34644 8812 34880
rect 9048 34644 9133 34880
rect 9369 34644 9454 34880
rect 9690 34644 9775 34880
rect 10011 34644 10096 34880
rect 10332 34644 10417 34880
rect 10653 34644 10738 34880
rect 10974 34644 11059 34880
rect 11295 34644 11380 34880
rect 11616 34644 11701 34880
rect 11937 34644 12022 34880
rect 12258 34644 12343 34880
rect 12579 34644 12664 34880
rect 12900 34644 12985 34880
rect 13221 34644 13306 34880
rect 13542 34644 13627 34880
rect 13863 34644 13948 34880
rect 14184 34644 14269 34880
rect 14505 34644 14590 34880
rect 14826 34644 14911 34880
rect 15147 34644 15232 34880
rect 15468 34644 15553 34880
rect 15789 34644 15874 34880
rect 16110 34644 16195 34880
rect 16431 34644 16516 34880
rect 16752 34644 16837 34880
rect 17073 34644 17158 34880
rect 17394 34644 17479 34880
rect 17715 34644 17800 34880
rect 18036 34644 18121 34880
rect 18357 34644 18442 34880
rect 18678 34644 18763 34880
rect 18999 34644 19084 34880
rect 19320 34644 19405 34880
rect 19641 34644 19726 34880
rect 19962 34644 20047 34880
rect 20283 34644 20368 34880
rect 20604 34644 20689 34880
rect 20925 34644 21010 34880
rect 21246 34644 21331 34880
rect 21567 34644 21652 34880
rect 21888 34644 21973 34880
rect 22209 34644 22294 34880
rect 22530 34644 22615 34880
rect 22851 34644 22936 34880
rect 23172 34644 23257 34880
rect 23493 34644 23578 34880
rect 23814 34644 23899 34880
rect 24135 34644 24220 34880
rect 24456 34644 24640 34880
rect -3360 34633 24640 34644
rect -3360 34608 -2720 34633
rect 24000 34608 24640 34633
rect -3360 18424 -2720 18451
rect 24000 18424 24640 18451
rect -3360 18423 24640 18424
rect -3360 18187 -3185 18423
rect -2949 18187 -2862 18423
rect -2626 18187 -2539 18423
rect -2303 18187 -2216 18423
rect -1980 18187 -1893 18423
rect -1657 18187 -1570 18423
rect -1334 18187 -1247 18423
rect -1011 18187 -924 18423
rect -688 18187 -601 18423
rect -365 18187 -278 18423
rect -42 18187 45 18423
rect 281 18187 368 18423
rect 604 18187 691 18423
rect 927 18187 1014 18423
rect 1250 18187 1337 18423
rect 1573 18187 1660 18423
rect 1896 18187 1983 18423
rect 2219 18187 2306 18423
rect 2542 18187 2629 18423
rect 2865 18187 2952 18423
rect 3188 18187 3275 18423
rect 3511 18187 3598 18423
rect 3834 18187 3921 18423
rect 4157 18187 4244 18423
rect 4480 18187 4567 18423
rect 4803 18187 4890 18423
rect 5126 18187 5213 18423
rect 5449 18187 5536 18423
rect 5772 18187 5859 18423
rect 6095 18187 6182 18423
rect 6418 18187 6505 18423
rect 6741 18187 6828 18423
rect 7064 18187 7150 18423
rect 7386 18187 7472 18423
rect 7708 18187 7794 18423
rect 8030 18187 8116 18423
rect 8352 18187 8438 18423
rect 8674 18187 8760 18423
rect 8996 18187 9082 18423
rect 9318 18187 9404 18423
rect 9640 18187 9726 18423
rect 9962 18187 10048 18423
rect 10284 18187 10370 18423
rect 10606 18187 10692 18423
rect 10928 18187 11014 18423
rect 11250 18187 11336 18423
rect 11572 18187 11658 18423
rect 11894 18187 11980 18423
rect 12216 18187 12302 18423
rect 12538 18187 12624 18423
rect 12860 18187 12946 18423
rect 13182 18187 13268 18423
rect 13504 18187 13590 18423
rect 13826 18187 13912 18423
rect 14148 18187 14234 18423
rect 14470 18187 14556 18423
rect 14792 18187 14878 18423
rect 15114 18187 15200 18423
rect 15436 18187 15522 18423
rect 15758 18187 15844 18423
rect 16080 18187 16166 18423
rect 16402 18187 16488 18423
rect 16724 18187 16810 18423
rect 17046 18187 17132 18423
rect 17368 18187 17454 18423
rect 17690 18187 17776 18423
rect 18012 18187 18098 18423
rect 18334 18187 18420 18423
rect 18656 18187 18742 18423
rect 18978 18187 19064 18423
rect 19300 18187 19386 18423
rect 19622 18187 19708 18423
rect 19944 18187 20030 18423
rect 20266 18187 20352 18423
rect 20588 18187 20674 18423
rect 20910 18187 20996 18423
rect 21232 18187 21318 18423
rect 21554 18187 21640 18423
rect 21876 18187 21962 18423
rect 22198 18187 22284 18423
rect 22520 18187 22606 18423
rect 22842 18187 22928 18423
rect 23164 18187 23250 18423
rect 23486 18187 23572 18423
rect 23808 18187 23894 18423
rect 24130 18187 24216 18423
rect 24452 18187 24640 18423
rect -3360 18087 24640 18187
rect -3360 17851 -3185 18087
rect -2949 17851 -2862 18087
rect -2626 17851 -2539 18087
rect -2303 17851 -2216 18087
rect -1980 17851 -1893 18087
rect -1657 17851 -1570 18087
rect -1334 17851 -1247 18087
rect -1011 17851 -924 18087
rect -688 17851 -601 18087
rect -365 17851 -278 18087
rect -42 17851 45 18087
rect 281 17851 368 18087
rect 604 17851 691 18087
rect 927 17851 1014 18087
rect 1250 17851 1337 18087
rect 1573 17851 1660 18087
rect 1896 17851 1983 18087
rect 2219 17851 2306 18087
rect 2542 17851 2629 18087
rect 2865 17851 2952 18087
rect 3188 17851 3275 18087
rect 3511 17851 3598 18087
rect 3834 17851 3921 18087
rect 4157 17851 4244 18087
rect 4480 17851 4567 18087
rect 4803 17851 4890 18087
rect 5126 17851 5213 18087
rect 5449 17851 5536 18087
rect 5772 17851 5859 18087
rect 6095 17851 6182 18087
rect 6418 17851 6505 18087
rect 6741 17851 6828 18087
rect 7064 17851 7150 18087
rect 7386 17851 7472 18087
rect 7708 17851 7794 18087
rect 8030 17851 8116 18087
rect 8352 17851 8438 18087
rect 8674 17851 8760 18087
rect 8996 17851 9082 18087
rect 9318 17851 9404 18087
rect 9640 17851 9726 18087
rect 9962 17851 10048 18087
rect 10284 17851 10370 18087
rect 10606 17851 10692 18087
rect 10928 17851 11014 18087
rect 11250 17851 11336 18087
rect 11572 17851 11658 18087
rect 11894 17851 11980 18087
rect 12216 17851 12302 18087
rect 12538 17851 12624 18087
rect 12860 17851 12946 18087
rect 13182 17851 13268 18087
rect 13504 17851 13590 18087
rect 13826 17851 13912 18087
rect 14148 17851 14234 18087
rect 14470 17851 14556 18087
rect 14792 17851 14878 18087
rect 15114 17851 15200 18087
rect 15436 17851 15522 18087
rect 15758 17851 15844 18087
rect 16080 17851 16166 18087
rect 16402 17851 16488 18087
rect 16724 17851 16810 18087
rect 17046 17851 17132 18087
rect 17368 17851 17454 18087
rect 17690 17851 17776 18087
rect 18012 17851 18098 18087
rect 18334 17851 18420 18087
rect 18656 17851 18742 18087
rect 18978 17851 19064 18087
rect 19300 17851 19386 18087
rect 19622 17851 19708 18087
rect 19944 17851 20030 18087
rect 20266 17851 20352 18087
rect 20588 17851 20674 18087
rect 20910 17851 20996 18087
rect 21232 17851 21318 18087
rect 21554 17851 21640 18087
rect 21876 17851 21962 18087
rect 22198 17851 22284 18087
rect 22520 17851 22606 18087
rect 22842 17851 22928 18087
rect 23164 17851 23250 18087
rect 23486 17851 23572 18087
rect 23808 17851 23894 18087
rect 24130 17851 24216 18087
rect 24452 17851 24640 18087
rect -3360 17751 24640 17851
rect -3360 17515 -3185 17751
rect -2949 17515 -2862 17751
rect -2626 17515 -2539 17751
rect -2303 17515 -2216 17751
rect -1980 17515 -1893 17751
rect -1657 17515 -1570 17751
rect -1334 17515 -1247 17751
rect -1011 17515 -924 17751
rect -688 17515 -601 17751
rect -365 17515 -278 17751
rect -42 17515 45 17751
rect 281 17515 368 17751
rect 604 17515 691 17751
rect 927 17515 1014 17751
rect 1250 17515 1337 17751
rect 1573 17515 1660 17751
rect 1896 17515 1983 17751
rect 2219 17515 2306 17751
rect 2542 17515 2629 17751
rect 2865 17515 2952 17751
rect 3188 17515 3275 17751
rect 3511 17515 3598 17751
rect 3834 17515 3921 17751
rect 4157 17515 4244 17751
rect 4480 17515 4567 17751
rect 4803 17515 4890 17751
rect 5126 17515 5213 17751
rect 5449 17515 5536 17751
rect 5772 17515 5859 17751
rect 6095 17515 6182 17751
rect 6418 17515 6505 17751
rect 6741 17515 6828 17751
rect 7064 17515 7150 17751
rect 7386 17515 7472 17751
rect 7708 17515 7794 17751
rect 8030 17515 8116 17751
rect 8352 17515 8438 17751
rect 8674 17515 8760 17751
rect 8996 17515 9082 17751
rect 9318 17515 9404 17751
rect 9640 17515 9726 17751
rect 9962 17515 10048 17751
rect 10284 17515 10370 17751
rect 10606 17515 10692 17751
rect 10928 17515 11014 17751
rect 11250 17515 11336 17751
rect 11572 17515 11658 17751
rect 11894 17515 11980 17751
rect 12216 17515 12302 17751
rect 12538 17515 12624 17751
rect 12860 17515 12946 17751
rect 13182 17515 13268 17751
rect 13504 17515 13590 17751
rect 13826 17515 13912 17751
rect 14148 17515 14234 17751
rect 14470 17515 14556 17751
rect 14792 17515 14878 17751
rect 15114 17515 15200 17751
rect 15436 17515 15522 17751
rect 15758 17515 15844 17751
rect 16080 17515 16166 17751
rect 16402 17515 16488 17751
rect 16724 17515 16810 17751
rect 17046 17515 17132 17751
rect 17368 17515 17454 17751
rect 17690 17515 17776 17751
rect 18012 17515 18098 17751
rect 18334 17515 18420 17751
rect 18656 17515 18742 17751
rect 18978 17515 19064 17751
rect 19300 17515 19386 17751
rect 19622 17515 19708 17751
rect 19944 17515 20030 17751
rect 20266 17515 20352 17751
rect 20588 17515 20674 17751
rect 20910 17515 20996 17751
rect 21232 17515 21318 17751
rect 21554 17515 21640 17751
rect 21876 17515 21962 17751
rect 22198 17515 22284 17751
rect 22520 17515 22606 17751
rect 22842 17515 22928 17751
rect 23164 17515 23250 17751
rect 23486 17515 23572 17751
rect 23808 17515 23894 17751
rect 24130 17515 24216 17751
rect 24452 17515 24640 17751
rect -3360 17415 24640 17515
rect -3360 17179 -3185 17415
rect -2949 17179 -2862 17415
rect -2626 17179 -2539 17415
rect -2303 17179 -2216 17415
rect -1980 17179 -1893 17415
rect -1657 17179 -1570 17415
rect -1334 17179 -1247 17415
rect -1011 17179 -924 17415
rect -688 17179 -601 17415
rect -365 17179 -278 17415
rect -42 17179 45 17415
rect 281 17179 368 17415
rect 604 17179 691 17415
rect 927 17179 1014 17415
rect 1250 17179 1337 17415
rect 1573 17179 1660 17415
rect 1896 17179 1983 17415
rect 2219 17179 2306 17415
rect 2542 17179 2629 17415
rect 2865 17179 2952 17415
rect 3188 17179 3275 17415
rect 3511 17179 3598 17415
rect 3834 17179 3921 17415
rect 4157 17179 4244 17415
rect 4480 17179 4567 17415
rect 4803 17179 4890 17415
rect 5126 17179 5213 17415
rect 5449 17179 5536 17415
rect 5772 17179 5859 17415
rect 6095 17179 6182 17415
rect 6418 17179 6505 17415
rect 6741 17179 6828 17415
rect 7064 17179 7150 17415
rect 7386 17179 7472 17415
rect 7708 17179 7794 17415
rect 8030 17179 8116 17415
rect 8352 17179 8438 17415
rect 8674 17179 8760 17415
rect 8996 17179 9082 17415
rect 9318 17179 9404 17415
rect 9640 17179 9726 17415
rect 9962 17179 10048 17415
rect 10284 17179 10370 17415
rect 10606 17179 10692 17415
rect 10928 17179 11014 17415
rect 11250 17179 11336 17415
rect 11572 17179 11658 17415
rect 11894 17179 11980 17415
rect 12216 17179 12302 17415
rect 12538 17179 12624 17415
rect 12860 17179 12946 17415
rect 13182 17179 13268 17415
rect 13504 17179 13590 17415
rect 13826 17179 13912 17415
rect 14148 17179 14234 17415
rect 14470 17179 14556 17415
rect 14792 17179 14878 17415
rect 15114 17179 15200 17415
rect 15436 17179 15522 17415
rect 15758 17179 15844 17415
rect 16080 17179 16166 17415
rect 16402 17179 16488 17415
rect 16724 17179 16810 17415
rect 17046 17179 17132 17415
rect 17368 17179 17454 17415
rect 17690 17179 17776 17415
rect 18012 17179 18098 17415
rect 18334 17179 18420 17415
rect 18656 17179 18742 17415
rect 18978 17179 19064 17415
rect 19300 17179 19386 17415
rect 19622 17179 19708 17415
rect 19944 17179 20030 17415
rect 20266 17179 20352 17415
rect 20588 17179 20674 17415
rect 20910 17179 20996 17415
rect 21232 17179 21318 17415
rect 21554 17179 21640 17415
rect 21876 17179 21962 17415
rect 22198 17179 22284 17415
rect 22520 17179 22606 17415
rect 22842 17179 22928 17415
rect 23164 17179 23250 17415
rect 23486 17179 23572 17415
rect 23808 17179 23894 17415
rect 24130 17179 24216 17415
rect 24452 17179 24640 17415
rect -3360 17079 24640 17179
rect -3360 16843 -3185 17079
rect -2949 16843 -2862 17079
rect -2626 16843 -2539 17079
rect -2303 16843 -2216 17079
rect -1980 16843 -1893 17079
rect -1657 16843 -1570 17079
rect -1334 16843 -1247 17079
rect -1011 16843 -924 17079
rect -688 16843 -601 17079
rect -365 16843 -278 17079
rect -42 16843 45 17079
rect 281 16843 368 17079
rect 604 16843 691 17079
rect 927 16843 1014 17079
rect 1250 16843 1337 17079
rect 1573 16843 1660 17079
rect 1896 16843 1983 17079
rect 2219 16843 2306 17079
rect 2542 16843 2629 17079
rect 2865 16843 2952 17079
rect 3188 16843 3275 17079
rect 3511 16843 3598 17079
rect 3834 16843 3921 17079
rect 4157 16843 4244 17079
rect 4480 16843 4567 17079
rect 4803 16843 4890 17079
rect 5126 16843 5213 17079
rect 5449 16843 5536 17079
rect 5772 16843 5859 17079
rect 6095 16843 6182 17079
rect 6418 16843 6505 17079
rect 6741 16843 6828 17079
rect 7064 16843 7150 17079
rect 7386 16843 7472 17079
rect 7708 16843 7794 17079
rect 8030 16843 8116 17079
rect 8352 16843 8438 17079
rect 8674 16843 8760 17079
rect 8996 16843 9082 17079
rect 9318 16843 9404 17079
rect 9640 16843 9726 17079
rect 9962 16843 10048 17079
rect 10284 16843 10370 17079
rect 10606 16843 10692 17079
rect 10928 16843 11014 17079
rect 11250 16843 11336 17079
rect 11572 16843 11658 17079
rect 11894 16843 11980 17079
rect 12216 16843 12302 17079
rect 12538 16843 12624 17079
rect 12860 16843 12946 17079
rect 13182 16843 13268 17079
rect 13504 16843 13590 17079
rect 13826 16843 13912 17079
rect 14148 16843 14234 17079
rect 14470 16843 14556 17079
rect 14792 16843 14878 17079
rect 15114 16843 15200 17079
rect 15436 16843 15522 17079
rect 15758 16843 15844 17079
rect 16080 16843 16166 17079
rect 16402 16843 16488 17079
rect 16724 16843 16810 17079
rect 17046 16843 17132 17079
rect 17368 16843 17454 17079
rect 17690 16843 17776 17079
rect 18012 16843 18098 17079
rect 18334 16843 18420 17079
rect 18656 16843 18742 17079
rect 18978 16843 19064 17079
rect 19300 16843 19386 17079
rect 19622 16843 19708 17079
rect 19944 16843 20030 17079
rect 20266 16843 20352 17079
rect 20588 16843 20674 17079
rect 20910 16843 20996 17079
rect 21232 16843 21318 17079
rect 21554 16843 21640 17079
rect 21876 16843 21962 17079
rect 22198 16843 22284 17079
rect 22520 16843 22606 17079
rect 22842 16843 22928 17079
rect 23164 16843 23250 17079
rect 23486 16843 23572 17079
rect 23808 16843 23894 17079
rect 24130 16843 24216 17079
rect 24452 16843 24640 17079
rect -3360 16743 24640 16843
rect -3360 16507 -3185 16743
rect -2949 16507 -2862 16743
rect -2626 16507 -2539 16743
rect -2303 16507 -2216 16743
rect -1980 16507 -1893 16743
rect -1657 16507 -1570 16743
rect -1334 16507 -1247 16743
rect -1011 16507 -924 16743
rect -688 16507 -601 16743
rect -365 16507 -278 16743
rect -42 16507 45 16743
rect 281 16507 368 16743
rect 604 16507 691 16743
rect 927 16507 1014 16743
rect 1250 16507 1337 16743
rect 1573 16507 1660 16743
rect 1896 16507 1983 16743
rect 2219 16507 2306 16743
rect 2542 16507 2629 16743
rect 2865 16507 2952 16743
rect 3188 16507 3275 16743
rect 3511 16507 3598 16743
rect 3834 16507 3921 16743
rect 4157 16507 4244 16743
rect 4480 16507 4567 16743
rect 4803 16507 4890 16743
rect 5126 16507 5213 16743
rect 5449 16507 5536 16743
rect 5772 16507 5859 16743
rect 6095 16507 6182 16743
rect 6418 16507 6505 16743
rect 6741 16507 6828 16743
rect 7064 16507 7150 16743
rect 7386 16507 7472 16743
rect 7708 16507 7794 16743
rect 8030 16507 8116 16743
rect 8352 16507 8438 16743
rect 8674 16507 8760 16743
rect 8996 16507 9082 16743
rect 9318 16507 9404 16743
rect 9640 16507 9726 16743
rect 9962 16507 10048 16743
rect 10284 16507 10370 16743
rect 10606 16507 10692 16743
rect 10928 16507 11014 16743
rect 11250 16507 11336 16743
rect 11572 16507 11658 16743
rect 11894 16507 11980 16743
rect 12216 16507 12302 16743
rect 12538 16507 12624 16743
rect 12860 16507 12946 16743
rect 13182 16507 13268 16743
rect 13504 16507 13590 16743
rect 13826 16507 13912 16743
rect 14148 16507 14234 16743
rect 14470 16507 14556 16743
rect 14792 16507 14878 16743
rect 15114 16507 15200 16743
rect 15436 16507 15522 16743
rect 15758 16507 15844 16743
rect 16080 16507 16166 16743
rect 16402 16507 16488 16743
rect 16724 16507 16810 16743
rect 17046 16507 17132 16743
rect 17368 16507 17454 16743
rect 17690 16507 17776 16743
rect 18012 16507 18098 16743
rect 18334 16507 18420 16743
rect 18656 16507 18742 16743
rect 18978 16507 19064 16743
rect 19300 16507 19386 16743
rect 19622 16507 19708 16743
rect 19944 16507 20030 16743
rect 20266 16507 20352 16743
rect 20588 16507 20674 16743
rect 20910 16507 20996 16743
rect 21232 16507 21318 16743
rect 21554 16507 21640 16743
rect 21876 16507 21962 16743
rect 22198 16507 22284 16743
rect 22520 16507 22606 16743
rect 22842 16507 22928 16743
rect 23164 16507 23250 16743
rect 23486 16507 23572 16743
rect 23808 16507 23894 16743
rect 24130 16507 24216 16743
rect 24452 16507 24640 16743
rect -3360 16407 24640 16507
rect -3360 16171 -3185 16407
rect -2949 16171 -2862 16407
rect -2626 16171 -2539 16407
rect -2303 16171 -2216 16407
rect -1980 16171 -1893 16407
rect -1657 16171 -1570 16407
rect -1334 16171 -1247 16407
rect -1011 16171 -924 16407
rect -688 16171 -601 16407
rect -365 16171 -278 16407
rect -42 16171 45 16407
rect 281 16171 368 16407
rect 604 16171 691 16407
rect 927 16171 1014 16407
rect 1250 16171 1337 16407
rect 1573 16171 1660 16407
rect 1896 16171 1983 16407
rect 2219 16171 2306 16407
rect 2542 16171 2629 16407
rect 2865 16171 2952 16407
rect 3188 16171 3275 16407
rect 3511 16171 3598 16407
rect 3834 16171 3921 16407
rect 4157 16171 4244 16407
rect 4480 16171 4567 16407
rect 4803 16171 4890 16407
rect 5126 16171 5213 16407
rect 5449 16171 5536 16407
rect 5772 16171 5859 16407
rect 6095 16171 6182 16407
rect 6418 16171 6505 16407
rect 6741 16171 6828 16407
rect 7064 16171 7150 16407
rect 7386 16171 7472 16407
rect 7708 16171 7794 16407
rect 8030 16171 8116 16407
rect 8352 16171 8438 16407
rect 8674 16171 8760 16407
rect 8996 16171 9082 16407
rect 9318 16171 9404 16407
rect 9640 16171 9726 16407
rect 9962 16171 10048 16407
rect 10284 16171 10370 16407
rect 10606 16171 10692 16407
rect 10928 16171 11014 16407
rect 11250 16171 11336 16407
rect 11572 16171 11658 16407
rect 11894 16171 11980 16407
rect 12216 16171 12302 16407
rect 12538 16171 12624 16407
rect 12860 16171 12946 16407
rect 13182 16171 13268 16407
rect 13504 16171 13590 16407
rect 13826 16171 13912 16407
rect 14148 16171 14234 16407
rect 14470 16171 14556 16407
rect 14792 16171 14878 16407
rect 15114 16171 15200 16407
rect 15436 16171 15522 16407
rect 15758 16171 15844 16407
rect 16080 16171 16166 16407
rect 16402 16171 16488 16407
rect 16724 16171 16810 16407
rect 17046 16171 17132 16407
rect 17368 16171 17454 16407
rect 17690 16171 17776 16407
rect 18012 16171 18098 16407
rect 18334 16171 18420 16407
rect 18656 16171 18742 16407
rect 18978 16171 19064 16407
rect 19300 16171 19386 16407
rect 19622 16171 19708 16407
rect 19944 16171 20030 16407
rect 20266 16171 20352 16407
rect 20588 16171 20674 16407
rect 20910 16171 20996 16407
rect 21232 16171 21318 16407
rect 21554 16171 21640 16407
rect 21876 16171 21962 16407
rect 22198 16171 22284 16407
rect 22520 16171 22606 16407
rect 22842 16171 22928 16407
rect 23164 16171 23250 16407
rect 23486 16171 23572 16407
rect 23808 16171 23894 16407
rect 24130 16171 24216 16407
rect 24452 16171 24640 16407
rect -3360 16071 24640 16171
rect -3360 15835 -3185 16071
rect -2949 15835 -2862 16071
rect -2626 15835 -2539 16071
rect -2303 15835 -2216 16071
rect -1980 15835 -1893 16071
rect -1657 15835 -1570 16071
rect -1334 15835 -1247 16071
rect -1011 15835 -924 16071
rect -688 15835 -601 16071
rect -365 15835 -278 16071
rect -42 15835 45 16071
rect 281 15835 368 16071
rect 604 15835 691 16071
rect 927 15835 1014 16071
rect 1250 15835 1337 16071
rect 1573 15835 1660 16071
rect 1896 15835 1983 16071
rect 2219 15835 2306 16071
rect 2542 15835 2629 16071
rect 2865 15835 2952 16071
rect 3188 15835 3275 16071
rect 3511 15835 3598 16071
rect 3834 15835 3921 16071
rect 4157 15835 4244 16071
rect 4480 15835 4567 16071
rect 4803 15835 4890 16071
rect 5126 15835 5213 16071
rect 5449 15835 5536 16071
rect 5772 15835 5859 16071
rect 6095 15835 6182 16071
rect 6418 15835 6505 16071
rect 6741 15835 6828 16071
rect 7064 15835 7150 16071
rect 7386 15835 7472 16071
rect 7708 15835 7794 16071
rect 8030 15835 8116 16071
rect 8352 15835 8438 16071
rect 8674 15835 8760 16071
rect 8996 15835 9082 16071
rect 9318 15835 9404 16071
rect 9640 15835 9726 16071
rect 9962 15835 10048 16071
rect 10284 15835 10370 16071
rect 10606 15835 10692 16071
rect 10928 15835 11014 16071
rect 11250 15835 11336 16071
rect 11572 15835 11658 16071
rect 11894 15835 11980 16071
rect 12216 15835 12302 16071
rect 12538 15835 12624 16071
rect 12860 15835 12946 16071
rect 13182 15835 13268 16071
rect 13504 15835 13590 16071
rect 13826 15835 13912 16071
rect 14148 15835 14234 16071
rect 14470 15835 14556 16071
rect 14792 15835 14878 16071
rect 15114 15835 15200 16071
rect 15436 15835 15522 16071
rect 15758 15835 15844 16071
rect 16080 15835 16166 16071
rect 16402 15835 16488 16071
rect 16724 15835 16810 16071
rect 17046 15835 17132 16071
rect 17368 15835 17454 16071
rect 17690 15835 17776 16071
rect 18012 15835 18098 16071
rect 18334 15835 18420 16071
rect 18656 15835 18742 16071
rect 18978 15835 19064 16071
rect 19300 15835 19386 16071
rect 19622 15835 19708 16071
rect 19944 15835 20030 16071
rect 20266 15835 20352 16071
rect 20588 15835 20674 16071
rect 20910 15835 20996 16071
rect 21232 15835 21318 16071
rect 21554 15835 21640 16071
rect 21876 15835 21962 16071
rect 22198 15835 22284 16071
rect 22520 15835 22606 16071
rect 22842 15835 22928 16071
rect 23164 15835 23250 16071
rect 23486 15835 23572 16071
rect 23808 15835 23894 16071
rect 24130 15835 24216 16071
rect 24452 15835 24640 16071
rect -3360 15735 24640 15835
rect -3360 15499 -3185 15735
rect -2949 15499 -2862 15735
rect -2626 15499 -2539 15735
rect -2303 15499 -2216 15735
rect -1980 15499 -1893 15735
rect -1657 15499 -1570 15735
rect -1334 15499 -1247 15735
rect -1011 15499 -924 15735
rect -688 15499 -601 15735
rect -365 15499 -278 15735
rect -42 15499 45 15735
rect 281 15499 368 15735
rect 604 15499 691 15735
rect 927 15499 1014 15735
rect 1250 15499 1337 15735
rect 1573 15499 1660 15735
rect 1896 15499 1983 15735
rect 2219 15499 2306 15735
rect 2542 15499 2629 15735
rect 2865 15499 2952 15735
rect 3188 15499 3275 15735
rect 3511 15499 3598 15735
rect 3834 15499 3921 15735
rect 4157 15499 4244 15735
rect 4480 15499 4567 15735
rect 4803 15499 4890 15735
rect 5126 15499 5213 15735
rect 5449 15499 5536 15735
rect 5772 15499 5859 15735
rect 6095 15499 6182 15735
rect 6418 15499 6505 15735
rect 6741 15499 6828 15735
rect 7064 15499 7150 15735
rect 7386 15499 7472 15735
rect 7708 15499 7794 15735
rect 8030 15499 8116 15735
rect 8352 15499 8438 15735
rect 8674 15499 8760 15735
rect 8996 15499 9082 15735
rect 9318 15499 9404 15735
rect 9640 15499 9726 15735
rect 9962 15499 10048 15735
rect 10284 15499 10370 15735
rect 10606 15499 10692 15735
rect 10928 15499 11014 15735
rect 11250 15499 11336 15735
rect 11572 15499 11658 15735
rect 11894 15499 11980 15735
rect 12216 15499 12302 15735
rect 12538 15499 12624 15735
rect 12860 15499 12946 15735
rect 13182 15499 13268 15735
rect 13504 15499 13590 15735
rect 13826 15499 13912 15735
rect 14148 15499 14234 15735
rect 14470 15499 14556 15735
rect 14792 15499 14878 15735
rect 15114 15499 15200 15735
rect 15436 15499 15522 15735
rect 15758 15499 15844 15735
rect 16080 15499 16166 15735
rect 16402 15499 16488 15735
rect 16724 15499 16810 15735
rect 17046 15499 17132 15735
rect 17368 15499 17454 15735
rect 17690 15499 17776 15735
rect 18012 15499 18098 15735
rect 18334 15499 18420 15735
rect 18656 15499 18742 15735
rect 18978 15499 19064 15735
rect 19300 15499 19386 15735
rect 19622 15499 19708 15735
rect 19944 15499 20030 15735
rect 20266 15499 20352 15735
rect 20588 15499 20674 15735
rect 20910 15499 20996 15735
rect 21232 15499 21318 15735
rect 21554 15499 21640 15735
rect 21876 15499 21962 15735
rect 22198 15499 22284 15735
rect 22520 15499 22606 15735
rect 22842 15499 22928 15735
rect 23164 15499 23250 15735
rect 23486 15499 23572 15735
rect 23808 15499 23894 15735
rect 24130 15499 24216 15735
rect 24452 15499 24640 15735
rect -3360 15399 24640 15499
rect -3360 15163 -3185 15399
rect -2949 15163 -2862 15399
rect -2626 15163 -2539 15399
rect -2303 15163 -2216 15399
rect -1980 15163 -1893 15399
rect -1657 15163 -1570 15399
rect -1334 15163 -1247 15399
rect -1011 15163 -924 15399
rect -688 15163 -601 15399
rect -365 15163 -278 15399
rect -42 15163 45 15399
rect 281 15163 368 15399
rect 604 15163 691 15399
rect 927 15163 1014 15399
rect 1250 15163 1337 15399
rect 1573 15163 1660 15399
rect 1896 15163 1983 15399
rect 2219 15163 2306 15399
rect 2542 15163 2629 15399
rect 2865 15163 2952 15399
rect 3188 15163 3275 15399
rect 3511 15163 3598 15399
rect 3834 15163 3921 15399
rect 4157 15163 4244 15399
rect 4480 15163 4567 15399
rect 4803 15163 4890 15399
rect 5126 15163 5213 15399
rect 5449 15163 5536 15399
rect 5772 15163 5859 15399
rect 6095 15163 6182 15399
rect 6418 15163 6505 15399
rect 6741 15163 6828 15399
rect 7064 15163 7150 15399
rect 7386 15163 7472 15399
rect 7708 15163 7794 15399
rect 8030 15163 8116 15399
rect 8352 15163 8438 15399
rect 8674 15163 8760 15399
rect 8996 15163 9082 15399
rect 9318 15163 9404 15399
rect 9640 15163 9726 15399
rect 9962 15163 10048 15399
rect 10284 15163 10370 15399
rect 10606 15163 10692 15399
rect 10928 15163 11014 15399
rect 11250 15163 11336 15399
rect 11572 15163 11658 15399
rect 11894 15163 11980 15399
rect 12216 15163 12302 15399
rect 12538 15163 12624 15399
rect 12860 15163 12946 15399
rect 13182 15163 13268 15399
rect 13504 15163 13590 15399
rect 13826 15163 13912 15399
rect 14148 15163 14234 15399
rect 14470 15163 14556 15399
rect 14792 15163 14878 15399
rect 15114 15163 15200 15399
rect 15436 15163 15522 15399
rect 15758 15163 15844 15399
rect 16080 15163 16166 15399
rect 16402 15163 16488 15399
rect 16724 15163 16810 15399
rect 17046 15163 17132 15399
rect 17368 15163 17454 15399
rect 17690 15163 17776 15399
rect 18012 15163 18098 15399
rect 18334 15163 18420 15399
rect 18656 15163 18742 15399
rect 18978 15163 19064 15399
rect 19300 15163 19386 15399
rect 19622 15163 19708 15399
rect 19944 15163 20030 15399
rect 20266 15163 20352 15399
rect 20588 15163 20674 15399
rect 20910 15163 20996 15399
rect 21232 15163 21318 15399
rect 21554 15163 21640 15399
rect 21876 15163 21962 15399
rect 22198 15163 22284 15399
rect 22520 15163 22606 15399
rect 22842 15163 22928 15399
rect 23164 15163 23250 15399
rect 23486 15163 23572 15399
rect 23808 15163 23894 15399
rect 24130 15163 24216 15399
rect 24452 15163 24640 15399
rect -3360 15063 24640 15163
rect -3360 14827 -3185 15063
rect -2949 14827 -2862 15063
rect -2626 14827 -2539 15063
rect -2303 14827 -2216 15063
rect -1980 14827 -1893 15063
rect -1657 14827 -1570 15063
rect -1334 14827 -1247 15063
rect -1011 14827 -924 15063
rect -688 14827 -601 15063
rect -365 14827 -278 15063
rect -42 14827 45 15063
rect 281 14827 368 15063
rect 604 14827 691 15063
rect 927 14827 1014 15063
rect 1250 14827 1337 15063
rect 1573 14827 1660 15063
rect 1896 14827 1983 15063
rect 2219 14827 2306 15063
rect 2542 14827 2629 15063
rect 2865 14827 2952 15063
rect 3188 14827 3275 15063
rect 3511 14827 3598 15063
rect 3834 14827 3921 15063
rect 4157 14827 4244 15063
rect 4480 14827 4567 15063
rect 4803 14827 4890 15063
rect 5126 14827 5213 15063
rect 5449 14827 5536 15063
rect 5772 14827 5859 15063
rect 6095 14827 6182 15063
rect 6418 14827 6505 15063
rect 6741 14827 6828 15063
rect 7064 14827 7150 15063
rect 7386 14827 7472 15063
rect 7708 14827 7794 15063
rect 8030 14827 8116 15063
rect 8352 14827 8438 15063
rect 8674 14827 8760 15063
rect 8996 14827 9082 15063
rect 9318 14827 9404 15063
rect 9640 14827 9726 15063
rect 9962 14827 10048 15063
rect 10284 14827 10370 15063
rect 10606 14827 10692 15063
rect 10928 14827 11014 15063
rect 11250 14827 11336 15063
rect 11572 14827 11658 15063
rect 11894 14827 11980 15063
rect 12216 14827 12302 15063
rect 12538 14827 12624 15063
rect 12860 14827 12946 15063
rect 13182 14827 13268 15063
rect 13504 14827 13590 15063
rect 13826 14827 13912 15063
rect 14148 14827 14234 15063
rect 14470 14827 14556 15063
rect 14792 14827 14878 15063
rect 15114 14827 15200 15063
rect 15436 14827 15522 15063
rect 15758 14827 15844 15063
rect 16080 14827 16166 15063
rect 16402 14827 16488 15063
rect 16724 14827 16810 15063
rect 17046 14827 17132 15063
rect 17368 14827 17454 15063
rect 17690 14827 17776 15063
rect 18012 14827 18098 15063
rect 18334 14827 18420 15063
rect 18656 14827 18742 15063
rect 18978 14827 19064 15063
rect 19300 14827 19386 15063
rect 19622 14827 19708 15063
rect 19944 14827 20030 15063
rect 20266 14827 20352 15063
rect 20588 14827 20674 15063
rect 20910 14827 20996 15063
rect 21232 14827 21318 15063
rect 21554 14827 21640 15063
rect 21876 14827 21962 15063
rect 22198 14827 22284 15063
rect 22520 14827 22606 15063
rect 22842 14827 22928 15063
rect 23164 14827 23250 15063
rect 23486 14827 23572 15063
rect 23808 14827 23894 15063
rect 24130 14827 24216 15063
rect 24452 14827 24640 15063
rect -3360 14727 24640 14827
rect -3360 14491 -3185 14727
rect -2949 14491 -2862 14727
rect -2626 14491 -2539 14727
rect -2303 14491 -2216 14727
rect -1980 14491 -1893 14727
rect -1657 14491 -1570 14727
rect -1334 14491 -1247 14727
rect -1011 14491 -924 14727
rect -688 14491 -601 14727
rect -365 14491 -278 14727
rect -42 14491 45 14727
rect 281 14491 368 14727
rect 604 14491 691 14727
rect 927 14491 1014 14727
rect 1250 14491 1337 14727
rect 1573 14491 1660 14727
rect 1896 14491 1983 14727
rect 2219 14491 2306 14727
rect 2542 14491 2629 14727
rect 2865 14491 2952 14727
rect 3188 14491 3275 14727
rect 3511 14491 3598 14727
rect 3834 14491 3921 14727
rect 4157 14491 4244 14727
rect 4480 14491 4567 14727
rect 4803 14491 4890 14727
rect 5126 14491 5213 14727
rect 5449 14491 5536 14727
rect 5772 14491 5859 14727
rect 6095 14491 6182 14727
rect 6418 14491 6505 14727
rect 6741 14491 6828 14727
rect 7064 14491 7150 14727
rect 7386 14491 7472 14727
rect 7708 14491 7794 14727
rect 8030 14491 8116 14727
rect 8352 14491 8438 14727
rect 8674 14491 8760 14727
rect 8996 14491 9082 14727
rect 9318 14491 9404 14727
rect 9640 14491 9726 14727
rect 9962 14491 10048 14727
rect 10284 14491 10370 14727
rect 10606 14491 10692 14727
rect 10928 14491 11014 14727
rect 11250 14491 11336 14727
rect 11572 14491 11658 14727
rect 11894 14491 11980 14727
rect 12216 14491 12302 14727
rect 12538 14491 12624 14727
rect 12860 14491 12946 14727
rect 13182 14491 13268 14727
rect 13504 14491 13590 14727
rect 13826 14491 13912 14727
rect 14148 14491 14234 14727
rect 14470 14491 14556 14727
rect 14792 14491 14878 14727
rect 15114 14491 15200 14727
rect 15436 14491 15522 14727
rect 15758 14491 15844 14727
rect 16080 14491 16166 14727
rect 16402 14491 16488 14727
rect 16724 14491 16810 14727
rect 17046 14491 17132 14727
rect 17368 14491 17454 14727
rect 17690 14491 17776 14727
rect 18012 14491 18098 14727
rect 18334 14491 18420 14727
rect 18656 14491 18742 14727
rect 18978 14491 19064 14727
rect 19300 14491 19386 14727
rect 19622 14491 19708 14727
rect 19944 14491 20030 14727
rect 20266 14491 20352 14727
rect 20588 14491 20674 14727
rect 20910 14491 20996 14727
rect 21232 14491 21318 14727
rect 21554 14491 21640 14727
rect 21876 14491 21962 14727
rect 22198 14491 22284 14727
rect 22520 14491 22606 14727
rect 22842 14491 22928 14727
rect 23164 14491 23250 14727
rect 23486 14491 23572 14727
rect 23808 14491 23894 14727
rect 24130 14491 24216 14727
rect 24452 14491 24640 14727
rect -3360 14391 24640 14491
rect -3360 14155 -3185 14391
rect -2949 14155 -2862 14391
rect -2626 14155 -2539 14391
rect -2303 14155 -2216 14391
rect -1980 14155 -1893 14391
rect -1657 14155 -1570 14391
rect -1334 14155 -1247 14391
rect -1011 14155 -924 14391
rect -688 14155 -601 14391
rect -365 14155 -278 14391
rect -42 14155 45 14391
rect 281 14155 368 14391
rect 604 14155 691 14391
rect 927 14155 1014 14391
rect 1250 14155 1337 14391
rect 1573 14155 1660 14391
rect 1896 14155 1983 14391
rect 2219 14155 2306 14391
rect 2542 14155 2629 14391
rect 2865 14155 2952 14391
rect 3188 14155 3275 14391
rect 3511 14155 3598 14391
rect 3834 14155 3921 14391
rect 4157 14155 4244 14391
rect 4480 14155 4567 14391
rect 4803 14155 4890 14391
rect 5126 14155 5213 14391
rect 5449 14155 5536 14391
rect 5772 14155 5859 14391
rect 6095 14155 6182 14391
rect 6418 14155 6505 14391
rect 6741 14155 6828 14391
rect 7064 14155 7150 14391
rect 7386 14155 7472 14391
rect 7708 14155 7794 14391
rect 8030 14155 8116 14391
rect 8352 14155 8438 14391
rect 8674 14155 8760 14391
rect 8996 14155 9082 14391
rect 9318 14155 9404 14391
rect 9640 14155 9726 14391
rect 9962 14155 10048 14391
rect 10284 14155 10370 14391
rect 10606 14155 10692 14391
rect 10928 14155 11014 14391
rect 11250 14155 11336 14391
rect 11572 14155 11658 14391
rect 11894 14155 11980 14391
rect 12216 14155 12302 14391
rect 12538 14155 12624 14391
rect 12860 14155 12946 14391
rect 13182 14155 13268 14391
rect 13504 14155 13590 14391
rect 13826 14155 13912 14391
rect 14148 14155 14234 14391
rect 14470 14155 14556 14391
rect 14792 14155 14878 14391
rect 15114 14155 15200 14391
rect 15436 14155 15522 14391
rect 15758 14155 15844 14391
rect 16080 14155 16166 14391
rect 16402 14155 16488 14391
rect 16724 14155 16810 14391
rect 17046 14155 17132 14391
rect 17368 14155 17454 14391
rect 17690 14155 17776 14391
rect 18012 14155 18098 14391
rect 18334 14155 18420 14391
rect 18656 14155 18742 14391
rect 18978 14155 19064 14391
rect 19300 14155 19386 14391
rect 19622 14155 19708 14391
rect 19944 14155 20030 14391
rect 20266 14155 20352 14391
rect 20588 14155 20674 14391
rect 20910 14155 20996 14391
rect 21232 14155 21318 14391
rect 21554 14155 21640 14391
rect 21876 14155 21962 14391
rect 22198 14155 22284 14391
rect 22520 14155 22606 14391
rect 22842 14155 22928 14391
rect 23164 14155 23250 14391
rect 23486 14155 23572 14391
rect 23808 14155 23894 14391
rect 24130 14155 24216 14391
rect 24452 14155 24640 14391
rect -3360 14055 24640 14155
rect -3360 13819 -3185 14055
rect -2949 13819 -2862 14055
rect -2626 13819 -2539 14055
rect -2303 13819 -2216 14055
rect -1980 13819 -1893 14055
rect -1657 13819 -1570 14055
rect -1334 13819 -1247 14055
rect -1011 13819 -924 14055
rect -688 13819 -601 14055
rect -365 13819 -278 14055
rect -42 13819 45 14055
rect 281 13819 368 14055
rect 604 13819 691 14055
rect 927 13819 1014 14055
rect 1250 13819 1337 14055
rect 1573 13819 1660 14055
rect 1896 13819 1983 14055
rect 2219 13819 2306 14055
rect 2542 13819 2629 14055
rect 2865 13819 2952 14055
rect 3188 13819 3275 14055
rect 3511 13819 3598 14055
rect 3834 13819 3921 14055
rect 4157 13819 4244 14055
rect 4480 13819 4567 14055
rect 4803 13819 4890 14055
rect 5126 13819 5213 14055
rect 5449 13819 5536 14055
rect 5772 13819 5859 14055
rect 6095 13819 6182 14055
rect 6418 13819 6505 14055
rect 6741 13819 6828 14055
rect 7064 13819 7150 14055
rect 7386 13819 7472 14055
rect 7708 13819 7794 14055
rect 8030 13819 8116 14055
rect 8352 13819 8438 14055
rect 8674 13819 8760 14055
rect 8996 13819 9082 14055
rect 9318 13819 9404 14055
rect 9640 13819 9726 14055
rect 9962 13819 10048 14055
rect 10284 13819 10370 14055
rect 10606 13819 10692 14055
rect 10928 13819 11014 14055
rect 11250 13819 11336 14055
rect 11572 13819 11658 14055
rect 11894 13819 11980 14055
rect 12216 13819 12302 14055
rect 12538 13819 12624 14055
rect 12860 13819 12946 14055
rect 13182 13819 13268 14055
rect 13504 13819 13590 14055
rect 13826 13819 13912 14055
rect 14148 13819 14234 14055
rect 14470 13819 14556 14055
rect 14792 13819 14878 14055
rect 15114 13819 15200 14055
rect 15436 13819 15522 14055
rect 15758 13819 15844 14055
rect 16080 13819 16166 14055
rect 16402 13819 16488 14055
rect 16724 13819 16810 14055
rect 17046 13819 17132 14055
rect 17368 13819 17454 14055
rect 17690 13819 17776 14055
rect 18012 13819 18098 14055
rect 18334 13819 18420 14055
rect 18656 13819 18742 14055
rect 18978 13819 19064 14055
rect 19300 13819 19386 14055
rect 19622 13819 19708 14055
rect 19944 13819 20030 14055
rect 20266 13819 20352 14055
rect 20588 13819 20674 14055
rect 20910 13819 20996 14055
rect 21232 13819 21318 14055
rect 21554 13819 21640 14055
rect 21876 13819 21962 14055
rect 22198 13819 22284 14055
rect 22520 13819 22606 14055
rect 22842 13819 22928 14055
rect 23164 13819 23250 14055
rect 23486 13819 23572 14055
rect 23808 13819 23894 14055
rect 24130 13819 24216 14055
rect 24452 13819 24640 14055
rect -3360 13719 24640 13819
rect -3360 13483 -3185 13719
rect -2949 13483 -2862 13719
rect -2626 13483 -2539 13719
rect -2303 13483 -2216 13719
rect -1980 13483 -1893 13719
rect -1657 13483 -1570 13719
rect -1334 13483 -1247 13719
rect -1011 13483 -924 13719
rect -688 13483 -601 13719
rect -365 13483 -278 13719
rect -42 13483 45 13719
rect 281 13483 368 13719
rect 604 13483 691 13719
rect 927 13483 1014 13719
rect 1250 13483 1337 13719
rect 1573 13483 1660 13719
rect 1896 13483 1983 13719
rect 2219 13483 2306 13719
rect 2542 13483 2629 13719
rect 2865 13483 2952 13719
rect 3188 13483 3275 13719
rect 3511 13483 3598 13719
rect 3834 13483 3921 13719
rect 4157 13483 4244 13719
rect 4480 13483 4567 13719
rect 4803 13483 4890 13719
rect 5126 13483 5213 13719
rect 5449 13483 5536 13719
rect 5772 13483 5859 13719
rect 6095 13483 6182 13719
rect 6418 13483 6505 13719
rect 6741 13483 6828 13719
rect 7064 13483 7150 13719
rect 7386 13483 7472 13719
rect 7708 13483 7794 13719
rect 8030 13483 8116 13719
rect 8352 13483 8438 13719
rect 8674 13483 8760 13719
rect 8996 13483 9082 13719
rect 9318 13483 9404 13719
rect 9640 13483 9726 13719
rect 9962 13483 10048 13719
rect 10284 13483 10370 13719
rect 10606 13483 10692 13719
rect 10928 13483 11014 13719
rect 11250 13483 11336 13719
rect 11572 13483 11658 13719
rect 11894 13483 11980 13719
rect 12216 13483 12302 13719
rect 12538 13483 12624 13719
rect 12860 13483 12946 13719
rect 13182 13483 13268 13719
rect 13504 13483 13590 13719
rect 13826 13483 13912 13719
rect 14148 13483 14234 13719
rect 14470 13483 14556 13719
rect 14792 13483 14878 13719
rect 15114 13483 15200 13719
rect 15436 13483 15522 13719
rect 15758 13483 15844 13719
rect 16080 13483 16166 13719
rect 16402 13483 16488 13719
rect 16724 13483 16810 13719
rect 17046 13483 17132 13719
rect 17368 13483 17454 13719
rect 17690 13483 17776 13719
rect 18012 13483 18098 13719
rect 18334 13483 18420 13719
rect 18656 13483 18742 13719
rect 18978 13483 19064 13719
rect 19300 13483 19386 13719
rect 19622 13483 19708 13719
rect 19944 13483 20030 13719
rect 20266 13483 20352 13719
rect 20588 13483 20674 13719
rect 20910 13483 20996 13719
rect 21232 13483 21318 13719
rect 21554 13483 21640 13719
rect 21876 13483 21962 13719
rect 22198 13483 22284 13719
rect 22520 13483 22606 13719
rect 22842 13483 22928 13719
rect 23164 13483 23250 13719
rect 23486 13483 23572 13719
rect 23808 13483 23894 13719
rect 24130 13483 24216 13719
rect 24452 13483 24640 13719
rect -3360 13482 24640 13483
rect -3360 13458 -2720 13482
rect 24000 13458 24640 13482
rect -3360 13114 -2720 13158
rect 24000 13114 24640 13158
rect -3360 12878 -3185 13114
rect -2949 12878 -2862 13114
rect -2626 12878 -2539 13114
rect -2303 12878 -2216 13114
rect -1980 12878 -1893 13114
rect -1657 12878 -1570 13114
rect -1334 12878 -1247 13114
rect -1011 12878 -924 13114
rect -688 12878 -601 13114
rect -365 12878 -278 13114
rect -42 12878 45 13114
rect 281 12878 368 13114
rect 604 12878 691 13114
rect 927 12878 1014 13114
rect 1250 12878 1337 13114
rect 1573 12878 1660 13114
rect 1896 12878 1983 13114
rect 2219 12878 2306 13114
rect 2542 12878 2629 13114
rect 2865 12878 2952 13114
rect 3188 12878 3275 13114
rect 3511 12878 3598 13114
rect 3834 12878 3921 13114
rect 4157 12878 4244 13114
rect 4480 12878 4567 13114
rect 4803 12878 4890 13114
rect 5126 12878 5213 13114
rect 5449 12878 5536 13114
rect 5772 12878 5859 13114
rect 6095 12878 6182 13114
rect 6418 12878 6504 13114
rect 6740 12878 6826 13114
rect 7062 12878 7148 13114
rect 7384 12878 7470 13114
rect 7706 12878 7792 13114
rect 8028 12878 8114 13114
rect 8350 12878 8436 13114
rect 8672 12878 8758 13114
rect 8994 12878 9080 13114
rect 9316 12878 9402 13114
rect 9638 12878 9724 13114
rect 9960 12878 10046 13114
rect 10282 12878 10368 13114
rect 10604 12878 10690 13114
rect 10926 12878 11012 13114
rect 11248 12878 11334 13114
rect 11570 12878 11656 13114
rect 11892 12878 11978 13114
rect 12214 12878 12300 13114
rect 12536 12878 12622 13114
rect 12858 12878 12944 13114
rect 13180 12878 13266 13114
rect 13502 12878 13588 13114
rect 13824 12878 13910 13114
rect 14146 12878 14232 13114
rect 14468 12878 14554 13114
rect 14790 12878 14876 13114
rect 15112 12878 15198 13114
rect 15434 12878 15520 13114
rect 15756 12878 15842 13114
rect 16078 12878 16164 13114
rect 16400 12878 16486 13114
rect 16722 12878 16808 13114
rect 17044 12878 17130 13114
rect 17366 12878 17452 13114
rect 17688 12878 17774 13114
rect 18010 12878 18096 13114
rect 18332 12878 18418 13114
rect 18654 12878 18740 13114
rect 18976 12878 19062 13114
rect 19298 12878 19384 13114
rect 19620 12878 19706 13114
rect 19942 12878 20028 13114
rect 20264 12878 20350 13114
rect 20586 12878 20672 13114
rect 20908 12878 20994 13114
rect 21230 12878 21316 13114
rect 21552 12878 21638 13114
rect 21874 12878 21960 13114
rect 22196 12878 22282 13114
rect 22518 12878 22604 13114
rect 22840 12878 22926 13114
rect 23162 12878 23248 13114
rect 23484 12878 23570 13114
rect 23806 12878 23892 13114
rect 24128 12878 24214 13114
rect 24450 12878 24640 13114
rect -3360 12548 24640 12878
rect -3360 12312 -3185 12548
rect -2949 12312 -2862 12548
rect -2626 12312 -2539 12548
rect -2303 12312 -2216 12548
rect -1980 12312 -1893 12548
rect -1657 12312 -1570 12548
rect -1334 12312 -1247 12548
rect -1011 12312 -924 12548
rect -688 12312 -601 12548
rect -365 12312 -278 12548
rect -42 12312 45 12548
rect 281 12312 368 12548
rect 604 12312 691 12548
rect 927 12312 1014 12548
rect 1250 12312 1337 12548
rect 1573 12312 1660 12548
rect 1896 12312 1983 12548
rect 2219 12312 2306 12548
rect 2542 12312 2629 12548
rect 2865 12312 2952 12548
rect 3188 12312 3275 12548
rect 3511 12312 3598 12548
rect 3834 12312 3921 12548
rect 4157 12312 4244 12548
rect 4480 12312 4567 12548
rect 4803 12312 4890 12548
rect 5126 12312 5213 12548
rect 5449 12312 5536 12548
rect 5772 12312 5859 12548
rect 6095 12312 6182 12548
rect 6418 12312 6504 12548
rect 6740 12312 6826 12548
rect 7062 12312 7148 12548
rect 7384 12312 7470 12548
rect 7706 12312 7792 12548
rect 8028 12312 8114 12548
rect 8350 12312 8436 12548
rect 8672 12312 8758 12548
rect 8994 12312 9080 12548
rect 9316 12312 9402 12548
rect 9638 12312 9724 12548
rect 9960 12312 10046 12548
rect 10282 12312 10368 12548
rect 10604 12312 10690 12548
rect 10926 12312 11012 12548
rect 11248 12312 11334 12548
rect 11570 12312 11656 12548
rect 11892 12312 11978 12548
rect 12214 12312 12300 12548
rect 12536 12312 12622 12548
rect 12858 12312 12944 12548
rect 13180 12312 13266 12548
rect 13502 12312 13588 12548
rect 13824 12312 13910 12548
rect 14146 12312 14232 12548
rect 14468 12312 14554 12548
rect 14790 12312 14876 12548
rect 15112 12312 15198 12548
rect 15434 12312 15520 12548
rect 15756 12312 15842 12548
rect 16078 12312 16164 12548
rect 16400 12312 16486 12548
rect 16722 12312 16808 12548
rect 17044 12312 17130 12548
rect 17366 12312 17452 12548
rect 17688 12312 17774 12548
rect 18010 12312 18096 12548
rect 18332 12312 18418 12548
rect 18654 12312 18740 12548
rect 18976 12312 19062 12548
rect 19298 12312 19384 12548
rect 19620 12312 19706 12548
rect 19942 12312 20028 12548
rect 20264 12312 20350 12548
rect 20586 12312 20672 12548
rect 20908 12312 20994 12548
rect 21230 12312 21316 12548
rect 21552 12312 21638 12548
rect 21874 12312 21960 12548
rect 22196 12312 22282 12548
rect 22518 12312 22604 12548
rect 22840 12312 22926 12548
rect 23162 12312 23248 12548
rect 23484 12312 23570 12548
rect 23806 12312 23892 12548
rect 24128 12312 24214 12548
rect 24450 12312 24640 12548
rect -3360 12268 -2720 12312
rect 24000 12268 24640 12312
rect -3360 11944 -2720 11988
rect 24000 11944 24640 11988
rect -3360 11708 -3185 11944
rect -2949 11708 -2862 11944
rect -2626 11708 -2539 11944
rect -2303 11708 -2216 11944
rect -1980 11708 -1893 11944
rect -1657 11708 -1570 11944
rect -1334 11708 -1247 11944
rect -1011 11708 -924 11944
rect -688 11708 -601 11944
rect -365 11708 -278 11944
rect -42 11708 45 11944
rect 281 11708 368 11944
rect 604 11708 691 11944
rect 927 11708 1014 11944
rect 1250 11708 1337 11944
rect 1573 11708 1660 11944
rect 1896 11708 1983 11944
rect 2219 11708 2306 11944
rect 2542 11708 2629 11944
rect 2865 11708 2952 11944
rect 3188 11708 3275 11944
rect 3511 11708 3598 11944
rect 3834 11708 3921 11944
rect 4157 11708 4244 11944
rect 4480 11708 4567 11944
rect 4803 11708 4890 11944
rect 5126 11708 5213 11944
rect 5449 11708 5536 11944
rect 5772 11708 5859 11944
rect 6095 11708 6182 11944
rect 6418 11708 6504 11944
rect 6740 11708 6826 11944
rect 7062 11708 7148 11944
rect 7384 11708 7470 11944
rect 7706 11708 7792 11944
rect 8028 11708 8114 11944
rect 8350 11708 8436 11944
rect 8672 11708 8758 11944
rect 8994 11708 9080 11944
rect 9316 11708 9402 11944
rect 9638 11708 9724 11944
rect 9960 11708 10046 11944
rect 10282 11708 10368 11944
rect 10604 11708 10690 11944
rect 10926 11708 11012 11944
rect 11248 11708 11334 11944
rect 11570 11708 11656 11944
rect 11892 11708 11978 11944
rect 12214 11708 12300 11944
rect 12536 11708 12622 11944
rect 12858 11708 12944 11944
rect 13180 11708 13266 11944
rect 13502 11708 13588 11944
rect 13824 11708 13910 11944
rect 14146 11708 14232 11944
rect 14468 11708 14554 11944
rect 14790 11708 14876 11944
rect 15112 11708 15198 11944
rect 15434 11708 15520 11944
rect 15756 11708 15842 11944
rect 16078 11708 16164 11944
rect 16400 11708 16486 11944
rect 16722 11708 16808 11944
rect 17044 11708 17130 11944
rect 17366 11708 17452 11944
rect 17688 11708 17774 11944
rect 18010 11708 18096 11944
rect 18332 11708 18418 11944
rect 18654 11708 18740 11944
rect 18976 11708 19062 11944
rect 19298 11708 19384 11944
rect 19620 11708 19706 11944
rect 19942 11708 20028 11944
rect 20264 11708 20350 11944
rect 20586 11708 20672 11944
rect 20908 11708 20994 11944
rect 21230 11708 21316 11944
rect 21552 11708 21638 11944
rect 21874 11708 21960 11944
rect 22196 11708 22282 11944
rect 22518 11708 22604 11944
rect 22840 11708 22926 11944
rect 23162 11708 23248 11944
rect 23484 11708 23570 11944
rect 23806 11708 23892 11944
rect 24128 11708 24214 11944
rect 24450 11708 24640 11944
rect -3360 11378 24640 11708
rect -3360 11142 -3185 11378
rect -2949 11142 -2862 11378
rect -2626 11142 -2539 11378
rect -2303 11142 -2216 11378
rect -1980 11142 -1893 11378
rect -1657 11142 -1570 11378
rect -1334 11142 -1247 11378
rect -1011 11142 -924 11378
rect -688 11142 -601 11378
rect -365 11142 -278 11378
rect -42 11142 45 11378
rect 281 11142 368 11378
rect 604 11142 691 11378
rect 927 11142 1014 11378
rect 1250 11142 1337 11378
rect 1573 11142 1660 11378
rect 1896 11142 1983 11378
rect 2219 11142 2306 11378
rect 2542 11142 2629 11378
rect 2865 11142 2952 11378
rect 3188 11142 3275 11378
rect 3511 11142 3598 11378
rect 3834 11142 3921 11378
rect 4157 11142 4244 11378
rect 4480 11142 4567 11378
rect 4803 11142 4890 11378
rect 5126 11142 5213 11378
rect 5449 11142 5536 11378
rect 5772 11142 5859 11378
rect 6095 11142 6182 11378
rect 6418 11142 6504 11378
rect 6740 11142 6826 11378
rect 7062 11142 7148 11378
rect 7384 11142 7470 11378
rect 7706 11142 7792 11378
rect 8028 11142 8114 11378
rect 8350 11142 8436 11378
rect 8672 11142 8758 11378
rect 8994 11142 9080 11378
rect 9316 11142 9402 11378
rect 9638 11142 9724 11378
rect 9960 11142 10046 11378
rect 10282 11142 10368 11378
rect 10604 11142 10690 11378
rect 10926 11142 11012 11378
rect 11248 11142 11334 11378
rect 11570 11142 11656 11378
rect 11892 11142 11978 11378
rect 12214 11142 12300 11378
rect 12536 11142 12622 11378
rect 12858 11142 12944 11378
rect 13180 11142 13266 11378
rect 13502 11142 13588 11378
rect 13824 11142 13910 11378
rect 14146 11142 14232 11378
rect 14468 11142 14554 11378
rect 14790 11142 14876 11378
rect 15112 11142 15198 11378
rect 15434 11142 15520 11378
rect 15756 11142 15842 11378
rect 16078 11142 16164 11378
rect 16400 11142 16486 11378
rect 16722 11142 16808 11378
rect 17044 11142 17130 11378
rect 17366 11142 17452 11378
rect 17688 11142 17774 11378
rect 18010 11142 18096 11378
rect 18332 11142 18418 11378
rect 18654 11142 18740 11378
rect 18976 11142 19062 11378
rect 19298 11142 19384 11378
rect 19620 11142 19706 11378
rect 19942 11142 20028 11378
rect 20264 11142 20350 11378
rect 20586 11142 20672 11378
rect 20908 11142 20994 11378
rect 21230 11142 21316 11378
rect 21552 11142 21638 11378
rect 21874 11142 21960 11378
rect 22196 11142 22282 11378
rect 22518 11142 22604 11378
rect 22840 11142 22926 11378
rect 23162 11142 23248 11378
rect 23484 11142 23570 11378
rect 23806 11142 23892 11378
rect 24128 11142 24214 11378
rect 24450 11142 24640 11378
rect -3360 11098 -2720 11142
rect 24000 11098 24640 11142
rect -3360 10732 -2720 10798
rect 24000 10732 24640 10798
rect -3360 10076 -2720 10672
rect 24000 10076 24640 10672
rect -3360 9780 -2720 10016
rect 24000 9780 24640 10016
rect -3360 9124 -2720 9720
rect 24000 9124 24640 9720
rect -3360 8998 -2720 9064
rect 24000 8998 24640 9064
rect -3360 8654 -2720 8698
rect 24000 8654 24640 8698
rect -3360 8418 -3185 8654
rect -2949 8418 -2862 8654
rect -2626 8418 -2539 8654
rect -2303 8418 -2216 8654
rect -1980 8418 -1893 8654
rect -1657 8418 -1570 8654
rect -1334 8418 -1247 8654
rect -1011 8418 -924 8654
rect -688 8418 -601 8654
rect -365 8418 -278 8654
rect -42 8418 45 8654
rect 281 8418 368 8654
rect 604 8418 691 8654
rect 927 8418 1014 8654
rect 1250 8418 1337 8654
rect 1573 8418 1660 8654
rect 1896 8418 1983 8654
rect 2219 8418 2306 8654
rect 2542 8418 2629 8654
rect 2865 8418 2952 8654
rect 3188 8418 3275 8654
rect 3511 8418 3598 8654
rect 3834 8418 3921 8654
rect 4157 8418 4244 8654
rect 4480 8418 4567 8654
rect 4803 8418 4890 8654
rect 5126 8418 5213 8654
rect 5449 8418 5536 8654
rect 5772 8418 5859 8654
rect 6095 8418 6182 8654
rect 6418 8418 6505 8654
rect 6741 8418 6828 8654
rect 7064 8418 7150 8654
rect 7386 8418 7472 8654
rect 7708 8418 7794 8654
rect 8030 8418 8116 8654
rect 8352 8418 8438 8654
rect 8674 8418 8760 8654
rect 8996 8418 9082 8654
rect 9318 8418 9404 8654
rect 9640 8418 9726 8654
rect 9962 8418 10048 8654
rect 10284 8418 10370 8654
rect 10606 8418 10692 8654
rect 10928 8418 11014 8654
rect 11250 8418 11336 8654
rect 11572 8418 11658 8654
rect 11894 8418 11980 8654
rect 12216 8418 12302 8654
rect 12538 8418 12624 8654
rect 12860 8418 12946 8654
rect 13182 8418 13268 8654
rect 13504 8418 13590 8654
rect 13826 8418 13912 8654
rect 14148 8418 14234 8654
rect 14470 8418 14556 8654
rect 14792 8418 14878 8654
rect 15114 8418 15200 8654
rect 15436 8418 15522 8654
rect 15758 8418 15844 8654
rect 16080 8418 16166 8654
rect 16402 8418 16488 8654
rect 16724 8418 16810 8654
rect 17046 8418 17132 8654
rect 17368 8418 17454 8654
rect 17690 8418 17776 8654
rect 18012 8418 18098 8654
rect 18334 8418 18420 8654
rect 18656 8418 18742 8654
rect 18978 8418 19064 8654
rect 19300 8418 19386 8654
rect 19622 8418 19708 8654
rect 19944 8418 20030 8654
rect 20266 8418 20352 8654
rect 20588 8418 20674 8654
rect 20910 8418 20996 8654
rect 21232 8418 21318 8654
rect 21554 8418 21640 8654
rect 21876 8418 21962 8654
rect 22198 8418 22284 8654
rect 22520 8418 22606 8654
rect 22842 8418 22928 8654
rect 23164 8418 23250 8654
rect 23486 8418 23572 8654
rect 23808 8418 23894 8654
rect 24130 8418 24216 8654
rect 24452 8418 24640 8654
rect -3360 8048 24640 8418
rect -3360 7812 -3185 8048
rect -2949 7812 -2862 8048
rect -2626 7812 -2539 8048
rect -2303 7812 -2216 8048
rect -1980 7812 -1893 8048
rect -1657 7812 -1570 8048
rect -1334 7812 -1247 8048
rect -1011 7812 -924 8048
rect -688 7812 -601 8048
rect -365 7812 -278 8048
rect -42 7812 45 8048
rect 281 7812 368 8048
rect 604 7812 691 8048
rect 927 7812 1014 8048
rect 1250 7812 1337 8048
rect 1573 7812 1660 8048
rect 1896 7812 1983 8048
rect 2219 7812 2306 8048
rect 2542 7812 2629 8048
rect 2865 7812 2952 8048
rect 3188 7812 3275 8048
rect 3511 7812 3598 8048
rect 3834 7812 3921 8048
rect 4157 7812 4244 8048
rect 4480 7812 4567 8048
rect 4803 7812 4890 8048
rect 5126 7812 5213 8048
rect 5449 7812 5536 8048
rect 5772 7812 5859 8048
rect 6095 7812 6182 8048
rect 6418 7812 6505 8048
rect 6741 7812 6828 8048
rect 7064 7812 7150 8048
rect 7386 7812 7472 8048
rect 7708 7812 7794 8048
rect 8030 7812 8116 8048
rect 8352 7812 8438 8048
rect 8674 7812 8760 8048
rect 8996 7812 9082 8048
rect 9318 7812 9404 8048
rect 9640 7812 9726 8048
rect 9962 7812 10048 8048
rect 10284 7812 10370 8048
rect 10606 7812 10692 8048
rect 10928 7812 11014 8048
rect 11250 7812 11336 8048
rect 11572 7812 11658 8048
rect 11894 7812 11980 8048
rect 12216 7812 12302 8048
rect 12538 7812 12624 8048
rect 12860 7812 12946 8048
rect 13182 7812 13268 8048
rect 13504 7812 13590 8048
rect 13826 7812 13912 8048
rect 14148 7812 14234 8048
rect 14470 7812 14556 8048
rect 14792 7812 14878 8048
rect 15114 7812 15200 8048
rect 15436 7812 15522 8048
rect 15758 7812 15844 8048
rect 16080 7812 16166 8048
rect 16402 7812 16488 8048
rect 16724 7812 16810 8048
rect 17046 7812 17132 8048
rect 17368 7812 17454 8048
rect 17690 7812 17776 8048
rect 18012 7812 18098 8048
rect 18334 7812 18420 8048
rect 18656 7812 18742 8048
rect 18978 7812 19064 8048
rect 19300 7812 19386 8048
rect 19622 7812 19708 8048
rect 19944 7812 20030 8048
rect 20266 7812 20352 8048
rect 20588 7812 20674 8048
rect 20910 7812 20996 8048
rect 21232 7812 21318 8048
rect 21554 7812 21640 8048
rect 21876 7812 21962 8048
rect 22198 7812 22284 8048
rect 22520 7812 22606 8048
rect 22842 7812 22928 8048
rect 23164 7812 23250 8048
rect 23486 7812 23572 8048
rect 23808 7812 23894 8048
rect 24130 7812 24216 8048
rect 24452 7812 24640 8048
rect -3360 7768 -2720 7812
rect 24000 7768 24640 7812
rect -3360 7444 -2720 7488
rect 24000 7444 24640 7488
rect -3360 7208 -3185 7444
rect -2949 7208 -2862 7444
rect -2626 7208 -2539 7444
rect -2303 7208 -2216 7444
rect -1980 7208 -1893 7444
rect -1657 7208 -1570 7444
rect -1334 7208 -1247 7444
rect -1011 7208 -924 7444
rect -688 7208 -601 7444
rect -365 7208 -278 7444
rect -42 7208 45 7444
rect 281 7208 368 7444
rect 604 7208 691 7444
rect 927 7208 1014 7444
rect 1250 7208 1337 7444
rect 1573 7208 1660 7444
rect 1896 7208 1983 7444
rect 2219 7208 2306 7444
rect 2542 7208 2629 7444
rect 2865 7208 2952 7444
rect 3188 7208 3275 7444
rect 3511 7208 3598 7444
rect 3834 7208 3921 7444
rect 4157 7208 4244 7444
rect 4480 7208 4567 7444
rect 4803 7208 4890 7444
rect 5126 7208 5213 7444
rect 5449 7208 5536 7444
rect 5772 7208 5859 7444
rect 6095 7208 6182 7444
rect 6418 7208 6505 7444
rect 6741 7208 6828 7444
rect 7064 7208 7150 7444
rect 7386 7208 7472 7444
rect 7708 7208 7794 7444
rect 8030 7208 8116 7444
rect 8352 7208 8438 7444
rect 8674 7208 8760 7444
rect 8996 7208 9082 7444
rect 9318 7208 9404 7444
rect 9640 7208 9726 7444
rect 9962 7208 10048 7444
rect 10284 7208 10370 7444
rect 10606 7208 10692 7444
rect 10928 7208 11014 7444
rect 11250 7208 11336 7444
rect 11572 7208 11658 7444
rect 11894 7208 11980 7444
rect 12216 7208 12302 7444
rect 12538 7208 12624 7444
rect 12860 7208 12946 7444
rect 13182 7208 13268 7444
rect 13504 7208 13590 7444
rect 13826 7208 13912 7444
rect 14148 7208 14234 7444
rect 14470 7208 14556 7444
rect 14792 7208 14878 7444
rect 15114 7208 15200 7444
rect 15436 7208 15522 7444
rect 15758 7208 15844 7444
rect 16080 7208 16166 7444
rect 16402 7208 16488 7444
rect 16724 7208 16810 7444
rect 17046 7208 17132 7444
rect 17368 7208 17454 7444
rect 17690 7208 17776 7444
rect 18012 7208 18098 7444
rect 18334 7208 18420 7444
rect 18656 7208 18742 7444
rect 18978 7208 19064 7444
rect 19300 7208 19386 7444
rect 19622 7208 19708 7444
rect 19944 7208 20030 7444
rect 20266 7208 20352 7444
rect 20588 7208 20674 7444
rect 20910 7208 20996 7444
rect 21232 7208 21318 7444
rect 21554 7208 21640 7444
rect 21876 7208 21962 7444
rect 22198 7208 22284 7444
rect 22520 7208 22606 7444
rect 22842 7208 22928 7444
rect 23164 7208 23250 7444
rect 23486 7208 23572 7444
rect 23808 7208 23894 7444
rect 24130 7208 24216 7444
rect 24452 7208 24640 7444
rect -3360 7078 24640 7208
rect -3360 6842 -3185 7078
rect -2949 6842 -2862 7078
rect -2626 6842 -2539 7078
rect -2303 6842 -2216 7078
rect -1980 6842 -1893 7078
rect -1657 6842 -1570 7078
rect -1334 6842 -1247 7078
rect -1011 6842 -924 7078
rect -688 6842 -601 7078
rect -365 6842 -278 7078
rect -42 6842 45 7078
rect 281 6842 368 7078
rect 604 6842 691 7078
rect 927 6842 1014 7078
rect 1250 6842 1337 7078
rect 1573 6842 1660 7078
rect 1896 6842 1983 7078
rect 2219 6842 2306 7078
rect 2542 6842 2629 7078
rect 2865 6842 2952 7078
rect 3188 6842 3275 7078
rect 3511 6842 3598 7078
rect 3834 6842 3921 7078
rect 4157 6842 4244 7078
rect 4480 6842 4567 7078
rect 4803 6842 4890 7078
rect 5126 6842 5213 7078
rect 5449 6842 5536 7078
rect 5772 6842 5859 7078
rect 6095 6842 6182 7078
rect 6418 6842 6505 7078
rect 6741 6842 6828 7078
rect 7064 6842 7150 7078
rect 7386 6842 7472 7078
rect 7708 6842 7794 7078
rect 8030 6842 8116 7078
rect 8352 6842 8438 7078
rect 8674 6842 8760 7078
rect 8996 6842 9082 7078
rect 9318 6842 9404 7078
rect 9640 6842 9726 7078
rect 9962 6842 10048 7078
rect 10284 6842 10370 7078
rect 10606 6842 10692 7078
rect 10928 6842 11014 7078
rect 11250 6842 11336 7078
rect 11572 6842 11658 7078
rect 11894 6842 11980 7078
rect 12216 6842 12302 7078
rect 12538 6842 12624 7078
rect 12860 6842 12946 7078
rect 13182 6842 13268 7078
rect 13504 6842 13590 7078
rect 13826 6842 13912 7078
rect 14148 6842 14234 7078
rect 14470 6842 14556 7078
rect 14792 6842 14878 7078
rect 15114 6842 15200 7078
rect 15436 6842 15522 7078
rect 15758 6842 15844 7078
rect 16080 6842 16166 7078
rect 16402 6842 16488 7078
rect 16724 6842 16810 7078
rect 17046 6842 17132 7078
rect 17368 6842 17454 7078
rect 17690 6842 17776 7078
rect 18012 6842 18098 7078
rect 18334 6842 18420 7078
rect 18656 6842 18742 7078
rect 18978 6842 19064 7078
rect 19300 6842 19386 7078
rect 19622 6842 19708 7078
rect 19944 6842 20030 7078
rect 20266 6842 20352 7078
rect 20588 6842 20674 7078
rect 20910 6842 20996 7078
rect 21232 6842 21318 7078
rect 21554 6842 21640 7078
rect 21876 6842 21962 7078
rect 22198 6842 22284 7078
rect 22520 6842 22606 7078
rect 22842 6842 22928 7078
rect 23164 6842 23250 7078
rect 23486 6842 23572 7078
rect 23808 6842 23894 7078
rect 24130 6842 24216 7078
rect 24452 6842 24640 7078
rect -3360 6798 -2720 6842
rect 24000 6798 24640 6842
rect -3360 6474 -2720 6518
rect 24000 6474 24640 6518
rect -3360 6238 -3185 6474
rect -2949 6238 -2862 6474
rect -2626 6238 -2539 6474
rect -2303 6238 -2216 6474
rect -1980 6238 -1893 6474
rect -1657 6238 -1570 6474
rect -1334 6238 -1247 6474
rect -1011 6238 -924 6474
rect -688 6238 -601 6474
rect -365 6238 -278 6474
rect -42 6238 45 6474
rect 281 6238 368 6474
rect 604 6238 691 6474
rect 927 6238 1014 6474
rect 1250 6238 1337 6474
rect 1573 6238 1660 6474
rect 1896 6238 1983 6474
rect 2219 6238 2306 6474
rect 2542 6238 2629 6474
rect 2865 6238 2952 6474
rect 3188 6238 3275 6474
rect 3511 6238 3598 6474
rect 3834 6238 3921 6474
rect 4157 6238 4244 6474
rect 4480 6238 4567 6474
rect 4803 6238 4890 6474
rect 5126 6238 5213 6474
rect 5449 6238 5536 6474
rect 5772 6238 5859 6474
rect 6095 6238 6182 6474
rect 6418 6238 6505 6474
rect 6741 6238 6828 6474
rect 7064 6238 7150 6474
rect 7386 6238 7472 6474
rect 7708 6238 7794 6474
rect 8030 6238 8116 6474
rect 8352 6238 8438 6474
rect 8674 6238 8760 6474
rect 8996 6238 9082 6474
rect 9318 6238 9404 6474
rect 9640 6238 9726 6474
rect 9962 6238 10048 6474
rect 10284 6238 10370 6474
rect 10606 6238 10692 6474
rect 10928 6238 11014 6474
rect 11250 6238 11336 6474
rect 11572 6238 11658 6474
rect 11894 6238 11980 6474
rect 12216 6238 12302 6474
rect 12538 6238 12624 6474
rect 12860 6238 12946 6474
rect 13182 6238 13268 6474
rect 13504 6238 13590 6474
rect 13826 6238 13912 6474
rect 14148 6238 14234 6474
rect 14470 6238 14556 6474
rect 14792 6238 14878 6474
rect 15114 6238 15200 6474
rect 15436 6238 15522 6474
rect 15758 6238 15844 6474
rect 16080 6238 16166 6474
rect 16402 6238 16488 6474
rect 16724 6238 16810 6474
rect 17046 6238 17132 6474
rect 17368 6238 17454 6474
rect 17690 6238 17776 6474
rect 18012 6238 18098 6474
rect 18334 6238 18420 6474
rect 18656 6238 18742 6474
rect 18978 6238 19064 6474
rect 19300 6238 19386 6474
rect 19622 6238 19708 6474
rect 19944 6238 20030 6474
rect 20266 6238 20352 6474
rect 20588 6238 20674 6474
rect 20910 6238 20996 6474
rect 21232 6238 21318 6474
rect 21554 6238 21640 6474
rect 21876 6238 21962 6474
rect 22198 6238 22284 6474
rect 22520 6238 22606 6474
rect 22842 6238 22928 6474
rect 23164 6238 23250 6474
rect 23486 6238 23572 6474
rect 23808 6238 23894 6474
rect 24130 6238 24216 6474
rect 24452 6238 24640 6474
rect -3360 6108 24640 6238
rect -3360 5872 -3185 6108
rect -2949 5872 -2862 6108
rect -2626 5872 -2539 6108
rect -2303 5872 -2216 6108
rect -1980 5872 -1893 6108
rect -1657 5872 -1570 6108
rect -1334 5872 -1247 6108
rect -1011 5872 -924 6108
rect -688 5872 -601 6108
rect -365 5872 -278 6108
rect -42 5872 45 6108
rect 281 5872 368 6108
rect 604 5872 691 6108
rect 927 5872 1014 6108
rect 1250 5872 1337 6108
rect 1573 5872 1660 6108
rect 1896 5872 1983 6108
rect 2219 5872 2306 6108
rect 2542 5872 2629 6108
rect 2865 5872 2952 6108
rect 3188 5872 3275 6108
rect 3511 5872 3598 6108
rect 3834 5872 3921 6108
rect 4157 5872 4244 6108
rect 4480 5872 4567 6108
rect 4803 5872 4890 6108
rect 5126 5872 5213 6108
rect 5449 5872 5536 6108
rect 5772 5872 5859 6108
rect 6095 5872 6182 6108
rect 6418 5872 6505 6108
rect 6741 5872 6828 6108
rect 7064 5872 7150 6108
rect 7386 5872 7472 6108
rect 7708 5872 7794 6108
rect 8030 5872 8116 6108
rect 8352 5872 8438 6108
rect 8674 5872 8760 6108
rect 8996 5872 9082 6108
rect 9318 5872 9404 6108
rect 9640 5872 9726 6108
rect 9962 5872 10048 6108
rect 10284 5872 10370 6108
rect 10606 5872 10692 6108
rect 10928 5872 11014 6108
rect 11250 5872 11336 6108
rect 11572 5872 11658 6108
rect 11894 5872 11980 6108
rect 12216 5872 12302 6108
rect 12538 5872 12624 6108
rect 12860 5872 12946 6108
rect 13182 5872 13268 6108
rect 13504 5872 13590 6108
rect 13826 5872 13912 6108
rect 14148 5872 14234 6108
rect 14470 5872 14556 6108
rect 14792 5872 14878 6108
rect 15114 5872 15200 6108
rect 15436 5872 15522 6108
rect 15758 5872 15844 6108
rect 16080 5872 16166 6108
rect 16402 5872 16488 6108
rect 16724 5872 16810 6108
rect 17046 5872 17132 6108
rect 17368 5872 17454 6108
rect 17690 5872 17776 6108
rect 18012 5872 18098 6108
rect 18334 5872 18420 6108
rect 18656 5872 18742 6108
rect 18978 5872 19064 6108
rect 19300 5872 19386 6108
rect 19622 5872 19708 6108
rect 19944 5872 20030 6108
rect 20266 5872 20352 6108
rect 20588 5872 20674 6108
rect 20910 5872 20996 6108
rect 21232 5872 21318 6108
rect 21554 5872 21640 6108
rect 21876 5872 21962 6108
rect 22198 5872 22284 6108
rect 22520 5872 22606 6108
rect 22842 5872 22928 6108
rect 23164 5872 23250 6108
rect 23486 5872 23572 6108
rect 23808 5872 23894 6108
rect 24130 5872 24216 6108
rect 24452 5872 24640 6108
rect -3360 5828 -2720 5872
rect 24000 5828 24640 5872
rect -3360 5504 -2720 5548
rect 24000 5504 24640 5548
rect -3360 5268 -3185 5504
rect -2949 5268 -2862 5504
rect -2626 5268 -2539 5504
rect -2303 5268 -2216 5504
rect -1980 5268 -1893 5504
rect -1657 5268 -1570 5504
rect -1334 5268 -1247 5504
rect -1011 5268 -924 5504
rect -688 5268 -601 5504
rect -365 5268 -278 5504
rect -42 5268 45 5504
rect 281 5268 368 5504
rect 604 5268 691 5504
rect 927 5268 1014 5504
rect 1250 5268 1337 5504
rect 1573 5268 1660 5504
rect 1896 5268 1983 5504
rect 2219 5268 2306 5504
rect 2542 5268 2629 5504
rect 2865 5268 2952 5504
rect 3188 5268 3275 5504
rect 3511 5268 3598 5504
rect 3834 5268 3921 5504
rect 4157 5268 4244 5504
rect 4480 5268 4567 5504
rect 4803 5268 4890 5504
rect 5126 5268 5213 5504
rect 5449 5268 5536 5504
rect 5772 5268 5859 5504
rect 6095 5268 6182 5504
rect 6418 5268 6505 5504
rect 6741 5268 6828 5504
rect 7064 5268 7150 5504
rect 7386 5268 7472 5504
rect 7708 5268 7794 5504
rect 8030 5268 8116 5504
rect 8352 5268 8438 5504
rect 8674 5268 8760 5504
rect 8996 5268 9082 5504
rect 9318 5268 9404 5504
rect 9640 5268 9726 5504
rect 9962 5268 10048 5504
rect 10284 5268 10370 5504
rect 10606 5268 10692 5504
rect 10928 5268 11014 5504
rect 11250 5268 11336 5504
rect 11572 5268 11658 5504
rect 11894 5268 11980 5504
rect 12216 5268 12302 5504
rect 12538 5268 12624 5504
rect 12860 5268 12946 5504
rect 13182 5268 13268 5504
rect 13504 5268 13590 5504
rect 13826 5268 13912 5504
rect 14148 5268 14234 5504
rect 14470 5268 14556 5504
rect 14792 5268 14878 5504
rect 15114 5268 15200 5504
rect 15436 5268 15522 5504
rect 15758 5268 15844 5504
rect 16080 5268 16166 5504
rect 16402 5268 16488 5504
rect 16724 5268 16810 5504
rect 17046 5268 17132 5504
rect 17368 5268 17454 5504
rect 17690 5268 17776 5504
rect 18012 5268 18098 5504
rect 18334 5268 18420 5504
rect 18656 5268 18742 5504
rect 18978 5268 19064 5504
rect 19300 5268 19386 5504
rect 19622 5268 19708 5504
rect 19944 5268 20030 5504
rect 20266 5268 20352 5504
rect 20588 5268 20674 5504
rect 20910 5268 20996 5504
rect 21232 5268 21318 5504
rect 21554 5268 21640 5504
rect 21876 5268 21962 5504
rect 22198 5268 22284 5504
rect 22520 5268 22606 5504
rect 22842 5268 22928 5504
rect 23164 5268 23250 5504
rect 23486 5268 23572 5504
rect 23808 5268 23894 5504
rect 24130 5268 24216 5504
rect 24452 5268 24640 5504
rect -3360 4898 24640 5268
rect -3360 4662 -3185 4898
rect -2949 4662 -2862 4898
rect -2626 4662 -2539 4898
rect -2303 4662 -2216 4898
rect -1980 4662 -1893 4898
rect -1657 4662 -1570 4898
rect -1334 4662 -1247 4898
rect -1011 4662 -924 4898
rect -688 4662 -601 4898
rect -365 4662 -278 4898
rect -42 4662 45 4898
rect 281 4662 368 4898
rect 604 4662 691 4898
rect 927 4662 1014 4898
rect 1250 4662 1337 4898
rect 1573 4662 1660 4898
rect 1896 4662 1983 4898
rect 2219 4662 2306 4898
rect 2542 4662 2629 4898
rect 2865 4662 2952 4898
rect 3188 4662 3275 4898
rect 3511 4662 3598 4898
rect 3834 4662 3921 4898
rect 4157 4662 4244 4898
rect 4480 4662 4567 4898
rect 4803 4662 4890 4898
rect 5126 4662 5213 4898
rect 5449 4662 5536 4898
rect 5772 4662 5859 4898
rect 6095 4662 6182 4898
rect 6418 4662 6505 4898
rect 6741 4662 6828 4898
rect 7064 4662 7150 4898
rect 7386 4662 7472 4898
rect 7708 4662 7794 4898
rect 8030 4662 8116 4898
rect 8352 4662 8438 4898
rect 8674 4662 8760 4898
rect 8996 4662 9082 4898
rect 9318 4662 9404 4898
rect 9640 4662 9726 4898
rect 9962 4662 10048 4898
rect 10284 4662 10370 4898
rect 10606 4662 10692 4898
rect 10928 4662 11014 4898
rect 11250 4662 11336 4898
rect 11572 4662 11658 4898
rect 11894 4662 11980 4898
rect 12216 4662 12302 4898
rect 12538 4662 12624 4898
rect 12860 4662 12946 4898
rect 13182 4662 13268 4898
rect 13504 4662 13590 4898
rect 13826 4662 13912 4898
rect 14148 4662 14234 4898
rect 14470 4662 14556 4898
rect 14792 4662 14878 4898
rect 15114 4662 15200 4898
rect 15436 4662 15522 4898
rect 15758 4662 15844 4898
rect 16080 4662 16166 4898
rect 16402 4662 16488 4898
rect 16724 4662 16810 4898
rect 17046 4662 17132 4898
rect 17368 4662 17454 4898
rect 17690 4662 17776 4898
rect 18012 4662 18098 4898
rect 18334 4662 18420 4898
rect 18656 4662 18742 4898
rect 18978 4662 19064 4898
rect 19300 4662 19386 4898
rect 19622 4662 19708 4898
rect 19944 4662 20030 4898
rect 20266 4662 20352 4898
rect 20588 4662 20674 4898
rect 20910 4662 20996 4898
rect 21232 4662 21318 4898
rect 21554 4662 21640 4898
rect 21876 4662 21962 4898
rect 22198 4662 22284 4898
rect 22520 4662 22606 4898
rect 22842 4662 22928 4898
rect 23164 4662 23250 4898
rect 23486 4662 23572 4898
rect 23808 4662 23894 4898
rect 24130 4662 24216 4898
rect 24452 4662 24640 4898
rect -3360 4618 -2720 4662
rect 24000 4618 24640 4662
rect -3360 4294 -2720 4338
rect 24000 4294 24640 4338
rect -3360 4058 -3185 4294
rect -2949 4058 -2862 4294
rect -2626 4058 -2539 4294
rect -2303 4058 -2216 4294
rect -1980 4058 -1893 4294
rect -1657 4058 -1570 4294
rect -1334 4058 -1247 4294
rect -1011 4058 -924 4294
rect -688 4058 -601 4294
rect -365 4058 -278 4294
rect -42 4058 45 4294
rect 281 4058 368 4294
rect 604 4058 691 4294
rect 927 4058 1014 4294
rect 1250 4058 1337 4294
rect 1573 4058 1660 4294
rect 1896 4058 1983 4294
rect 2219 4058 2306 4294
rect 2542 4058 2629 4294
rect 2865 4058 2952 4294
rect 3188 4058 3275 4294
rect 3511 4058 3598 4294
rect 3834 4058 3921 4294
rect 4157 4058 4244 4294
rect 4480 4058 4567 4294
rect 4803 4058 4890 4294
rect 5126 4058 5213 4294
rect 5449 4058 5536 4294
rect 5772 4058 5859 4294
rect 6095 4058 6182 4294
rect 6418 4058 6505 4294
rect 6741 4058 6828 4294
rect 7064 4058 7150 4294
rect 7386 4058 7472 4294
rect 7708 4058 7794 4294
rect 8030 4058 8116 4294
rect 8352 4058 8438 4294
rect 8674 4058 8760 4294
rect 8996 4058 9082 4294
rect 9318 4058 9404 4294
rect 9640 4058 9726 4294
rect 9962 4058 10048 4294
rect 10284 4058 10370 4294
rect 10606 4058 10692 4294
rect 10928 4058 11014 4294
rect 11250 4058 11336 4294
rect 11572 4058 11658 4294
rect 11894 4058 11980 4294
rect 12216 4058 12302 4294
rect 12538 4058 12624 4294
rect 12860 4058 12946 4294
rect 13182 4058 13268 4294
rect 13504 4058 13590 4294
rect 13826 4058 13912 4294
rect 14148 4058 14234 4294
rect 14470 4058 14556 4294
rect 14792 4058 14878 4294
rect 15114 4058 15200 4294
rect 15436 4058 15522 4294
rect 15758 4058 15844 4294
rect 16080 4058 16166 4294
rect 16402 4058 16488 4294
rect 16724 4058 16810 4294
rect 17046 4058 17132 4294
rect 17368 4058 17454 4294
rect 17690 4058 17776 4294
rect 18012 4058 18098 4294
rect 18334 4058 18420 4294
rect 18656 4058 18742 4294
rect 18978 4058 19064 4294
rect 19300 4058 19386 4294
rect 19622 4058 19708 4294
rect 19944 4058 20030 4294
rect 20266 4058 20352 4294
rect 20588 4058 20674 4294
rect 20910 4058 20996 4294
rect 21232 4058 21318 4294
rect 21554 4058 21640 4294
rect 21876 4058 21962 4294
rect 22198 4058 22284 4294
rect 22520 4058 22606 4294
rect 22842 4058 22928 4294
rect 23164 4058 23250 4294
rect 23486 4058 23572 4294
rect 23808 4058 23894 4294
rect 24130 4058 24216 4294
rect 24452 4058 24640 4294
rect -3360 3688 24640 4058
rect -3360 3452 -3185 3688
rect -2949 3452 -2862 3688
rect -2626 3452 -2539 3688
rect -2303 3452 -2216 3688
rect -1980 3452 -1893 3688
rect -1657 3452 -1570 3688
rect -1334 3452 -1247 3688
rect -1011 3452 -924 3688
rect -688 3452 -601 3688
rect -365 3452 -278 3688
rect -42 3452 45 3688
rect 281 3452 368 3688
rect 604 3452 691 3688
rect 927 3452 1014 3688
rect 1250 3452 1337 3688
rect 1573 3452 1660 3688
rect 1896 3452 1983 3688
rect 2219 3452 2306 3688
rect 2542 3452 2629 3688
rect 2865 3452 2952 3688
rect 3188 3452 3275 3688
rect 3511 3452 3598 3688
rect 3834 3452 3921 3688
rect 4157 3452 4244 3688
rect 4480 3452 4567 3688
rect 4803 3452 4890 3688
rect 5126 3452 5213 3688
rect 5449 3452 5536 3688
rect 5772 3452 5859 3688
rect 6095 3452 6182 3688
rect 6418 3452 6505 3688
rect 6741 3452 6828 3688
rect 7064 3452 7150 3688
rect 7386 3452 7472 3688
rect 7708 3452 7794 3688
rect 8030 3452 8116 3688
rect 8352 3452 8438 3688
rect 8674 3452 8760 3688
rect 8996 3452 9082 3688
rect 9318 3452 9404 3688
rect 9640 3452 9726 3688
rect 9962 3452 10048 3688
rect 10284 3452 10370 3688
rect 10606 3452 10692 3688
rect 10928 3452 11014 3688
rect 11250 3452 11336 3688
rect 11572 3452 11658 3688
rect 11894 3452 11980 3688
rect 12216 3452 12302 3688
rect 12538 3452 12624 3688
rect 12860 3452 12946 3688
rect 13182 3452 13268 3688
rect 13504 3452 13590 3688
rect 13826 3452 13912 3688
rect 14148 3452 14234 3688
rect 14470 3452 14556 3688
rect 14792 3452 14878 3688
rect 15114 3452 15200 3688
rect 15436 3452 15522 3688
rect 15758 3452 15844 3688
rect 16080 3452 16166 3688
rect 16402 3452 16488 3688
rect 16724 3452 16810 3688
rect 17046 3452 17132 3688
rect 17368 3452 17454 3688
rect 17690 3452 17776 3688
rect 18012 3452 18098 3688
rect 18334 3452 18420 3688
rect 18656 3452 18742 3688
rect 18978 3452 19064 3688
rect 19300 3452 19386 3688
rect 19622 3452 19708 3688
rect 19944 3452 20030 3688
rect 20266 3452 20352 3688
rect 20588 3452 20674 3688
rect 20910 3452 20996 3688
rect 21232 3452 21318 3688
rect 21554 3452 21640 3688
rect 21876 3452 21962 3688
rect 22198 3452 22284 3688
rect 22520 3452 22606 3688
rect 22842 3452 22928 3688
rect 23164 3452 23250 3688
rect 23486 3452 23572 3688
rect 23808 3452 23894 3688
rect 24130 3452 24216 3688
rect 24452 3452 24640 3688
rect -3360 3408 -2720 3452
rect 24000 3408 24640 3452
rect -3360 3084 -2720 3128
rect 24000 3084 24640 3128
rect -3360 2848 -3185 3084
rect -2949 2848 -2862 3084
rect -2626 2848 -2539 3084
rect -2303 2848 -2216 3084
rect -1980 2848 -1893 3084
rect -1657 2848 -1570 3084
rect -1334 2848 -1247 3084
rect -1011 2848 -924 3084
rect -688 2848 -601 3084
rect -365 2848 -278 3084
rect -42 2848 45 3084
rect 281 2848 368 3084
rect 604 2848 691 3084
rect 927 2848 1014 3084
rect 1250 2848 1337 3084
rect 1573 2848 1660 3084
rect 1896 2848 1983 3084
rect 2219 2848 2306 3084
rect 2542 2848 2629 3084
rect 2865 2848 2952 3084
rect 3188 2848 3275 3084
rect 3511 2848 3598 3084
rect 3834 2848 3921 3084
rect 4157 2848 4244 3084
rect 4480 2848 4567 3084
rect 4803 2848 4890 3084
rect 5126 2848 5213 3084
rect 5449 2848 5536 3084
rect 5772 2848 5859 3084
rect 6095 2848 6182 3084
rect 6418 2848 6505 3084
rect 6741 2848 6828 3084
rect 7064 2848 7150 3084
rect 7386 2848 7472 3084
rect 7708 2848 7794 3084
rect 8030 2848 8116 3084
rect 8352 2848 8438 3084
rect 8674 2848 8760 3084
rect 8996 2848 9082 3084
rect 9318 2848 9404 3084
rect 9640 2848 9726 3084
rect 9962 2848 10048 3084
rect 10284 2848 10370 3084
rect 10606 2848 10692 3084
rect 10928 2848 11014 3084
rect 11250 2848 11336 3084
rect 11572 2848 11658 3084
rect 11894 2848 11980 3084
rect 12216 2848 12302 3084
rect 12538 2848 12624 3084
rect 12860 2848 12946 3084
rect 13182 2848 13268 3084
rect 13504 2848 13590 3084
rect 13826 2848 13912 3084
rect 14148 2848 14234 3084
rect 14470 2848 14556 3084
rect 14792 2848 14878 3084
rect 15114 2848 15200 3084
rect 15436 2848 15522 3084
rect 15758 2848 15844 3084
rect 16080 2848 16166 3084
rect 16402 2848 16488 3084
rect 16724 2848 16810 3084
rect 17046 2848 17132 3084
rect 17368 2848 17454 3084
rect 17690 2848 17776 3084
rect 18012 2848 18098 3084
rect 18334 2848 18420 3084
rect 18656 2848 18742 3084
rect 18978 2848 19064 3084
rect 19300 2848 19386 3084
rect 19622 2848 19708 3084
rect 19944 2848 20030 3084
rect 20266 2848 20352 3084
rect 20588 2848 20674 3084
rect 20910 2848 20996 3084
rect 21232 2848 21318 3084
rect 21554 2848 21640 3084
rect 21876 2848 21962 3084
rect 22198 2848 22284 3084
rect 22520 2848 22606 3084
rect 22842 2848 22928 3084
rect 23164 2848 23250 3084
rect 23486 2848 23572 3084
rect 23808 2848 23894 3084
rect 24130 2848 24216 3084
rect 24452 2848 24640 3084
rect -3360 2718 24640 2848
rect -3360 2482 -3185 2718
rect -2949 2482 -2862 2718
rect -2626 2482 -2539 2718
rect -2303 2482 -2216 2718
rect -1980 2482 -1893 2718
rect -1657 2482 -1570 2718
rect -1334 2482 -1247 2718
rect -1011 2482 -924 2718
rect -688 2482 -601 2718
rect -365 2482 -278 2718
rect -42 2482 45 2718
rect 281 2482 368 2718
rect 604 2482 691 2718
rect 927 2482 1014 2718
rect 1250 2482 1337 2718
rect 1573 2482 1660 2718
rect 1896 2482 1983 2718
rect 2219 2482 2306 2718
rect 2542 2482 2629 2718
rect 2865 2482 2952 2718
rect 3188 2482 3275 2718
rect 3511 2482 3598 2718
rect 3834 2482 3921 2718
rect 4157 2482 4244 2718
rect 4480 2482 4567 2718
rect 4803 2482 4890 2718
rect 5126 2482 5213 2718
rect 5449 2482 5536 2718
rect 5772 2482 5859 2718
rect 6095 2482 6182 2718
rect 6418 2482 6505 2718
rect 6741 2482 6828 2718
rect 7064 2482 7150 2718
rect 7386 2482 7472 2718
rect 7708 2482 7794 2718
rect 8030 2482 8116 2718
rect 8352 2482 8438 2718
rect 8674 2482 8760 2718
rect 8996 2482 9082 2718
rect 9318 2482 9404 2718
rect 9640 2482 9726 2718
rect 9962 2482 10048 2718
rect 10284 2482 10370 2718
rect 10606 2482 10692 2718
rect 10928 2482 11014 2718
rect 11250 2482 11336 2718
rect 11572 2482 11658 2718
rect 11894 2482 11980 2718
rect 12216 2482 12302 2718
rect 12538 2482 12624 2718
rect 12860 2482 12946 2718
rect 13182 2482 13268 2718
rect 13504 2482 13590 2718
rect 13826 2482 13912 2718
rect 14148 2482 14234 2718
rect 14470 2482 14556 2718
rect 14792 2482 14878 2718
rect 15114 2482 15200 2718
rect 15436 2482 15522 2718
rect 15758 2482 15844 2718
rect 16080 2482 16166 2718
rect 16402 2482 16488 2718
rect 16724 2482 16810 2718
rect 17046 2482 17132 2718
rect 17368 2482 17454 2718
rect 17690 2482 17776 2718
rect 18012 2482 18098 2718
rect 18334 2482 18420 2718
rect 18656 2482 18742 2718
rect 18978 2482 19064 2718
rect 19300 2482 19386 2718
rect 19622 2482 19708 2718
rect 19944 2482 20030 2718
rect 20266 2482 20352 2718
rect 20588 2482 20674 2718
rect 20910 2482 20996 2718
rect 21232 2482 21318 2718
rect 21554 2482 21640 2718
rect 21876 2482 21962 2718
rect 22198 2482 22284 2718
rect 22520 2482 22606 2718
rect 22842 2482 22928 2718
rect 23164 2482 23250 2718
rect 23486 2482 23572 2718
rect 23808 2482 23894 2718
rect 24130 2482 24216 2718
rect 24452 2482 24640 2718
rect -3360 2438 -2720 2482
rect 24000 2438 24640 2482
rect -3360 2114 -2720 2158
rect 24000 2114 24640 2158
rect -3360 1878 -3185 2114
rect -2949 1878 -2862 2114
rect -2626 1878 -2539 2114
rect -2303 1878 -2216 2114
rect -1980 1878 -1893 2114
rect -1657 1878 -1570 2114
rect -1334 1878 -1247 2114
rect -1011 1878 -924 2114
rect -688 1878 -601 2114
rect -365 1878 -278 2114
rect -42 1878 45 2114
rect 281 1878 368 2114
rect 604 1878 691 2114
rect 927 1878 1014 2114
rect 1250 1878 1337 2114
rect 1573 1878 1660 2114
rect 1896 1878 1983 2114
rect 2219 1878 2306 2114
rect 2542 1878 2629 2114
rect 2865 1878 2952 2114
rect 3188 1878 3275 2114
rect 3511 1878 3598 2114
rect 3834 1878 3921 2114
rect 4157 1878 4244 2114
rect 4480 1878 4567 2114
rect 4803 1878 4890 2114
rect 5126 1878 5213 2114
rect 5449 1878 5536 2114
rect 5772 1878 5859 2114
rect 6095 1878 6182 2114
rect 6418 1878 6505 2114
rect 6741 1878 6828 2114
rect 7064 1878 7150 2114
rect 7386 1878 7472 2114
rect 7708 1878 7794 2114
rect 8030 1878 8116 2114
rect 8352 1878 8438 2114
rect 8674 1878 8760 2114
rect 8996 1878 9082 2114
rect 9318 1878 9404 2114
rect 9640 1878 9726 2114
rect 9962 1878 10048 2114
rect 10284 1878 10370 2114
rect 10606 1878 10692 2114
rect 10928 1878 11014 2114
rect 11250 1878 11336 2114
rect 11572 1878 11658 2114
rect 11894 1878 11980 2114
rect 12216 1878 12302 2114
rect 12538 1878 12624 2114
rect 12860 1878 12946 2114
rect 13182 1878 13268 2114
rect 13504 1878 13590 2114
rect 13826 1878 13912 2114
rect 14148 1878 14234 2114
rect 14470 1878 14556 2114
rect 14792 1878 14878 2114
rect 15114 1878 15200 2114
rect 15436 1878 15522 2114
rect 15758 1878 15844 2114
rect 16080 1878 16166 2114
rect 16402 1878 16488 2114
rect 16724 1878 16810 2114
rect 17046 1878 17132 2114
rect 17368 1878 17454 2114
rect 17690 1878 17776 2114
rect 18012 1878 18098 2114
rect 18334 1878 18420 2114
rect 18656 1878 18742 2114
rect 18978 1878 19064 2114
rect 19300 1878 19386 2114
rect 19622 1878 19708 2114
rect 19944 1878 20030 2114
rect 20266 1878 20352 2114
rect 20588 1878 20674 2114
rect 20910 1878 20996 2114
rect 21232 1878 21318 2114
rect 21554 1878 21640 2114
rect 21876 1878 21962 2114
rect 22198 1878 22284 2114
rect 22520 1878 22606 2114
rect 22842 1878 22928 2114
rect 23164 1878 23250 2114
rect 23486 1878 23572 2114
rect 23808 1878 23894 2114
rect 24130 1878 24216 2114
rect 24452 1878 24640 2114
rect -3360 1508 24640 1878
rect -3360 1272 -3185 1508
rect -2949 1272 -2862 1508
rect -2626 1272 -2539 1508
rect -2303 1272 -2216 1508
rect -1980 1272 -1893 1508
rect -1657 1272 -1570 1508
rect -1334 1272 -1247 1508
rect -1011 1272 -924 1508
rect -688 1272 -601 1508
rect -365 1272 -278 1508
rect -42 1272 45 1508
rect 281 1272 368 1508
rect 604 1272 691 1508
rect 927 1272 1014 1508
rect 1250 1272 1337 1508
rect 1573 1272 1660 1508
rect 1896 1272 1983 1508
rect 2219 1272 2306 1508
rect 2542 1272 2629 1508
rect 2865 1272 2952 1508
rect 3188 1272 3275 1508
rect 3511 1272 3598 1508
rect 3834 1272 3921 1508
rect 4157 1272 4244 1508
rect 4480 1272 4567 1508
rect 4803 1272 4890 1508
rect 5126 1272 5213 1508
rect 5449 1272 5536 1508
rect 5772 1272 5859 1508
rect 6095 1272 6182 1508
rect 6418 1272 6505 1508
rect 6741 1272 6828 1508
rect 7064 1272 7150 1508
rect 7386 1272 7472 1508
rect 7708 1272 7794 1508
rect 8030 1272 8116 1508
rect 8352 1272 8438 1508
rect 8674 1272 8760 1508
rect 8996 1272 9082 1508
rect 9318 1272 9404 1508
rect 9640 1272 9726 1508
rect 9962 1272 10048 1508
rect 10284 1272 10370 1508
rect 10606 1272 10692 1508
rect 10928 1272 11014 1508
rect 11250 1272 11336 1508
rect 11572 1272 11658 1508
rect 11894 1272 11980 1508
rect 12216 1272 12302 1508
rect 12538 1272 12624 1508
rect 12860 1272 12946 1508
rect 13182 1272 13268 1508
rect 13504 1272 13590 1508
rect 13826 1272 13912 1508
rect 14148 1272 14234 1508
rect 14470 1272 14556 1508
rect 14792 1272 14878 1508
rect 15114 1272 15200 1508
rect 15436 1272 15522 1508
rect 15758 1272 15844 1508
rect 16080 1272 16166 1508
rect 16402 1272 16488 1508
rect 16724 1272 16810 1508
rect 17046 1272 17132 1508
rect 17368 1272 17454 1508
rect 17690 1272 17776 1508
rect 18012 1272 18098 1508
rect 18334 1272 18420 1508
rect 18656 1272 18742 1508
rect 18978 1272 19064 1508
rect 19300 1272 19386 1508
rect 19622 1272 19708 1508
rect 19944 1272 20030 1508
rect 20266 1272 20352 1508
rect 20588 1272 20674 1508
rect 20910 1272 20996 1508
rect 21232 1272 21318 1508
rect 21554 1272 21640 1508
rect 21876 1272 21962 1508
rect 22198 1272 22284 1508
rect 22520 1272 22606 1508
rect 22842 1272 22928 1508
rect 23164 1272 23250 1508
rect 23486 1272 23572 1508
rect 23808 1272 23894 1508
rect 24130 1272 24216 1508
rect 24452 1272 24640 1508
rect -3360 1228 -2720 1272
rect 24000 1228 24640 1272
rect -3360 904 -2720 948
rect 24000 904 24640 948
rect -3360 903 24640 904
rect -3360 667 -3185 903
rect -2949 667 -2862 903
rect -2626 667 -2539 903
rect -2303 667 -2216 903
rect -1980 667 -1893 903
rect -1657 667 -1570 903
rect -1334 667 -1247 903
rect -1011 667 -924 903
rect -688 667 -601 903
rect -365 667 -278 903
rect -42 667 45 903
rect 281 667 368 903
rect 604 667 691 903
rect 927 667 1014 903
rect 1250 667 1337 903
rect 1573 667 1660 903
rect 1896 667 1983 903
rect 2219 667 2306 903
rect 2542 667 2629 903
rect 2865 667 2952 903
rect 3188 667 3275 903
rect 3511 667 3598 903
rect 3834 667 3921 903
rect 4157 667 4244 903
rect 4480 667 4567 903
rect 4803 667 4890 903
rect 5126 667 5213 903
rect 5449 667 5536 903
rect 5772 667 5859 903
rect 6095 667 6182 903
rect 6418 667 6505 903
rect 6741 667 6828 903
rect 7064 667 7150 903
rect 7386 667 7472 903
rect 7708 667 7794 903
rect 8030 667 8116 903
rect 8352 667 8438 903
rect 8674 667 8760 903
rect 8996 667 9082 903
rect 9318 667 9404 903
rect 9640 667 9726 903
rect 9962 667 10048 903
rect 10284 667 10370 903
rect 10606 667 10692 903
rect 10928 667 11014 903
rect 11250 667 11336 903
rect 11572 667 11658 903
rect 11894 667 11980 903
rect 12216 667 12302 903
rect 12538 667 12624 903
rect 12860 667 12946 903
rect 13182 667 13268 903
rect 13504 667 13590 903
rect 13826 667 13912 903
rect 14148 667 14234 903
rect 14470 667 14556 903
rect 14792 667 14878 903
rect 15114 667 15200 903
rect 15436 667 15522 903
rect 15758 667 15844 903
rect 16080 667 16166 903
rect 16402 667 16488 903
rect 16724 667 16810 903
rect 17046 667 17132 903
rect 17368 667 17454 903
rect 17690 667 17776 903
rect 18012 667 18098 903
rect 18334 667 18420 903
rect 18656 667 18742 903
rect 18978 667 19064 903
rect 19300 667 19386 903
rect 19622 667 19708 903
rect 19944 667 20030 903
rect 20266 667 20352 903
rect 20588 667 20674 903
rect 20910 667 20996 903
rect 21232 667 21318 903
rect 21554 667 21640 903
rect 21876 667 21962 903
rect 22198 667 22284 903
rect 22520 667 22606 903
rect 22842 667 22928 903
rect 23164 667 23250 903
rect 23486 667 23572 903
rect 23808 667 23894 903
rect 24130 667 24216 903
rect 24452 667 24640 903
rect -3360 521 24640 667
rect -3360 285 -3185 521
rect -2949 285 -2862 521
rect -2626 285 -2539 521
rect -2303 285 -2216 521
rect -1980 285 -1893 521
rect -1657 285 -1570 521
rect -1334 285 -1247 521
rect -1011 285 -924 521
rect -688 285 -601 521
rect -365 285 -278 521
rect -42 285 45 521
rect 281 285 368 521
rect 604 285 691 521
rect 927 285 1014 521
rect 1250 285 1337 521
rect 1573 285 1660 521
rect 1896 285 1983 521
rect 2219 285 2306 521
rect 2542 285 2629 521
rect 2865 285 2952 521
rect 3188 285 3275 521
rect 3511 285 3598 521
rect 3834 285 3921 521
rect 4157 285 4244 521
rect 4480 285 4567 521
rect 4803 285 4890 521
rect 5126 285 5213 521
rect 5449 285 5536 521
rect 5772 285 5859 521
rect 6095 285 6182 521
rect 6418 285 6505 521
rect 6741 285 6828 521
rect 7064 285 7150 521
rect 7386 285 7472 521
rect 7708 285 7794 521
rect 8030 285 8116 521
rect 8352 285 8438 521
rect 8674 285 8760 521
rect 8996 285 9082 521
rect 9318 285 9404 521
rect 9640 285 9726 521
rect 9962 285 10048 521
rect 10284 285 10370 521
rect 10606 285 10692 521
rect 10928 285 11014 521
rect 11250 285 11336 521
rect 11572 285 11658 521
rect 11894 285 11980 521
rect 12216 285 12302 521
rect 12538 285 12624 521
rect 12860 285 12946 521
rect 13182 285 13268 521
rect 13504 285 13590 521
rect 13826 285 13912 521
rect 14148 285 14234 521
rect 14470 285 14556 521
rect 14792 285 14878 521
rect 15114 285 15200 521
rect 15436 285 15522 521
rect 15758 285 15844 521
rect 16080 285 16166 521
rect 16402 285 16488 521
rect 16724 285 16810 521
rect 17046 285 17132 521
rect 17368 285 17454 521
rect 17690 285 17776 521
rect 18012 285 18098 521
rect 18334 285 18420 521
rect 18656 285 18742 521
rect 18978 285 19064 521
rect 19300 285 19386 521
rect 19622 285 19708 521
rect 19944 285 20030 521
rect 20266 285 20352 521
rect 20588 285 20674 521
rect 20910 285 20996 521
rect 21232 285 21318 521
rect 21554 285 21640 521
rect 21876 285 21962 521
rect 22198 285 22284 521
rect 22520 285 22606 521
rect 22842 285 22928 521
rect 23164 285 23250 521
rect 23486 285 23572 521
rect 23808 285 23894 521
rect 24130 285 24216 521
rect 24452 285 24640 521
rect -3360 139 24640 285
rect -3360 -97 -3185 139
rect -2949 -97 -2862 139
rect -2626 -97 -2539 139
rect -2303 -97 -2216 139
rect -1980 -97 -1893 139
rect -1657 -97 -1570 139
rect -1334 -97 -1247 139
rect -1011 -97 -924 139
rect -688 -97 -601 139
rect -365 -97 -278 139
rect -42 -97 45 139
rect 281 -97 368 139
rect 604 -97 691 139
rect 927 -97 1014 139
rect 1250 -97 1337 139
rect 1573 -97 1660 139
rect 1896 -97 1983 139
rect 2219 -97 2306 139
rect 2542 -97 2629 139
rect 2865 -97 2952 139
rect 3188 -97 3275 139
rect 3511 -97 3598 139
rect 3834 -97 3921 139
rect 4157 -97 4244 139
rect 4480 -97 4567 139
rect 4803 -97 4890 139
rect 5126 -97 5213 139
rect 5449 -97 5536 139
rect 5772 -97 5859 139
rect 6095 -97 6182 139
rect 6418 -97 6505 139
rect 6741 -97 6828 139
rect 7064 -97 7150 139
rect 7386 -97 7472 139
rect 7708 -97 7794 139
rect 8030 -97 8116 139
rect 8352 -97 8438 139
rect 8674 -97 8760 139
rect 8996 -97 9082 139
rect 9318 -97 9404 139
rect 9640 -97 9726 139
rect 9962 -97 10048 139
rect 10284 -97 10370 139
rect 10606 -97 10692 139
rect 10928 -97 11014 139
rect 11250 -97 11336 139
rect 11572 -97 11658 139
rect 11894 -97 11980 139
rect 12216 -97 12302 139
rect 12538 -97 12624 139
rect 12860 -97 12946 139
rect 13182 -97 13268 139
rect 13504 -97 13590 139
rect 13826 -97 13912 139
rect 14148 -97 14234 139
rect 14470 -97 14556 139
rect 14792 -97 14878 139
rect 15114 -97 15200 139
rect 15436 -97 15522 139
rect 15758 -97 15844 139
rect 16080 -97 16166 139
rect 16402 -97 16488 139
rect 16724 -97 16810 139
rect 17046 -97 17132 139
rect 17368 -97 17454 139
rect 17690 -97 17776 139
rect 18012 -97 18098 139
rect 18334 -97 18420 139
rect 18656 -97 18742 139
rect 18978 -97 19064 139
rect 19300 -97 19386 139
rect 19622 -97 19708 139
rect 19944 -97 20030 139
rect 20266 -97 20352 139
rect 20588 -97 20674 139
rect 20910 -97 20996 139
rect 21232 -97 21318 139
rect 21554 -97 21640 139
rect 21876 -97 21962 139
rect 22198 -97 22284 139
rect 22520 -97 22606 139
rect 22842 -97 22928 139
rect 23164 -97 23250 139
rect 23486 -97 23572 139
rect 23808 -97 23894 139
rect 24130 -97 24216 139
rect 24452 -97 24640 139
rect -3360 -98 24640 -97
rect -3360 -142 -2720 -98
rect 24000 -142 24640 -98
<< via4 >>
rect -3087 39180 -2851 39416
rect -2765 39180 -2529 39416
rect -2443 39180 -2207 39416
rect -2121 39180 -1885 39416
rect -1799 39180 -1563 39416
rect -1477 39180 -1241 39416
rect -1155 39180 -919 39416
rect -833 39180 -597 39416
rect -511 39180 -275 39416
rect -189 39180 47 39416
rect 133 39180 369 39416
rect 455 39180 691 39416
rect 777 39180 1013 39416
rect 1099 39180 1335 39416
rect 1421 39180 1657 39416
rect 1743 39180 1979 39416
rect 2065 39180 2301 39416
rect 2387 39180 2623 39416
rect 2709 39180 2945 39416
rect 3031 39180 3267 39416
rect 3353 39180 3589 39416
rect 3675 39180 3911 39416
rect 3997 39180 4233 39416
rect 4318 39180 4554 39416
rect 4639 39180 4875 39416
rect 4960 39180 5196 39416
rect 5281 39180 5517 39416
rect 5602 39180 5838 39416
rect 5923 39180 6159 39416
rect 6244 39180 6480 39416
rect 6565 39180 6801 39416
rect 6886 39180 7122 39416
rect 7207 39180 7443 39416
rect 7528 39180 7764 39416
rect 7849 39180 8085 39416
rect 8170 39180 8406 39416
rect 8491 39180 8727 39416
rect 8812 39180 9048 39416
rect 9133 39180 9369 39416
rect 9454 39180 9690 39416
rect 9775 39180 10011 39416
rect 10096 39180 10332 39416
rect 10417 39180 10653 39416
rect 10738 39180 10974 39416
rect 11059 39180 11295 39416
rect 11380 39180 11616 39416
rect 11701 39180 11937 39416
rect 12022 39180 12258 39416
rect 12343 39180 12579 39416
rect 12664 39180 12900 39416
rect 12985 39180 13221 39416
rect 13306 39180 13542 39416
rect 13627 39180 13863 39416
rect 13948 39180 14184 39416
rect 14269 39180 14505 39416
rect 14590 39180 14826 39416
rect 14911 39180 15147 39416
rect 15232 39180 15468 39416
rect 15553 39180 15789 39416
rect 15874 39180 16110 39416
rect 16195 39180 16431 39416
rect 16516 39180 16752 39416
rect 16837 39180 17073 39416
rect 17158 39180 17394 39416
rect 17479 39180 17715 39416
rect 17800 39180 18036 39416
rect 18121 39180 18357 39416
rect 18442 39180 18678 39416
rect 18763 39180 18999 39416
rect 19084 39180 19320 39416
rect 19405 39180 19641 39416
rect 19726 39180 19962 39416
rect 20047 39180 20283 39416
rect 20368 39180 20604 39416
rect 20689 39180 20925 39416
rect 21010 39180 21246 39416
rect 21331 39180 21567 39416
rect 21652 39180 21888 39416
rect 21973 39180 22209 39416
rect 22294 39180 22530 39416
rect 22615 39180 22851 39416
rect 22936 39180 23172 39416
rect 23257 39180 23493 39416
rect 23578 39180 23814 39416
rect 23899 39180 24135 39416
rect 24220 39180 24456 39416
rect -3087 38856 -2851 39092
rect -2765 38856 -2529 39092
rect -2443 38856 -2207 39092
rect -2121 38856 -1885 39092
rect -1799 38856 -1563 39092
rect -1477 38856 -1241 39092
rect -1155 38856 -919 39092
rect -833 38856 -597 39092
rect -511 38856 -275 39092
rect -189 38856 47 39092
rect 133 38856 369 39092
rect 455 38856 691 39092
rect 777 38856 1013 39092
rect 1099 38856 1335 39092
rect 1421 38856 1657 39092
rect 1743 38856 1979 39092
rect 2065 38856 2301 39092
rect 2387 38856 2623 39092
rect 2709 38856 2945 39092
rect 3031 38856 3267 39092
rect 3353 38856 3589 39092
rect 3675 38856 3911 39092
rect 3997 38856 4233 39092
rect 4318 38856 4554 39092
rect 4639 38856 4875 39092
rect 4960 38856 5196 39092
rect 5281 38856 5517 39092
rect 5602 38856 5838 39092
rect 5923 38856 6159 39092
rect 6244 38856 6480 39092
rect 6565 38856 6801 39092
rect 6886 38856 7122 39092
rect 7207 38856 7443 39092
rect 7528 38856 7764 39092
rect 7849 38856 8085 39092
rect 8170 38856 8406 39092
rect 8491 38856 8727 39092
rect 8812 38856 9048 39092
rect 9133 38856 9369 39092
rect 9454 38856 9690 39092
rect 9775 38856 10011 39092
rect 10096 38856 10332 39092
rect 10417 38856 10653 39092
rect 10738 38856 10974 39092
rect 11059 38856 11295 39092
rect 11380 38856 11616 39092
rect 11701 38856 11937 39092
rect 12022 38856 12258 39092
rect 12343 38856 12579 39092
rect 12664 38856 12900 39092
rect 12985 38856 13221 39092
rect 13306 38856 13542 39092
rect 13627 38856 13863 39092
rect 13948 38856 14184 39092
rect 14269 38856 14505 39092
rect 14590 38856 14826 39092
rect 14911 38856 15147 39092
rect 15232 38856 15468 39092
rect 15553 38856 15789 39092
rect 15874 38856 16110 39092
rect 16195 38856 16431 39092
rect 16516 38856 16752 39092
rect 16837 38856 17073 39092
rect 17158 38856 17394 39092
rect 17479 38856 17715 39092
rect 17800 38856 18036 39092
rect 18121 38856 18357 39092
rect 18442 38856 18678 39092
rect 18763 38856 18999 39092
rect 19084 38856 19320 39092
rect 19405 38856 19641 39092
rect 19726 38856 19962 39092
rect 20047 38856 20283 39092
rect 20368 38856 20604 39092
rect 20689 38856 20925 39092
rect 21010 38856 21246 39092
rect 21331 38856 21567 39092
rect 21652 38856 21888 39092
rect 21973 38856 22209 39092
rect 22294 38856 22530 39092
rect 22615 38856 22851 39092
rect 22936 38856 23172 39092
rect 23257 38856 23493 39092
rect 23578 38856 23814 39092
rect 23899 38856 24135 39092
rect 24220 38856 24456 39092
rect -3087 38532 -2851 38768
rect -2765 38532 -2529 38768
rect -2443 38532 -2207 38768
rect -2121 38532 -1885 38768
rect -1799 38532 -1563 38768
rect -1477 38532 -1241 38768
rect -1155 38532 -919 38768
rect -833 38532 -597 38768
rect -511 38532 -275 38768
rect -189 38532 47 38768
rect 133 38532 369 38768
rect 455 38532 691 38768
rect 777 38532 1013 38768
rect 1099 38532 1335 38768
rect 1421 38532 1657 38768
rect 1743 38532 1979 38768
rect 2065 38532 2301 38768
rect 2387 38532 2623 38768
rect 2709 38532 2945 38768
rect 3031 38532 3267 38768
rect 3353 38532 3589 38768
rect 3675 38532 3911 38768
rect 3997 38532 4233 38768
rect 4318 38532 4554 38768
rect 4639 38532 4875 38768
rect 4960 38532 5196 38768
rect 5281 38532 5517 38768
rect 5602 38532 5838 38768
rect 5923 38532 6159 38768
rect 6244 38532 6480 38768
rect 6565 38532 6801 38768
rect 6886 38532 7122 38768
rect 7207 38532 7443 38768
rect 7528 38532 7764 38768
rect 7849 38532 8085 38768
rect 8170 38532 8406 38768
rect 8491 38532 8727 38768
rect 8812 38532 9048 38768
rect 9133 38532 9369 38768
rect 9454 38532 9690 38768
rect 9775 38532 10011 38768
rect 10096 38532 10332 38768
rect 10417 38532 10653 38768
rect 10738 38532 10974 38768
rect 11059 38532 11295 38768
rect 11380 38532 11616 38768
rect 11701 38532 11937 38768
rect 12022 38532 12258 38768
rect 12343 38532 12579 38768
rect 12664 38532 12900 38768
rect 12985 38532 13221 38768
rect 13306 38532 13542 38768
rect 13627 38532 13863 38768
rect 13948 38532 14184 38768
rect 14269 38532 14505 38768
rect 14590 38532 14826 38768
rect 14911 38532 15147 38768
rect 15232 38532 15468 38768
rect 15553 38532 15789 38768
rect 15874 38532 16110 38768
rect 16195 38532 16431 38768
rect 16516 38532 16752 38768
rect 16837 38532 17073 38768
rect 17158 38532 17394 38768
rect 17479 38532 17715 38768
rect 17800 38532 18036 38768
rect 18121 38532 18357 38768
rect 18442 38532 18678 38768
rect 18763 38532 18999 38768
rect 19084 38532 19320 38768
rect 19405 38532 19641 38768
rect 19726 38532 19962 38768
rect 20047 38532 20283 38768
rect 20368 38532 20604 38768
rect 20689 38532 20925 38768
rect 21010 38532 21246 38768
rect 21331 38532 21567 38768
rect 21652 38532 21888 38768
rect 21973 38532 22209 38768
rect 22294 38532 22530 38768
rect 22615 38532 22851 38768
rect 22936 38532 23172 38768
rect 23257 38532 23493 38768
rect 23578 38532 23814 38768
rect 23899 38532 24135 38768
rect 24220 38532 24456 38768
rect -3087 38208 -2851 38444
rect -2765 38208 -2529 38444
rect -2443 38208 -2207 38444
rect -2121 38208 -1885 38444
rect -1799 38208 -1563 38444
rect -1477 38208 -1241 38444
rect -1155 38208 -919 38444
rect -833 38208 -597 38444
rect -511 38208 -275 38444
rect -189 38208 47 38444
rect 133 38208 369 38444
rect 455 38208 691 38444
rect 777 38208 1013 38444
rect 1099 38208 1335 38444
rect 1421 38208 1657 38444
rect 1743 38208 1979 38444
rect 2065 38208 2301 38444
rect 2387 38208 2623 38444
rect 2709 38208 2945 38444
rect 3031 38208 3267 38444
rect 3353 38208 3589 38444
rect 3675 38208 3911 38444
rect 3997 38208 4233 38444
rect 4318 38208 4554 38444
rect 4639 38208 4875 38444
rect 4960 38208 5196 38444
rect 5281 38208 5517 38444
rect 5602 38208 5838 38444
rect 5923 38208 6159 38444
rect 6244 38208 6480 38444
rect 6565 38208 6801 38444
rect 6886 38208 7122 38444
rect 7207 38208 7443 38444
rect 7528 38208 7764 38444
rect 7849 38208 8085 38444
rect 8170 38208 8406 38444
rect 8491 38208 8727 38444
rect 8812 38208 9048 38444
rect 9133 38208 9369 38444
rect 9454 38208 9690 38444
rect 9775 38208 10011 38444
rect 10096 38208 10332 38444
rect 10417 38208 10653 38444
rect 10738 38208 10974 38444
rect 11059 38208 11295 38444
rect 11380 38208 11616 38444
rect 11701 38208 11937 38444
rect 12022 38208 12258 38444
rect 12343 38208 12579 38444
rect 12664 38208 12900 38444
rect 12985 38208 13221 38444
rect 13306 38208 13542 38444
rect 13627 38208 13863 38444
rect 13948 38208 14184 38444
rect 14269 38208 14505 38444
rect 14590 38208 14826 38444
rect 14911 38208 15147 38444
rect 15232 38208 15468 38444
rect 15553 38208 15789 38444
rect 15874 38208 16110 38444
rect 16195 38208 16431 38444
rect 16516 38208 16752 38444
rect 16837 38208 17073 38444
rect 17158 38208 17394 38444
rect 17479 38208 17715 38444
rect 17800 38208 18036 38444
rect 18121 38208 18357 38444
rect 18442 38208 18678 38444
rect 18763 38208 18999 38444
rect 19084 38208 19320 38444
rect 19405 38208 19641 38444
rect 19726 38208 19962 38444
rect 20047 38208 20283 38444
rect 20368 38208 20604 38444
rect 20689 38208 20925 38444
rect 21010 38208 21246 38444
rect 21331 38208 21567 38444
rect 21652 38208 21888 38444
rect 21973 38208 22209 38444
rect 22294 38208 22530 38444
rect 22615 38208 22851 38444
rect 22936 38208 23172 38444
rect 23257 38208 23493 38444
rect 23578 38208 23814 38444
rect 23899 38208 24135 38444
rect 24220 38208 24456 38444
rect -3087 37884 -2851 38120
rect -2765 37884 -2529 38120
rect -2443 37884 -2207 38120
rect -2121 37884 -1885 38120
rect -1799 37884 -1563 38120
rect -1477 37884 -1241 38120
rect -1155 37884 -919 38120
rect -833 37884 -597 38120
rect -511 37884 -275 38120
rect -189 37884 47 38120
rect 133 37884 369 38120
rect 455 37884 691 38120
rect 777 37884 1013 38120
rect 1099 37884 1335 38120
rect 1421 37884 1657 38120
rect 1743 37884 1979 38120
rect 2065 37884 2301 38120
rect 2387 37884 2623 38120
rect 2709 37884 2945 38120
rect 3031 37884 3267 38120
rect 3353 37884 3589 38120
rect 3675 37884 3911 38120
rect 3997 37884 4233 38120
rect 4318 37884 4554 38120
rect 4639 37884 4875 38120
rect 4960 37884 5196 38120
rect 5281 37884 5517 38120
rect 5602 37884 5838 38120
rect 5923 37884 6159 38120
rect 6244 37884 6480 38120
rect 6565 37884 6801 38120
rect 6886 37884 7122 38120
rect 7207 37884 7443 38120
rect 7528 37884 7764 38120
rect 7849 37884 8085 38120
rect 8170 37884 8406 38120
rect 8491 37884 8727 38120
rect 8812 37884 9048 38120
rect 9133 37884 9369 38120
rect 9454 37884 9690 38120
rect 9775 37884 10011 38120
rect 10096 37884 10332 38120
rect 10417 37884 10653 38120
rect 10738 37884 10974 38120
rect 11059 37884 11295 38120
rect 11380 37884 11616 38120
rect 11701 37884 11937 38120
rect 12022 37884 12258 38120
rect 12343 37884 12579 38120
rect 12664 37884 12900 38120
rect 12985 37884 13221 38120
rect 13306 37884 13542 38120
rect 13627 37884 13863 38120
rect 13948 37884 14184 38120
rect 14269 37884 14505 38120
rect 14590 37884 14826 38120
rect 14911 37884 15147 38120
rect 15232 37884 15468 38120
rect 15553 37884 15789 38120
rect 15874 37884 16110 38120
rect 16195 37884 16431 38120
rect 16516 37884 16752 38120
rect 16837 37884 17073 38120
rect 17158 37884 17394 38120
rect 17479 37884 17715 38120
rect 17800 37884 18036 38120
rect 18121 37884 18357 38120
rect 18442 37884 18678 38120
rect 18763 37884 18999 38120
rect 19084 37884 19320 38120
rect 19405 37884 19641 38120
rect 19726 37884 19962 38120
rect 20047 37884 20283 38120
rect 20368 37884 20604 38120
rect 20689 37884 20925 38120
rect 21010 37884 21246 38120
rect 21331 37884 21567 38120
rect 21652 37884 21888 38120
rect 21973 37884 22209 38120
rect 22294 37884 22530 38120
rect 22615 37884 22851 38120
rect 22936 37884 23172 38120
rect 23257 37884 23493 38120
rect 23578 37884 23814 38120
rect 23899 37884 24135 38120
rect 24220 37884 24456 38120
rect -3087 37560 -2851 37796
rect -2765 37560 -2529 37796
rect -2443 37560 -2207 37796
rect -2121 37560 -1885 37796
rect -1799 37560 -1563 37796
rect -1477 37560 -1241 37796
rect -1155 37560 -919 37796
rect -833 37560 -597 37796
rect -511 37560 -275 37796
rect -189 37560 47 37796
rect 133 37560 369 37796
rect 455 37560 691 37796
rect 777 37560 1013 37796
rect 1099 37560 1335 37796
rect 1421 37560 1657 37796
rect 1743 37560 1979 37796
rect 2065 37560 2301 37796
rect 2387 37560 2623 37796
rect 2709 37560 2945 37796
rect 3031 37560 3267 37796
rect 3353 37560 3589 37796
rect 3675 37560 3911 37796
rect 3997 37560 4233 37796
rect 4318 37560 4554 37796
rect 4639 37560 4875 37796
rect 4960 37560 5196 37796
rect 5281 37560 5517 37796
rect 5602 37560 5838 37796
rect 5923 37560 6159 37796
rect 6244 37560 6480 37796
rect 6565 37560 6801 37796
rect 6886 37560 7122 37796
rect 7207 37560 7443 37796
rect 7528 37560 7764 37796
rect 7849 37560 8085 37796
rect 8170 37560 8406 37796
rect 8491 37560 8727 37796
rect 8812 37560 9048 37796
rect 9133 37560 9369 37796
rect 9454 37560 9690 37796
rect 9775 37560 10011 37796
rect 10096 37560 10332 37796
rect 10417 37560 10653 37796
rect 10738 37560 10974 37796
rect 11059 37560 11295 37796
rect 11380 37560 11616 37796
rect 11701 37560 11937 37796
rect 12022 37560 12258 37796
rect 12343 37560 12579 37796
rect 12664 37560 12900 37796
rect 12985 37560 13221 37796
rect 13306 37560 13542 37796
rect 13627 37560 13863 37796
rect 13948 37560 14184 37796
rect 14269 37560 14505 37796
rect 14590 37560 14826 37796
rect 14911 37560 15147 37796
rect 15232 37560 15468 37796
rect 15553 37560 15789 37796
rect 15874 37560 16110 37796
rect 16195 37560 16431 37796
rect 16516 37560 16752 37796
rect 16837 37560 17073 37796
rect 17158 37560 17394 37796
rect 17479 37560 17715 37796
rect 17800 37560 18036 37796
rect 18121 37560 18357 37796
rect 18442 37560 18678 37796
rect 18763 37560 18999 37796
rect 19084 37560 19320 37796
rect 19405 37560 19641 37796
rect 19726 37560 19962 37796
rect 20047 37560 20283 37796
rect 20368 37560 20604 37796
rect 20689 37560 20925 37796
rect 21010 37560 21246 37796
rect 21331 37560 21567 37796
rect 21652 37560 21888 37796
rect 21973 37560 22209 37796
rect 22294 37560 22530 37796
rect 22615 37560 22851 37796
rect 22936 37560 23172 37796
rect 23257 37560 23493 37796
rect 23578 37560 23814 37796
rect 23899 37560 24135 37796
rect 24220 37560 24456 37796
rect -3087 37236 -2851 37472
rect -2765 37236 -2529 37472
rect -2443 37236 -2207 37472
rect -2121 37236 -1885 37472
rect -1799 37236 -1563 37472
rect -1477 37236 -1241 37472
rect -1155 37236 -919 37472
rect -833 37236 -597 37472
rect -511 37236 -275 37472
rect -189 37236 47 37472
rect 133 37236 369 37472
rect 455 37236 691 37472
rect 777 37236 1013 37472
rect 1099 37236 1335 37472
rect 1421 37236 1657 37472
rect 1743 37236 1979 37472
rect 2065 37236 2301 37472
rect 2387 37236 2623 37472
rect 2709 37236 2945 37472
rect 3031 37236 3267 37472
rect 3353 37236 3589 37472
rect 3675 37236 3911 37472
rect 3997 37236 4233 37472
rect 4318 37236 4554 37472
rect 4639 37236 4875 37472
rect 4960 37236 5196 37472
rect 5281 37236 5517 37472
rect 5602 37236 5838 37472
rect 5923 37236 6159 37472
rect 6244 37236 6480 37472
rect 6565 37236 6801 37472
rect 6886 37236 7122 37472
rect 7207 37236 7443 37472
rect 7528 37236 7764 37472
rect 7849 37236 8085 37472
rect 8170 37236 8406 37472
rect 8491 37236 8727 37472
rect 8812 37236 9048 37472
rect 9133 37236 9369 37472
rect 9454 37236 9690 37472
rect 9775 37236 10011 37472
rect 10096 37236 10332 37472
rect 10417 37236 10653 37472
rect 10738 37236 10974 37472
rect 11059 37236 11295 37472
rect 11380 37236 11616 37472
rect 11701 37236 11937 37472
rect 12022 37236 12258 37472
rect 12343 37236 12579 37472
rect 12664 37236 12900 37472
rect 12985 37236 13221 37472
rect 13306 37236 13542 37472
rect 13627 37236 13863 37472
rect 13948 37236 14184 37472
rect 14269 37236 14505 37472
rect 14590 37236 14826 37472
rect 14911 37236 15147 37472
rect 15232 37236 15468 37472
rect 15553 37236 15789 37472
rect 15874 37236 16110 37472
rect 16195 37236 16431 37472
rect 16516 37236 16752 37472
rect 16837 37236 17073 37472
rect 17158 37236 17394 37472
rect 17479 37236 17715 37472
rect 17800 37236 18036 37472
rect 18121 37236 18357 37472
rect 18442 37236 18678 37472
rect 18763 37236 18999 37472
rect 19084 37236 19320 37472
rect 19405 37236 19641 37472
rect 19726 37236 19962 37472
rect 20047 37236 20283 37472
rect 20368 37236 20604 37472
rect 20689 37236 20925 37472
rect 21010 37236 21246 37472
rect 21331 37236 21567 37472
rect 21652 37236 21888 37472
rect 21973 37236 22209 37472
rect 22294 37236 22530 37472
rect 22615 37236 22851 37472
rect 22936 37236 23172 37472
rect 23257 37236 23493 37472
rect 23578 37236 23814 37472
rect 23899 37236 24135 37472
rect 24220 37236 24456 37472
rect -3087 36912 -2851 37148
rect -2765 36912 -2529 37148
rect -2443 36912 -2207 37148
rect -2121 36912 -1885 37148
rect -1799 36912 -1563 37148
rect -1477 36912 -1241 37148
rect -1155 36912 -919 37148
rect -833 36912 -597 37148
rect -511 36912 -275 37148
rect -189 36912 47 37148
rect 133 36912 369 37148
rect 455 36912 691 37148
rect 777 36912 1013 37148
rect 1099 36912 1335 37148
rect 1421 36912 1657 37148
rect 1743 36912 1979 37148
rect 2065 36912 2301 37148
rect 2387 36912 2623 37148
rect 2709 36912 2945 37148
rect 3031 36912 3267 37148
rect 3353 36912 3589 37148
rect 3675 36912 3911 37148
rect 3997 36912 4233 37148
rect 4318 36912 4554 37148
rect 4639 36912 4875 37148
rect 4960 36912 5196 37148
rect 5281 36912 5517 37148
rect 5602 36912 5838 37148
rect 5923 36912 6159 37148
rect 6244 36912 6480 37148
rect 6565 36912 6801 37148
rect 6886 36912 7122 37148
rect 7207 36912 7443 37148
rect 7528 36912 7764 37148
rect 7849 36912 8085 37148
rect 8170 36912 8406 37148
rect 8491 36912 8727 37148
rect 8812 36912 9048 37148
rect 9133 36912 9369 37148
rect 9454 36912 9690 37148
rect 9775 36912 10011 37148
rect 10096 36912 10332 37148
rect 10417 36912 10653 37148
rect 10738 36912 10974 37148
rect 11059 36912 11295 37148
rect 11380 36912 11616 37148
rect 11701 36912 11937 37148
rect 12022 36912 12258 37148
rect 12343 36912 12579 37148
rect 12664 36912 12900 37148
rect 12985 36912 13221 37148
rect 13306 36912 13542 37148
rect 13627 36912 13863 37148
rect 13948 36912 14184 37148
rect 14269 36912 14505 37148
rect 14590 36912 14826 37148
rect 14911 36912 15147 37148
rect 15232 36912 15468 37148
rect 15553 36912 15789 37148
rect 15874 36912 16110 37148
rect 16195 36912 16431 37148
rect 16516 36912 16752 37148
rect 16837 36912 17073 37148
rect 17158 36912 17394 37148
rect 17479 36912 17715 37148
rect 17800 36912 18036 37148
rect 18121 36912 18357 37148
rect 18442 36912 18678 37148
rect 18763 36912 18999 37148
rect 19084 36912 19320 37148
rect 19405 36912 19641 37148
rect 19726 36912 19962 37148
rect 20047 36912 20283 37148
rect 20368 36912 20604 37148
rect 20689 36912 20925 37148
rect 21010 36912 21246 37148
rect 21331 36912 21567 37148
rect 21652 36912 21888 37148
rect 21973 36912 22209 37148
rect 22294 36912 22530 37148
rect 22615 36912 22851 37148
rect 22936 36912 23172 37148
rect 23257 36912 23493 37148
rect 23578 36912 23814 37148
rect 23899 36912 24135 37148
rect 24220 36912 24456 37148
rect -3087 36588 -2851 36824
rect -2765 36588 -2529 36824
rect -2443 36588 -2207 36824
rect -2121 36588 -1885 36824
rect -1799 36588 -1563 36824
rect -1477 36588 -1241 36824
rect -1155 36588 -919 36824
rect -833 36588 -597 36824
rect -511 36588 -275 36824
rect -189 36588 47 36824
rect 133 36588 369 36824
rect 455 36588 691 36824
rect 777 36588 1013 36824
rect 1099 36588 1335 36824
rect 1421 36588 1657 36824
rect 1743 36588 1979 36824
rect 2065 36588 2301 36824
rect 2387 36588 2623 36824
rect 2709 36588 2945 36824
rect 3031 36588 3267 36824
rect 3353 36588 3589 36824
rect 3675 36588 3911 36824
rect 3997 36588 4233 36824
rect 4318 36588 4554 36824
rect 4639 36588 4875 36824
rect 4960 36588 5196 36824
rect 5281 36588 5517 36824
rect 5602 36588 5838 36824
rect 5923 36588 6159 36824
rect 6244 36588 6480 36824
rect 6565 36588 6801 36824
rect 6886 36588 7122 36824
rect 7207 36588 7443 36824
rect 7528 36588 7764 36824
rect 7849 36588 8085 36824
rect 8170 36588 8406 36824
rect 8491 36588 8727 36824
rect 8812 36588 9048 36824
rect 9133 36588 9369 36824
rect 9454 36588 9690 36824
rect 9775 36588 10011 36824
rect 10096 36588 10332 36824
rect 10417 36588 10653 36824
rect 10738 36588 10974 36824
rect 11059 36588 11295 36824
rect 11380 36588 11616 36824
rect 11701 36588 11937 36824
rect 12022 36588 12258 36824
rect 12343 36588 12579 36824
rect 12664 36588 12900 36824
rect 12985 36588 13221 36824
rect 13306 36588 13542 36824
rect 13627 36588 13863 36824
rect 13948 36588 14184 36824
rect 14269 36588 14505 36824
rect 14590 36588 14826 36824
rect 14911 36588 15147 36824
rect 15232 36588 15468 36824
rect 15553 36588 15789 36824
rect 15874 36588 16110 36824
rect 16195 36588 16431 36824
rect 16516 36588 16752 36824
rect 16837 36588 17073 36824
rect 17158 36588 17394 36824
rect 17479 36588 17715 36824
rect 17800 36588 18036 36824
rect 18121 36588 18357 36824
rect 18442 36588 18678 36824
rect 18763 36588 18999 36824
rect 19084 36588 19320 36824
rect 19405 36588 19641 36824
rect 19726 36588 19962 36824
rect 20047 36588 20283 36824
rect 20368 36588 20604 36824
rect 20689 36588 20925 36824
rect 21010 36588 21246 36824
rect 21331 36588 21567 36824
rect 21652 36588 21888 36824
rect 21973 36588 22209 36824
rect 22294 36588 22530 36824
rect 22615 36588 22851 36824
rect 22936 36588 23172 36824
rect 23257 36588 23493 36824
rect 23578 36588 23814 36824
rect 23899 36588 24135 36824
rect 24220 36588 24456 36824
rect -3087 36264 -2851 36500
rect -2765 36264 -2529 36500
rect -2443 36264 -2207 36500
rect -2121 36264 -1885 36500
rect -1799 36264 -1563 36500
rect -1477 36264 -1241 36500
rect -1155 36264 -919 36500
rect -833 36264 -597 36500
rect -511 36264 -275 36500
rect -189 36264 47 36500
rect 133 36264 369 36500
rect 455 36264 691 36500
rect 777 36264 1013 36500
rect 1099 36264 1335 36500
rect 1421 36264 1657 36500
rect 1743 36264 1979 36500
rect 2065 36264 2301 36500
rect 2387 36264 2623 36500
rect 2709 36264 2945 36500
rect 3031 36264 3267 36500
rect 3353 36264 3589 36500
rect 3675 36264 3911 36500
rect 3997 36264 4233 36500
rect 4318 36264 4554 36500
rect 4639 36264 4875 36500
rect 4960 36264 5196 36500
rect 5281 36264 5517 36500
rect 5602 36264 5838 36500
rect 5923 36264 6159 36500
rect 6244 36264 6480 36500
rect 6565 36264 6801 36500
rect 6886 36264 7122 36500
rect 7207 36264 7443 36500
rect 7528 36264 7764 36500
rect 7849 36264 8085 36500
rect 8170 36264 8406 36500
rect 8491 36264 8727 36500
rect 8812 36264 9048 36500
rect 9133 36264 9369 36500
rect 9454 36264 9690 36500
rect 9775 36264 10011 36500
rect 10096 36264 10332 36500
rect 10417 36264 10653 36500
rect 10738 36264 10974 36500
rect 11059 36264 11295 36500
rect 11380 36264 11616 36500
rect 11701 36264 11937 36500
rect 12022 36264 12258 36500
rect 12343 36264 12579 36500
rect 12664 36264 12900 36500
rect 12985 36264 13221 36500
rect 13306 36264 13542 36500
rect 13627 36264 13863 36500
rect 13948 36264 14184 36500
rect 14269 36264 14505 36500
rect 14590 36264 14826 36500
rect 14911 36264 15147 36500
rect 15232 36264 15468 36500
rect 15553 36264 15789 36500
rect 15874 36264 16110 36500
rect 16195 36264 16431 36500
rect 16516 36264 16752 36500
rect 16837 36264 17073 36500
rect 17158 36264 17394 36500
rect 17479 36264 17715 36500
rect 17800 36264 18036 36500
rect 18121 36264 18357 36500
rect 18442 36264 18678 36500
rect 18763 36264 18999 36500
rect 19084 36264 19320 36500
rect 19405 36264 19641 36500
rect 19726 36264 19962 36500
rect 20047 36264 20283 36500
rect 20368 36264 20604 36500
rect 20689 36264 20925 36500
rect 21010 36264 21246 36500
rect 21331 36264 21567 36500
rect 21652 36264 21888 36500
rect 21973 36264 22209 36500
rect 22294 36264 22530 36500
rect 22615 36264 22851 36500
rect 22936 36264 23172 36500
rect 23257 36264 23493 36500
rect 23578 36264 23814 36500
rect 23899 36264 24135 36500
rect 24220 36264 24456 36500
rect -3087 35940 -2851 36176
rect -2765 35940 -2529 36176
rect -2443 35940 -2207 36176
rect -2121 35940 -1885 36176
rect -1799 35940 -1563 36176
rect -1477 35940 -1241 36176
rect -1155 35940 -919 36176
rect -833 35940 -597 36176
rect -511 35940 -275 36176
rect -189 35940 47 36176
rect 133 35940 369 36176
rect 455 35940 691 36176
rect 777 35940 1013 36176
rect 1099 35940 1335 36176
rect 1421 35940 1657 36176
rect 1743 35940 1979 36176
rect 2065 35940 2301 36176
rect 2387 35940 2623 36176
rect 2709 35940 2945 36176
rect 3031 35940 3267 36176
rect 3353 35940 3589 36176
rect 3675 35940 3911 36176
rect 3997 35940 4233 36176
rect 4318 35940 4554 36176
rect 4639 35940 4875 36176
rect 4960 35940 5196 36176
rect 5281 35940 5517 36176
rect 5602 35940 5838 36176
rect 5923 35940 6159 36176
rect 6244 35940 6480 36176
rect 6565 35940 6801 36176
rect 6886 35940 7122 36176
rect 7207 35940 7443 36176
rect 7528 35940 7764 36176
rect 7849 35940 8085 36176
rect 8170 35940 8406 36176
rect 8491 35940 8727 36176
rect 8812 35940 9048 36176
rect 9133 35940 9369 36176
rect 9454 35940 9690 36176
rect 9775 35940 10011 36176
rect 10096 35940 10332 36176
rect 10417 35940 10653 36176
rect 10738 35940 10974 36176
rect 11059 35940 11295 36176
rect 11380 35940 11616 36176
rect 11701 35940 11937 36176
rect 12022 35940 12258 36176
rect 12343 35940 12579 36176
rect 12664 35940 12900 36176
rect 12985 35940 13221 36176
rect 13306 35940 13542 36176
rect 13627 35940 13863 36176
rect 13948 35940 14184 36176
rect 14269 35940 14505 36176
rect 14590 35940 14826 36176
rect 14911 35940 15147 36176
rect 15232 35940 15468 36176
rect 15553 35940 15789 36176
rect 15874 35940 16110 36176
rect 16195 35940 16431 36176
rect 16516 35940 16752 36176
rect 16837 35940 17073 36176
rect 17158 35940 17394 36176
rect 17479 35940 17715 36176
rect 17800 35940 18036 36176
rect 18121 35940 18357 36176
rect 18442 35940 18678 36176
rect 18763 35940 18999 36176
rect 19084 35940 19320 36176
rect 19405 35940 19641 36176
rect 19726 35940 19962 36176
rect 20047 35940 20283 36176
rect 20368 35940 20604 36176
rect 20689 35940 20925 36176
rect 21010 35940 21246 36176
rect 21331 35940 21567 36176
rect 21652 35940 21888 36176
rect 21973 35940 22209 36176
rect 22294 35940 22530 36176
rect 22615 35940 22851 36176
rect 22936 35940 23172 36176
rect 23257 35940 23493 36176
rect 23578 35940 23814 36176
rect 23899 35940 24135 36176
rect 24220 35940 24456 36176
rect -3087 35616 -2851 35852
rect -2765 35616 -2529 35852
rect -2443 35616 -2207 35852
rect -2121 35616 -1885 35852
rect -1799 35616 -1563 35852
rect -1477 35616 -1241 35852
rect -1155 35616 -919 35852
rect -833 35616 -597 35852
rect -511 35616 -275 35852
rect -189 35616 47 35852
rect 133 35616 369 35852
rect 455 35616 691 35852
rect 777 35616 1013 35852
rect 1099 35616 1335 35852
rect 1421 35616 1657 35852
rect 1743 35616 1979 35852
rect 2065 35616 2301 35852
rect 2387 35616 2623 35852
rect 2709 35616 2945 35852
rect 3031 35616 3267 35852
rect 3353 35616 3589 35852
rect 3675 35616 3911 35852
rect 3997 35616 4233 35852
rect 4318 35616 4554 35852
rect 4639 35616 4875 35852
rect 4960 35616 5196 35852
rect 5281 35616 5517 35852
rect 5602 35616 5838 35852
rect 5923 35616 6159 35852
rect 6244 35616 6480 35852
rect 6565 35616 6801 35852
rect 6886 35616 7122 35852
rect 7207 35616 7443 35852
rect 7528 35616 7764 35852
rect 7849 35616 8085 35852
rect 8170 35616 8406 35852
rect 8491 35616 8727 35852
rect 8812 35616 9048 35852
rect 9133 35616 9369 35852
rect 9454 35616 9690 35852
rect 9775 35616 10011 35852
rect 10096 35616 10332 35852
rect 10417 35616 10653 35852
rect 10738 35616 10974 35852
rect 11059 35616 11295 35852
rect 11380 35616 11616 35852
rect 11701 35616 11937 35852
rect 12022 35616 12258 35852
rect 12343 35616 12579 35852
rect 12664 35616 12900 35852
rect 12985 35616 13221 35852
rect 13306 35616 13542 35852
rect 13627 35616 13863 35852
rect 13948 35616 14184 35852
rect 14269 35616 14505 35852
rect 14590 35616 14826 35852
rect 14911 35616 15147 35852
rect 15232 35616 15468 35852
rect 15553 35616 15789 35852
rect 15874 35616 16110 35852
rect 16195 35616 16431 35852
rect 16516 35616 16752 35852
rect 16837 35616 17073 35852
rect 17158 35616 17394 35852
rect 17479 35616 17715 35852
rect 17800 35616 18036 35852
rect 18121 35616 18357 35852
rect 18442 35616 18678 35852
rect 18763 35616 18999 35852
rect 19084 35616 19320 35852
rect 19405 35616 19641 35852
rect 19726 35616 19962 35852
rect 20047 35616 20283 35852
rect 20368 35616 20604 35852
rect 20689 35616 20925 35852
rect 21010 35616 21246 35852
rect 21331 35616 21567 35852
rect 21652 35616 21888 35852
rect 21973 35616 22209 35852
rect 22294 35616 22530 35852
rect 22615 35616 22851 35852
rect 22936 35616 23172 35852
rect 23257 35616 23493 35852
rect 23578 35616 23814 35852
rect 23899 35616 24135 35852
rect 24220 35616 24456 35852
rect -3087 35292 -2851 35528
rect -2765 35292 -2529 35528
rect -2443 35292 -2207 35528
rect -2121 35292 -1885 35528
rect -1799 35292 -1563 35528
rect -1477 35292 -1241 35528
rect -1155 35292 -919 35528
rect -833 35292 -597 35528
rect -511 35292 -275 35528
rect -189 35292 47 35528
rect 133 35292 369 35528
rect 455 35292 691 35528
rect 777 35292 1013 35528
rect 1099 35292 1335 35528
rect 1421 35292 1657 35528
rect 1743 35292 1979 35528
rect 2065 35292 2301 35528
rect 2387 35292 2623 35528
rect 2709 35292 2945 35528
rect 3031 35292 3267 35528
rect 3353 35292 3589 35528
rect 3675 35292 3911 35528
rect 3997 35292 4233 35528
rect 4318 35292 4554 35528
rect 4639 35292 4875 35528
rect 4960 35292 5196 35528
rect 5281 35292 5517 35528
rect 5602 35292 5838 35528
rect 5923 35292 6159 35528
rect 6244 35292 6480 35528
rect 6565 35292 6801 35528
rect 6886 35292 7122 35528
rect 7207 35292 7443 35528
rect 7528 35292 7764 35528
rect 7849 35292 8085 35528
rect 8170 35292 8406 35528
rect 8491 35292 8727 35528
rect 8812 35292 9048 35528
rect 9133 35292 9369 35528
rect 9454 35292 9690 35528
rect 9775 35292 10011 35528
rect 10096 35292 10332 35528
rect 10417 35292 10653 35528
rect 10738 35292 10974 35528
rect 11059 35292 11295 35528
rect 11380 35292 11616 35528
rect 11701 35292 11937 35528
rect 12022 35292 12258 35528
rect 12343 35292 12579 35528
rect 12664 35292 12900 35528
rect 12985 35292 13221 35528
rect 13306 35292 13542 35528
rect 13627 35292 13863 35528
rect 13948 35292 14184 35528
rect 14269 35292 14505 35528
rect 14590 35292 14826 35528
rect 14911 35292 15147 35528
rect 15232 35292 15468 35528
rect 15553 35292 15789 35528
rect 15874 35292 16110 35528
rect 16195 35292 16431 35528
rect 16516 35292 16752 35528
rect 16837 35292 17073 35528
rect 17158 35292 17394 35528
rect 17479 35292 17715 35528
rect 17800 35292 18036 35528
rect 18121 35292 18357 35528
rect 18442 35292 18678 35528
rect 18763 35292 18999 35528
rect 19084 35292 19320 35528
rect 19405 35292 19641 35528
rect 19726 35292 19962 35528
rect 20047 35292 20283 35528
rect 20368 35292 20604 35528
rect 20689 35292 20925 35528
rect 21010 35292 21246 35528
rect 21331 35292 21567 35528
rect 21652 35292 21888 35528
rect 21973 35292 22209 35528
rect 22294 35292 22530 35528
rect 22615 35292 22851 35528
rect 22936 35292 23172 35528
rect 23257 35292 23493 35528
rect 23578 35292 23814 35528
rect 23899 35292 24135 35528
rect 24220 35292 24456 35528
rect -3087 34968 -2851 35204
rect -2765 34968 -2529 35204
rect -2443 34968 -2207 35204
rect -2121 34968 -1885 35204
rect -1799 34968 -1563 35204
rect -1477 34968 -1241 35204
rect -1155 34968 -919 35204
rect -833 34968 -597 35204
rect -511 34968 -275 35204
rect -189 34968 47 35204
rect 133 34968 369 35204
rect 455 34968 691 35204
rect 777 34968 1013 35204
rect 1099 34968 1335 35204
rect 1421 34968 1657 35204
rect 1743 34968 1979 35204
rect 2065 34968 2301 35204
rect 2387 34968 2623 35204
rect 2709 34968 2945 35204
rect 3031 34968 3267 35204
rect 3353 34968 3589 35204
rect 3675 34968 3911 35204
rect 3997 34968 4233 35204
rect 4318 34968 4554 35204
rect 4639 34968 4875 35204
rect 4960 34968 5196 35204
rect 5281 34968 5517 35204
rect 5602 34968 5838 35204
rect 5923 34968 6159 35204
rect 6244 34968 6480 35204
rect 6565 34968 6801 35204
rect 6886 34968 7122 35204
rect 7207 34968 7443 35204
rect 7528 34968 7764 35204
rect 7849 34968 8085 35204
rect 8170 34968 8406 35204
rect 8491 34968 8727 35204
rect 8812 34968 9048 35204
rect 9133 34968 9369 35204
rect 9454 34968 9690 35204
rect 9775 34968 10011 35204
rect 10096 34968 10332 35204
rect 10417 34968 10653 35204
rect 10738 34968 10974 35204
rect 11059 34968 11295 35204
rect 11380 34968 11616 35204
rect 11701 34968 11937 35204
rect 12022 34968 12258 35204
rect 12343 34968 12579 35204
rect 12664 34968 12900 35204
rect 12985 34968 13221 35204
rect 13306 34968 13542 35204
rect 13627 34968 13863 35204
rect 13948 34968 14184 35204
rect 14269 34968 14505 35204
rect 14590 34968 14826 35204
rect 14911 34968 15147 35204
rect 15232 34968 15468 35204
rect 15553 34968 15789 35204
rect 15874 34968 16110 35204
rect 16195 34968 16431 35204
rect 16516 34968 16752 35204
rect 16837 34968 17073 35204
rect 17158 34968 17394 35204
rect 17479 34968 17715 35204
rect 17800 34968 18036 35204
rect 18121 34968 18357 35204
rect 18442 34968 18678 35204
rect 18763 34968 18999 35204
rect 19084 34968 19320 35204
rect 19405 34968 19641 35204
rect 19726 34968 19962 35204
rect 20047 34968 20283 35204
rect 20368 34968 20604 35204
rect 20689 34968 20925 35204
rect 21010 34968 21246 35204
rect 21331 34968 21567 35204
rect 21652 34968 21888 35204
rect 21973 34968 22209 35204
rect 22294 34968 22530 35204
rect 22615 34968 22851 35204
rect 22936 34968 23172 35204
rect 23257 34968 23493 35204
rect 23578 34968 23814 35204
rect 23899 34968 24135 35204
rect 24220 34968 24456 35204
rect -3087 34644 -2851 34880
rect -2765 34644 -2529 34880
rect -2443 34644 -2207 34880
rect -2121 34644 -1885 34880
rect -1799 34644 -1563 34880
rect -1477 34644 -1241 34880
rect -1155 34644 -919 34880
rect -833 34644 -597 34880
rect -511 34644 -275 34880
rect -189 34644 47 34880
rect 133 34644 369 34880
rect 455 34644 691 34880
rect 777 34644 1013 34880
rect 1099 34644 1335 34880
rect 1421 34644 1657 34880
rect 1743 34644 1979 34880
rect 2065 34644 2301 34880
rect 2387 34644 2623 34880
rect 2709 34644 2945 34880
rect 3031 34644 3267 34880
rect 3353 34644 3589 34880
rect 3675 34644 3911 34880
rect 3997 34644 4233 34880
rect 4318 34644 4554 34880
rect 4639 34644 4875 34880
rect 4960 34644 5196 34880
rect 5281 34644 5517 34880
rect 5602 34644 5838 34880
rect 5923 34644 6159 34880
rect 6244 34644 6480 34880
rect 6565 34644 6801 34880
rect 6886 34644 7122 34880
rect 7207 34644 7443 34880
rect 7528 34644 7764 34880
rect 7849 34644 8085 34880
rect 8170 34644 8406 34880
rect 8491 34644 8727 34880
rect 8812 34644 9048 34880
rect 9133 34644 9369 34880
rect 9454 34644 9690 34880
rect 9775 34644 10011 34880
rect 10096 34644 10332 34880
rect 10417 34644 10653 34880
rect 10738 34644 10974 34880
rect 11059 34644 11295 34880
rect 11380 34644 11616 34880
rect 11701 34644 11937 34880
rect 12022 34644 12258 34880
rect 12343 34644 12579 34880
rect 12664 34644 12900 34880
rect 12985 34644 13221 34880
rect 13306 34644 13542 34880
rect 13627 34644 13863 34880
rect 13948 34644 14184 34880
rect 14269 34644 14505 34880
rect 14590 34644 14826 34880
rect 14911 34644 15147 34880
rect 15232 34644 15468 34880
rect 15553 34644 15789 34880
rect 15874 34644 16110 34880
rect 16195 34644 16431 34880
rect 16516 34644 16752 34880
rect 16837 34644 17073 34880
rect 17158 34644 17394 34880
rect 17479 34644 17715 34880
rect 17800 34644 18036 34880
rect 18121 34644 18357 34880
rect 18442 34644 18678 34880
rect 18763 34644 18999 34880
rect 19084 34644 19320 34880
rect 19405 34644 19641 34880
rect 19726 34644 19962 34880
rect 20047 34644 20283 34880
rect 20368 34644 20604 34880
rect 20689 34644 20925 34880
rect 21010 34644 21246 34880
rect 21331 34644 21567 34880
rect 21652 34644 21888 34880
rect 21973 34644 22209 34880
rect 22294 34644 22530 34880
rect 22615 34644 22851 34880
rect 22936 34644 23172 34880
rect 23257 34644 23493 34880
rect 23578 34644 23814 34880
rect 23899 34644 24135 34880
rect 24220 34644 24456 34880
rect -3185 18187 -2949 18423
rect -2862 18187 -2626 18423
rect -2539 18187 -2303 18423
rect -2216 18187 -1980 18423
rect -1893 18187 -1657 18423
rect -1570 18187 -1334 18423
rect -1247 18187 -1011 18423
rect -924 18187 -688 18423
rect -601 18187 -365 18423
rect -278 18187 -42 18423
rect 45 18187 281 18423
rect 368 18187 604 18423
rect 691 18187 927 18423
rect 1014 18187 1250 18423
rect 1337 18187 1573 18423
rect 1660 18187 1896 18423
rect 1983 18187 2219 18423
rect 2306 18187 2542 18423
rect 2629 18187 2865 18423
rect 2952 18187 3188 18423
rect 3275 18187 3511 18423
rect 3598 18187 3834 18423
rect 3921 18187 4157 18423
rect 4244 18187 4480 18423
rect 4567 18187 4803 18423
rect 4890 18187 5126 18423
rect 5213 18187 5449 18423
rect 5536 18187 5772 18423
rect 5859 18187 6095 18423
rect 6182 18187 6418 18423
rect 6505 18187 6741 18423
rect 6828 18187 7064 18423
rect 7150 18187 7386 18423
rect 7472 18187 7708 18423
rect 7794 18187 8030 18423
rect 8116 18187 8352 18423
rect 8438 18187 8674 18423
rect 8760 18187 8996 18423
rect 9082 18187 9318 18423
rect 9404 18187 9640 18423
rect 9726 18187 9962 18423
rect 10048 18187 10284 18423
rect 10370 18187 10606 18423
rect 10692 18187 10928 18423
rect 11014 18187 11250 18423
rect 11336 18187 11572 18423
rect 11658 18187 11894 18423
rect 11980 18187 12216 18423
rect 12302 18187 12538 18423
rect 12624 18187 12860 18423
rect 12946 18187 13182 18423
rect 13268 18187 13504 18423
rect 13590 18187 13826 18423
rect 13912 18187 14148 18423
rect 14234 18187 14470 18423
rect 14556 18187 14792 18423
rect 14878 18187 15114 18423
rect 15200 18187 15436 18423
rect 15522 18187 15758 18423
rect 15844 18187 16080 18423
rect 16166 18187 16402 18423
rect 16488 18187 16724 18423
rect 16810 18187 17046 18423
rect 17132 18187 17368 18423
rect 17454 18187 17690 18423
rect 17776 18187 18012 18423
rect 18098 18187 18334 18423
rect 18420 18187 18656 18423
rect 18742 18187 18978 18423
rect 19064 18187 19300 18423
rect 19386 18187 19622 18423
rect 19708 18187 19944 18423
rect 20030 18187 20266 18423
rect 20352 18187 20588 18423
rect 20674 18187 20910 18423
rect 20996 18187 21232 18423
rect 21318 18187 21554 18423
rect 21640 18187 21876 18423
rect 21962 18187 22198 18423
rect 22284 18187 22520 18423
rect 22606 18187 22842 18423
rect 22928 18187 23164 18423
rect 23250 18187 23486 18423
rect 23572 18187 23808 18423
rect 23894 18187 24130 18423
rect 24216 18187 24452 18423
rect -3185 17851 -2949 18087
rect -2862 17851 -2626 18087
rect -2539 17851 -2303 18087
rect -2216 17851 -1980 18087
rect -1893 17851 -1657 18087
rect -1570 17851 -1334 18087
rect -1247 17851 -1011 18087
rect -924 17851 -688 18087
rect -601 17851 -365 18087
rect -278 17851 -42 18087
rect 45 17851 281 18087
rect 368 17851 604 18087
rect 691 17851 927 18087
rect 1014 17851 1250 18087
rect 1337 17851 1573 18087
rect 1660 17851 1896 18087
rect 1983 17851 2219 18087
rect 2306 17851 2542 18087
rect 2629 17851 2865 18087
rect 2952 17851 3188 18087
rect 3275 17851 3511 18087
rect 3598 17851 3834 18087
rect 3921 17851 4157 18087
rect 4244 17851 4480 18087
rect 4567 17851 4803 18087
rect 4890 17851 5126 18087
rect 5213 17851 5449 18087
rect 5536 17851 5772 18087
rect 5859 17851 6095 18087
rect 6182 17851 6418 18087
rect 6505 17851 6741 18087
rect 6828 17851 7064 18087
rect 7150 17851 7386 18087
rect 7472 17851 7708 18087
rect 7794 17851 8030 18087
rect 8116 17851 8352 18087
rect 8438 17851 8674 18087
rect 8760 17851 8996 18087
rect 9082 17851 9318 18087
rect 9404 17851 9640 18087
rect 9726 17851 9962 18087
rect 10048 17851 10284 18087
rect 10370 17851 10606 18087
rect 10692 17851 10928 18087
rect 11014 17851 11250 18087
rect 11336 17851 11572 18087
rect 11658 17851 11894 18087
rect 11980 17851 12216 18087
rect 12302 17851 12538 18087
rect 12624 17851 12860 18087
rect 12946 17851 13182 18087
rect 13268 17851 13504 18087
rect 13590 17851 13826 18087
rect 13912 17851 14148 18087
rect 14234 17851 14470 18087
rect 14556 17851 14792 18087
rect 14878 17851 15114 18087
rect 15200 17851 15436 18087
rect 15522 17851 15758 18087
rect 15844 17851 16080 18087
rect 16166 17851 16402 18087
rect 16488 17851 16724 18087
rect 16810 17851 17046 18087
rect 17132 17851 17368 18087
rect 17454 17851 17690 18087
rect 17776 17851 18012 18087
rect 18098 17851 18334 18087
rect 18420 17851 18656 18087
rect 18742 17851 18978 18087
rect 19064 17851 19300 18087
rect 19386 17851 19622 18087
rect 19708 17851 19944 18087
rect 20030 17851 20266 18087
rect 20352 17851 20588 18087
rect 20674 17851 20910 18087
rect 20996 17851 21232 18087
rect 21318 17851 21554 18087
rect 21640 17851 21876 18087
rect 21962 17851 22198 18087
rect 22284 17851 22520 18087
rect 22606 17851 22842 18087
rect 22928 17851 23164 18087
rect 23250 17851 23486 18087
rect 23572 17851 23808 18087
rect 23894 17851 24130 18087
rect 24216 17851 24452 18087
rect -3185 17515 -2949 17751
rect -2862 17515 -2626 17751
rect -2539 17515 -2303 17751
rect -2216 17515 -1980 17751
rect -1893 17515 -1657 17751
rect -1570 17515 -1334 17751
rect -1247 17515 -1011 17751
rect -924 17515 -688 17751
rect -601 17515 -365 17751
rect -278 17515 -42 17751
rect 45 17515 281 17751
rect 368 17515 604 17751
rect 691 17515 927 17751
rect 1014 17515 1250 17751
rect 1337 17515 1573 17751
rect 1660 17515 1896 17751
rect 1983 17515 2219 17751
rect 2306 17515 2542 17751
rect 2629 17515 2865 17751
rect 2952 17515 3188 17751
rect 3275 17515 3511 17751
rect 3598 17515 3834 17751
rect 3921 17515 4157 17751
rect 4244 17515 4480 17751
rect 4567 17515 4803 17751
rect 4890 17515 5126 17751
rect 5213 17515 5449 17751
rect 5536 17515 5772 17751
rect 5859 17515 6095 17751
rect 6182 17515 6418 17751
rect 6505 17515 6741 17751
rect 6828 17515 7064 17751
rect 7150 17515 7386 17751
rect 7472 17515 7708 17751
rect 7794 17515 8030 17751
rect 8116 17515 8352 17751
rect 8438 17515 8674 17751
rect 8760 17515 8996 17751
rect 9082 17515 9318 17751
rect 9404 17515 9640 17751
rect 9726 17515 9962 17751
rect 10048 17515 10284 17751
rect 10370 17515 10606 17751
rect 10692 17515 10928 17751
rect 11014 17515 11250 17751
rect 11336 17515 11572 17751
rect 11658 17515 11894 17751
rect 11980 17515 12216 17751
rect 12302 17515 12538 17751
rect 12624 17515 12860 17751
rect 12946 17515 13182 17751
rect 13268 17515 13504 17751
rect 13590 17515 13826 17751
rect 13912 17515 14148 17751
rect 14234 17515 14470 17751
rect 14556 17515 14792 17751
rect 14878 17515 15114 17751
rect 15200 17515 15436 17751
rect 15522 17515 15758 17751
rect 15844 17515 16080 17751
rect 16166 17515 16402 17751
rect 16488 17515 16724 17751
rect 16810 17515 17046 17751
rect 17132 17515 17368 17751
rect 17454 17515 17690 17751
rect 17776 17515 18012 17751
rect 18098 17515 18334 17751
rect 18420 17515 18656 17751
rect 18742 17515 18978 17751
rect 19064 17515 19300 17751
rect 19386 17515 19622 17751
rect 19708 17515 19944 17751
rect 20030 17515 20266 17751
rect 20352 17515 20588 17751
rect 20674 17515 20910 17751
rect 20996 17515 21232 17751
rect 21318 17515 21554 17751
rect 21640 17515 21876 17751
rect 21962 17515 22198 17751
rect 22284 17515 22520 17751
rect 22606 17515 22842 17751
rect 22928 17515 23164 17751
rect 23250 17515 23486 17751
rect 23572 17515 23808 17751
rect 23894 17515 24130 17751
rect 24216 17515 24452 17751
rect -3185 17179 -2949 17415
rect -2862 17179 -2626 17415
rect -2539 17179 -2303 17415
rect -2216 17179 -1980 17415
rect -1893 17179 -1657 17415
rect -1570 17179 -1334 17415
rect -1247 17179 -1011 17415
rect -924 17179 -688 17415
rect -601 17179 -365 17415
rect -278 17179 -42 17415
rect 45 17179 281 17415
rect 368 17179 604 17415
rect 691 17179 927 17415
rect 1014 17179 1250 17415
rect 1337 17179 1573 17415
rect 1660 17179 1896 17415
rect 1983 17179 2219 17415
rect 2306 17179 2542 17415
rect 2629 17179 2865 17415
rect 2952 17179 3188 17415
rect 3275 17179 3511 17415
rect 3598 17179 3834 17415
rect 3921 17179 4157 17415
rect 4244 17179 4480 17415
rect 4567 17179 4803 17415
rect 4890 17179 5126 17415
rect 5213 17179 5449 17415
rect 5536 17179 5772 17415
rect 5859 17179 6095 17415
rect 6182 17179 6418 17415
rect 6505 17179 6741 17415
rect 6828 17179 7064 17415
rect 7150 17179 7386 17415
rect 7472 17179 7708 17415
rect 7794 17179 8030 17415
rect 8116 17179 8352 17415
rect 8438 17179 8674 17415
rect 8760 17179 8996 17415
rect 9082 17179 9318 17415
rect 9404 17179 9640 17415
rect 9726 17179 9962 17415
rect 10048 17179 10284 17415
rect 10370 17179 10606 17415
rect 10692 17179 10928 17415
rect 11014 17179 11250 17415
rect 11336 17179 11572 17415
rect 11658 17179 11894 17415
rect 11980 17179 12216 17415
rect 12302 17179 12538 17415
rect 12624 17179 12860 17415
rect 12946 17179 13182 17415
rect 13268 17179 13504 17415
rect 13590 17179 13826 17415
rect 13912 17179 14148 17415
rect 14234 17179 14470 17415
rect 14556 17179 14792 17415
rect 14878 17179 15114 17415
rect 15200 17179 15436 17415
rect 15522 17179 15758 17415
rect 15844 17179 16080 17415
rect 16166 17179 16402 17415
rect 16488 17179 16724 17415
rect 16810 17179 17046 17415
rect 17132 17179 17368 17415
rect 17454 17179 17690 17415
rect 17776 17179 18012 17415
rect 18098 17179 18334 17415
rect 18420 17179 18656 17415
rect 18742 17179 18978 17415
rect 19064 17179 19300 17415
rect 19386 17179 19622 17415
rect 19708 17179 19944 17415
rect 20030 17179 20266 17415
rect 20352 17179 20588 17415
rect 20674 17179 20910 17415
rect 20996 17179 21232 17415
rect 21318 17179 21554 17415
rect 21640 17179 21876 17415
rect 21962 17179 22198 17415
rect 22284 17179 22520 17415
rect 22606 17179 22842 17415
rect 22928 17179 23164 17415
rect 23250 17179 23486 17415
rect 23572 17179 23808 17415
rect 23894 17179 24130 17415
rect 24216 17179 24452 17415
rect -3185 16843 -2949 17079
rect -2862 16843 -2626 17079
rect -2539 16843 -2303 17079
rect -2216 16843 -1980 17079
rect -1893 16843 -1657 17079
rect -1570 16843 -1334 17079
rect -1247 16843 -1011 17079
rect -924 16843 -688 17079
rect -601 16843 -365 17079
rect -278 16843 -42 17079
rect 45 16843 281 17079
rect 368 16843 604 17079
rect 691 16843 927 17079
rect 1014 16843 1250 17079
rect 1337 16843 1573 17079
rect 1660 16843 1896 17079
rect 1983 16843 2219 17079
rect 2306 16843 2542 17079
rect 2629 16843 2865 17079
rect 2952 16843 3188 17079
rect 3275 16843 3511 17079
rect 3598 16843 3834 17079
rect 3921 16843 4157 17079
rect 4244 16843 4480 17079
rect 4567 16843 4803 17079
rect 4890 16843 5126 17079
rect 5213 16843 5449 17079
rect 5536 16843 5772 17079
rect 5859 16843 6095 17079
rect 6182 16843 6418 17079
rect 6505 16843 6741 17079
rect 6828 16843 7064 17079
rect 7150 16843 7386 17079
rect 7472 16843 7708 17079
rect 7794 16843 8030 17079
rect 8116 16843 8352 17079
rect 8438 16843 8674 17079
rect 8760 16843 8996 17079
rect 9082 16843 9318 17079
rect 9404 16843 9640 17079
rect 9726 16843 9962 17079
rect 10048 16843 10284 17079
rect 10370 16843 10606 17079
rect 10692 16843 10928 17079
rect 11014 16843 11250 17079
rect 11336 16843 11572 17079
rect 11658 16843 11894 17079
rect 11980 16843 12216 17079
rect 12302 16843 12538 17079
rect 12624 16843 12860 17079
rect 12946 16843 13182 17079
rect 13268 16843 13504 17079
rect 13590 16843 13826 17079
rect 13912 16843 14148 17079
rect 14234 16843 14470 17079
rect 14556 16843 14792 17079
rect 14878 16843 15114 17079
rect 15200 16843 15436 17079
rect 15522 16843 15758 17079
rect 15844 16843 16080 17079
rect 16166 16843 16402 17079
rect 16488 16843 16724 17079
rect 16810 16843 17046 17079
rect 17132 16843 17368 17079
rect 17454 16843 17690 17079
rect 17776 16843 18012 17079
rect 18098 16843 18334 17079
rect 18420 16843 18656 17079
rect 18742 16843 18978 17079
rect 19064 16843 19300 17079
rect 19386 16843 19622 17079
rect 19708 16843 19944 17079
rect 20030 16843 20266 17079
rect 20352 16843 20588 17079
rect 20674 16843 20910 17079
rect 20996 16843 21232 17079
rect 21318 16843 21554 17079
rect 21640 16843 21876 17079
rect 21962 16843 22198 17079
rect 22284 16843 22520 17079
rect 22606 16843 22842 17079
rect 22928 16843 23164 17079
rect 23250 16843 23486 17079
rect 23572 16843 23808 17079
rect 23894 16843 24130 17079
rect 24216 16843 24452 17079
rect -3185 16507 -2949 16743
rect -2862 16507 -2626 16743
rect -2539 16507 -2303 16743
rect -2216 16507 -1980 16743
rect -1893 16507 -1657 16743
rect -1570 16507 -1334 16743
rect -1247 16507 -1011 16743
rect -924 16507 -688 16743
rect -601 16507 -365 16743
rect -278 16507 -42 16743
rect 45 16507 281 16743
rect 368 16507 604 16743
rect 691 16507 927 16743
rect 1014 16507 1250 16743
rect 1337 16507 1573 16743
rect 1660 16507 1896 16743
rect 1983 16507 2219 16743
rect 2306 16507 2542 16743
rect 2629 16507 2865 16743
rect 2952 16507 3188 16743
rect 3275 16507 3511 16743
rect 3598 16507 3834 16743
rect 3921 16507 4157 16743
rect 4244 16507 4480 16743
rect 4567 16507 4803 16743
rect 4890 16507 5126 16743
rect 5213 16507 5449 16743
rect 5536 16507 5772 16743
rect 5859 16507 6095 16743
rect 6182 16507 6418 16743
rect 6505 16507 6741 16743
rect 6828 16507 7064 16743
rect 7150 16507 7386 16743
rect 7472 16507 7708 16743
rect 7794 16507 8030 16743
rect 8116 16507 8352 16743
rect 8438 16507 8674 16743
rect 8760 16507 8996 16743
rect 9082 16507 9318 16743
rect 9404 16507 9640 16743
rect 9726 16507 9962 16743
rect 10048 16507 10284 16743
rect 10370 16507 10606 16743
rect 10692 16507 10928 16743
rect 11014 16507 11250 16743
rect 11336 16507 11572 16743
rect 11658 16507 11894 16743
rect 11980 16507 12216 16743
rect 12302 16507 12538 16743
rect 12624 16507 12860 16743
rect 12946 16507 13182 16743
rect 13268 16507 13504 16743
rect 13590 16507 13826 16743
rect 13912 16507 14148 16743
rect 14234 16507 14470 16743
rect 14556 16507 14792 16743
rect 14878 16507 15114 16743
rect 15200 16507 15436 16743
rect 15522 16507 15758 16743
rect 15844 16507 16080 16743
rect 16166 16507 16402 16743
rect 16488 16507 16724 16743
rect 16810 16507 17046 16743
rect 17132 16507 17368 16743
rect 17454 16507 17690 16743
rect 17776 16507 18012 16743
rect 18098 16507 18334 16743
rect 18420 16507 18656 16743
rect 18742 16507 18978 16743
rect 19064 16507 19300 16743
rect 19386 16507 19622 16743
rect 19708 16507 19944 16743
rect 20030 16507 20266 16743
rect 20352 16507 20588 16743
rect 20674 16507 20910 16743
rect 20996 16507 21232 16743
rect 21318 16507 21554 16743
rect 21640 16507 21876 16743
rect 21962 16507 22198 16743
rect 22284 16507 22520 16743
rect 22606 16507 22842 16743
rect 22928 16507 23164 16743
rect 23250 16507 23486 16743
rect 23572 16507 23808 16743
rect 23894 16507 24130 16743
rect 24216 16507 24452 16743
rect -3185 16171 -2949 16407
rect -2862 16171 -2626 16407
rect -2539 16171 -2303 16407
rect -2216 16171 -1980 16407
rect -1893 16171 -1657 16407
rect -1570 16171 -1334 16407
rect -1247 16171 -1011 16407
rect -924 16171 -688 16407
rect -601 16171 -365 16407
rect -278 16171 -42 16407
rect 45 16171 281 16407
rect 368 16171 604 16407
rect 691 16171 927 16407
rect 1014 16171 1250 16407
rect 1337 16171 1573 16407
rect 1660 16171 1896 16407
rect 1983 16171 2219 16407
rect 2306 16171 2542 16407
rect 2629 16171 2865 16407
rect 2952 16171 3188 16407
rect 3275 16171 3511 16407
rect 3598 16171 3834 16407
rect 3921 16171 4157 16407
rect 4244 16171 4480 16407
rect 4567 16171 4803 16407
rect 4890 16171 5126 16407
rect 5213 16171 5449 16407
rect 5536 16171 5772 16407
rect 5859 16171 6095 16407
rect 6182 16171 6418 16407
rect 6505 16171 6741 16407
rect 6828 16171 7064 16407
rect 7150 16171 7386 16407
rect 7472 16171 7708 16407
rect 7794 16171 8030 16407
rect 8116 16171 8352 16407
rect 8438 16171 8674 16407
rect 8760 16171 8996 16407
rect 9082 16171 9318 16407
rect 9404 16171 9640 16407
rect 9726 16171 9962 16407
rect 10048 16171 10284 16407
rect 10370 16171 10606 16407
rect 10692 16171 10928 16407
rect 11014 16171 11250 16407
rect 11336 16171 11572 16407
rect 11658 16171 11894 16407
rect 11980 16171 12216 16407
rect 12302 16171 12538 16407
rect 12624 16171 12860 16407
rect 12946 16171 13182 16407
rect 13268 16171 13504 16407
rect 13590 16171 13826 16407
rect 13912 16171 14148 16407
rect 14234 16171 14470 16407
rect 14556 16171 14792 16407
rect 14878 16171 15114 16407
rect 15200 16171 15436 16407
rect 15522 16171 15758 16407
rect 15844 16171 16080 16407
rect 16166 16171 16402 16407
rect 16488 16171 16724 16407
rect 16810 16171 17046 16407
rect 17132 16171 17368 16407
rect 17454 16171 17690 16407
rect 17776 16171 18012 16407
rect 18098 16171 18334 16407
rect 18420 16171 18656 16407
rect 18742 16171 18978 16407
rect 19064 16171 19300 16407
rect 19386 16171 19622 16407
rect 19708 16171 19944 16407
rect 20030 16171 20266 16407
rect 20352 16171 20588 16407
rect 20674 16171 20910 16407
rect 20996 16171 21232 16407
rect 21318 16171 21554 16407
rect 21640 16171 21876 16407
rect 21962 16171 22198 16407
rect 22284 16171 22520 16407
rect 22606 16171 22842 16407
rect 22928 16171 23164 16407
rect 23250 16171 23486 16407
rect 23572 16171 23808 16407
rect 23894 16171 24130 16407
rect 24216 16171 24452 16407
rect -3185 15835 -2949 16071
rect -2862 15835 -2626 16071
rect -2539 15835 -2303 16071
rect -2216 15835 -1980 16071
rect -1893 15835 -1657 16071
rect -1570 15835 -1334 16071
rect -1247 15835 -1011 16071
rect -924 15835 -688 16071
rect -601 15835 -365 16071
rect -278 15835 -42 16071
rect 45 15835 281 16071
rect 368 15835 604 16071
rect 691 15835 927 16071
rect 1014 15835 1250 16071
rect 1337 15835 1573 16071
rect 1660 15835 1896 16071
rect 1983 15835 2219 16071
rect 2306 15835 2542 16071
rect 2629 15835 2865 16071
rect 2952 15835 3188 16071
rect 3275 15835 3511 16071
rect 3598 15835 3834 16071
rect 3921 15835 4157 16071
rect 4244 15835 4480 16071
rect 4567 15835 4803 16071
rect 4890 15835 5126 16071
rect 5213 15835 5449 16071
rect 5536 15835 5772 16071
rect 5859 15835 6095 16071
rect 6182 15835 6418 16071
rect 6505 15835 6741 16071
rect 6828 15835 7064 16071
rect 7150 15835 7386 16071
rect 7472 15835 7708 16071
rect 7794 15835 8030 16071
rect 8116 15835 8352 16071
rect 8438 15835 8674 16071
rect 8760 15835 8996 16071
rect 9082 15835 9318 16071
rect 9404 15835 9640 16071
rect 9726 15835 9962 16071
rect 10048 15835 10284 16071
rect 10370 15835 10606 16071
rect 10692 15835 10928 16071
rect 11014 15835 11250 16071
rect 11336 15835 11572 16071
rect 11658 15835 11894 16071
rect 11980 15835 12216 16071
rect 12302 15835 12538 16071
rect 12624 15835 12860 16071
rect 12946 15835 13182 16071
rect 13268 15835 13504 16071
rect 13590 15835 13826 16071
rect 13912 15835 14148 16071
rect 14234 15835 14470 16071
rect 14556 15835 14792 16071
rect 14878 15835 15114 16071
rect 15200 15835 15436 16071
rect 15522 15835 15758 16071
rect 15844 15835 16080 16071
rect 16166 15835 16402 16071
rect 16488 15835 16724 16071
rect 16810 15835 17046 16071
rect 17132 15835 17368 16071
rect 17454 15835 17690 16071
rect 17776 15835 18012 16071
rect 18098 15835 18334 16071
rect 18420 15835 18656 16071
rect 18742 15835 18978 16071
rect 19064 15835 19300 16071
rect 19386 15835 19622 16071
rect 19708 15835 19944 16071
rect 20030 15835 20266 16071
rect 20352 15835 20588 16071
rect 20674 15835 20910 16071
rect 20996 15835 21232 16071
rect 21318 15835 21554 16071
rect 21640 15835 21876 16071
rect 21962 15835 22198 16071
rect 22284 15835 22520 16071
rect 22606 15835 22842 16071
rect 22928 15835 23164 16071
rect 23250 15835 23486 16071
rect 23572 15835 23808 16071
rect 23894 15835 24130 16071
rect 24216 15835 24452 16071
rect -3185 15499 -2949 15735
rect -2862 15499 -2626 15735
rect -2539 15499 -2303 15735
rect -2216 15499 -1980 15735
rect -1893 15499 -1657 15735
rect -1570 15499 -1334 15735
rect -1247 15499 -1011 15735
rect -924 15499 -688 15735
rect -601 15499 -365 15735
rect -278 15499 -42 15735
rect 45 15499 281 15735
rect 368 15499 604 15735
rect 691 15499 927 15735
rect 1014 15499 1250 15735
rect 1337 15499 1573 15735
rect 1660 15499 1896 15735
rect 1983 15499 2219 15735
rect 2306 15499 2542 15735
rect 2629 15499 2865 15735
rect 2952 15499 3188 15735
rect 3275 15499 3511 15735
rect 3598 15499 3834 15735
rect 3921 15499 4157 15735
rect 4244 15499 4480 15735
rect 4567 15499 4803 15735
rect 4890 15499 5126 15735
rect 5213 15499 5449 15735
rect 5536 15499 5772 15735
rect 5859 15499 6095 15735
rect 6182 15499 6418 15735
rect 6505 15499 6741 15735
rect 6828 15499 7064 15735
rect 7150 15499 7386 15735
rect 7472 15499 7708 15735
rect 7794 15499 8030 15735
rect 8116 15499 8352 15735
rect 8438 15499 8674 15735
rect 8760 15499 8996 15735
rect 9082 15499 9318 15735
rect 9404 15499 9640 15735
rect 9726 15499 9962 15735
rect 10048 15499 10284 15735
rect 10370 15499 10606 15735
rect 10692 15499 10928 15735
rect 11014 15499 11250 15735
rect 11336 15499 11572 15735
rect 11658 15499 11894 15735
rect 11980 15499 12216 15735
rect 12302 15499 12538 15735
rect 12624 15499 12860 15735
rect 12946 15499 13182 15735
rect 13268 15499 13504 15735
rect 13590 15499 13826 15735
rect 13912 15499 14148 15735
rect 14234 15499 14470 15735
rect 14556 15499 14792 15735
rect 14878 15499 15114 15735
rect 15200 15499 15436 15735
rect 15522 15499 15758 15735
rect 15844 15499 16080 15735
rect 16166 15499 16402 15735
rect 16488 15499 16724 15735
rect 16810 15499 17046 15735
rect 17132 15499 17368 15735
rect 17454 15499 17690 15735
rect 17776 15499 18012 15735
rect 18098 15499 18334 15735
rect 18420 15499 18656 15735
rect 18742 15499 18978 15735
rect 19064 15499 19300 15735
rect 19386 15499 19622 15735
rect 19708 15499 19944 15735
rect 20030 15499 20266 15735
rect 20352 15499 20588 15735
rect 20674 15499 20910 15735
rect 20996 15499 21232 15735
rect 21318 15499 21554 15735
rect 21640 15499 21876 15735
rect 21962 15499 22198 15735
rect 22284 15499 22520 15735
rect 22606 15499 22842 15735
rect 22928 15499 23164 15735
rect 23250 15499 23486 15735
rect 23572 15499 23808 15735
rect 23894 15499 24130 15735
rect 24216 15499 24452 15735
rect -3185 15163 -2949 15399
rect -2862 15163 -2626 15399
rect -2539 15163 -2303 15399
rect -2216 15163 -1980 15399
rect -1893 15163 -1657 15399
rect -1570 15163 -1334 15399
rect -1247 15163 -1011 15399
rect -924 15163 -688 15399
rect -601 15163 -365 15399
rect -278 15163 -42 15399
rect 45 15163 281 15399
rect 368 15163 604 15399
rect 691 15163 927 15399
rect 1014 15163 1250 15399
rect 1337 15163 1573 15399
rect 1660 15163 1896 15399
rect 1983 15163 2219 15399
rect 2306 15163 2542 15399
rect 2629 15163 2865 15399
rect 2952 15163 3188 15399
rect 3275 15163 3511 15399
rect 3598 15163 3834 15399
rect 3921 15163 4157 15399
rect 4244 15163 4480 15399
rect 4567 15163 4803 15399
rect 4890 15163 5126 15399
rect 5213 15163 5449 15399
rect 5536 15163 5772 15399
rect 5859 15163 6095 15399
rect 6182 15163 6418 15399
rect 6505 15163 6741 15399
rect 6828 15163 7064 15399
rect 7150 15163 7386 15399
rect 7472 15163 7708 15399
rect 7794 15163 8030 15399
rect 8116 15163 8352 15399
rect 8438 15163 8674 15399
rect 8760 15163 8996 15399
rect 9082 15163 9318 15399
rect 9404 15163 9640 15399
rect 9726 15163 9962 15399
rect 10048 15163 10284 15399
rect 10370 15163 10606 15399
rect 10692 15163 10928 15399
rect 11014 15163 11250 15399
rect 11336 15163 11572 15399
rect 11658 15163 11894 15399
rect 11980 15163 12216 15399
rect 12302 15163 12538 15399
rect 12624 15163 12860 15399
rect 12946 15163 13182 15399
rect 13268 15163 13504 15399
rect 13590 15163 13826 15399
rect 13912 15163 14148 15399
rect 14234 15163 14470 15399
rect 14556 15163 14792 15399
rect 14878 15163 15114 15399
rect 15200 15163 15436 15399
rect 15522 15163 15758 15399
rect 15844 15163 16080 15399
rect 16166 15163 16402 15399
rect 16488 15163 16724 15399
rect 16810 15163 17046 15399
rect 17132 15163 17368 15399
rect 17454 15163 17690 15399
rect 17776 15163 18012 15399
rect 18098 15163 18334 15399
rect 18420 15163 18656 15399
rect 18742 15163 18978 15399
rect 19064 15163 19300 15399
rect 19386 15163 19622 15399
rect 19708 15163 19944 15399
rect 20030 15163 20266 15399
rect 20352 15163 20588 15399
rect 20674 15163 20910 15399
rect 20996 15163 21232 15399
rect 21318 15163 21554 15399
rect 21640 15163 21876 15399
rect 21962 15163 22198 15399
rect 22284 15163 22520 15399
rect 22606 15163 22842 15399
rect 22928 15163 23164 15399
rect 23250 15163 23486 15399
rect 23572 15163 23808 15399
rect 23894 15163 24130 15399
rect 24216 15163 24452 15399
rect -3185 14827 -2949 15063
rect -2862 14827 -2626 15063
rect -2539 14827 -2303 15063
rect -2216 14827 -1980 15063
rect -1893 14827 -1657 15063
rect -1570 14827 -1334 15063
rect -1247 14827 -1011 15063
rect -924 14827 -688 15063
rect -601 14827 -365 15063
rect -278 14827 -42 15063
rect 45 14827 281 15063
rect 368 14827 604 15063
rect 691 14827 927 15063
rect 1014 14827 1250 15063
rect 1337 14827 1573 15063
rect 1660 14827 1896 15063
rect 1983 14827 2219 15063
rect 2306 14827 2542 15063
rect 2629 14827 2865 15063
rect 2952 14827 3188 15063
rect 3275 14827 3511 15063
rect 3598 14827 3834 15063
rect 3921 14827 4157 15063
rect 4244 14827 4480 15063
rect 4567 14827 4803 15063
rect 4890 14827 5126 15063
rect 5213 14827 5449 15063
rect 5536 14827 5772 15063
rect 5859 14827 6095 15063
rect 6182 14827 6418 15063
rect 6505 14827 6741 15063
rect 6828 14827 7064 15063
rect 7150 14827 7386 15063
rect 7472 14827 7708 15063
rect 7794 14827 8030 15063
rect 8116 14827 8352 15063
rect 8438 14827 8674 15063
rect 8760 14827 8996 15063
rect 9082 14827 9318 15063
rect 9404 14827 9640 15063
rect 9726 14827 9962 15063
rect 10048 14827 10284 15063
rect 10370 14827 10606 15063
rect 10692 14827 10928 15063
rect 11014 14827 11250 15063
rect 11336 14827 11572 15063
rect 11658 14827 11894 15063
rect 11980 14827 12216 15063
rect 12302 14827 12538 15063
rect 12624 14827 12860 15063
rect 12946 14827 13182 15063
rect 13268 14827 13504 15063
rect 13590 14827 13826 15063
rect 13912 14827 14148 15063
rect 14234 14827 14470 15063
rect 14556 14827 14792 15063
rect 14878 14827 15114 15063
rect 15200 14827 15436 15063
rect 15522 14827 15758 15063
rect 15844 14827 16080 15063
rect 16166 14827 16402 15063
rect 16488 14827 16724 15063
rect 16810 14827 17046 15063
rect 17132 14827 17368 15063
rect 17454 14827 17690 15063
rect 17776 14827 18012 15063
rect 18098 14827 18334 15063
rect 18420 14827 18656 15063
rect 18742 14827 18978 15063
rect 19064 14827 19300 15063
rect 19386 14827 19622 15063
rect 19708 14827 19944 15063
rect 20030 14827 20266 15063
rect 20352 14827 20588 15063
rect 20674 14827 20910 15063
rect 20996 14827 21232 15063
rect 21318 14827 21554 15063
rect 21640 14827 21876 15063
rect 21962 14827 22198 15063
rect 22284 14827 22520 15063
rect 22606 14827 22842 15063
rect 22928 14827 23164 15063
rect 23250 14827 23486 15063
rect 23572 14827 23808 15063
rect 23894 14827 24130 15063
rect 24216 14827 24452 15063
rect -3185 14491 -2949 14727
rect -2862 14491 -2626 14727
rect -2539 14491 -2303 14727
rect -2216 14491 -1980 14727
rect -1893 14491 -1657 14727
rect -1570 14491 -1334 14727
rect -1247 14491 -1011 14727
rect -924 14491 -688 14727
rect -601 14491 -365 14727
rect -278 14491 -42 14727
rect 45 14491 281 14727
rect 368 14491 604 14727
rect 691 14491 927 14727
rect 1014 14491 1250 14727
rect 1337 14491 1573 14727
rect 1660 14491 1896 14727
rect 1983 14491 2219 14727
rect 2306 14491 2542 14727
rect 2629 14491 2865 14727
rect 2952 14491 3188 14727
rect 3275 14491 3511 14727
rect 3598 14491 3834 14727
rect 3921 14491 4157 14727
rect 4244 14491 4480 14727
rect 4567 14491 4803 14727
rect 4890 14491 5126 14727
rect 5213 14491 5449 14727
rect 5536 14491 5772 14727
rect 5859 14491 6095 14727
rect 6182 14491 6418 14727
rect 6505 14491 6741 14727
rect 6828 14491 7064 14727
rect 7150 14491 7386 14727
rect 7472 14491 7708 14727
rect 7794 14491 8030 14727
rect 8116 14491 8352 14727
rect 8438 14491 8674 14727
rect 8760 14491 8996 14727
rect 9082 14491 9318 14727
rect 9404 14491 9640 14727
rect 9726 14491 9962 14727
rect 10048 14491 10284 14727
rect 10370 14491 10606 14727
rect 10692 14491 10928 14727
rect 11014 14491 11250 14727
rect 11336 14491 11572 14727
rect 11658 14491 11894 14727
rect 11980 14491 12216 14727
rect 12302 14491 12538 14727
rect 12624 14491 12860 14727
rect 12946 14491 13182 14727
rect 13268 14491 13504 14727
rect 13590 14491 13826 14727
rect 13912 14491 14148 14727
rect 14234 14491 14470 14727
rect 14556 14491 14792 14727
rect 14878 14491 15114 14727
rect 15200 14491 15436 14727
rect 15522 14491 15758 14727
rect 15844 14491 16080 14727
rect 16166 14491 16402 14727
rect 16488 14491 16724 14727
rect 16810 14491 17046 14727
rect 17132 14491 17368 14727
rect 17454 14491 17690 14727
rect 17776 14491 18012 14727
rect 18098 14491 18334 14727
rect 18420 14491 18656 14727
rect 18742 14491 18978 14727
rect 19064 14491 19300 14727
rect 19386 14491 19622 14727
rect 19708 14491 19944 14727
rect 20030 14491 20266 14727
rect 20352 14491 20588 14727
rect 20674 14491 20910 14727
rect 20996 14491 21232 14727
rect 21318 14491 21554 14727
rect 21640 14491 21876 14727
rect 21962 14491 22198 14727
rect 22284 14491 22520 14727
rect 22606 14491 22842 14727
rect 22928 14491 23164 14727
rect 23250 14491 23486 14727
rect 23572 14491 23808 14727
rect 23894 14491 24130 14727
rect 24216 14491 24452 14727
rect -3185 14155 -2949 14391
rect -2862 14155 -2626 14391
rect -2539 14155 -2303 14391
rect -2216 14155 -1980 14391
rect -1893 14155 -1657 14391
rect -1570 14155 -1334 14391
rect -1247 14155 -1011 14391
rect -924 14155 -688 14391
rect -601 14155 -365 14391
rect -278 14155 -42 14391
rect 45 14155 281 14391
rect 368 14155 604 14391
rect 691 14155 927 14391
rect 1014 14155 1250 14391
rect 1337 14155 1573 14391
rect 1660 14155 1896 14391
rect 1983 14155 2219 14391
rect 2306 14155 2542 14391
rect 2629 14155 2865 14391
rect 2952 14155 3188 14391
rect 3275 14155 3511 14391
rect 3598 14155 3834 14391
rect 3921 14155 4157 14391
rect 4244 14155 4480 14391
rect 4567 14155 4803 14391
rect 4890 14155 5126 14391
rect 5213 14155 5449 14391
rect 5536 14155 5772 14391
rect 5859 14155 6095 14391
rect 6182 14155 6418 14391
rect 6505 14155 6741 14391
rect 6828 14155 7064 14391
rect 7150 14155 7386 14391
rect 7472 14155 7708 14391
rect 7794 14155 8030 14391
rect 8116 14155 8352 14391
rect 8438 14155 8674 14391
rect 8760 14155 8996 14391
rect 9082 14155 9318 14391
rect 9404 14155 9640 14391
rect 9726 14155 9962 14391
rect 10048 14155 10284 14391
rect 10370 14155 10606 14391
rect 10692 14155 10928 14391
rect 11014 14155 11250 14391
rect 11336 14155 11572 14391
rect 11658 14155 11894 14391
rect 11980 14155 12216 14391
rect 12302 14155 12538 14391
rect 12624 14155 12860 14391
rect 12946 14155 13182 14391
rect 13268 14155 13504 14391
rect 13590 14155 13826 14391
rect 13912 14155 14148 14391
rect 14234 14155 14470 14391
rect 14556 14155 14792 14391
rect 14878 14155 15114 14391
rect 15200 14155 15436 14391
rect 15522 14155 15758 14391
rect 15844 14155 16080 14391
rect 16166 14155 16402 14391
rect 16488 14155 16724 14391
rect 16810 14155 17046 14391
rect 17132 14155 17368 14391
rect 17454 14155 17690 14391
rect 17776 14155 18012 14391
rect 18098 14155 18334 14391
rect 18420 14155 18656 14391
rect 18742 14155 18978 14391
rect 19064 14155 19300 14391
rect 19386 14155 19622 14391
rect 19708 14155 19944 14391
rect 20030 14155 20266 14391
rect 20352 14155 20588 14391
rect 20674 14155 20910 14391
rect 20996 14155 21232 14391
rect 21318 14155 21554 14391
rect 21640 14155 21876 14391
rect 21962 14155 22198 14391
rect 22284 14155 22520 14391
rect 22606 14155 22842 14391
rect 22928 14155 23164 14391
rect 23250 14155 23486 14391
rect 23572 14155 23808 14391
rect 23894 14155 24130 14391
rect 24216 14155 24452 14391
rect -3185 13819 -2949 14055
rect -2862 13819 -2626 14055
rect -2539 13819 -2303 14055
rect -2216 13819 -1980 14055
rect -1893 13819 -1657 14055
rect -1570 13819 -1334 14055
rect -1247 13819 -1011 14055
rect -924 13819 -688 14055
rect -601 13819 -365 14055
rect -278 13819 -42 14055
rect 45 13819 281 14055
rect 368 13819 604 14055
rect 691 13819 927 14055
rect 1014 13819 1250 14055
rect 1337 13819 1573 14055
rect 1660 13819 1896 14055
rect 1983 13819 2219 14055
rect 2306 13819 2542 14055
rect 2629 13819 2865 14055
rect 2952 13819 3188 14055
rect 3275 13819 3511 14055
rect 3598 13819 3834 14055
rect 3921 13819 4157 14055
rect 4244 13819 4480 14055
rect 4567 13819 4803 14055
rect 4890 13819 5126 14055
rect 5213 13819 5449 14055
rect 5536 13819 5772 14055
rect 5859 13819 6095 14055
rect 6182 13819 6418 14055
rect 6505 13819 6741 14055
rect 6828 13819 7064 14055
rect 7150 13819 7386 14055
rect 7472 13819 7708 14055
rect 7794 13819 8030 14055
rect 8116 13819 8352 14055
rect 8438 13819 8674 14055
rect 8760 13819 8996 14055
rect 9082 13819 9318 14055
rect 9404 13819 9640 14055
rect 9726 13819 9962 14055
rect 10048 13819 10284 14055
rect 10370 13819 10606 14055
rect 10692 13819 10928 14055
rect 11014 13819 11250 14055
rect 11336 13819 11572 14055
rect 11658 13819 11894 14055
rect 11980 13819 12216 14055
rect 12302 13819 12538 14055
rect 12624 13819 12860 14055
rect 12946 13819 13182 14055
rect 13268 13819 13504 14055
rect 13590 13819 13826 14055
rect 13912 13819 14148 14055
rect 14234 13819 14470 14055
rect 14556 13819 14792 14055
rect 14878 13819 15114 14055
rect 15200 13819 15436 14055
rect 15522 13819 15758 14055
rect 15844 13819 16080 14055
rect 16166 13819 16402 14055
rect 16488 13819 16724 14055
rect 16810 13819 17046 14055
rect 17132 13819 17368 14055
rect 17454 13819 17690 14055
rect 17776 13819 18012 14055
rect 18098 13819 18334 14055
rect 18420 13819 18656 14055
rect 18742 13819 18978 14055
rect 19064 13819 19300 14055
rect 19386 13819 19622 14055
rect 19708 13819 19944 14055
rect 20030 13819 20266 14055
rect 20352 13819 20588 14055
rect 20674 13819 20910 14055
rect 20996 13819 21232 14055
rect 21318 13819 21554 14055
rect 21640 13819 21876 14055
rect 21962 13819 22198 14055
rect 22284 13819 22520 14055
rect 22606 13819 22842 14055
rect 22928 13819 23164 14055
rect 23250 13819 23486 14055
rect 23572 13819 23808 14055
rect 23894 13819 24130 14055
rect 24216 13819 24452 14055
rect -3185 13483 -2949 13719
rect -2862 13483 -2626 13719
rect -2539 13483 -2303 13719
rect -2216 13483 -1980 13719
rect -1893 13483 -1657 13719
rect -1570 13483 -1334 13719
rect -1247 13483 -1011 13719
rect -924 13483 -688 13719
rect -601 13483 -365 13719
rect -278 13483 -42 13719
rect 45 13483 281 13719
rect 368 13483 604 13719
rect 691 13483 927 13719
rect 1014 13483 1250 13719
rect 1337 13483 1573 13719
rect 1660 13483 1896 13719
rect 1983 13483 2219 13719
rect 2306 13483 2542 13719
rect 2629 13483 2865 13719
rect 2952 13483 3188 13719
rect 3275 13483 3511 13719
rect 3598 13483 3834 13719
rect 3921 13483 4157 13719
rect 4244 13483 4480 13719
rect 4567 13483 4803 13719
rect 4890 13483 5126 13719
rect 5213 13483 5449 13719
rect 5536 13483 5772 13719
rect 5859 13483 6095 13719
rect 6182 13483 6418 13719
rect 6505 13483 6741 13719
rect 6828 13483 7064 13719
rect 7150 13483 7386 13719
rect 7472 13483 7708 13719
rect 7794 13483 8030 13719
rect 8116 13483 8352 13719
rect 8438 13483 8674 13719
rect 8760 13483 8996 13719
rect 9082 13483 9318 13719
rect 9404 13483 9640 13719
rect 9726 13483 9962 13719
rect 10048 13483 10284 13719
rect 10370 13483 10606 13719
rect 10692 13483 10928 13719
rect 11014 13483 11250 13719
rect 11336 13483 11572 13719
rect 11658 13483 11894 13719
rect 11980 13483 12216 13719
rect 12302 13483 12538 13719
rect 12624 13483 12860 13719
rect 12946 13483 13182 13719
rect 13268 13483 13504 13719
rect 13590 13483 13826 13719
rect 13912 13483 14148 13719
rect 14234 13483 14470 13719
rect 14556 13483 14792 13719
rect 14878 13483 15114 13719
rect 15200 13483 15436 13719
rect 15522 13483 15758 13719
rect 15844 13483 16080 13719
rect 16166 13483 16402 13719
rect 16488 13483 16724 13719
rect 16810 13483 17046 13719
rect 17132 13483 17368 13719
rect 17454 13483 17690 13719
rect 17776 13483 18012 13719
rect 18098 13483 18334 13719
rect 18420 13483 18656 13719
rect 18742 13483 18978 13719
rect 19064 13483 19300 13719
rect 19386 13483 19622 13719
rect 19708 13483 19944 13719
rect 20030 13483 20266 13719
rect 20352 13483 20588 13719
rect 20674 13483 20910 13719
rect 20996 13483 21232 13719
rect 21318 13483 21554 13719
rect 21640 13483 21876 13719
rect 21962 13483 22198 13719
rect 22284 13483 22520 13719
rect 22606 13483 22842 13719
rect 22928 13483 23164 13719
rect 23250 13483 23486 13719
rect 23572 13483 23808 13719
rect 23894 13483 24130 13719
rect 24216 13483 24452 13719
rect -3185 12878 -2949 13114
rect -2862 12878 -2626 13114
rect -2539 12878 -2303 13114
rect -2216 12878 -1980 13114
rect -1893 12878 -1657 13114
rect -1570 12878 -1334 13114
rect -1247 12878 -1011 13114
rect -924 12878 -688 13114
rect -601 12878 -365 13114
rect -278 12878 -42 13114
rect 45 12878 281 13114
rect 368 12878 604 13114
rect 691 12878 927 13114
rect 1014 12878 1250 13114
rect 1337 12878 1573 13114
rect 1660 12878 1896 13114
rect 1983 12878 2219 13114
rect 2306 12878 2542 13114
rect 2629 12878 2865 13114
rect 2952 12878 3188 13114
rect 3275 12878 3511 13114
rect 3598 12878 3834 13114
rect 3921 12878 4157 13114
rect 4244 12878 4480 13114
rect 4567 12878 4803 13114
rect 4890 12878 5126 13114
rect 5213 12878 5449 13114
rect 5536 12878 5772 13114
rect 5859 12878 6095 13114
rect 6182 12878 6418 13114
rect 6504 12878 6740 13114
rect 6826 12878 7062 13114
rect 7148 12878 7384 13114
rect 7470 12878 7706 13114
rect 7792 12878 8028 13114
rect 8114 12878 8350 13114
rect 8436 12878 8672 13114
rect 8758 12878 8994 13114
rect 9080 12878 9316 13114
rect 9402 12878 9638 13114
rect 9724 12878 9960 13114
rect 10046 12878 10282 13114
rect 10368 12878 10604 13114
rect 10690 12878 10926 13114
rect 11012 12878 11248 13114
rect 11334 12878 11570 13114
rect 11656 12878 11892 13114
rect 11978 12878 12214 13114
rect 12300 12878 12536 13114
rect 12622 12878 12858 13114
rect 12944 12878 13180 13114
rect 13266 12878 13502 13114
rect 13588 12878 13824 13114
rect 13910 12878 14146 13114
rect 14232 12878 14468 13114
rect 14554 12878 14790 13114
rect 14876 12878 15112 13114
rect 15198 12878 15434 13114
rect 15520 12878 15756 13114
rect 15842 12878 16078 13114
rect 16164 12878 16400 13114
rect 16486 12878 16722 13114
rect 16808 12878 17044 13114
rect 17130 12878 17366 13114
rect 17452 12878 17688 13114
rect 17774 12878 18010 13114
rect 18096 12878 18332 13114
rect 18418 12878 18654 13114
rect 18740 12878 18976 13114
rect 19062 12878 19298 13114
rect 19384 12878 19620 13114
rect 19706 12878 19942 13114
rect 20028 12878 20264 13114
rect 20350 12878 20586 13114
rect 20672 12878 20908 13114
rect 20994 12878 21230 13114
rect 21316 12878 21552 13114
rect 21638 12878 21874 13114
rect 21960 12878 22196 13114
rect 22282 12878 22518 13114
rect 22604 12878 22840 13114
rect 22926 12878 23162 13114
rect 23248 12878 23484 13114
rect 23570 12878 23806 13114
rect 23892 12878 24128 13114
rect 24214 12878 24450 13114
rect -3185 12312 -2949 12548
rect -2862 12312 -2626 12548
rect -2539 12312 -2303 12548
rect -2216 12312 -1980 12548
rect -1893 12312 -1657 12548
rect -1570 12312 -1334 12548
rect -1247 12312 -1011 12548
rect -924 12312 -688 12548
rect -601 12312 -365 12548
rect -278 12312 -42 12548
rect 45 12312 281 12548
rect 368 12312 604 12548
rect 691 12312 927 12548
rect 1014 12312 1250 12548
rect 1337 12312 1573 12548
rect 1660 12312 1896 12548
rect 1983 12312 2219 12548
rect 2306 12312 2542 12548
rect 2629 12312 2865 12548
rect 2952 12312 3188 12548
rect 3275 12312 3511 12548
rect 3598 12312 3834 12548
rect 3921 12312 4157 12548
rect 4244 12312 4480 12548
rect 4567 12312 4803 12548
rect 4890 12312 5126 12548
rect 5213 12312 5449 12548
rect 5536 12312 5772 12548
rect 5859 12312 6095 12548
rect 6182 12312 6418 12548
rect 6504 12312 6740 12548
rect 6826 12312 7062 12548
rect 7148 12312 7384 12548
rect 7470 12312 7706 12548
rect 7792 12312 8028 12548
rect 8114 12312 8350 12548
rect 8436 12312 8672 12548
rect 8758 12312 8994 12548
rect 9080 12312 9316 12548
rect 9402 12312 9638 12548
rect 9724 12312 9960 12548
rect 10046 12312 10282 12548
rect 10368 12312 10604 12548
rect 10690 12312 10926 12548
rect 11012 12312 11248 12548
rect 11334 12312 11570 12548
rect 11656 12312 11892 12548
rect 11978 12312 12214 12548
rect 12300 12312 12536 12548
rect 12622 12312 12858 12548
rect 12944 12312 13180 12548
rect 13266 12312 13502 12548
rect 13588 12312 13824 12548
rect 13910 12312 14146 12548
rect 14232 12312 14468 12548
rect 14554 12312 14790 12548
rect 14876 12312 15112 12548
rect 15198 12312 15434 12548
rect 15520 12312 15756 12548
rect 15842 12312 16078 12548
rect 16164 12312 16400 12548
rect 16486 12312 16722 12548
rect 16808 12312 17044 12548
rect 17130 12312 17366 12548
rect 17452 12312 17688 12548
rect 17774 12312 18010 12548
rect 18096 12312 18332 12548
rect 18418 12312 18654 12548
rect 18740 12312 18976 12548
rect 19062 12312 19298 12548
rect 19384 12312 19620 12548
rect 19706 12312 19942 12548
rect 20028 12312 20264 12548
rect 20350 12312 20586 12548
rect 20672 12312 20908 12548
rect 20994 12312 21230 12548
rect 21316 12312 21552 12548
rect 21638 12312 21874 12548
rect 21960 12312 22196 12548
rect 22282 12312 22518 12548
rect 22604 12312 22840 12548
rect 22926 12312 23162 12548
rect 23248 12312 23484 12548
rect 23570 12312 23806 12548
rect 23892 12312 24128 12548
rect 24214 12312 24450 12548
rect -3185 11708 -2949 11944
rect -2862 11708 -2626 11944
rect -2539 11708 -2303 11944
rect -2216 11708 -1980 11944
rect -1893 11708 -1657 11944
rect -1570 11708 -1334 11944
rect -1247 11708 -1011 11944
rect -924 11708 -688 11944
rect -601 11708 -365 11944
rect -278 11708 -42 11944
rect 45 11708 281 11944
rect 368 11708 604 11944
rect 691 11708 927 11944
rect 1014 11708 1250 11944
rect 1337 11708 1573 11944
rect 1660 11708 1896 11944
rect 1983 11708 2219 11944
rect 2306 11708 2542 11944
rect 2629 11708 2865 11944
rect 2952 11708 3188 11944
rect 3275 11708 3511 11944
rect 3598 11708 3834 11944
rect 3921 11708 4157 11944
rect 4244 11708 4480 11944
rect 4567 11708 4803 11944
rect 4890 11708 5126 11944
rect 5213 11708 5449 11944
rect 5536 11708 5772 11944
rect 5859 11708 6095 11944
rect 6182 11708 6418 11944
rect 6504 11708 6740 11944
rect 6826 11708 7062 11944
rect 7148 11708 7384 11944
rect 7470 11708 7706 11944
rect 7792 11708 8028 11944
rect 8114 11708 8350 11944
rect 8436 11708 8672 11944
rect 8758 11708 8994 11944
rect 9080 11708 9316 11944
rect 9402 11708 9638 11944
rect 9724 11708 9960 11944
rect 10046 11708 10282 11944
rect 10368 11708 10604 11944
rect 10690 11708 10926 11944
rect 11012 11708 11248 11944
rect 11334 11708 11570 11944
rect 11656 11708 11892 11944
rect 11978 11708 12214 11944
rect 12300 11708 12536 11944
rect 12622 11708 12858 11944
rect 12944 11708 13180 11944
rect 13266 11708 13502 11944
rect 13588 11708 13824 11944
rect 13910 11708 14146 11944
rect 14232 11708 14468 11944
rect 14554 11708 14790 11944
rect 14876 11708 15112 11944
rect 15198 11708 15434 11944
rect 15520 11708 15756 11944
rect 15842 11708 16078 11944
rect 16164 11708 16400 11944
rect 16486 11708 16722 11944
rect 16808 11708 17044 11944
rect 17130 11708 17366 11944
rect 17452 11708 17688 11944
rect 17774 11708 18010 11944
rect 18096 11708 18332 11944
rect 18418 11708 18654 11944
rect 18740 11708 18976 11944
rect 19062 11708 19298 11944
rect 19384 11708 19620 11944
rect 19706 11708 19942 11944
rect 20028 11708 20264 11944
rect 20350 11708 20586 11944
rect 20672 11708 20908 11944
rect 20994 11708 21230 11944
rect 21316 11708 21552 11944
rect 21638 11708 21874 11944
rect 21960 11708 22196 11944
rect 22282 11708 22518 11944
rect 22604 11708 22840 11944
rect 22926 11708 23162 11944
rect 23248 11708 23484 11944
rect 23570 11708 23806 11944
rect 23892 11708 24128 11944
rect 24214 11708 24450 11944
rect -3185 11142 -2949 11378
rect -2862 11142 -2626 11378
rect -2539 11142 -2303 11378
rect -2216 11142 -1980 11378
rect -1893 11142 -1657 11378
rect -1570 11142 -1334 11378
rect -1247 11142 -1011 11378
rect -924 11142 -688 11378
rect -601 11142 -365 11378
rect -278 11142 -42 11378
rect 45 11142 281 11378
rect 368 11142 604 11378
rect 691 11142 927 11378
rect 1014 11142 1250 11378
rect 1337 11142 1573 11378
rect 1660 11142 1896 11378
rect 1983 11142 2219 11378
rect 2306 11142 2542 11378
rect 2629 11142 2865 11378
rect 2952 11142 3188 11378
rect 3275 11142 3511 11378
rect 3598 11142 3834 11378
rect 3921 11142 4157 11378
rect 4244 11142 4480 11378
rect 4567 11142 4803 11378
rect 4890 11142 5126 11378
rect 5213 11142 5449 11378
rect 5536 11142 5772 11378
rect 5859 11142 6095 11378
rect 6182 11142 6418 11378
rect 6504 11142 6740 11378
rect 6826 11142 7062 11378
rect 7148 11142 7384 11378
rect 7470 11142 7706 11378
rect 7792 11142 8028 11378
rect 8114 11142 8350 11378
rect 8436 11142 8672 11378
rect 8758 11142 8994 11378
rect 9080 11142 9316 11378
rect 9402 11142 9638 11378
rect 9724 11142 9960 11378
rect 10046 11142 10282 11378
rect 10368 11142 10604 11378
rect 10690 11142 10926 11378
rect 11012 11142 11248 11378
rect 11334 11142 11570 11378
rect 11656 11142 11892 11378
rect 11978 11142 12214 11378
rect 12300 11142 12536 11378
rect 12622 11142 12858 11378
rect 12944 11142 13180 11378
rect 13266 11142 13502 11378
rect 13588 11142 13824 11378
rect 13910 11142 14146 11378
rect 14232 11142 14468 11378
rect 14554 11142 14790 11378
rect 14876 11142 15112 11378
rect 15198 11142 15434 11378
rect 15520 11142 15756 11378
rect 15842 11142 16078 11378
rect 16164 11142 16400 11378
rect 16486 11142 16722 11378
rect 16808 11142 17044 11378
rect 17130 11142 17366 11378
rect 17452 11142 17688 11378
rect 17774 11142 18010 11378
rect 18096 11142 18332 11378
rect 18418 11142 18654 11378
rect 18740 11142 18976 11378
rect 19062 11142 19298 11378
rect 19384 11142 19620 11378
rect 19706 11142 19942 11378
rect 20028 11142 20264 11378
rect 20350 11142 20586 11378
rect 20672 11142 20908 11378
rect 20994 11142 21230 11378
rect 21316 11142 21552 11378
rect 21638 11142 21874 11378
rect 21960 11142 22196 11378
rect 22282 11142 22518 11378
rect 22604 11142 22840 11378
rect 22926 11142 23162 11378
rect 23248 11142 23484 11378
rect 23570 11142 23806 11378
rect 23892 11142 24128 11378
rect 24214 11142 24450 11378
rect -3185 8418 -2949 8654
rect -2862 8418 -2626 8654
rect -2539 8418 -2303 8654
rect -2216 8418 -1980 8654
rect -1893 8418 -1657 8654
rect -1570 8418 -1334 8654
rect -1247 8418 -1011 8654
rect -924 8418 -688 8654
rect -601 8418 -365 8654
rect -278 8418 -42 8654
rect 45 8418 281 8654
rect 368 8418 604 8654
rect 691 8418 927 8654
rect 1014 8418 1250 8654
rect 1337 8418 1573 8654
rect 1660 8418 1896 8654
rect 1983 8418 2219 8654
rect 2306 8418 2542 8654
rect 2629 8418 2865 8654
rect 2952 8418 3188 8654
rect 3275 8418 3511 8654
rect 3598 8418 3834 8654
rect 3921 8418 4157 8654
rect 4244 8418 4480 8654
rect 4567 8418 4803 8654
rect 4890 8418 5126 8654
rect 5213 8418 5449 8654
rect 5536 8418 5772 8654
rect 5859 8418 6095 8654
rect 6182 8418 6418 8654
rect 6505 8418 6741 8654
rect 6828 8418 7064 8654
rect 7150 8418 7386 8654
rect 7472 8418 7708 8654
rect 7794 8418 8030 8654
rect 8116 8418 8352 8654
rect 8438 8418 8674 8654
rect 8760 8418 8996 8654
rect 9082 8418 9318 8654
rect 9404 8418 9640 8654
rect 9726 8418 9962 8654
rect 10048 8418 10284 8654
rect 10370 8418 10606 8654
rect 10692 8418 10928 8654
rect 11014 8418 11250 8654
rect 11336 8418 11572 8654
rect 11658 8418 11894 8654
rect 11980 8418 12216 8654
rect 12302 8418 12538 8654
rect 12624 8418 12860 8654
rect 12946 8418 13182 8654
rect 13268 8418 13504 8654
rect 13590 8418 13826 8654
rect 13912 8418 14148 8654
rect 14234 8418 14470 8654
rect 14556 8418 14792 8654
rect 14878 8418 15114 8654
rect 15200 8418 15436 8654
rect 15522 8418 15758 8654
rect 15844 8418 16080 8654
rect 16166 8418 16402 8654
rect 16488 8418 16724 8654
rect 16810 8418 17046 8654
rect 17132 8418 17368 8654
rect 17454 8418 17690 8654
rect 17776 8418 18012 8654
rect 18098 8418 18334 8654
rect 18420 8418 18656 8654
rect 18742 8418 18978 8654
rect 19064 8418 19300 8654
rect 19386 8418 19622 8654
rect 19708 8418 19944 8654
rect 20030 8418 20266 8654
rect 20352 8418 20588 8654
rect 20674 8418 20910 8654
rect 20996 8418 21232 8654
rect 21318 8418 21554 8654
rect 21640 8418 21876 8654
rect 21962 8418 22198 8654
rect 22284 8418 22520 8654
rect 22606 8418 22842 8654
rect 22928 8418 23164 8654
rect 23250 8418 23486 8654
rect 23572 8418 23808 8654
rect 23894 8418 24130 8654
rect 24216 8418 24452 8654
rect -3185 7812 -2949 8048
rect -2862 7812 -2626 8048
rect -2539 7812 -2303 8048
rect -2216 7812 -1980 8048
rect -1893 7812 -1657 8048
rect -1570 7812 -1334 8048
rect -1247 7812 -1011 8048
rect -924 7812 -688 8048
rect -601 7812 -365 8048
rect -278 7812 -42 8048
rect 45 7812 281 8048
rect 368 7812 604 8048
rect 691 7812 927 8048
rect 1014 7812 1250 8048
rect 1337 7812 1573 8048
rect 1660 7812 1896 8048
rect 1983 7812 2219 8048
rect 2306 7812 2542 8048
rect 2629 7812 2865 8048
rect 2952 7812 3188 8048
rect 3275 7812 3511 8048
rect 3598 7812 3834 8048
rect 3921 7812 4157 8048
rect 4244 7812 4480 8048
rect 4567 7812 4803 8048
rect 4890 7812 5126 8048
rect 5213 7812 5449 8048
rect 5536 7812 5772 8048
rect 5859 7812 6095 8048
rect 6182 7812 6418 8048
rect 6505 7812 6741 8048
rect 6828 7812 7064 8048
rect 7150 7812 7386 8048
rect 7472 7812 7708 8048
rect 7794 7812 8030 8048
rect 8116 7812 8352 8048
rect 8438 7812 8674 8048
rect 8760 7812 8996 8048
rect 9082 7812 9318 8048
rect 9404 7812 9640 8048
rect 9726 7812 9962 8048
rect 10048 7812 10284 8048
rect 10370 7812 10606 8048
rect 10692 7812 10928 8048
rect 11014 7812 11250 8048
rect 11336 7812 11572 8048
rect 11658 7812 11894 8048
rect 11980 7812 12216 8048
rect 12302 7812 12538 8048
rect 12624 7812 12860 8048
rect 12946 7812 13182 8048
rect 13268 7812 13504 8048
rect 13590 7812 13826 8048
rect 13912 7812 14148 8048
rect 14234 7812 14470 8048
rect 14556 7812 14792 8048
rect 14878 7812 15114 8048
rect 15200 7812 15436 8048
rect 15522 7812 15758 8048
rect 15844 7812 16080 8048
rect 16166 7812 16402 8048
rect 16488 7812 16724 8048
rect 16810 7812 17046 8048
rect 17132 7812 17368 8048
rect 17454 7812 17690 8048
rect 17776 7812 18012 8048
rect 18098 7812 18334 8048
rect 18420 7812 18656 8048
rect 18742 7812 18978 8048
rect 19064 7812 19300 8048
rect 19386 7812 19622 8048
rect 19708 7812 19944 8048
rect 20030 7812 20266 8048
rect 20352 7812 20588 8048
rect 20674 7812 20910 8048
rect 20996 7812 21232 8048
rect 21318 7812 21554 8048
rect 21640 7812 21876 8048
rect 21962 7812 22198 8048
rect 22284 7812 22520 8048
rect 22606 7812 22842 8048
rect 22928 7812 23164 8048
rect 23250 7812 23486 8048
rect 23572 7812 23808 8048
rect 23894 7812 24130 8048
rect 24216 7812 24452 8048
rect -3185 7208 -2949 7444
rect -2862 7208 -2626 7444
rect -2539 7208 -2303 7444
rect -2216 7208 -1980 7444
rect -1893 7208 -1657 7444
rect -1570 7208 -1334 7444
rect -1247 7208 -1011 7444
rect -924 7208 -688 7444
rect -601 7208 -365 7444
rect -278 7208 -42 7444
rect 45 7208 281 7444
rect 368 7208 604 7444
rect 691 7208 927 7444
rect 1014 7208 1250 7444
rect 1337 7208 1573 7444
rect 1660 7208 1896 7444
rect 1983 7208 2219 7444
rect 2306 7208 2542 7444
rect 2629 7208 2865 7444
rect 2952 7208 3188 7444
rect 3275 7208 3511 7444
rect 3598 7208 3834 7444
rect 3921 7208 4157 7444
rect 4244 7208 4480 7444
rect 4567 7208 4803 7444
rect 4890 7208 5126 7444
rect 5213 7208 5449 7444
rect 5536 7208 5772 7444
rect 5859 7208 6095 7444
rect 6182 7208 6418 7444
rect 6505 7208 6741 7444
rect 6828 7208 7064 7444
rect 7150 7208 7386 7444
rect 7472 7208 7708 7444
rect 7794 7208 8030 7444
rect 8116 7208 8352 7444
rect 8438 7208 8674 7444
rect 8760 7208 8996 7444
rect 9082 7208 9318 7444
rect 9404 7208 9640 7444
rect 9726 7208 9962 7444
rect 10048 7208 10284 7444
rect 10370 7208 10606 7444
rect 10692 7208 10928 7444
rect 11014 7208 11250 7444
rect 11336 7208 11572 7444
rect 11658 7208 11894 7444
rect 11980 7208 12216 7444
rect 12302 7208 12538 7444
rect 12624 7208 12860 7444
rect 12946 7208 13182 7444
rect 13268 7208 13504 7444
rect 13590 7208 13826 7444
rect 13912 7208 14148 7444
rect 14234 7208 14470 7444
rect 14556 7208 14792 7444
rect 14878 7208 15114 7444
rect 15200 7208 15436 7444
rect 15522 7208 15758 7444
rect 15844 7208 16080 7444
rect 16166 7208 16402 7444
rect 16488 7208 16724 7444
rect 16810 7208 17046 7444
rect 17132 7208 17368 7444
rect 17454 7208 17690 7444
rect 17776 7208 18012 7444
rect 18098 7208 18334 7444
rect 18420 7208 18656 7444
rect 18742 7208 18978 7444
rect 19064 7208 19300 7444
rect 19386 7208 19622 7444
rect 19708 7208 19944 7444
rect 20030 7208 20266 7444
rect 20352 7208 20588 7444
rect 20674 7208 20910 7444
rect 20996 7208 21232 7444
rect 21318 7208 21554 7444
rect 21640 7208 21876 7444
rect 21962 7208 22198 7444
rect 22284 7208 22520 7444
rect 22606 7208 22842 7444
rect 22928 7208 23164 7444
rect 23250 7208 23486 7444
rect 23572 7208 23808 7444
rect 23894 7208 24130 7444
rect 24216 7208 24452 7444
rect -3185 6842 -2949 7078
rect -2862 6842 -2626 7078
rect -2539 6842 -2303 7078
rect -2216 6842 -1980 7078
rect -1893 6842 -1657 7078
rect -1570 6842 -1334 7078
rect -1247 6842 -1011 7078
rect -924 6842 -688 7078
rect -601 6842 -365 7078
rect -278 6842 -42 7078
rect 45 6842 281 7078
rect 368 6842 604 7078
rect 691 6842 927 7078
rect 1014 6842 1250 7078
rect 1337 6842 1573 7078
rect 1660 6842 1896 7078
rect 1983 6842 2219 7078
rect 2306 6842 2542 7078
rect 2629 6842 2865 7078
rect 2952 6842 3188 7078
rect 3275 6842 3511 7078
rect 3598 6842 3834 7078
rect 3921 6842 4157 7078
rect 4244 6842 4480 7078
rect 4567 6842 4803 7078
rect 4890 6842 5126 7078
rect 5213 6842 5449 7078
rect 5536 6842 5772 7078
rect 5859 6842 6095 7078
rect 6182 6842 6418 7078
rect 6505 6842 6741 7078
rect 6828 6842 7064 7078
rect 7150 6842 7386 7078
rect 7472 6842 7708 7078
rect 7794 6842 8030 7078
rect 8116 6842 8352 7078
rect 8438 6842 8674 7078
rect 8760 6842 8996 7078
rect 9082 6842 9318 7078
rect 9404 6842 9640 7078
rect 9726 6842 9962 7078
rect 10048 6842 10284 7078
rect 10370 6842 10606 7078
rect 10692 6842 10928 7078
rect 11014 6842 11250 7078
rect 11336 6842 11572 7078
rect 11658 6842 11894 7078
rect 11980 6842 12216 7078
rect 12302 6842 12538 7078
rect 12624 6842 12860 7078
rect 12946 6842 13182 7078
rect 13268 6842 13504 7078
rect 13590 6842 13826 7078
rect 13912 6842 14148 7078
rect 14234 6842 14470 7078
rect 14556 6842 14792 7078
rect 14878 6842 15114 7078
rect 15200 6842 15436 7078
rect 15522 6842 15758 7078
rect 15844 6842 16080 7078
rect 16166 6842 16402 7078
rect 16488 6842 16724 7078
rect 16810 6842 17046 7078
rect 17132 6842 17368 7078
rect 17454 6842 17690 7078
rect 17776 6842 18012 7078
rect 18098 6842 18334 7078
rect 18420 6842 18656 7078
rect 18742 6842 18978 7078
rect 19064 6842 19300 7078
rect 19386 6842 19622 7078
rect 19708 6842 19944 7078
rect 20030 6842 20266 7078
rect 20352 6842 20588 7078
rect 20674 6842 20910 7078
rect 20996 6842 21232 7078
rect 21318 6842 21554 7078
rect 21640 6842 21876 7078
rect 21962 6842 22198 7078
rect 22284 6842 22520 7078
rect 22606 6842 22842 7078
rect 22928 6842 23164 7078
rect 23250 6842 23486 7078
rect 23572 6842 23808 7078
rect 23894 6842 24130 7078
rect 24216 6842 24452 7078
rect -3185 6238 -2949 6474
rect -2862 6238 -2626 6474
rect -2539 6238 -2303 6474
rect -2216 6238 -1980 6474
rect -1893 6238 -1657 6474
rect -1570 6238 -1334 6474
rect -1247 6238 -1011 6474
rect -924 6238 -688 6474
rect -601 6238 -365 6474
rect -278 6238 -42 6474
rect 45 6238 281 6474
rect 368 6238 604 6474
rect 691 6238 927 6474
rect 1014 6238 1250 6474
rect 1337 6238 1573 6474
rect 1660 6238 1896 6474
rect 1983 6238 2219 6474
rect 2306 6238 2542 6474
rect 2629 6238 2865 6474
rect 2952 6238 3188 6474
rect 3275 6238 3511 6474
rect 3598 6238 3834 6474
rect 3921 6238 4157 6474
rect 4244 6238 4480 6474
rect 4567 6238 4803 6474
rect 4890 6238 5126 6474
rect 5213 6238 5449 6474
rect 5536 6238 5772 6474
rect 5859 6238 6095 6474
rect 6182 6238 6418 6474
rect 6505 6238 6741 6474
rect 6828 6238 7064 6474
rect 7150 6238 7386 6474
rect 7472 6238 7708 6474
rect 7794 6238 8030 6474
rect 8116 6238 8352 6474
rect 8438 6238 8674 6474
rect 8760 6238 8996 6474
rect 9082 6238 9318 6474
rect 9404 6238 9640 6474
rect 9726 6238 9962 6474
rect 10048 6238 10284 6474
rect 10370 6238 10606 6474
rect 10692 6238 10928 6474
rect 11014 6238 11250 6474
rect 11336 6238 11572 6474
rect 11658 6238 11894 6474
rect 11980 6238 12216 6474
rect 12302 6238 12538 6474
rect 12624 6238 12860 6474
rect 12946 6238 13182 6474
rect 13268 6238 13504 6474
rect 13590 6238 13826 6474
rect 13912 6238 14148 6474
rect 14234 6238 14470 6474
rect 14556 6238 14792 6474
rect 14878 6238 15114 6474
rect 15200 6238 15436 6474
rect 15522 6238 15758 6474
rect 15844 6238 16080 6474
rect 16166 6238 16402 6474
rect 16488 6238 16724 6474
rect 16810 6238 17046 6474
rect 17132 6238 17368 6474
rect 17454 6238 17690 6474
rect 17776 6238 18012 6474
rect 18098 6238 18334 6474
rect 18420 6238 18656 6474
rect 18742 6238 18978 6474
rect 19064 6238 19300 6474
rect 19386 6238 19622 6474
rect 19708 6238 19944 6474
rect 20030 6238 20266 6474
rect 20352 6238 20588 6474
rect 20674 6238 20910 6474
rect 20996 6238 21232 6474
rect 21318 6238 21554 6474
rect 21640 6238 21876 6474
rect 21962 6238 22198 6474
rect 22284 6238 22520 6474
rect 22606 6238 22842 6474
rect 22928 6238 23164 6474
rect 23250 6238 23486 6474
rect 23572 6238 23808 6474
rect 23894 6238 24130 6474
rect 24216 6238 24452 6474
rect -3185 5872 -2949 6108
rect -2862 5872 -2626 6108
rect -2539 5872 -2303 6108
rect -2216 5872 -1980 6108
rect -1893 5872 -1657 6108
rect -1570 5872 -1334 6108
rect -1247 5872 -1011 6108
rect -924 5872 -688 6108
rect -601 5872 -365 6108
rect -278 5872 -42 6108
rect 45 5872 281 6108
rect 368 5872 604 6108
rect 691 5872 927 6108
rect 1014 5872 1250 6108
rect 1337 5872 1573 6108
rect 1660 5872 1896 6108
rect 1983 5872 2219 6108
rect 2306 5872 2542 6108
rect 2629 5872 2865 6108
rect 2952 5872 3188 6108
rect 3275 5872 3511 6108
rect 3598 5872 3834 6108
rect 3921 5872 4157 6108
rect 4244 5872 4480 6108
rect 4567 5872 4803 6108
rect 4890 5872 5126 6108
rect 5213 5872 5449 6108
rect 5536 5872 5772 6108
rect 5859 5872 6095 6108
rect 6182 5872 6418 6108
rect 6505 5872 6741 6108
rect 6828 5872 7064 6108
rect 7150 5872 7386 6108
rect 7472 5872 7708 6108
rect 7794 5872 8030 6108
rect 8116 5872 8352 6108
rect 8438 5872 8674 6108
rect 8760 5872 8996 6108
rect 9082 5872 9318 6108
rect 9404 5872 9640 6108
rect 9726 5872 9962 6108
rect 10048 5872 10284 6108
rect 10370 5872 10606 6108
rect 10692 5872 10928 6108
rect 11014 5872 11250 6108
rect 11336 5872 11572 6108
rect 11658 5872 11894 6108
rect 11980 5872 12216 6108
rect 12302 5872 12538 6108
rect 12624 5872 12860 6108
rect 12946 5872 13182 6108
rect 13268 5872 13504 6108
rect 13590 5872 13826 6108
rect 13912 5872 14148 6108
rect 14234 5872 14470 6108
rect 14556 5872 14792 6108
rect 14878 5872 15114 6108
rect 15200 5872 15436 6108
rect 15522 5872 15758 6108
rect 15844 5872 16080 6108
rect 16166 5872 16402 6108
rect 16488 5872 16724 6108
rect 16810 5872 17046 6108
rect 17132 5872 17368 6108
rect 17454 5872 17690 6108
rect 17776 5872 18012 6108
rect 18098 5872 18334 6108
rect 18420 5872 18656 6108
rect 18742 5872 18978 6108
rect 19064 5872 19300 6108
rect 19386 5872 19622 6108
rect 19708 5872 19944 6108
rect 20030 5872 20266 6108
rect 20352 5872 20588 6108
rect 20674 5872 20910 6108
rect 20996 5872 21232 6108
rect 21318 5872 21554 6108
rect 21640 5872 21876 6108
rect 21962 5872 22198 6108
rect 22284 5872 22520 6108
rect 22606 5872 22842 6108
rect 22928 5872 23164 6108
rect 23250 5872 23486 6108
rect 23572 5872 23808 6108
rect 23894 5872 24130 6108
rect 24216 5872 24452 6108
rect -3185 5268 -2949 5504
rect -2862 5268 -2626 5504
rect -2539 5268 -2303 5504
rect -2216 5268 -1980 5504
rect -1893 5268 -1657 5504
rect -1570 5268 -1334 5504
rect -1247 5268 -1011 5504
rect -924 5268 -688 5504
rect -601 5268 -365 5504
rect -278 5268 -42 5504
rect 45 5268 281 5504
rect 368 5268 604 5504
rect 691 5268 927 5504
rect 1014 5268 1250 5504
rect 1337 5268 1573 5504
rect 1660 5268 1896 5504
rect 1983 5268 2219 5504
rect 2306 5268 2542 5504
rect 2629 5268 2865 5504
rect 2952 5268 3188 5504
rect 3275 5268 3511 5504
rect 3598 5268 3834 5504
rect 3921 5268 4157 5504
rect 4244 5268 4480 5504
rect 4567 5268 4803 5504
rect 4890 5268 5126 5504
rect 5213 5268 5449 5504
rect 5536 5268 5772 5504
rect 5859 5268 6095 5504
rect 6182 5268 6418 5504
rect 6505 5268 6741 5504
rect 6828 5268 7064 5504
rect 7150 5268 7386 5504
rect 7472 5268 7708 5504
rect 7794 5268 8030 5504
rect 8116 5268 8352 5504
rect 8438 5268 8674 5504
rect 8760 5268 8996 5504
rect 9082 5268 9318 5504
rect 9404 5268 9640 5504
rect 9726 5268 9962 5504
rect 10048 5268 10284 5504
rect 10370 5268 10606 5504
rect 10692 5268 10928 5504
rect 11014 5268 11250 5504
rect 11336 5268 11572 5504
rect 11658 5268 11894 5504
rect 11980 5268 12216 5504
rect 12302 5268 12538 5504
rect 12624 5268 12860 5504
rect 12946 5268 13182 5504
rect 13268 5268 13504 5504
rect 13590 5268 13826 5504
rect 13912 5268 14148 5504
rect 14234 5268 14470 5504
rect 14556 5268 14792 5504
rect 14878 5268 15114 5504
rect 15200 5268 15436 5504
rect 15522 5268 15758 5504
rect 15844 5268 16080 5504
rect 16166 5268 16402 5504
rect 16488 5268 16724 5504
rect 16810 5268 17046 5504
rect 17132 5268 17368 5504
rect 17454 5268 17690 5504
rect 17776 5268 18012 5504
rect 18098 5268 18334 5504
rect 18420 5268 18656 5504
rect 18742 5268 18978 5504
rect 19064 5268 19300 5504
rect 19386 5268 19622 5504
rect 19708 5268 19944 5504
rect 20030 5268 20266 5504
rect 20352 5268 20588 5504
rect 20674 5268 20910 5504
rect 20996 5268 21232 5504
rect 21318 5268 21554 5504
rect 21640 5268 21876 5504
rect 21962 5268 22198 5504
rect 22284 5268 22520 5504
rect 22606 5268 22842 5504
rect 22928 5268 23164 5504
rect 23250 5268 23486 5504
rect 23572 5268 23808 5504
rect 23894 5268 24130 5504
rect 24216 5268 24452 5504
rect -3185 4662 -2949 4898
rect -2862 4662 -2626 4898
rect -2539 4662 -2303 4898
rect -2216 4662 -1980 4898
rect -1893 4662 -1657 4898
rect -1570 4662 -1334 4898
rect -1247 4662 -1011 4898
rect -924 4662 -688 4898
rect -601 4662 -365 4898
rect -278 4662 -42 4898
rect 45 4662 281 4898
rect 368 4662 604 4898
rect 691 4662 927 4898
rect 1014 4662 1250 4898
rect 1337 4662 1573 4898
rect 1660 4662 1896 4898
rect 1983 4662 2219 4898
rect 2306 4662 2542 4898
rect 2629 4662 2865 4898
rect 2952 4662 3188 4898
rect 3275 4662 3511 4898
rect 3598 4662 3834 4898
rect 3921 4662 4157 4898
rect 4244 4662 4480 4898
rect 4567 4662 4803 4898
rect 4890 4662 5126 4898
rect 5213 4662 5449 4898
rect 5536 4662 5772 4898
rect 5859 4662 6095 4898
rect 6182 4662 6418 4898
rect 6505 4662 6741 4898
rect 6828 4662 7064 4898
rect 7150 4662 7386 4898
rect 7472 4662 7708 4898
rect 7794 4662 8030 4898
rect 8116 4662 8352 4898
rect 8438 4662 8674 4898
rect 8760 4662 8996 4898
rect 9082 4662 9318 4898
rect 9404 4662 9640 4898
rect 9726 4662 9962 4898
rect 10048 4662 10284 4898
rect 10370 4662 10606 4898
rect 10692 4662 10928 4898
rect 11014 4662 11250 4898
rect 11336 4662 11572 4898
rect 11658 4662 11894 4898
rect 11980 4662 12216 4898
rect 12302 4662 12538 4898
rect 12624 4662 12860 4898
rect 12946 4662 13182 4898
rect 13268 4662 13504 4898
rect 13590 4662 13826 4898
rect 13912 4662 14148 4898
rect 14234 4662 14470 4898
rect 14556 4662 14792 4898
rect 14878 4662 15114 4898
rect 15200 4662 15436 4898
rect 15522 4662 15758 4898
rect 15844 4662 16080 4898
rect 16166 4662 16402 4898
rect 16488 4662 16724 4898
rect 16810 4662 17046 4898
rect 17132 4662 17368 4898
rect 17454 4662 17690 4898
rect 17776 4662 18012 4898
rect 18098 4662 18334 4898
rect 18420 4662 18656 4898
rect 18742 4662 18978 4898
rect 19064 4662 19300 4898
rect 19386 4662 19622 4898
rect 19708 4662 19944 4898
rect 20030 4662 20266 4898
rect 20352 4662 20588 4898
rect 20674 4662 20910 4898
rect 20996 4662 21232 4898
rect 21318 4662 21554 4898
rect 21640 4662 21876 4898
rect 21962 4662 22198 4898
rect 22284 4662 22520 4898
rect 22606 4662 22842 4898
rect 22928 4662 23164 4898
rect 23250 4662 23486 4898
rect 23572 4662 23808 4898
rect 23894 4662 24130 4898
rect 24216 4662 24452 4898
rect -3185 4058 -2949 4294
rect -2862 4058 -2626 4294
rect -2539 4058 -2303 4294
rect -2216 4058 -1980 4294
rect -1893 4058 -1657 4294
rect -1570 4058 -1334 4294
rect -1247 4058 -1011 4294
rect -924 4058 -688 4294
rect -601 4058 -365 4294
rect -278 4058 -42 4294
rect 45 4058 281 4294
rect 368 4058 604 4294
rect 691 4058 927 4294
rect 1014 4058 1250 4294
rect 1337 4058 1573 4294
rect 1660 4058 1896 4294
rect 1983 4058 2219 4294
rect 2306 4058 2542 4294
rect 2629 4058 2865 4294
rect 2952 4058 3188 4294
rect 3275 4058 3511 4294
rect 3598 4058 3834 4294
rect 3921 4058 4157 4294
rect 4244 4058 4480 4294
rect 4567 4058 4803 4294
rect 4890 4058 5126 4294
rect 5213 4058 5449 4294
rect 5536 4058 5772 4294
rect 5859 4058 6095 4294
rect 6182 4058 6418 4294
rect 6505 4058 6741 4294
rect 6828 4058 7064 4294
rect 7150 4058 7386 4294
rect 7472 4058 7708 4294
rect 7794 4058 8030 4294
rect 8116 4058 8352 4294
rect 8438 4058 8674 4294
rect 8760 4058 8996 4294
rect 9082 4058 9318 4294
rect 9404 4058 9640 4294
rect 9726 4058 9962 4294
rect 10048 4058 10284 4294
rect 10370 4058 10606 4294
rect 10692 4058 10928 4294
rect 11014 4058 11250 4294
rect 11336 4058 11572 4294
rect 11658 4058 11894 4294
rect 11980 4058 12216 4294
rect 12302 4058 12538 4294
rect 12624 4058 12860 4294
rect 12946 4058 13182 4294
rect 13268 4058 13504 4294
rect 13590 4058 13826 4294
rect 13912 4058 14148 4294
rect 14234 4058 14470 4294
rect 14556 4058 14792 4294
rect 14878 4058 15114 4294
rect 15200 4058 15436 4294
rect 15522 4058 15758 4294
rect 15844 4058 16080 4294
rect 16166 4058 16402 4294
rect 16488 4058 16724 4294
rect 16810 4058 17046 4294
rect 17132 4058 17368 4294
rect 17454 4058 17690 4294
rect 17776 4058 18012 4294
rect 18098 4058 18334 4294
rect 18420 4058 18656 4294
rect 18742 4058 18978 4294
rect 19064 4058 19300 4294
rect 19386 4058 19622 4294
rect 19708 4058 19944 4294
rect 20030 4058 20266 4294
rect 20352 4058 20588 4294
rect 20674 4058 20910 4294
rect 20996 4058 21232 4294
rect 21318 4058 21554 4294
rect 21640 4058 21876 4294
rect 21962 4058 22198 4294
rect 22284 4058 22520 4294
rect 22606 4058 22842 4294
rect 22928 4058 23164 4294
rect 23250 4058 23486 4294
rect 23572 4058 23808 4294
rect 23894 4058 24130 4294
rect 24216 4058 24452 4294
rect -3185 3452 -2949 3688
rect -2862 3452 -2626 3688
rect -2539 3452 -2303 3688
rect -2216 3452 -1980 3688
rect -1893 3452 -1657 3688
rect -1570 3452 -1334 3688
rect -1247 3452 -1011 3688
rect -924 3452 -688 3688
rect -601 3452 -365 3688
rect -278 3452 -42 3688
rect 45 3452 281 3688
rect 368 3452 604 3688
rect 691 3452 927 3688
rect 1014 3452 1250 3688
rect 1337 3452 1573 3688
rect 1660 3452 1896 3688
rect 1983 3452 2219 3688
rect 2306 3452 2542 3688
rect 2629 3452 2865 3688
rect 2952 3452 3188 3688
rect 3275 3452 3511 3688
rect 3598 3452 3834 3688
rect 3921 3452 4157 3688
rect 4244 3452 4480 3688
rect 4567 3452 4803 3688
rect 4890 3452 5126 3688
rect 5213 3452 5449 3688
rect 5536 3452 5772 3688
rect 5859 3452 6095 3688
rect 6182 3452 6418 3688
rect 6505 3452 6741 3688
rect 6828 3452 7064 3688
rect 7150 3452 7386 3688
rect 7472 3452 7708 3688
rect 7794 3452 8030 3688
rect 8116 3452 8352 3688
rect 8438 3452 8674 3688
rect 8760 3452 8996 3688
rect 9082 3452 9318 3688
rect 9404 3452 9640 3688
rect 9726 3452 9962 3688
rect 10048 3452 10284 3688
rect 10370 3452 10606 3688
rect 10692 3452 10928 3688
rect 11014 3452 11250 3688
rect 11336 3452 11572 3688
rect 11658 3452 11894 3688
rect 11980 3452 12216 3688
rect 12302 3452 12538 3688
rect 12624 3452 12860 3688
rect 12946 3452 13182 3688
rect 13268 3452 13504 3688
rect 13590 3452 13826 3688
rect 13912 3452 14148 3688
rect 14234 3452 14470 3688
rect 14556 3452 14792 3688
rect 14878 3452 15114 3688
rect 15200 3452 15436 3688
rect 15522 3452 15758 3688
rect 15844 3452 16080 3688
rect 16166 3452 16402 3688
rect 16488 3452 16724 3688
rect 16810 3452 17046 3688
rect 17132 3452 17368 3688
rect 17454 3452 17690 3688
rect 17776 3452 18012 3688
rect 18098 3452 18334 3688
rect 18420 3452 18656 3688
rect 18742 3452 18978 3688
rect 19064 3452 19300 3688
rect 19386 3452 19622 3688
rect 19708 3452 19944 3688
rect 20030 3452 20266 3688
rect 20352 3452 20588 3688
rect 20674 3452 20910 3688
rect 20996 3452 21232 3688
rect 21318 3452 21554 3688
rect 21640 3452 21876 3688
rect 21962 3452 22198 3688
rect 22284 3452 22520 3688
rect 22606 3452 22842 3688
rect 22928 3452 23164 3688
rect 23250 3452 23486 3688
rect 23572 3452 23808 3688
rect 23894 3452 24130 3688
rect 24216 3452 24452 3688
rect -3185 2848 -2949 3084
rect -2862 2848 -2626 3084
rect -2539 2848 -2303 3084
rect -2216 2848 -1980 3084
rect -1893 2848 -1657 3084
rect -1570 2848 -1334 3084
rect -1247 2848 -1011 3084
rect -924 2848 -688 3084
rect -601 2848 -365 3084
rect -278 2848 -42 3084
rect 45 2848 281 3084
rect 368 2848 604 3084
rect 691 2848 927 3084
rect 1014 2848 1250 3084
rect 1337 2848 1573 3084
rect 1660 2848 1896 3084
rect 1983 2848 2219 3084
rect 2306 2848 2542 3084
rect 2629 2848 2865 3084
rect 2952 2848 3188 3084
rect 3275 2848 3511 3084
rect 3598 2848 3834 3084
rect 3921 2848 4157 3084
rect 4244 2848 4480 3084
rect 4567 2848 4803 3084
rect 4890 2848 5126 3084
rect 5213 2848 5449 3084
rect 5536 2848 5772 3084
rect 5859 2848 6095 3084
rect 6182 2848 6418 3084
rect 6505 2848 6741 3084
rect 6828 2848 7064 3084
rect 7150 2848 7386 3084
rect 7472 2848 7708 3084
rect 7794 2848 8030 3084
rect 8116 2848 8352 3084
rect 8438 2848 8674 3084
rect 8760 2848 8996 3084
rect 9082 2848 9318 3084
rect 9404 2848 9640 3084
rect 9726 2848 9962 3084
rect 10048 2848 10284 3084
rect 10370 2848 10606 3084
rect 10692 2848 10928 3084
rect 11014 2848 11250 3084
rect 11336 2848 11572 3084
rect 11658 2848 11894 3084
rect 11980 2848 12216 3084
rect 12302 2848 12538 3084
rect 12624 2848 12860 3084
rect 12946 2848 13182 3084
rect 13268 2848 13504 3084
rect 13590 2848 13826 3084
rect 13912 2848 14148 3084
rect 14234 2848 14470 3084
rect 14556 2848 14792 3084
rect 14878 2848 15114 3084
rect 15200 2848 15436 3084
rect 15522 2848 15758 3084
rect 15844 2848 16080 3084
rect 16166 2848 16402 3084
rect 16488 2848 16724 3084
rect 16810 2848 17046 3084
rect 17132 2848 17368 3084
rect 17454 2848 17690 3084
rect 17776 2848 18012 3084
rect 18098 2848 18334 3084
rect 18420 2848 18656 3084
rect 18742 2848 18978 3084
rect 19064 2848 19300 3084
rect 19386 2848 19622 3084
rect 19708 2848 19944 3084
rect 20030 2848 20266 3084
rect 20352 2848 20588 3084
rect 20674 2848 20910 3084
rect 20996 2848 21232 3084
rect 21318 2848 21554 3084
rect 21640 2848 21876 3084
rect 21962 2848 22198 3084
rect 22284 2848 22520 3084
rect 22606 2848 22842 3084
rect 22928 2848 23164 3084
rect 23250 2848 23486 3084
rect 23572 2848 23808 3084
rect 23894 2848 24130 3084
rect 24216 2848 24452 3084
rect -3185 2482 -2949 2718
rect -2862 2482 -2626 2718
rect -2539 2482 -2303 2718
rect -2216 2482 -1980 2718
rect -1893 2482 -1657 2718
rect -1570 2482 -1334 2718
rect -1247 2482 -1011 2718
rect -924 2482 -688 2718
rect -601 2482 -365 2718
rect -278 2482 -42 2718
rect 45 2482 281 2718
rect 368 2482 604 2718
rect 691 2482 927 2718
rect 1014 2482 1250 2718
rect 1337 2482 1573 2718
rect 1660 2482 1896 2718
rect 1983 2482 2219 2718
rect 2306 2482 2542 2718
rect 2629 2482 2865 2718
rect 2952 2482 3188 2718
rect 3275 2482 3511 2718
rect 3598 2482 3834 2718
rect 3921 2482 4157 2718
rect 4244 2482 4480 2718
rect 4567 2482 4803 2718
rect 4890 2482 5126 2718
rect 5213 2482 5449 2718
rect 5536 2482 5772 2718
rect 5859 2482 6095 2718
rect 6182 2482 6418 2718
rect 6505 2482 6741 2718
rect 6828 2482 7064 2718
rect 7150 2482 7386 2718
rect 7472 2482 7708 2718
rect 7794 2482 8030 2718
rect 8116 2482 8352 2718
rect 8438 2482 8674 2718
rect 8760 2482 8996 2718
rect 9082 2482 9318 2718
rect 9404 2482 9640 2718
rect 9726 2482 9962 2718
rect 10048 2482 10284 2718
rect 10370 2482 10606 2718
rect 10692 2482 10928 2718
rect 11014 2482 11250 2718
rect 11336 2482 11572 2718
rect 11658 2482 11894 2718
rect 11980 2482 12216 2718
rect 12302 2482 12538 2718
rect 12624 2482 12860 2718
rect 12946 2482 13182 2718
rect 13268 2482 13504 2718
rect 13590 2482 13826 2718
rect 13912 2482 14148 2718
rect 14234 2482 14470 2718
rect 14556 2482 14792 2718
rect 14878 2482 15114 2718
rect 15200 2482 15436 2718
rect 15522 2482 15758 2718
rect 15844 2482 16080 2718
rect 16166 2482 16402 2718
rect 16488 2482 16724 2718
rect 16810 2482 17046 2718
rect 17132 2482 17368 2718
rect 17454 2482 17690 2718
rect 17776 2482 18012 2718
rect 18098 2482 18334 2718
rect 18420 2482 18656 2718
rect 18742 2482 18978 2718
rect 19064 2482 19300 2718
rect 19386 2482 19622 2718
rect 19708 2482 19944 2718
rect 20030 2482 20266 2718
rect 20352 2482 20588 2718
rect 20674 2482 20910 2718
rect 20996 2482 21232 2718
rect 21318 2482 21554 2718
rect 21640 2482 21876 2718
rect 21962 2482 22198 2718
rect 22284 2482 22520 2718
rect 22606 2482 22842 2718
rect 22928 2482 23164 2718
rect 23250 2482 23486 2718
rect 23572 2482 23808 2718
rect 23894 2482 24130 2718
rect 24216 2482 24452 2718
rect -3185 1878 -2949 2114
rect -2862 1878 -2626 2114
rect -2539 1878 -2303 2114
rect -2216 1878 -1980 2114
rect -1893 1878 -1657 2114
rect -1570 1878 -1334 2114
rect -1247 1878 -1011 2114
rect -924 1878 -688 2114
rect -601 1878 -365 2114
rect -278 1878 -42 2114
rect 45 1878 281 2114
rect 368 1878 604 2114
rect 691 1878 927 2114
rect 1014 1878 1250 2114
rect 1337 1878 1573 2114
rect 1660 1878 1896 2114
rect 1983 1878 2219 2114
rect 2306 1878 2542 2114
rect 2629 1878 2865 2114
rect 2952 1878 3188 2114
rect 3275 1878 3511 2114
rect 3598 1878 3834 2114
rect 3921 1878 4157 2114
rect 4244 1878 4480 2114
rect 4567 1878 4803 2114
rect 4890 1878 5126 2114
rect 5213 1878 5449 2114
rect 5536 1878 5772 2114
rect 5859 1878 6095 2114
rect 6182 1878 6418 2114
rect 6505 1878 6741 2114
rect 6828 1878 7064 2114
rect 7150 1878 7386 2114
rect 7472 1878 7708 2114
rect 7794 1878 8030 2114
rect 8116 1878 8352 2114
rect 8438 1878 8674 2114
rect 8760 1878 8996 2114
rect 9082 1878 9318 2114
rect 9404 1878 9640 2114
rect 9726 1878 9962 2114
rect 10048 1878 10284 2114
rect 10370 1878 10606 2114
rect 10692 1878 10928 2114
rect 11014 1878 11250 2114
rect 11336 1878 11572 2114
rect 11658 1878 11894 2114
rect 11980 1878 12216 2114
rect 12302 1878 12538 2114
rect 12624 1878 12860 2114
rect 12946 1878 13182 2114
rect 13268 1878 13504 2114
rect 13590 1878 13826 2114
rect 13912 1878 14148 2114
rect 14234 1878 14470 2114
rect 14556 1878 14792 2114
rect 14878 1878 15114 2114
rect 15200 1878 15436 2114
rect 15522 1878 15758 2114
rect 15844 1878 16080 2114
rect 16166 1878 16402 2114
rect 16488 1878 16724 2114
rect 16810 1878 17046 2114
rect 17132 1878 17368 2114
rect 17454 1878 17690 2114
rect 17776 1878 18012 2114
rect 18098 1878 18334 2114
rect 18420 1878 18656 2114
rect 18742 1878 18978 2114
rect 19064 1878 19300 2114
rect 19386 1878 19622 2114
rect 19708 1878 19944 2114
rect 20030 1878 20266 2114
rect 20352 1878 20588 2114
rect 20674 1878 20910 2114
rect 20996 1878 21232 2114
rect 21318 1878 21554 2114
rect 21640 1878 21876 2114
rect 21962 1878 22198 2114
rect 22284 1878 22520 2114
rect 22606 1878 22842 2114
rect 22928 1878 23164 2114
rect 23250 1878 23486 2114
rect 23572 1878 23808 2114
rect 23894 1878 24130 2114
rect 24216 1878 24452 2114
rect -3185 1272 -2949 1508
rect -2862 1272 -2626 1508
rect -2539 1272 -2303 1508
rect -2216 1272 -1980 1508
rect -1893 1272 -1657 1508
rect -1570 1272 -1334 1508
rect -1247 1272 -1011 1508
rect -924 1272 -688 1508
rect -601 1272 -365 1508
rect -278 1272 -42 1508
rect 45 1272 281 1508
rect 368 1272 604 1508
rect 691 1272 927 1508
rect 1014 1272 1250 1508
rect 1337 1272 1573 1508
rect 1660 1272 1896 1508
rect 1983 1272 2219 1508
rect 2306 1272 2542 1508
rect 2629 1272 2865 1508
rect 2952 1272 3188 1508
rect 3275 1272 3511 1508
rect 3598 1272 3834 1508
rect 3921 1272 4157 1508
rect 4244 1272 4480 1508
rect 4567 1272 4803 1508
rect 4890 1272 5126 1508
rect 5213 1272 5449 1508
rect 5536 1272 5772 1508
rect 5859 1272 6095 1508
rect 6182 1272 6418 1508
rect 6505 1272 6741 1508
rect 6828 1272 7064 1508
rect 7150 1272 7386 1508
rect 7472 1272 7708 1508
rect 7794 1272 8030 1508
rect 8116 1272 8352 1508
rect 8438 1272 8674 1508
rect 8760 1272 8996 1508
rect 9082 1272 9318 1508
rect 9404 1272 9640 1508
rect 9726 1272 9962 1508
rect 10048 1272 10284 1508
rect 10370 1272 10606 1508
rect 10692 1272 10928 1508
rect 11014 1272 11250 1508
rect 11336 1272 11572 1508
rect 11658 1272 11894 1508
rect 11980 1272 12216 1508
rect 12302 1272 12538 1508
rect 12624 1272 12860 1508
rect 12946 1272 13182 1508
rect 13268 1272 13504 1508
rect 13590 1272 13826 1508
rect 13912 1272 14148 1508
rect 14234 1272 14470 1508
rect 14556 1272 14792 1508
rect 14878 1272 15114 1508
rect 15200 1272 15436 1508
rect 15522 1272 15758 1508
rect 15844 1272 16080 1508
rect 16166 1272 16402 1508
rect 16488 1272 16724 1508
rect 16810 1272 17046 1508
rect 17132 1272 17368 1508
rect 17454 1272 17690 1508
rect 17776 1272 18012 1508
rect 18098 1272 18334 1508
rect 18420 1272 18656 1508
rect 18742 1272 18978 1508
rect 19064 1272 19300 1508
rect 19386 1272 19622 1508
rect 19708 1272 19944 1508
rect 20030 1272 20266 1508
rect 20352 1272 20588 1508
rect 20674 1272 20910 1508
rect 20996 1272 21232 1508
rect 21318 1272 21554 1508
rect 21640 1272 21876 1508
rect 21962 1272 22198 1508
rect 22284 1272 22520 1508
rect 22606 1272 22842 1508
rect 22928 1272 23164 1508
rect 23250 1272 23486 1508
rect 23572 1272 23808 1508
rect 23894 1272 24130 1508
rect 24216 1272 24452 1508
rect -3185 667 -2949 903
rect -2862 667 -2626 903
rect -2539 667 -2303 903
rect -2216 667 -1980 903
rect -1893 667 -1657 903
rect -1570 667 -1334 903
rect -1247 667 -1011 903
rect -924 667 -688 903
rect -601 667 -365 903
rect -278 667 -42 903
rect 45 667 281 903
rect 368 667 604 903
rect 691 667 927 903
rect 1014 667 1250 903
rect 1337 667 1573 903
rect 1660 667 1896 903
rect 1983 667 2219 903
rect 2306 667 2542 903
rect 2629 667 2865 903
rect 2952 667 3188 903
rect 3275 667 3511 903
rect 3598 667 3834 903
rect 3921 667 4157 903
rect 4244 667 4480 903
rect 4567 667 4803 903
rect 4890 667 5126 903
rect 5213 667 5449 903
rect 5536 667 5772 903
rect 5859 667 6095 903
rect 6182 667 6418 903
rect 6505 667 6741 903
rect 6828 667 7064 903
rect 7150 667 7386 903
rect 7472 667 7708 903
rect 7794 667 8030 903
rect 8116 667 8352 903
rect 8438 667 8674 903
rect 8760 667 8996 903
rect 9082 667 9318 903
rect 9404 667 9640 903
rect 9726 667 9962 903
rect 10048 667 10284 903
rect 10370 667 10606 903
rect 10692 667 10928 903
rect 11014 667 11250 903
rect 11336 667 11572 903
rect 11658 667 11894 903
rect 11980 667 12216 903
rect 12302 667 12538 903
rect 12624 667 12860 903
rect 12946 667 13182 903
rect 13268 667 13504 903
rect 13590 667 13826 903
rect 13912 667 14148 903
rect 14234 667 14470 903
rect 14556 667 14792 903
rect 14878 667 15114 903
rect 15200 667 15436 903
rect 15522 667 15758 903
rect 15844 667 16080 903
rect 16166 667 16402 903
rect 16488 667 16724 903
rect 16810 667 17046 903
rect 17132 667 17368 903
rect 17454 667 17690 903
rect 17776 667 18012 903
rect 18098 667 18334 903
rect 18420 667 18656 903
rect 18742 667 18978 903
rect 19064 667 19300 903
rect 19386 667 19622 903
rect 19708 667 19944 903
rect 20030 667 20266 903
rect 20352 667 20588 903
rect 20674 667 20910 903
rect 20996 667 21232 903
rect 21318 667 21554 903
rect 21640 667 21876 903
rect 21962 667 22198 903
rect 22284 667 22520 903
rect 22606 667 22842 903
rect 22928 667 23164 903
rect 23250 667 23486 903
rect 23572 667 23808 903
rect 23894 667 24130 903
rect 24216 667 24452 903
rect -3185 285 -2949 521
rect -2862 285 -2626 521
rect -2539 285 -2303 521
rect -2216 285 -1980 521
rect -1893 285 -1657 521
rect -1570 285 -1334 521
rect -1247 285 -1011 521
rect -924 285 -688 521
rect -601 285 -365 521
rect -278 285 -42 521
rect 45 285 281 521
rect 368 285 604 521
rect 691 285 927 521
rect 1014 285 1250 521
rect 1337 285 1573 521
rect 1660 285 1896 521
rect 1983 285 2219 521
rect 2306 285 2542 521
rect 2629 285 2865 521
rect 2952 285 3188 521
rect 3275 285 3511 521
rect 3598 285 3834 521
rect 3921 285 4157 521
rect 4244 285 4480 521
rect 4567 285 4803 521
rect 4890 285 5126 521
rect 5213 285 5449 521
rect 5536 285 5772 521
rect 5859 285 6095 521
rect 6182 285 6418 521
rect 6505 285 6741 521
rect 6828 285 7064 521
rect 7150 285 7386 521
rect 7472 285 7708 521
rect 7794 285 8030 521
rect 8116 285 8352 521
rect 8438 285 8674 521
rect 8760 285 8996 521
rect 9082 285 9318 521
rect 9404 285 9640 521
rect 9726 285 9962 521
rect 10048 285 10284 521
rect 10370 285 10606 521
rect 10692 285 10928 521
rect 11014 285 11250 521
rect 11336 285 11572 521
rect 11658 285 11894 521
rect 11980 285 12216 521
rect 12302 285 12538 521
rect 12624 285 12860 521
rect 12946 285 13182 521
rect 13268 285 13504 521
rect 13590 285 13826 521
rect 13912 285 14148 521
rect 14234 285 14470 521
rect 14556 285 14792 521
rect 14878 285 15114 521
rect 15200 285 15436 521
rect 15522 285 15758 521
rect 15844 285 16080 521
rect 16166 285 16402 521
rect 16488 285 16724 521
rect 16810 285 17046 521
rect 17132 285 17368 521
rect 17454 285 17690 521
rect 17776 285 18012 521
rect 18098 285 18334 521
rect 18420 285 18656 521
rect 18742 285 18978 521
rect 19064 285 19300 521
rect 19386 285 19622 521
rect 19708 285 19944 521
rect 20030 285 20266 521
rect 20352 285 20588 521
rect 20674 285 20910 521
rect 20996 285 21232 521
rect 21318 285 21554 521
rect 21640 285 21876 521
rect 21962 285 22198 521
rect 22284 285 22520 521
rect 22606 285 22842 521
rect 22928 285 23164 521
rect 23250 285 23486 521
rect 23572 285 23808 521
rect 23894 285 24130 521
rect 24216 285 24452 521
rect -3185 -97 -2949 139
rect -2862 -97 -2626 139
rect -2539 -97 -2303 139
rect -2216 -97 -1980 139
rect -1893 -97 -1657 139
rect -1570 -97 -1334 139
rect -1247 -97 -1011 139
rect -924 -97 -688 139
rect -601 -97 -365 139
rect -278 -97 -42 139
rect 45 -97 281 139
rect 368 -97 604 139
rect 691 -97 927 139
rect 1014 -97 1250 139
rect 1337 -97 1573 139
rect 1660 -97 1896 139
rect 1983 -97 2219 139
rect 2306 -97 2542 139
rect 2629 -97 2865 139
rect 2952 -97 3188 139
rect 3275 -97 3511 139
rect 3598 -97 3834 139
rect 3921 -97 4157 139
rect 4244 -97 4480 139
rect 4567 -97 4803 139
rect 4890 -97 5126 139
rect 5213 -97 5449 139
rect 5536 -97 5772 139
rect 5859 -97 6095 139
rect 6182 -97 6418 139
rect 6505 -97 6741 139
rect 6828 -97 7064 139
rect 7150 -97 7386 139
rect 7472 -97 7708 139
rect 7794 -97 8030 139
rect 8116 -97 8352 139
rect 8438 -97 8674 139
rect 8760 -97 8996 139
rect 9082 -97 9318 139
rect 9404 -97 9640 139
rect 9726 -97 9962 139
rect 10048 -97 10284 139
rect 10370 -97 10606 139
rect 10692 -97 10928 139
rect 11014 -97 11250 139
rect 11336 -97 11572 139
rect 11658 -97 11894 139
rect 11980 -97 12216 139
rect 12302 -97 12538 139
rect 12624 -97 12860 139
rect 12946 -97 13182 139
rect 13268 -97 13504 139
rect 13590 -97 13826 139
rect 13912 -97 14148 139
rect 14234 -97 14470 139
rect 14556 -97 14792 139
rect 14878 -97 15114 139
rect 15200 -97 15436 139
rect 15522 -97 15758 139
rect 15844 -97 16080 139
rect 16166 -97 16402 139
rect 16488 -97 16724 139
rect 16810 -97 17046 139
rect 17132 -97 17368 139
rect 17454 -97 17690 139
rect 17776 -97 18012 139
rect 18098 -97 18334 139
rect 18420 -97 18656 139
rect 18742 -97 18978 139
rect 19064 -97 19300 139
rect 19386 -97 19622 139
rect 19708 -97 19944 139
rect 20030 -97 20266 139
rect 20352 -97 20588 139
rect 20674 -97 20910 139
rect 20996 -97 21232 139
rect 21318 -97 21554 139
rect 21640 -97 21876 139
rect 21962 -97 22198 139
rect 22284 -97 22520 139
rect 22606 -97 22842 139
rect 22928 -97 23164 139
rect 23250 -97 23486 139
rect 23572 -97 23808 139
rect 23894 -97 24130 139
rect 24216 -97 24452 139
<< metal5 >>
rect -3360 39416 24640 39451
rect -3360 39180 -3087 39416
rect -2851 39180 -2765 39416
rect -2529 39180 -2443 39416
rect -2207 39180 -2121 39416
rect -1885 39180 -1799 39416
rect -1563 39180 -1477 39416
rect -1241 39180 -1155 39416
rect -919 39180 -833 39416
rect -597 39180 -511 39416
rect -275 39180 -189 39416
rect 47 39180 133 39416
rect 369 39180 455 39416
rect 691 39180 777 39416
rect 1013 39180 1099 39416
rect 1335 39180 1421 39416
rect 1657 39180 1743 39416
rect 1979 39180 2065 39416
rect 2301 39180 2387 39416
rect 2623 39180 2709 39416
rect 2945 39180 3031 39416
rect 3267 39180 3353 39416
rect 3589 39180 3675 39416
rect 3911 39180 3997 39416
rect 4233 39180 4318 39416
rect 4554 39180 4639 39416
rect 4875 39180 4960 39416
rect 5196 39180 5281 39416
rect 5517 39180 5602 39416
rect 5838 39180 5923 39416
rect 6159 39180 6244 39416
rect 6480 39180 6565 39416
rect 6801 39180 6886 39416
rect 7122 39180 7207 39416
rect 7443 39180 7528 39416
rect 7764 39180 7849 39416
rect 8085 39180 8170 39416
rect 8406 39180 8491 39416
rect 8727 39180 8812 39416
rect 9048 39180 9133 39416
rect 9369 39180 9454 39416
rect 9690 39180 9775 39416
rect 10011 39180 10096 39416
rect 10332 39180 10417 39416
rect 10653 39180 10738 39416
rect 10974 39180 11059 39416
rect 11295 39180 11380 39416
rect 11616 39180 11701 39416
rect 11937 39180 12022 39416
rect 12258 39180 12343 39416
rect 12579 39180 12664 39416
rect 12900 39180 12985 39416
rect 13221 39180 13306 39416
rect 13542 39180 13627 39416
rect 13863 39180 13948 39416
rect 14184 39180 14269 39416
rect 14505 39180 14590 39416
rect 14826 39180 14911 39416
rect 15147 39180 15232 39416
rect 15468 39180 15553 39416
rect 15789 39180 15874 39416
rect 16110 39180 16195 39416
rect 16431 39180 16516 39416
rect 16752 39180 16837 39416
rect 17073 39180 17158 39416
rect 17394 39180 17479 39416
rect 17715 39180 17800 39416
rect 18036 39180 18121 39416
rect 18357 39180 18442 39416
rect 18678 39180 18763 39416
rect 18999 39180 19084 39416
rect 19320 39180 19405 39416
rect 19641 39180 19726 39416
rect 19962 39180 20047 39416
rect 20283 39180 20368 39416
rect 20604 39180 20689 39416
rect 20925 39180 21010 39416
rect 21246 39180 21331 39416
rect 21567 39180 21652 39416
rect 21888 39180 21973 39416
rect 22209 39180 22294 39416
rect 22530 39180 22615 39416
rect 22851 39180 22936 39416
rect 23172 39180 23257 39416
rect 23493 39180 23578 39416
rect 23814 39180 23899 39416
rect 24135 39180 24220 39416
rect 24456 39180 24640 39416
rect -3360 39092 24640 39180
rect -3360 38856 -3087 39092
rect -2851 38856 -2765 39092
rect -2529 38856 -2443 39092
rect -2207 38856 -2121 39092
rect -1885 38856 -1799 39092
rect -1563 38856 -1477 39092
rect -1241 38856 -1155 39092
rect -919 38856 -833 39092
rect -597 38856 -511 39092
rect -275 38856 -189 39092
rect 47 38856 133 39092
rect 369 38856 455 39092
rect 691 38856 777 39092
rect 1013 38856 1099 39092
rect 1335 38856 1421 39092
rect 1657 38856 1743 39092
rect 1979 38856 2065 39092
rect 2301 38856 2387 39092
rect 2623 38856 2709 39092
rect 2945 38856 3031 39092
rect 3267 38856 3353 39092
rect 3589 38856 3675 39092
rect 3911 38856 3997 39092
rect 4233 38856 4318 39092
rect 4554 38856 4639 39092
rect 4875 38856 4960 39092
rect 5196 38856 5281 39092
rect 5517 38856 5602 39092
rect 5838 38856 5923 39092
rect 6159 38856 6244 39092
rect 6480 38856 6565 39092
rect 6801 38856 6886 39092
rect 7122 38856 7207 39092
rect 7443 38856 7528 39092
rect 7764 38856 7849 39092
rect 8085 38856 8170 39092
rect 8406 38856 8491 39092
rect 8727 38856 8812 39092
rect 9048 38856 9133 39092
rect 9369 38856 9454 39092
rect 9690 38856 9775 39092
rect 10011 38856 10096 39092
rect 10332 38856 10417 39092
rect 10653 38856 10738 39092
rect 10974 38856 11059 39092
rect 11295 38856 11380 39092
rect 11616 38856 11701 39092
rect 11937 38856 12022 39092
rect 12258 38856 12343 39092
rect 12579 38856 12664 39092
rect 12900 38856 12985 39092
rect 13221 38856 13306 39092
rect 13542 38856 13627 39092
rect 13863 38856 13948 39092
rect 14184 38856 14269 39092
rect 14505 38856 14590 39092
rect 14826 38856 14911 39092
rect 15147 38856 15232 39092
rect 15468 38856 15553 39092
rect 15789 38856 15874 39092
rect 16110 38856 16195 39092
rect 16431 38856 16516 39092
rect 16752 38856 16837 39092
rect 17073 38856 17158 39092
rect 17394 38856 17479 39092
rect 17715 38856 17800 39092
rect 18036 38856 18121 39092
rect 18357 38856 18442 39092
rect 18678 38856 18763 39092
rect 18999 38856 19084 39092
rect 19320 38856 19405 39092
rect 19641 38856 19726 39092
rect 19962 38856 20047 39092
rect 20283 38856 20368 39092
rect 20604 38856 20689 39092
rect 20925 38856 21010 39092
rect 21246 38856 21331 39092
rect 21567 38856 21652 39092
rect 21888 38856 21973 39092
rect 22209 38856 22294 39092
rect 22530 38856 22615 39092
rect 22851 38856 22936 39092
rect 23172 38856 23257 39092
rect 23493 38856 23578 39092
rect 23814 38856 23899 39092
rect 24135 38856 24220 39092
rect 24456 38856 24640 39092
rect -3360 38768 24640 38856
rect -3360 38532 -3087 38768
rect -2851 38532 -2765 38768
rect -2529 38532 -2443 38768
rect -2207 38532 -2121 38768
rect -1885 38532 -1799 38768
rect -1563 38532 -1477 38768
rect -1241 38532 -1155 38768
rect -919 38532 -833 38768
rect -597 38532 -511 38768
rect -275 38532 -189 38768
rect 47 38532 133 38768
rect 369 38532 455 38768
rect 691 38532 777 38768
rect 1013 38532 1099 38768
rect 1335 38532 1421 38768
rect 1657 38532 1743 38768
rect 1979 38532 2065 38768
rect 2301 38532 2387 38768
rect 2623 38532 2709 38768
rect 2945 38532 3031 38768
rect 3267 38532 3353 38768
rect 3589 38532 3675 38768
rect 3911 38532 3997 38768
rect 4233 38532 4318 38768
rect 4554 38532 4639 38768
rect 4875 38532 4960 38768
rect 5196 38532 5281 38768
rect 5517 38532 5602 38768
rect 5838 38532 5923 38768
rect 6159 38532 6244 38768
rect 6480 38532 6565 38768
rect 6801 38532 6886 38768
rect 7122 38532 7207 38768
rect 7443 38532 7528 38768
rect 7764 38532 7849 38768
rect 8085 38532 8170 38768
rect 8406 38532 8491 38768
rect 8727 38532 8812 38768
rect 9048 38532 9133 38768
rect 9369 38532 9454 38768
rect 9690 38532 9775 38768
rect 10011 38532 10096 38768
rect 10332 38532 10417 38768
rect 10653 38532 10738 38768
rect 10974 38532 11059 38768
rect 11295 38532 11380 38768
rect 11616 38532 11701 38768
rect 11937 38532 12022 38768
rect 12258 38532 12343 38768
rect 12579 38532 12664 38768
rect 12900 38532 12985 38768
rect 13221 38532 13306 38768
rect 13542 38532 13627 38768
rect 13863 38532 13948 38768
rect 14184 38532 14269 38768
rect 14505 38532 14590 38768
rect 14826 38532 14911 38768
rect 15147 38532 15232 38768
rect 15468 38532 15553 38768
rect 15789 38532 15874 38768
rect 16110 38532 16195 38768
rect 16431 38532 16516 38768
rect 16752 38532 16837 38768
rect 17073 38532 17158 38768
rect 17394 38532 17479 38768
rect 17715 38532 17800 38768
rect 18036 38532 18121 38768
rect 18357 38532 18442 38768
rect 18678 38532 18763 38768
rect 18999 38532 19084 38768
rect 19320 38532 19405 38768
rect 19641 38532 19726 38768
rect 19962 38532 20047 38768
rect 20283 38532 20368 38768
rect 20604 38532 20689 38768
rect 20925 38532 21010 38768
rect 21246 38532 21331 38768
rect 21567 38532 21652 38768
rect 21888 38532 21973 38768
rect 22209 38532 22294 38768
rect 22530 38532 22615 38768
rect 22851 38532 22936 38768
rect 23172 38532 23257 38768
rect 23493 38532 23578 38768
rect 23814 38532 23899 38768
rect 24135 38532 24220 38768
rect 24456 38532 24640 38768
rect -3360 38444 24640 38532
rect -3360 38208 -3087 38444
rect -2851 38208 -2765 38444
rect -2529 38208 -2443 38444
rect -2207 38208 -2121 38444
rect -1885 38208 -1799 38444
rect -1563 38208 -1477 38444
rect -1241 38208 -1155 38444
rect -919 38208 -833 38444
rect -597 38208 -511 38444
rect -275 38208 -189 38444
rect 47 38208 133 38444
rect 369 38208 455 38444
rect 691 38208 777 38444
rect 1013 38208 1099 38444
rect 1335 38208 1421 38444
rect 1657 38208 1743 38444
rect 1979 38208 2065 38444
rect 2301 38208 2387 38444
rect 2623 38208 2709 38444
rect 2945 38208 3031 38444
rect 3267 38208 3353 38444
rect 3589 38208 3675 38444
rect 3911 38208 3997 38444
rect 4233 38208 4318 38444
rect 4554 38208 4639 38444
rect 4875 38208 4960 38444
rect 5196 38208 5281 38444
rect 5517 38208 5602 38444
rect 5838 38208 5923 38444
rect 6159 38208 6244 38444
rect 6480 38208 6565 38444
rect 6801 38208 6886 38444
rect 7122 38208 7207 38444
rect 7443 38208 7528 38444
rect 7764 38208 7849 38444
rect 8085 38208 8170 38444
rect 8406 38208 8491 38444
rect 8727 38208 8812 38444
rect 9048 38208 9133 38444
rect 9369 38208 9454 38444
rect 9690 38208 9775 38444
rect 10011 38208 10096 38444
rect 10332 38208 10417 38444
rect 10653 38208 10738 38444
rect 10974 38208 11059 38444
rect 11295 38208 11380 38444
rect 11616 38208 11701 38444
rect 11937 38208 12022 38444
rect 12258 38208 12343 38444
rect 12579 38208 12664 38444
rect 12900 38208 12985 38444
rect 13221 38208 13306 38444
rect 13542 38208 13627 38444
rect 13863 38208 13948 38444
rect 14184 38208 14269 38444
rect 14505 38208 14590 38444
rect 14826 38208 14911 38444
rect 15147 38208 15232 38444
rect 15468 38208 15553 38444
rect 15789 38208 15874 38444
rect 16110 38208 16195 38444
rect 16431 38208 16516 38444
rect 16752 38208 16837 38444
rect 17073 38208 17158 38444
rect 17394 38208 17479 38444
rect 17715 38208 17800 38444
rect 18036 38208 18121 38444
rect 18357 38208 18442 38444
rect 18678 38208 18763 38444
rect 18999 38208 19084 38444
rect 19320 38208 19405 38444
rect 19641 38208 19726 38444
rect 19962 38208 20047 38444
rect 20283 38208 20368 38444
rect 20604 38208 20689 38444
rect 20925 38208 21010 38444
rect 21246 38208 21331 38444
rect 21567 38208 21652 38444
rect 21888 38208 21973 38444
rect 22209 38208 22294 38444
rect 22530 38208 22615 38444
rect 22851 38208 22936 38444
rect 23172 38208 23257 38444
rect 23493 38208 23578 38444
rect 23814 38208 23899 38444
rect 24135 38208 24220 38444
rect 24456 38208 24640 38444
rect -3360 38120 24640 38208
rect -3360 37884 -3087 38120
rect -2851 37884 -2765 38120
rect -2529 37884 -2443 38120
rect -2207 37884 -2121 38120
rect -1885 37884 -1799 38120
rect -1563 37884 -1477 38120
rect -1241 37884 -1155 38120
rect -919 37884 -833 38120
rect -597 37884 -511 38120
rect -275 37884 -189 38120
rect 47 37884 133 38120
rect 369 37884 455 38120
rect 691 37884 777 38120
rect 1013 37884 1099 38120
rect 1335 37884 1421 38120
rect 1657 37884 1743 38120
rect 1979 37884 2065 38120
rect 2301 37884 2387 38120
rect 2623 37884 2709 38120
rect 2945 37884 3031 38120
rect 3267 37884 3353 38120
rect 3589 37884 3675 38120
rect 3911 37884 3997 38120
rect 4233 37884 4318 38120
rect 4554 37884 4639 38120
rect 4875 37884 4960 38120
rect 5196 37884 5281 38120
rect 5517 37884 5602 38120
rect 5838 37884 5923 38120
rect 6159 37884 6244 38120
rect 6480 37884 6565 38120
rect 6801 37884 6886 38120
rect 7122 37884 7207 38120
rect 7443 37884 7528 38120
rect 7764 37884 7849 38120
rect 8085 37884 8170 38120
rect 8406 37884 8491 38120
rect 8727 37884 8812 38120
rect 9048 37884 9133 38120
rect 9369 37884 9454 38120
rect 9690 37884 9775 38120
rect 10011 37884 10096 38120
rect 10332 37884 10417 38120
rect 10653 37884 10738 38120
rect 10974 37884 11059 38120
rect 11295 37884 11380 38120
rect 11616 37884 11701 38120
rect 11937 37884 12022 38120
rect 12258 37884 12343 38120
rect 12579 37884 12664 38120
rect 12900 37884 12985 38120
rect 13221 37884 13306 38120
rect 13542 37884 13627 38120
rect 13863 37884 13948 38120
rect 14184 37884 14269 38120
rect 14505 37884 14590 38120
rect 14826 37884 14911 38120
rect 15147 37884 15232 38120
rect 15468 37884 15553 38120
rect 15789 37884 15874 38120
rect 16110 37884 16195 38120
rect 16431 37884 16516 38120
rect 16752 37884 16837 38120
rect 17073 37884 17158 38120
rect 17394 37884 17479 38120
rect 17715 37884 17800 38120
rect 18036 37884 18121 38120
rect 18357 37884 18442 38120
rect 18678 37884 18763 38120
rect 18999 37884 19084 38120
rect 19320 37884 19405 38120
rect 19641 37884 19726 38120
rect 19962 37884 20047 38120
rect 20283 37884 20368 38120
rect 20604 37884 20689 38120
rect 20925 37884 21010 38120
rect 21246 37884 21331 38120
rect 21567 37884 21652 38120
rect 21888 37884 21973 38120
rect 22209 37884 22294 38120
rect 22530 37884 22615 38120
rect 22851 37884 22936 38120
rect 23172 37884 23257 38120
rect 23493 37884 23578 38120
rect 23814 37884 23899 38120
rect 24135 37884 24220 38120
rect 24456 37884 24640 38120
rect -3360 37796 24640 37884
rect -3360 37560 -3087 37796
rect -2851 37560 -2765 37796
rect -2529 37560 -2443 37796
rect -2207 37560 -2121 37796
rect -1885 37560 -1799 37796
rect -1563 37560 -1477 37796
rect -1241 37560 -1155 37796
rect -919 37560 -833 37796
rect -597 37560 -511 37796
rect -275 37560 -189 37796
rect 47 37560 133 37796
rect 369 37560 455 37796
rect 691 37560 777 37796
rect 1013 37560 1099 37796
rect 1335 37560 1421 37796
rect 1657 37560 1743 37796
rect 1979 37560 2065 37796
rect 2301 37560 2387 37796
rect 2623 37560 2709 37796
rect 2945 37560 3031 37796
rect 3267 37560 3353 37796
rect 3589 37560 3675 37796
rect 3911 37560 3997 37796
rect 4233 37560 4318 37796
rect 4554 37560 4639 37796
rect 4875 37560 4960 37796
rect 5196 37560 5281 37796
rect 5517 37560 5602 37796
rect 5838 37560 5923 37796
rect 6159 37560 6244 37796
rect 6480 37560 6565 37796
rect 6801 37560 6886 37796
rect 7122 37560 7207 37796
rect 7443 37560 7528 37796
rect 7764 37560 7849 37796
rect 8085 37560 8170 37796
rect 8406 37560 8491 37796
rect 8727 37560 8812 37796
rect 9048 37560 9133 37796
rect 9369 37560 9454 37796
rect 9690 37560 9775 37796
rect 10011 37560 10096 37796
rect 10332 37560 10417 37796
rect 10653 37560 10738 37796
rect 10974 37560 11059 37796
rect 11295 37560 11380 37796
rect 11616 37560 11701 37796
rect 11937 37560 12022 37796
rect 12258 37560 12343 37796
rect 12579 37560 12664 37796
rect 12900 37560 12985 37796
rect 13221 37560 13306 37796
rect 13542 37560 13627 37796
rect 13863 37560 13948 37796
rect 14184 37560 14269 37796
rect 14505 37560 14590 37796
rect 14826 37560 14911 37796
rect 15147 37560 15232 37796
rect 15468 37560 15553 37796
rect 15789 37560 15874 37796
rect 16110 37560 16195 37796
rect 16431 37560 16516 37796
rect 16752 37560 16837 37796
rect 17073 37560 17158 37796
rect 17394 37560 17479 37796
rect 17715 37560 17800 37796
rect 18036 37560 18121 37796
rect 18357 37560 18442 37796
rect 18678 37560 18763 37796
rect 18999 37560 19084 37796
rect 19320 37560 19405 37796
rect 19641 37560 19726 37796
rect 19962 37560 20047 37796
rect 20283 37560 20368 37796
rect 20604 37560 20689 37796
rect 20925 37560 21010 37796
rect 21246 37560 21331 37796
rect 21567 37560 21652 37796
rect 21888 37560 21973 37796
rect 22209 37560 22294 37796
rect 22530 37560 22615 37796
rect 22851 37560 22936 37796
rect 23172 37560 23257 37796
rect 23493 37560 23578 37796
rect 23814 37560 23899 37796
rect 24135 37560 24220 37796
rect 24456 37560 24640 37796
rect -3360 37472 24640 37560
rect -3360 37236 -3087 37472
rect -2851 37236 -2765 37472
rect -2529 37236 -2443 37472
rect -2207 37236 -2121 37472
rect -1885 37236 -1799 37472
rect -1563 37236 -1477 37472
rect -1241 37236 -1155 37472
rect -919 37236 -833 37472
rect -597 37236 -511 37472
rect -275 37236 -189 37472
rect 47 37236 133 37472
rect 369 37236 455 37472
rect 691 37236 777 37472
rect 1013 37236 1099 37472
rect 1335 37236 1421 37472
rect 1657 37236 1743 37472
rect 1979 37236 2065 37472
rect 2301 37236 2387 37472
rect 2623 37236 2709 37472
rect 2945 37236 3031 37472
rect 3267 37236 3353 37472
rect 3589 37236 3675 37472
rect 3911 37236 3997 37472
rect 4233 37236 4318 37472
rect 4554 37236 4639 37472
rect 4875 37236 4960 37472
rect 5196 37236 5281 37472
rect 5517 37236 5602 37472
rect 5838 37236 5923 37472
rect 6159 37236 6244 37472
rect 6480 37236 6565 37472
rect 6801 37236 6886 37472
rect 7122 37236 7207 37472
rect 7443 37236 7528 37472
rect 7764 37236 7849 37472
rect 8085 37236 8170 37472
rect 8406 37236 8491 37472
rect 8727 37236 8812 37472
rect 9048 37236 9133 37472
rect 9369 37236 9454 37472
rect 9690 37236 9775 37472
rect 10011 37236 10096 37472
rect 10332 37236 10417 37472
rect 10653 37236 10738 37472
rect 10974 37236 11059 37472
rect 11295 37236 11380 37472
rect 11616 37236 11701 37472
rect 11937 37236 12022 37472
rect 12258 37236 12343 37472
rect 12579 37236 12664 37472
rect 12900 37236 12985 37472
rect 13221 37236 13306 37472
rect 13542 37236 13627 37472
rect 13863 37236 13948 37472
rect 14184 37236 14269 37472
rect 14505 37236 14590 37472
rect 14826 37236 14911 37472
rect 15147 37236 15232 37472
rect 15468 37236 15553 37472
rect 15789 37236 15874 37472
rect 16110 37236 16195 37472
rect 16431 37236 16516 37472
rect 16752 37236 16837 37472
rect 17073 37236 17158 37472
rect 17394 37236 17479 37472
rect 17715 37236 17800 37472
rect 18036 37236 18121 37472
rect 18357 37236 18442 37472
rect 18678 37236 18763 37472
rect 18999 37236 19084 37472
rect 19320 37236 19405 37472
rect 19641 37236 19726 37472
rect 19962 37236 20047 37472
rect 20283 37236 20368 37472
rect 20604 37236 20689 37472
rect 20925 37236 21010 37472
rect 21246 37236 21331 37472
rect 21567 37236 21652 37472
rect 21888 37236 21973 37472
rect 22209 37236 22294 37472
rect 22530 37236 22615 37472
rect 22851 37236 22936 37472
rect 23172 37236 23257 37472
rect 23493 37236 23578 37472
rect 23814 37236 23899 37472
rect 24135 37236 24220 37472
rect 24456 37236 24640 37472
rect -3360 37148 24640 37236
rect -3360 36912 -3087 37148
rect -2851 36912 -2765 37148
rect -2529 36912 -2443 37148
rect -2207 36912 -2121 37148
rect -1885 36912 -1799 37148
rect -1563 36912 -1477 37148
rect -1241 36912 -1155 37148
rect -919 36912 -833 37148
rect -597 36912 -511 37148
rect -275 36912 -189 37148
rect 47 36912 133 37148
rect 369 36912 455 37148
rect 691 36912 777 37148
rect 1013 36912 1099 37148
rect 1335 36912 1421 37148
rect 1657 36912 1743 37148
rect 1979 36912 2065 37148
rect 2301 36912 2387 37148
rect 2623 36912 2709 37148
rect 2945 36912 3031 37148
rect 3267 36912 3353 37148
rect 3589 36912 3675 37148
rect 3911 36912 3997 37148
rect 4233 36912 4318 37148
rect 4554 36912 4639 37148
rect 4875 36912 4960 37148
rect 5196 36912 5281 37148
rect 5517 36912 5602 37148
rect 5838 36912 5923 37148
rect 6159 36912 6244 37148
rect 6480 36912 6565 37148
rect 6801 36912 6886 37148
rect 7122 36912 7207 37148
rect 7443 36912 7528 37148
rect 7764 36912 7849 37148
rect 8085 36912 8170 37148
rect 8406 36912 8491 37148
rect 8727 36912 8812 37148
rect 9048 36912 9133 37148
rect 9369 36912 9454 37148
rect 9690 36912 9775 37148
rect 10011 36912 10096 37148
rect 10332 36912 10417 37148
rect 10653 36912 10738 37148
rect 10974 36912 11059 37148
rect 11295 36912 11380 37148
rect 11616 36912 11701 37148
rect 11937 36912 12022 37148
rect 12258 36912 12343 37148
rect 12579 36912 12664 37148
rect 12900 36912 12985 37148
rect 13221 36912 13306 37148
rect 13542 36912 13627 37148
rect 13863 36912 13948 37148
rect 14184 36912 14269 37148
rect 14505 36912 14590 37148
rect 14826 36912 14911 37148
rect 15147 36912 15232 37148
rect 15468 36912 15553 37148
rect 15789 36912 15874 37148
rect 16110 36912 16195 37148
rect 16431 36912 16516 37148
rect 16752 36912 16837 37148
rect 17073 36912 17158 37148
rect 17394 36912 17479 37148
rect 17715 36912 17800 37148
rect 18036 36912 18121 37148
rect 18357 36912 18442 37148
rect 18678 36912 18763 37148
rect 18999 36912 19084 37148
rect 19320 36912 19405 37148
rect 19641 36912 19726 37148
rect 19962 36912 20047 37148
rect 20283 36912 20368 37148
rect 20604 36912 20689 37148
rect 20925 36912 21010 37148
rect 21246 36912 21331 37148
rect 21567 36912 21652 37148
rect 21888 36912 21973 37148
rect 22209 36912 22294 37148
rect 22530 36912 22615 37148
rect 22851 36912 22936 37148
rect 23172 36912 23257 37148
rect 23493 36912 23578 37148
rect 23814 36912 23899 37148
rect 24135 36912 24220 37148
rect 24456 36912 24640 37148
rect -3360 36824 24640 36912
rect -3360 36588 -3087 36824
rect -2851 36588 -2765 36824
rect -2529 36588 -2443 36824
rect -2207 36588 -2121 36824
rect -1885 36588 -1799 36824
rect -1563 36588 -1477 36824
rect -1241 36588 -1155 36824
rect -919 36588 -833 36824
rect -597 36588 -511 36824
rect -275 36588 -189 36824
rect 47 36588 133 36824
rect 369 36588 455 36824
rect 691 36588 777 36824
rect 1013 36588 1099 36824
rect 1335 36588 1421 36824
rect 1657 36588 1743 36824
rect 1979 36588 2065 36824
rect 2301 36588 2387 36824
rect 2623 36588 2709 36824
rect 2945 36588 3031 36824
rect 3267 36588 3353 36824
rect 3589 36588 3675 36824
rect 3911 36588 3997 36824
rect 4233 36588 4318 36824
rect 4554 36588 4639 36824
rect 4875 36588 4960 36824
rect 5196 36588 5281 36824
rect 5517 36588 5602 36824
rect 5838 36588 5923 36824
rect 6159 36588 6244 36824
rect 6480 36588 6565 36824
rect 6801 36588 6886 36824
rect 7122 36588 7207 36824
rect 7443 36588 7528 36824
rect 7764 36588 7849 36824
rect 8085 36588 8170 36824
rect 8406 36588 8491 36824
rect 8727 36588 8812 36824
rect 9048 36588 9133 36824
rect 9369 36588 9454 36824
rect 9690 36588 9775 36824
rect 10011 36588 10096 36824
rect 10332 36588 10417 36824
rect 10653 36588 10738 36824
rect 10974 36588 11059 36824
rect 11295 36588 11380 36824
rect 11616 36588 11701 36824
rect 11937 36588 12022 36824
rect 12258 36588 12343 36824
rect 12579 36588 12664 36824
rect 12900 36588 12985 36824
rect 13221 36588 13306 36824
rect 13542 36588 13627 36824
rect 13863 36588 13948 36824
rect 14184 36588 14269 36824
rect 14505 36588 14590 36824
rect 14826 36588 14911 36824
rect 15147 36588 15232 36824
rect 15468 36588 15553 36824
rect 15789 36588 15874 36824
rect 16110 36588 16195 36824
rect 16431 36588 16516 36824
rect 16752 36588 16837 36824
rect 17073 36588 17158 36824
rect 17394 36588 17479 36824
rect 17715 36588 17800 36824
rect 18036 36588 18121 36824
rect 18357 36588 18442 36824
rect 18678 36588 18763 36824
rect 18999 36588 19084 36824
rect 19320 36588 19405 36824
rect 19641 36588 19726 36824
rect 19962 36588 20047 36824
rect 20283 36588 20368 36824
rect 20604 36588 20689 36824
rect 20925 36588 21010 36824
rect 21246 36588 21331 36824
rect 21567 36588 21652 36824
rect 21888 36588 21973 36824
rect 22209 36588 22294 36824
rect 22530 36588 22615 36824
rect 22851 36588 22936 36824
rect 23172 36588 23257 36824
rect 23493 36588 23578 36824
rect 23814 36588 23899 36824
rect 24135 36588 24220 36824
rect 24456 36588 24640 36824
rect -3360 36500 24640 36588
rect -3360 36264 -3087 36500
rect -2851 36264 -2765 36500
rect -2529 36264 -2443 36500
rect -2207 36264 -2121 36500
rect -1885 36264 -1799 36500
rect -1563 36264 -1477 36500
rect -1241 36264 -1155 36500
rect -919 36264 -833 36500
rect -597 36264 -511 36500
rect -275 36264 -189 36500
rect 47 36264 133 36500
rect 369 36264 455 36500
rect 691 36264 777 36500
rect 1013 36264 1099 36500
rect 1335 36264 1421 36500
rect 1657 36264 1743 36500
rect 1979 36264 2065 36500
rect 2301 36264 2387 36500
rect 2623 36264 2709 36500
rect 2945 36264 3031 36500
rect 3267 36264 3353 36500
rect 3589 36264 3675 36500
rect 3911 36264 3997 36500
rect 4233 36264 4318 36500
rect 4554 36264 4639 36500
rect 4875 36264 4960 36500
rect 5196 36264 5281 36500
rect 5517 36264 5602 36500
rect 5838 36264 5923 36500
rect 6159 36264 6244 36500
rect 6480 36264 6565 36500
rect 6801 36264 6886 36500
rect 7122 36264 7207 36500
rect 7443 36264 7528 36500
rect 7764 36264 7849 36500
rect 8085 36264 8170 36500
rect 8406 36264 8491 36500
rect 8727 36264 8812 36500
rect 9048 36264 9133 36500
rect 9369 36264 9454 36500
rect 9690 36264 9775 36500
rect 10011 36264 10096 36500
rect 10332 36264 10417 36500
rect 10653 36264 10738 36500
rect 10974 36264 11059 36500
rect 11295 36264 11380 36500
rect 11616 36264 11701 36500
rect 11937 36264 12022 36500
rect 12258 36264 12343 36500
rect 12579 36264 12664 36500
rect 12900 36264 12985 36500
rect 13221 36264 13306 36500
rect 13542 36264 13627 36500
rect 13863 36264 13948 36500
rect 14184 36264 14269 36500
rect 14505 36264 14590 36500
rect 14826 36264 14911 36500
rect 15147 36264 15232 36500
rect 15468 36264 15553 36500
rect 15789 36264 15874 36500
rect 16110 36264 16195 36500
rect 16431 36264 16516 36500
rect 16752 36264 16837 36500
rect 17073 36264 17158 36500
rect 17394 36264 17479 36500
rect 17715 36264 17800 36500
rect 18036 36264 18121 36500
rect 18357 36264 18442 36500
rect 18678 36264 18763 36500
rect 18999 36264 19084 36500
rect 19320 36264 19405 36500
rect 19641 36264 19726 36500
rect 19962 36264 20047 36500
rect 20283 36264 20368 36500
rect 20604 36264 20689 36500
rect 20925 36264 21010 36500
rect 21246 36264 21331 36500
rect 21567 36264 21652 36500
rect 21888 36264 21973 36500
rect 22209 36264 22294 36500
rect 22530 36264 22615 36500
rect 22851 36264 22936 36500
rect 23172 36264 23257 36500
rect 23493 36264 23578 36500
rect 23814 36264 23899 36500
rect 24135 36264 24220 36500
rect 24456 36264 24640 36500
rect -3360 36176 24640 36264
rect -3360 35940 -3087 36176
rect -2851 35940 -2765 36176
rect -2529 35940 -2443 36176
rect -2207 35940 -2121 36176
rect -1885 35940 -1799 36176
rect -1563 35940 -1477 36176
rect -1241 35940 -1155 36176
rect -919 35940 -833 36176
rect -597 35940 -511 36176
rect -275 35940 -189 36176
rect 47 35940 133 36176
rect 369 35940 455 36176
rect 691 35940 777 36176
rect 1013 35940 1099 36176
rect 1335 35940 1421 36176
rect 1657 35940 1743 36176
rect 1979 35940 2065 36176
rect 2301 35940 2387 36176
rect 2623 35940 2709 36176
rect 2945 35940 3031 36176
rect 3267 35940 3353 36176
rect 3589 35940 3675 36176
rect 3911 35940 3997 36176
rect 4233 35940 4318 36176
rect 4554 35940 4639 36176
rect 4875 35940 4960 36176
rect 5196 35940 5281 36176
rect 5517 35940 5602 36176
rect 5838 35940 5923 36176
rect 6159 35940 6244 36176
rect 6480 35940 6565 36176
rect 6801 35940 6886 36176
rect 7122 35940 7207 36176
rect 7443 35940 7528 36176
rect 7764 35940 7849 36176
rect 8085 35940 8170 36176
rect 8406 35940 8491 36176
rect 8727 35940 8812 36176
rect 9048 35940 9133 36176
rect 9369 35940 9454 36176
rect 9690 35940 9775 36176
rect 10011 35940 10096 36176
rect 10332 35940 10417 36176
rect 10653 35940 10738 36176
rect 10974 35940 11059 36176
rect 11295 35940 11380 36176
rect 11616 35940 11701 36176
rect 11937 35940 12022 36176
rect 12258 35940 12343 36176
rect 12579 35940 12664 36176
rect 12900 35940 12985 36176
rect 13221 35940 13306 36176
rect 13542 35940 13627 36176
rect 13863 35940 13948 36176
rect 14184 35940 14269 36176
rect 14505 35940 14590 36176
rect 14826 35940 14911 36176
rect 15147 35940 15232 36176
rect 15468 35940 15553 36176
rect 15789 35940 15874 36176
rect 16110 35940 16195 36176
rect 16431 35940 16516 36176
rect 16752 35940 16837 36176
rect 17073 35940 17158 36176
rect 17394 35940 17479 36176
rect 17715 35940 17800 36176
rect 18036 35940 18121 36176
rect 18357 35940 18442 36176
rect 18678 35940 18763 36176
rect 18999 35940 19084 36176
rect 19320 35940 19405 36176
rect 19641 35940 19726 36176
rect 19962 35940 20047 36176
rect 20283 35940 20368 36176
rect 20604 35940 20689 36176
rect 20925 35940 21010 36176
rect 21246 35940 21331 36176
rect 21567 35940 21652 36176
rect 21888 35940 21973 36176
rect 22209 35940 22294 36176
rect 22530 35940 22615 36176
rect 22851 35940 22936 36176
rect 23172 35940 23257 36176
rect 23493 35940 23578 36176
rect 23814 35940 23899 36176
rect 24135 35940 24220 36176
rect 24456 35940 24640 36176
rect -3360 35852 24640 35940
rect -3360 35616 -3087 35852
rect -2851 35616 -2765 35852
rect -2529 35616 -2443 35852
rect -2207 35616 -2121 35852
rect -1885 35616 -1799 35852
rect -1563 35616 -1477 35852
rect -1241 35616 -1155 35852
rect -919 35616 -833 35852
rect -597 35616 -511 35852
rect -275 35616 -189 35852
rect 47 35616 133 35852
rect 369 35616 455 35852
rect 691 35616 777 35852
rect 1013 35616 1099 35852
rect 1335 35616 1421 35852
rect 1657 35616 1743 35852
rect 1979 35616 2065 35852
rect 2301 35616 2387 35852
rect 2623 35616 2709 35852
rect 2945 35616 3031 35852
rect 3267 35616 3353 35852
rect 3589 35616 3675 35852
rect 3911 35616 3997 35852
rect 4233 35616 4318 35852
rect 4554 35616 4639 35852
rect 4875 35616 4960 35852
rect 5196 35616 5281 35852
rect 5517 35616 5602 35852
rect 5838 35616 5923 35852
rect 6159 35616 6244 35852
rect 6480 35616 6565 35852
rect 6801 35616 6886 35852
rect 7122 35616 7207 35852
rect 7443 35616 7528 35852
rect 7764 35616 7849 35852
rect 8085 35616 8170 35852
rect 8406 35616 8491 35852
rect 8727 35616 8812 35852
rect 9048 35616 9133 35852
rect 9369 35616 9454 35852
rect 9690 35616 9775 35852
rect 10011 35616 10096 35852
rect 10332 35616 10417 35852
rect 10653 35616 10738 35852
rect 10974 35616 11059 35852
rect 11295 35616 11380 35852
rect 11616 35616 11701 35852
rect 11937 35616 12022 35852
rect 12258 35616 12343 35852
rect 12579 35616 12664 35852
rect 12900 35616 12985 35852
rect 13221 35616 13306 35852
rect 13542 35616 13627 35852
rect 13863 35616 13948 35852
rect 14184 35616 14269 35852
rect 14505 35616 14590 35852
rect 14826 35616 14911 35852
rect 15147 35616 15232 35852
rect 15468 35616 15553 35852
rect 15789 35616 15874 35852
rect 16110 35616 16195 35852
rect 16431 35616 16516 35852
rect 16752 35616 16837 35852
rect 17073 35616 17158 35852
rect 17394 35616 17479 35852
rect 17715 35616 17800 35852
rect 18036 35616 18121 35852
rect 18357 35616 18442 35852
rect 18678 35616 18763 35852
rect 18999 35616 19084 35852
rect 19320 35616 19405 35852
rect 19641 35616 19726 35852
rect 19962 35616 20047 35852
rect 20283 35616 20368 35852
rect 20604 35616 20689 35852
rect 20925 35616 21010 35852
rect 21246 35616 21331 35852
rect 21567 35616 21652 35852
rect 21888 35616 21973 35852
rect 22209 35616 22294 35852
rect 22530 35616 22615 35852
rect 22851 35616 22936 35852
rect 23172 35616 23257 35852
rect 23493 35616 23578 35852
rect 23814 35616 23899 35852
rect 24135 35616 24220 35852
rect 24456 35616 24640 35852
rect -3360 35528 24640 35616
rect -3360 35292 -3087 35528
rect -2851 35292 -2765 35528
rect -2529 35292 -2443 35528
rect -2207 35292 -2121 35528
rect -1885 35292 -1799 35528
rect -1563 35292 -1477 35528
rect -1241 35292 -1155 35528
rect -919 35292 -833 35528
rect -597 35292 -511 35528
rect -275 35292 -189 35528
rect 47 35292 133 35528
rect 369 35292 455 35528
rect 691 35292 777 35528
rect 1013 35292 1099 35528
rect 1335 35292 1421 35528
rect 1657 35292 1743 35528
rect 1979 35292 2065 35528
rect 2301 35292 2387 35528
rect 2623 35292 2709 35528
rect 2945 35292 3031 35528
rect 3267 35292 3353 35528
rect 3589 35292 3675 35528
rect 3911 35292 3997 35528
rect 4233 35292 4318 35528
rect 4554 35292 4639 35528
rect 4875 35292 4960 35528
rect 5196 35292 5281 35528
rect 5517 35292 5602 35528
rect 5838 35292 5923 35528
rect 6159 35292 6244 35528
rect 6480 35292 6565 35528
rect 6801 35292 6886 35528
rect 7122 35292 7207 35528
rect 7443 35292 7528 35528
rect 7764 35292 7849 35528
rect 8085 35292 8170 35528
rect 8406 35292 8491 35528
rect 8727 35292 8812 35528
rect 9048 35292 9133 35528
rect 9369 35292 9454 35528
rect 9690 35292 9775 35528
rect 10011 35292 10096 35528
rect 10332 35292 10417 35528
rect 10653 35292 10738 35528
rect 10974 35292 11059 35528
rect 11295 35292 11380 35528
rect 11616 35292 11701 35528
rect 11937 35292 12022 35528
rect 12258 35292 12343 35528
rect 12579 35292 12664 35528
rect 12900 35292 12985 35528
rect 13221 35292 13306 35528
rect 13542 35292 13627 35528
rect 13863 35292 13948 35528
rect 14184 35292 14269 35528
rect 14505 35292 14590 35528
rect 14826 35292 14911 35528
rect 15147 35292 15232 35528
rect 15468 35292 15553 35528
rect 15789 35292 15874 35528
rect 16110 35292 16195 35528
rect 16431 35292 16516 35528
rect 16752 35292 16837 35528
rect 17073 35292 17158 35528
rect 17394 35292 17479 35528
rect 17715 35292 17800 35528
rect 18036 35292 18121 35528
rect 18357 35292 18442 35528
rect 18678 35292 18763 35528
rect 18999 35292 19084 35528
rect 19320 35292 19405 35528
rect 19641 35292 19726 35528
rect 19962 35292 20047 35528
rect 20283 35292 20368 35528
rect 20604 35292 20689 35528
rect 20925 35292 21010 35528
rect 21246 35292 21331 35528
rect 21567 35292 21652 35528
rect 21888 35292 21973 35528
rect 22209 35292 22294 35528
rect 22530 35292 22615 35528
rect 22851 35292 22936 35528
rect 23172 35292 23257 35528
rect 23493 35292 23578 35528
rect 23814 35292 23899 35528
rect 24135 35292 24220 35528
rect 24456 35292 24640 35528
rect -3360 35204 24640 35292
rect -3360 34968 -3087 35204
rect -2851 34968 -2765 35204
rect -2529 34968 -2443 35204
rect -2207 34968 -2121 35204
rect -1885 34968 -1799 35204
rect -1563 34968 -1477 35204
rect -1241 34968 -1155 35204
rect -919 34968 -833 35204
rect -597 34968 -511 35204
rect -275 34968 -189 35204
rect 47 34968 133 35204
rect 369 34968 455 35204
rect 691 34968 777 35204
rect 1013 34968 1099 35204
rect 1335 34968 1421 35204
rect 1657 34968 1743 35204
rect 1979 34968 2065 35204
rect 2301 34968 2387 35204
rect 2623 34968 2709 35204
rect 2945 34968 3031 35204
rect 3267 34968 3353 35204
rect 3589 34968 3675 35204
rect 3911 34968 3997 35204
rect 4233 34968 4318 35204
rect 4554 34968 4639 35204
rect 4875 34968 4960 35204
rect 5196 34968 5281 35204
rect 5517 34968 5602 35204
rect 5838 34968 5923 35204
rect 6159 34968 6244 35204
rect 6480 34968 6565 35204
rect 6801 34968 6886 35204
rect 7122 34968 7207 35204
rect 7443 34968 7528 35204
rect 7764 34968 7849 35204
rect 8085 34968 8170 35204
rect 8406 34968 8491 35204
rect 8727 34968 8812 35204
rect 9048 34968 9133 35204
rect 9369 34968 9454 35204
rect 9690 34968 9775 35204
rect 10011 34968 10096 35204
rect 10332 34968 10417 35204
rect 10653 34968 10738 35204
rect 10974 34968 11059 35204
rect 11295 34968 11380 35204
rect 11616 34968 11701 35204
rect 11937 34968 12022 35204
rect 12258 34968 12343 35204
rect 12579 34968 12664 35204
rect 12900 34968 12985 35204
rect 13221 34968 13306 35204
rect 13542 34968 13627 35204
rect 13863 34968 13948 35204
rect 14184 34968 14269 35204
rect 14505 34968 14590 35204
rect 14826 34968 14911 35204
rect 15147 34968 15232 35204
rect 15468 34968 15553 35204
rect 15789 34968 15874 35204
rect 16110 34968 16195 35204
rect 16431 34968 16516 35204
rect 16752 34968 16837 35204
rect 17073 34968 17158 35204
rect 17394 34968 17479 35204
rect 17715 34968 17800 35204
rect 18036 34968 18121 35204
rect 18357 34968 18442 35204
rect 18678 34968 18763 35204
rect 18999 34968 19084 35204
rect 19320 34968 19405 35204
rect 19641 34968 19726 35204
rect 19962 34968 20047 35204
rect 20283 34968 20368 35204
rect 20604 34968 20689 35204
rect 20925 34968 21010 35204
rect 21246 34968 21331 35204
rect 21567 34968 21652 35204
rect 21888 34968 21973 35204
rect 22209 34968 22294 35204
rect 22530 34968 22615 35204
rect 22851 34968 22936 35204
rect 23172 34968 23257 35204
rect 23493 34968 23578 35204
rect 23814 34968 23899 35204
rect 24135 34968 24220 35204
rect 24456 34968 24640 35204
rect -3360 34880 24640 34968
rect -3360 34644 -3087 34880
rect -2851 34644 -2765 34880
rect -2529 34644 -2443 34880
rect -2207 34644 -2121 34880
rect -1885 34644 -1799 34880
rect -1563 34644 -1477 34880
rect -1241 34644 -1155 34880
rect -919 34644 -833 34880
rect -597 34644 -511 34880
rect -275 34644 -189 34880
rect 47 34644 133 34880
rect 369 34644 455 34880
rect 691 34644 777 34880
rect 1013 34644 1099 34880
rect 1335 34644 1421 34880
rect 1657 34644 1743 34880
rect 1979 34644 2065 34880
rect 2301 34644 2387 34880
rect 2623 34644 2709 34880
rect 2945 34644 3031 34880
rect 3267 34644 3353 34880
rect 3589 34644 3675 34880
rect 3911 34644 3997 34880
rect 4233 34644 4318 34880
rect 4554 34644 4639 34880
rect 4875 34644 4960 34880
rect 5196 34644 5281 34880
rect 5517 34644 5602 34880
rect 5838 34644 5923 34880
rect 6159 34644 6244 34880
rect 6480 34644 6565 34880
rect 6801 34644 6886 34880
rect 7122 34644 7207 34880
rect 7443 34644 7528 34880
rect 7764 34644 7849 34880
rect 8085 34644 8170 34880
rect 8406 34644 8491 34880
rect 8727 34644 8812 34880
rect 9048 34644 9133 34880
rect 9369 34644 9454 34880
rect 9690 34644 9775 34880
rect 10011 34644 10096 34880
rect 10332 34644 10417 34880
rect 10653 34644 10738 34880
rect 10974 34644 11059 34880
rect 11295 34644 11380 34880
rect 11616 34644 11701 34880
rect 11937 34644 12022 34880
rect 12258 34644 12343 34880
rect 12579 34644 12664 34880
rect 12900 34644 12985 34880
rect 13221 34644 13306 34880
rect 13542 34644 13627 34880
rect 13863 34644 13948 34880
rect 14184 34644 14269 34880
rect 14505 34644 14590 34880
rect 14826 34644 14911 34880
rect 15147 34644 15232 34880
rect 15468 34644 15553 34880
rect 15789 34644 15874 34880
rect 16110 34644 16195 34880
rect 16431 34644 16516 34880
rect 16752 34644 16837 34880
rect 17073 34644 17158 34880
rect 17394 34644 17479 34880
rect 17715 34644 17800 34880
rect 18036 34644 18121 34880
rect 18357 34644 18442 34880
rect 18678 34644 18763 34880
rect 18999 34644 19084 34880
rect 19320 34644 19405 34880
rect 19641 34644 19726 34880
rect 19962 34644 20047 34880
rect 20283 34644 20368 34880
rect 20604 34644 20689 34880
rect 20925 34644 21010 34880
rect 21246 34644 21331 34880
rect 21567 34644 21652 34880
rect 21888 34644 21973 34880
rect 22209 34644 22294 34880
rect 22530 34644 22615 34880
rect 22851 34644 22936 34880
rect 23172 34644 23257 34880
rect 23493 34644 23578 34880
rect 23814 34644 23899 34880
rect 24135 34644 24220 34880
rect 24456 34644 24640 34880
rect -3360 34609 24640 34644
rect -3360 34608 -2720 34609
rect 24000 34608 24640 34609
rect -3360 18423 24640 18448
rect -3360 18187 -3185 18423
rect -2949 18187 -2862 18423
rect -2626 18187 -2539 18423
rect -2303 18187 -2216 18423
rect -1980 18187 -1893 18423
rect -1657 18187 -1570 18423
rect -1334 18187 -1247 18423
rect -1011 18187 -924 18423
rect -688 18187 -601 18423
rect -365 18187 -278 18423
rect -42 18187 45 18423
rect 281 18187 368 18423
rect 604 18187 691 18423
rect 927 18187 1014 18423
rect 1250 18187 1337 18423
rect 1573 18187 1660 18423
rect 1896 18187 1983 18423
rect 2219 18187 2306 18423
rect 2542 18187 2629 18423
rect 2865 18187 2952 18423
rect 3188 18187 3275 18423
rect 3511 18187 3598 18423
rect 3834 18187 3921 18423
rect 4157 18187 4244 18423
rect 4480 18187 4567 18423
rect 4803 18187 4890 18423
rect 5126 18187 5213 18423
rect 5449 18187 5536 18423
rect 5772 18187 5859 18423
rect 6095 18187 6182 18423
rect 6418 18187 6505 18423
rect 6741 18187 6828 18423
rect 7064 18187 7150 18423
rect 7386 18187 7472 18423
rect 7708 18187 7794 18423
rect 8030 18187 8116 18423
rect 8352 18187 8438 18423
rect 8674 18187 8760 18423
rect 8996 18187 9082 18423
rect 9318 18187 9404 18423
rect 9640 18187 9726 18423
rect 9962 18187 10048 18423
rect 10284 18187 10370 18423
rect 10606 18187 10692 18423
rect 10928 18187 11014 18423
rect 11250 18187 11336 18423
rect 11572 18187 11658 18423
rect 11894 18187 11980 18423
rect 12216 18187 12302 18423
rect 12538 18187 12624 18423
rect 12860 18187 12946 18423
rect 13182 18187 13268 18423
rect 13504 18187 13590 18423
rect 13826 18187 13912 18423
rect 14148 18187 14234 18423
rect 14470 18187 14556 18423
rect 14792 18187 14878 18423
rect 15114 18187 15200 18423
rect 15436 18187 15522 18423
rect 15758 18187 15844 18423
rect 16080 18187 16166 18423
rect 16402 18187 16488 18423
rect 16724 18187 16810 18423
rect 17046 18187 17132 18423
rect 17368 18187 17454 18423
rect 17690 18187 17776 18423
rect 18012 18187 18098 18423
rect 18334 18187 18420 18423
rect 18656 18187 18742 18423
rect 18978 18187 19064 18423
rect 19300 18187 19386 18423
rect 19622 18187 19708 18423
rect 19944 18187 20030 18423
rect 20266 18187 20352 18423
rect 20588 18187 20674 18423
rect 20910 18187 20996 18423
rect 21232 18187 21318 18423
rect 21554 18187 21640 18423
rect 21876 18187 21962 18423
rect 22198 18187 22284 18423
rect 22520 18187 22606 18423
rect 22842 18187 22928 18423
rect 23164 18187 23250 18423
rect 23486 18187 23572 18423
rect 23808 18187 23894 18423
rect 24130 18187 24216 18423
rect 24452 18187 24640 18423
rect -3360 18087 24640 18187
rect -3360 17851 -3185 18087
rect -2949 17851 -2862 18087
rect -2626 17851 -2539 18087
rect -2303 17851 -2216 18087
rect -1980 17851 -1893 18087
rect -1657 17851 -1570 18087
rect -1334 17851 -1247 18087
rect -1011 17851 -924 18087
rect -688 17851 -601 18087
rect -365 17851 -278 18087
rect -42 17851 45 18087
rect 281 17851 368 18087
rect 604 17851 691 18087
rect 927 17851 1014 18087
rect 1250 17851 1337 18087
rect 1573 17851 1660 18087
rect 1896 17851 1983 18087
rect 2219 17851 2306 18087
rect 2542 17851 2629 18087
rect 2865 17851 2952 18087
rect 3188 17851 3275 18087
rect 3511 17851 3598 18087
rect 3834 17851 3921 18087
rect 4157 17851 4244 18087
rect 4480 17851 4567 18087
rect 4803 17851 4890 18087
rect 5126 17851 5213 18087
rect 5449 17851 5536 18087
rect 5772 17851 5859 18087
rect 6095 17851 6182 18087
rect 6418 17851 6505 18087
rect 6741 17851 6828 18087
rect 7064 17851 7150 18087
rect 7386 17851 7472 18087
rect 7708 17851 7794 18087
rect 8030 17851 8116 18087
rect 8352 17851 8438 18087
rect 8674 17851 8760 18087
rect 8996 17851 9082 18087
rect 9318 17851 9404 18087
rect 9640 17851 9726 18087
rect 9962 17851 10048 18087
rect 10284 17851 10370 18087
rect 10606 17851 10692 18087
rect 10928 17851 11014 18087
rect 11250 17851 11336 18087
rect 11572 17851 11658 18087
rect 11894 17851 11980 18087
rect 12216 17851 12302 18087
rect 12538 17851 12624 18087
rect 12860 17851 12946 18087
rect 13182 17851 13268 18087
rect 13504 17851 13590 18087
rect 13826 17851 13912 18087
rect 14148 17851 14234 18087
rect 14470 17851 14556 18087
rect 14792 17851 14878 18087
rect 15114 17851 15200 18087
rect 15436 17851 15522 18087
rect 15758 17851 15844 18087
rect 16080 17851 16166 18087
rect 16402 17851 16488 18087
rect 16724 17851 16810 18087
rect 17046 17851 17132 18087
rect 17368 17851 17454 18087
rect 17690 17851 17776 18087
rect 18012 17851 18098 18087
rect 18334 17851 18420 18087
rect 18656 17851 18742 18087
rect 18978 17851 19064 18087
rect 19300 17851 19386 18087
rect 19622 17851 19708 18087
rect 19944 17851 20030 18087
rect 20266 17851 20352 18087
rect 20588 17851 20674 18087
rect 20910 17851 20996 18087
rect 21232 17851 21318 18087
rect 21554 17851 21640 18087
rect 21876 17851 21962 18087
rect 22198 17851 22284 18087
rect 22520 17851 22606 18087
rect 22842 17851 22928 18087
rect 23164 17851 23250 18087
rect 23486 17851 23572 18087
rect 23808 17851 23894 18087
rect 24130 17851 24216 18087
rect 24452 17851 24640 18087
rect -3360 17751 24640 17851
rect -3360 17515 -3185 17751
rect -2949 17515 -2862 17751
rect -2626 17515 -2539 17751
rect -2303 17515 -2216 17751
rect -1980 17515 -1893 17751
rect -1657 17515 -1570 17751
rect -1334 17515 -1247 17751
rect -1011 17515 -924 17751
rect -688 17515 -601 17751
rect -365 17515 -278 17751
rect -42 17515 45 17751
rect 281 17515 368 17751
rect 604 17515 691 17751
rect 927 17515 1014 17751
rect 1250 17515 1337 17751
rect 1573 17515 1660 17751
rect 1896 17515 1983 17751
rect 2219 17515 2306 17751
rect 2542 17515 2629 17751
rect 2865 17515 2952 17751
rect 3188 17515 3275 17751
rect 3511 17515 3598 17751
rect 3834 17515 3921 17751
rect 4157 17515 4244 17751
rect 4480 17515 4567 17751
rect 4803 17515 4890 17751
rect 5126 17515 5213 17751
rect 5449 17515 5536 17751
rect 5772 17515 5859 17751
rect 6095 17515 6182 17751
rect 6418 17515 6505 17751
rect 6741 17515 6828 17751
rect 7064 17515 7150 17751
rect 7386 17515 7472 17751
rect 7708 17515 7794 17751
rect 8030 17515 8116 17751
rect 8352 17515 8438 17751
rect 8674 17515 8760 17751
rect 8996 17515 9082 17751
rect 9318 17515 9404 17751
rect 9640 17515 9726 17751
rect 9962 17515 10048 17751
rect 10284 17515 10370 17751
rect 10606 17515 10692 17751
rect 10928 17515 11014 17751
rect 11250 17515 11336 17751
rect 11572 17515 11658 17751
rect 11894 17515 11980 17751
rect 12216 17515 12302 17751
rect 12538 17515 12624 17751
rect 12860 17515 12946 17751
rect 13182 17515 13268 17751
rect 13504 17515 13590 17751
rect 13826 17515 13912 17751
rect 14148 17515 14234 17751
rect 14470 17515 14556 17751
rect 14792 17515 14878 17751
rect 15114 17515 15200 17751
rect 15436 17515 15522 17751
rect 15758 17515 15844 17751
rect 16080 17515 16166 17751
rect 16402 17515 16488 17751
rect 16724 17515 16810 17751
rect 17046 17515 17132 17751
rect 17368 17515 17454 17751
rect 17690 17515 17776 17751
rect 18012 17515 18098 17751
rect 18334 17515 18420 17751
rect 18656 17515 18742 17751
rect 18978 17515 19064 17751
rect 19300 17515 19386 17751
rect 19622 17515 19708 17751
rect 19944 17515 20030 17751
rect 20266 17515 20352 17751
rect 20588 17515 20674 17751
rect 20910 17515 20996 17751
rect 21232 17515 21318 17751
rect 21554 17515 21640 17751
rect 21876 17515 21962 17751
rect 22198 17515 22284 17751
rect 22520 17515 22606 17751
rect 22842 17515 22928 17751
rect 23164 17515 23250 17751
rect 23486 17515 23572 17751
rect 23808 17515 23894 17751
rect 24130 17515 24216 17751
rect 24452 17515 24640 17751
rect -3360 17415 24640 17515
rect -3360 17179 -3185 17415
rect -2949 17179 -2862 17415
rect -2626 17179 -2539 17415
rect -2303 17179 -2216 17415
rect -1980 17179 -1893 17415
rect -1657 17179 -1570 17415
rect -1334 17179 -1247 17415
rect -1011 17179 -924 17415
rect -688 17179 -601 17415
rect -365 17179 -278 17415
rect -42 17179 45 17415
rect 281 17179 368 17415
rect 604 17179 691 17415
rect 927 17179 1014 17415
rect 1250 17179 1337 17415
rect 1573 17179 1660 17415
rect 1896 17179 1983 17415
rect 2219 17179 2306 17415
rect 2542 17179 2629 17415
rect 2865 17179 2952 17415
rect 3188 17179 3275 17415
rect 3511 17179 3598 17415
rect 3834 17179 3921 17415
rect 4157 17179 4244 17415
rect 4480 17179 4567 17415
rect 4803 17179 4890 17415
rect 5126 17179 5213 17415
rect 5449 17179 5536 17415
rect 5772 17179 5859 17415
rect 6095 17179 6182 17415
rect 6418 17179 6505 17415
rect 6741 17179 6828 17415
rect 7064 17179 7150 17415
rect 7386 17179 7472 17415
rect 7708 17179 7794 17415
rect 8030 17179 8116 17415
rect 8352 17179 8438 17415
rect 8674 17179 8760 17415
rect 8996 17179 9082 17415
rect 9318 17179 9404 17415
rect 9640 17179 9726 17415
rect 9962 17179 10048 17415
rect 10284 17179 10370 17415
rect 10606 17179 10692 17415
rect 10928 17179 11014 17415
rect 11250 17179 11336 17415
rect 11572 17179 11658 17415
rect 11894 17179 11980 17415
rect 12216 17179 12302 17415
rect 12538 17179 12624 17415
rect 12860 17179 12946 17415
rect 13182 17179 13268 17415
rect 13504 17179 13590 17415
rect 13826 17179 13912 17415
rect 14148 17179 14234 17415
rect 14470 17179 14556 17415
rect 14792 17179 14878 17415
rect 15114 17179 15200 17415
rect 15436 17179 15522 17415
rect 15758 17179 15844 17415
rect 16080 17179 16166 17415
rect 16402 17179 16488 17415
rect 16724 17179 16810 17415
rect 17046 17179 17132 17415
rect 17368 17179 17454 17415
rect 17690 17179 17776 17415
rect 18012 17179 18098 17415
rect 18334 17179 18420 17415
rect 18656 17179 18742 17415
rect 18978 17179 19064 17415
rect 19300 17179 19386 17415
rect 19622 17179 19708 17415
rect 19944 17179 20030 17415
rect 20266 17179 20352 17415
rect 20588 17179 20674 17415
rect 20910 17179 20996 17415
rect 21232 17179 21318 17415
rect 21554 17179 21640 17415
rect 21876 17179 21962 17415
rect 22198 17179 22284 17415
rect 22520 17179 22606 17415
rect 22842 17179 22928 17415
rect 23164 17179 23250 17415
rect 23486 17179 23572 17415
rect 23808 17179 23894 17415
rect 24130 17179 24216 17415
rect 24452 17179 24640 17415
rect -3360 17079 24640 17179
rect -3360 16843 -3185 17079
rect -2949 16843 -2862 17079
rect -2626 16843 -2539 17079
rect -2303 16843 -2216 17079
rect -1980 16843 -1893 17079
rect -1657 16843 -1570 17079
rect -1334 16843 -1247 17079
rect -1011 16843 -924 17079
rect -688 16843 -601 17079
rect -365 16843 -278 17079
rect -42 16843 45 17079
rect 281 16843 368 17079
rect 604 16843 691 17079
rect 927 16843 1014 17079
rect 1250 16843 1337 17079
rect 1573 16843 1660 17079
rect 1896 16843 1983 17079
rect 2219 16843 2306 17079
rect 2542 16843 2629 17079
rect 2865 16843 2952 17079
rect 3188 16843 3275 17079
rect 3511 16843 3598 17079
rect 3834 16843 3921 17079
rect 4157 16843 4244 17079
rect 4480 16843 4567 17079
rect 4803 16843 4890 17079
rect 5126 16843 5213 17079
rect 5449 16843 5536 17079
rect 5772 16843 5859 17079
rect 6095 16843 6182 17079
rect 6418 16843 6505 17079
rect 6741 16843 6828 17079
rect 7064 16843 7150 17079
rect 7386 16843 7472 17079
rect 7708 16843 7794 17079
rect 8030 16843 8116 17079
rect 8352 16843 8438 17079
rect 8674 16843 8760 17079
rect 8996 16843 9082 17079
rect 9318 16843 9404 17079
rect 9640 16843 9726 17079
rect 9962 16843 10048 17079
rect 10284 16843 10370 17079
rect 10606 16843 10692 17079
rect 10928 16843 11014 17079
rect 11250 16843 11336 17079
rect 11572 16843 11658 17079
rect 11894 16843 11980 17079
rect 12216 16843 12302 17079
rect 12538 16843 12624 17079
rect 12860 16843 12946 17079
rect 13182 16843 13268 17079
rect 13504 16843 13590 17079
rect 13826 16843 13912 17079
rect 14148 16843 14234 17079
rect 14470 16843 14556 17079
rect 14792 16843 14878 17079
rect 15114 16843 15200 17079
rect 15436 16843 15522 17079
rect 15758 16843 15844 17079
rect 16080 16843 16166 17079
rect 16402 16843 16488 17079
rect 16724 16843 16810 17079
rect 17046 16843 17132 17079
rect 17368 16843 17454 17079
rect 17690 16843 17776 17079
rect 18012 16843 18098 17079
rect 18334 16843 18420 17079
rect 18656 16843 18742 17079
rect 18978 16843 19064 17079
rect 19300 16843 19386 17079
rect 19622 16843 19708 17079
rect 19944 16843 20030 17079
rect 20266 16843 20352 17079
rect 20588 16843 20674 17079
rect 20910 16843 20996 17079
rect 21232 16843 21318 17079
rect 21554 16843 21640 17079
rect 21876 16843 21962 17079
rect 22198 16843 22284 17079
rect 22520 16843 22606 17079
rect 22842 16843 22928 17079
rect 23164 16843 23250 17079
rect 23486 16843 23572 17079
rect 23808 16843 23894 17079
rect 24130 16843 24216 17079
rect 24452 16843 24640 17079
rect -3360 16743 24640 16843
rect -3360 16507 -3185 16743
rect -2949 16507 -2862 16743
rect -2626 16507 -2539 16743
rect -2303 16507 -2216 16743
rect -1980 16507 -1893 16743
rect -1657 16507 -1570 16743
rect -1334 16507 -1247 16743
rect -1011 16507 -924 16743
rect -688 16507 -601 16743
rect -365 16507 -278 16743
rect -42 16507 45 16743
rect 281 16507 368 16743
rect 604 16507 691 16743
rect 927 16507 1014 16743
rect 1250 16507 1337 16743
rect 1573 16507 1660 16743
rect 1896 16507 1983 16743
rect 2219 16507 2306 16743
rect 2542 16507 2629 16743
rect 2865 16507 2952 16743
rect 3188 16507 3275 16743
rect 3511 16507 3598 16743
rect 3834 16507 3921 16743
rect 4157 16507 4244 16743
rect 4480 16507 4567 16743
rect 4803 16507 4890 16743
rect 5126 16507 5213 16743
rect 5449 16507 5536 16743
rect 5772 16507 5859 16743
rect 6095 16507 6182 16743
rect 6418 16507 6505 16743
rect 6741 16507 6828 16743
rect 7064 16507 7150 16743
rect 7386 16507 7472 16743
rect 7708 16507 7794 16743
rect 8030 16507 8116 16743
rect 8352 16507 8438 16743
rect 8674 16507 8760 16743
rect 8996 16507 9082 16743
rect 9318 16507 9404 16743
rect 9640 16507 9726 16743
rect 9962 16507 10048 16743
rect 10284 16507 10370 16743
rect 10606 16507 10692 16743
rect 10928 16507 11014 16743
rect 11250 16507 11336 16743
rect 11572 16507 11658 16743
rect 11894 16507 11980 16743
rect 12216 16507 12302 16743
rect 12538 16507 12624 16743
rect 12860 16507 12946 16743
rect 13182 16507 13268 16743
rect 13504 16507 13590 16743
rect 13826 16507 13912 16743
rect 14148 16507 14234 16743
rect 14470 16507 14556 16743
rect 14792 16507 14878 16743
rect 15114 16507 15200 16743
rect 15436 16507 15522 16743
rect 15758 16507 15844 16743
rect 16080 16507 16166 16743
rect 16402 16507 16488 16743
rect 16724 16507 16810 16743
rect 17046 16507 17132 16743
rect 17368 16507 17454 16743
rect 17690 16507 17776 16743
rect 18012 16507 18098 16743
rect 18334 16507 18420 16743
rect 18656 16507 18742 16743
rect 18978 16507 19064 16743
rect 19300 16507 19386 16743
rect 19622 16507 19708 16743
rect 19944 16507 20030 16743
rect 20266 16507 20352 16743
rect 20588 16507 20674 16743
rect 20910 16507 20996 16743
rect 21232 16507 21318 16743
rect 21554 16507 21640 16743
rect 21876 16507 21962 16743
rect 22198 16507 22284 16743
rect 22520 16507 22606 16743
rect 22842 16507 22928 16743
rect 23164 16507 23250 16743
rect 23486 16507 23572 16743
rect 23808 16507 23894 16743
rect 24130 16507 24216 16743
rect 24452 16507 24640 16743
rect -3360 16407 24640 16507
rect -3360 16171 -3185 16407
rect -2949 16171 -2862 16407
rect -2626 16171 -2539 16407
rect -2303 16171 -2216 16407
rect -1980 16171 -1893 16407
rect -1657 16171 -1570 16407
rect -1334 16171 -1247 16407
rect -1011 16171 -924 16407
rect -688 16171 -601 16407
rect -365 16171 -278 16407
rect -42 16171 45 16407
rect 281 16171 368 16407
rect 604 16171 691 16407
rect 927 16171 1014 16407
rect 1250 16171 1337 16407
rect 1573 16171 1660 16407
rect 1896 16171 1983 16407
rect 2219 16171 2306 16407
rect 2542 16171 2629 16407
rect 2865 16171 2952 16407
rect 3188 16171 3275 16407
rect 3511 16171 3598 16407
rect 3834 16171 3921 16407
rect 4157 16171 4244 16407
rect 4480 16171 4567 16407
rect 4803 16171 4890 16407
rect 5126 16171 5213 16407
rect 5449 16171 5536 16407
rect 5772 16171 5859 16407
rect 6095 16171 6182 16407
rect 6418 16171 6505 16407
rect 6741 16171 6828 16407
rect 7064 16171 7150 16407
rect 7386 16171 7472 16407
rect 7708 16171 7794 16407
rect 8030 16171 8116 16407
rect 8352 16171 8438 16407
rect 8674 16171 8760 16407
rect 8996 16171 9082 16407
rect 9318 16171 9404 16407
rect 9640 16171 9726 16407
rect 9962 16171 10048 16407
rect 10284 16171 10370 16407
rect 10606 16171 10692 16407
rect 10928 16171 11014 16407
rect 11250 16171 11336 16407
rect 11572 16171 11658 16407
rect 11894 16171 11980 16407
rect 12216 16171 12302 16407
rect 12538 16171 12624 16407
rect 12860 16171 12946 16407
rect 13182 16171 13268 16407
rect 13504 16171 13590 16407
rect 13826 16171 13912 16407
rect 14148 16171 14234 16407
rect 14470 16171 14556 16407
rect 14792 16171 14878 16407
rect 15114 16171 15200 16407
rect 15436 16171 15522 16407
rect 15758 16171 15844 16407
rect 16080 16171 16166 16407
rect 16402 16171 16488 16407
rect 16724 16171 16810 16407
rect 17046 16171 17132 16407
rect 17368 16171 17454 16407
rect 17690 16171 17776 16407
rect 18012 16171 18098 16407
rect 18334 16171 18420 16407
rect 18656 16171 18742 16407
rect 18978 16171 19064 16407
rect 19300 16171 19386 16407
rect 19622 16171 19708 16407
rect 19944 16171 20030 16407
rect 20266 16171 20352 16407
rect 20588 16171 20674 16407
rect 20910 16171 20996 16407
rect 21232 16171 21318 16407
rect 21554 16171 21640 16407
rect 21876 16171 21962 16407
rect 22198 16171 22284 16407
rect 22520 16171 22606 16407
rect 22842 16171 22928 16407
rect 23164 16171 23250 16407
rect 23486 16171 23572 16407
rect 23808 16171 23894 16407
rect 24130 16171 24216 16407
rect 24452 16171 24640 16407
rect -3360 16071 24640 16171
rect -3360 15835 -3185 16071
rect -2949 15835 -2862 16071
rect -2626 15835 -2539 16071
rect -2303 15835 -2216 16071
rect -1980 15835 -1893 16071
rect -1657 15835 -1570 16071
rect -1334 15835 -1247 16071
rect -1011 15835 -924 16071
rect -688 15835 -601 16071
rect -365 15835 -278 16071
rect -42 15835 45 16071
rect 281 15835 368 16071
rect 604 15835 691 16071
rect 927 15835 1014 16071
rect 1250 15835 1337 16071
rect 1573 15835 1660 16071
rect 1896 15835 1983 16071
rect 2219 15835 2306 16071
rect 2542 15835 2629 16071
rect 2865 15835 2952 16071
rect 3188 15835 3275 16071
rect 3511 15835 3598 16071
rect 3834 15835 3921 16071
rect 4157 15835 4244 16071
rect 4480 15835 4567 16071
rect 4803 15835 4890 16071
rect 5126 15835 5213 16071
rect 5449 15835 5536 16071
rect 5772 15835 5859 16071
rect 6095 15835 6182 16071
rect 6418 15835 6505 16071
rect 6741 15835 6828 16071
rect 7064 15835 7150 16071
rect 7386 15835 7472 16071
rect 7708 15835 7794 16071
rect 8030 15835 8116 16071
rect 8352 15835 8438 16071
rect 8674 15835 8760 16071
rect 8996 15835 9082 16071
rect 9318 15835 9404 16071
rect 9640 15835 9726 16071
rect 9962 15835 10048 16071
rect 10284 15835 10370 16071
rect 10606 15835 10692 16071
rect 10928 15835 11014 16071
rect 11250 15835 11336 16071
rect 11572 15835 11658 16071
rect 11894 15835 11980 16071
rect 12216 15835 12302 16071
rect 12538 15835 12624 16071
rect 12860 15835 12946 16071
rect 13182 15835 13268 16071
rect 13504 15835 13590 16071
rect 13826 15835 13912 16071
rect 14148 15835 14234 16071
rect 14470 15835 14556 16071
rect 14792 15835 14878 16071
rect 15114 15835 15200 16071
rect 15436 15835 15522 16071
rect 15758 15835 15844 16071
rect 16080 15835 16166 16071
rect 16402 15835 16488 16071
rect 16724 15835 16810 16071
rect 17046 15835 17132 16071
rect 17368 15835 17454 16071
rect 17690 15835 17776 16071
rect 18012 15835 18098 16071
rect 18334 15835 18420 16071
rect 18656 15835 18742 16071
rect 18978 15835 19064 16071
rect 19300 15835 19386 16071
rect 19622 15835 19708 16071
rect 19944 15835 20030 16071
rect 20266 15835 20352 16071
rect 20588 15835 20674 16071
rect 20910 15835 20996 16071
rect 21232 15835 21318 16071
rect 21554 15835 21640 16071
rect 21876 15835 21962 16071
rect 22198 15835 22284 16071
rect 22520 15835 22606 16071
rect 22842 15835 22928 16071
rect 23164 15835 23250 16071
rect 23486 15835 23572 16071
rect 23808 15835 23894 16071
rect 24130 15835 24216 16071
rect 24452 15835 24640 16071
rect -3360 15735 24640 15835
rect -3360 15499 -3185 15735
rect -2949 15499 -2862 15735
rect -2626 15499 -2539 15735
rect -2303 15499 -2216 15735
rect -1980 15499 -1893 15735
rect -1657 15499 -1570 15735
rect -1334 15499 -1247 15735
rect -1011 15499 -924 15735
rect -688 15499 -601 15735
rect -365 15499 -278 15735
rect -42 15499 45 15735
rect 281 15499 368 15735
rect 604 15499 691 15735
rect 927 15499 1014 15735
rect 1250 15499 1337 15735
rect 1573 15499 1660 15735
rect 1896 15499 1983 15735
rect 2219 15499 2306 15735
rect 2542 15499 2629 15735
rect 2865 15499 2952 15735
rect 3188 15499 3275 15735
rect 3511 15499 3598 15735
rect 3834 15499 3921 15735
rect 4157 15499 4244 15735
rect 4480 15499 4567 15735
rect 4803 15499 4890 15735
rect 5126 15499 5213 15735
rect 5449 15499 5536 15735
rect 5772 15499 5859 15735
rect 6095 15499 6182 15735
rect 6418 15499 6505 15735
rect 6741 15499 6828 15735
rect 7064 15499 7150 15735
rect 7386 15499 7472 15735
rect 7708 15499 7794 15735
rect 8030 15499 8116 15735
rect 8352 15499 8438 15735
rect 8674 15499 8760 15735
rect 8996 15499 9082 15735
rect 9318 15499 9404 15735
rect 9640 15499 9726 15735
rect 9962 15499 10048 15735
rect 10284 15499 10370 15735
rect 10606 15499 10692 15735
rect 10928 15499 11014 15735
rect 11250 15499 11336 15735
rect 11572 15499 11658 15735
rect 11894 15499 11980 15735
rect 12216 15499 12302 15735
rect 12538 15499 12624 15735
rect 12860 15499 12946 15735
rect 13182 15499 13268 15735
rect 13504 15499 13590 15735
rect 13826 15499 13912 15735
rect 14148 15499 14234 15735
rect 14470 15499 14556 15735
rect 14792 15499 14878 15735
rect 15114 15499 15200 15735
rect 15436 15499 15522 15735
rect 15758 15499 15844 15735
rect 16080 15499 16166 15735
rect 16402 15499 16488 15735
rect 16724 15499 16810 15735
rect 17046 15499 17132 15735
rect 17368 15499 17454 15735
rect 17690 15499 17776 15735
rect 18012 15499 18098 15735
rect 18334 15499 18420 15735
rect 18656 15499 18742 15735
rect 18978 15499 19064 15735
rect 19300 15499 19386 15735
rect 19622 15499 19708 15735
rect 19944 15499 20030 15735
rect 20266 15499 20352 15735
rect 20588 15499 20674 15735
rect 20910 15499 20996 15735
rect 21232 15499 21318 15735
rect 21554 15499 21640 15735
rect 21876 15499 21962 15735
rect 22198 15499 22284 15735
rect 22520 15499 22606 15735
rect 22842 15499 22928 15735
rect 23164 15499 23250 15735
rect 23486 15499 23572 15735
rect 23808 15499 23894 15735
rect 24130 15499 24216 15735
rect 24452 15499 24640 15735
rect -3360 15399 24640 15499
rect -3360 15163 -3185 15399
rect -2949 15163 -2862 15399
rect -2626 15163 -2539 15399
rect -2303 15163 -2216 15399
rect -1980 15163 -1893 15399
rect -1657 15163 -1570 15399
rect -1334 15163 -1247 15399
rect -1011 15163 -924 15399
rect -688 15163 -601 15399
rect -365 15163 -278 15399
rect -42 15163 45 15399
rect 281 15163 368 15399
rect 604 15163 691 15399
rect 927 15163 1014 15399
rect 1250 15163 1337 15399
rect 1573 15163 1660 15399
rect 1896 15163 1983 15399
rect 2219 15163 2306 15399
rect 2542 15163 2629 15399
rect 2865 15163 2952 15399
rect 3188 15163 3275 15399
rect 3511 15163 3598 15399
rect 3834 15163 3921 15399
rect 4157 15163 4244 15399
rect 4480 15163 4567 15399
rect 4803 15163 4890 15399
rect 5126 15163 5213 15399
rect 5449 15163 5536 15399
rect 5772 15163 5859 15399
rect 6095 15163 6182 15399
rect 6418 15163 6505 15399
rect 6741 15163 6828 15399
rect 7064 15163 7150 15399
rect 7386 15163 7472 15399
rect 7708 15163 7794 15399
rect 8030 15163 8116 15399
rect 8352 15163 8438 15399
rect 8674 15163 8760 15399
rect 8996 15163 9082 15399
rect 9318 15163 9404 15399
rect 9640 15163 9726 15399
rect 9962 15163 10048 15399
rect 10284 15163 10370 15399
rect 10606 15163 10692 15399
rect 10928 15163 11014 15399
rect 11250 15163 11336 15399
rect 11572 15163 11658 15399
rect 11894 15163 11980 15399
rect 12216 15163 12302 15399
rect 12538 15163 12624 15399
rect 12860 15163 12946 15399
rect 13182 15163 13268 15399
rect 13504 15163 13590 15399
rect 13826 15163 13912 15399
rect 14148 15163 14234 15399
rect 14470 15163 14556 15399
rect 14792 15163 14878 15399
rect 15114 15163 15200 15399
rect 15436 15163 15522 15399
rect 15758 15163 15844 15399
rect 16080 15163 16166 15399
rect 16402 15163 16488 15399
rect 16724 15163 16810 15399
rect 17046 15163 17132 15399
rect 17368 15163 17454 15399
rect 17690 15163 17776 15399
rect 18012 15163 18098 15399
rect 18334 15163 18420 15399
rect 18656 15163 18742 15399
rect 18978 15163 19064 15399
rect 19300 15163 19386 15399
rect 19622 15163 19708 15399
rect 19944 15163 20030 15399
rect 20266 15163 20352 15399
rect 20588 15163 20674 15399
rect 20910 15163 20996 15399
rect 21232 15163 21318 15399
rect 21554 15163 21640 15399
rect 21876 15163 21962 15399
rect 22198 15163 22284 15399
rect 22520 15163 22606 15399
rect 22842 15163 22928 15399
rect 23164 15163 23250 15399
rect 23486 15163 23572 15399
rect 23808 15163 23894 15399
rect 24130 15163 24216 15399
rect 24452 15163 24640 15399
rect -3360 15063 24640 15163
rect -3360 14827 -3185 15063
rect -2949 14827 -2862 15063
rect -2626 14827 -2539 15063
rect -2303 14827 -2216 15063
rect -1980 14827 -1893 15063
rect -1657 14827 -1570 15063
rect -1334 14827 -1247 15063
rect -1011 14827 -924 15063
rect -688 14827 -601 15063
rect -365 14827 -278 15063
rect -42 14827 45 15063
rect 281 14827 368 15063
rect 604 14827 691 15063
rect 927 14827 1014 15063
rect 1250 14827 1337 15063
rect 1573 14827 1660 15063
rect 1896 14827 1983 15063
rect 2219 14827 2306 15063
rect 2542 14827 2629 15063
rect 2865 14827 2952 15063
rect 3188 14827 3275 15063
rect 3511 14827 3598 15063
rect 3834 14827 3921 15063
rect 4157 14827 4244 15063
rect 4480 14827 4567 15063
rect 4803 14827 4890 15063
rect 5126 14827 5213 15063
rect 5449 14827 5536 15063
rect 5772 14827 5859 15063
rect 6095 14827 6182 15063
rect 6418 14827 6505 15063
rect 6741 14827 6828 15063
rect 7064 14827 7150 15063
rect 7386 14827 7472 15063
rect 7708 14827 7794 15063
rect 8030 14827 8116 15063
rect 8352 14827 8438 15063
rect 8674 14827 8760 15063
rect 8996 14827 9082 15063
rect 9318 14827 9404 15063
rect 9640 14827 9726 15063
rect 9962 14827 10048 15063
rect 10284 14827 10370 15063
rect 10606 14827 10692 15063
rect 10928 14827 11014 15063
rect 11250 14827 11336 15063
rect 11572 14827 11658 15063
rect 11894 14827 11980 15063
rect 12216 14827 12302 15063
rect 12538 14827 12624 15063
rect 12860 14827 12946 15063
rect 13182 14827 13268 15063
rect 13504 14827 13590 15063
rect 13826 14827 13912 15063
rect 14148 14827 14234 15063
rect 14470 14827 14556 15063
rect 14792 14827 14878 15063
rect 15114 14827 15200 15063
rect 15436 14827 15522 15063
rect 15758 14827 15844 15063
rect 16080 14827 16166 15063
rect 16402 14827 16488 15063
rect 16724 14827 16810 15063
rect 17046 14827 17132 15063
rect 17368 14827 17454 15063
rect 17690 14827 17776 15063
rect 18012 14827 18098 15063
rect 18334 14827 18420 15063
rect 18656 14827 18742 15063
rect 18978 14827 19064 15063
rect 19300 14827 19386 15063
rect 19622 14827 19708 15063
rect 19944 14827 20030 15063
rect 20266 14827 20352 15063
rect 20588 14827 20674 15063
rect 20910 14827 20996 15063
rect 21232 14827 21318 15063
rect 21554 14827 21640 15063
rect 21876 14827 21962 15063
rect 22198 14827 22284 15063
rect 22520 14827 22606 15063
rect 22842 14827 22928 15063
rect 23164 14827 23250 15063
rect 23486 14827 23572 15063
rect 23808 14827 23894 15063
rect 24130 14827 24216 15063
rect 24452 14827 24640 15063
rect -3360 14727 24640 14827
rect -3360 14491 -3185 14727
rect -2949 14491 -2862 14727
rect -2626 14491 -2539 14727
rect -2303 14491 -2216 14727
rect -1980 14491 -1893 14727
rect -1657 14491 -1570 14727
rect -1334 14491 -1247 14727
rect -1011 14491 -924 14727
rect -688 14491 -601 14727
rect -365 14491 -278 14727
rect -42 14491 45 14727
rect 281 14491 368 14727
rect 604 14491 691 14727
rect 927 14491 1014 14727
rect 1250 14491 1337 14727
rect 1573 14491 1660 14727
rect 1896 14491 1983 14727
rect 2219 14491 2306 14727
rect 2542 14491 2629 14727
rect 2865 14491 2952 14727
rect 3188 14491 3275 14727
rect 3511 14491 3598 14727
rect 3834 14491 3921 14727
rect 4157 14491 4244 14727
rect 4480 14491 4567 14727
rect 4803 14491 4890 14727
rect 5126 14491 5213 14727
rect 5449 14491 5536 14727
rect 5772 14491 5859 14727
rect 6095 14491 6182 14727
rect 6418 14491 6505 14727
rect 6741 14491 6828 14727
rect 7064 14491 7150 14727
rect 7386 14491 7472 14727
rect 7708 14491 7794 14727
rect 8030 14491 8116 14727
rect 8352 14491 8438 14727
rect 8674 14491 8760 14727
rect 8996 14491 9082 14727
rect 9318 14491 9404 14727
rect 9640 14491 9726 14727
rect 9962 14491 10048 14727
rect 10284 14491 10370 14727
rect 10606 14491 10692 14727
rect 10928 14491 11014 14727
rect 11250 14491 11336 14727
rect 11572 14491 11658 14727
rect 11894 14491 11980 14727
rect 12216 14491 12302 14727
rect 12538 14491 12624 14727
rect 12860 14491 12946 14727
rect 13182 14491 13268 14727
rect 13504 14491 13590 14727
rect 13826 14491 13912 14727
rect 14148 14491 14234 14727
rect 14470 14491 14556 14727
rect 14792 14491 14878 14727
rect 15114 14491 15200 14727
rect 15436 14491 15522 14727
rect 15758 14491 15844 14727
rect 16080 14491 16166 14727
rect 16402 14491 16488 14727
rect 16724 14491 16810 14727
rect 17046 14491 17132 14727
rect 17368 14491 17454 14727
rect 17690 14491 17776 14727
rect 18012 14491 18098 14727
rect 18334 14491 18420 14727
rect 18656 14491 18742 14727
rect 18978 14491 19064 14727
rect 19300 14491 19386 14727
rect 19622 14491 19708 14727
rect 19944 14491 20030 14727
rect 20266 14491 20352 14727
rect 20588 14491 20674 14727
rect 20910 14491 20996 14727
rect 21232 14491 21318 14727
rect 21554 14491 21640 14727
rect 21876 14491 21962 14727
rect 22198 14491 22284 14727
rect 22520 14491 22606 14727
rect 22842 14491 22928 14727
rect 23164 14491 23250 14727
rect 23486 14491 23572 14727
rect 23808 14491 23894 14727
rect 24130 14491 24216 14727
rect 24452 14491 24640 14727
rect -3360 14391 24640 14491
rect -3360 14155 -3185 14391
rect -2949 14155 -2862 14391
rect -2626 14155 -2539 14391
rect -2303 14155 -2216 14391
rect -1980 14155 -1893 14391
rect -1657 14155 -1570 14391
rect -1334 14155 -1247 14391
rect -1011 14155 -924 14391
rect -688 14155 -601 14391
rect -365 14155 -278 14391
rect -42 14155 45 14391
rect 281 14155 368 14391
rect 604 14155 691 14391
rect 927 14155 1014 14391
rect 1250 14155 1337 14391
rect 1573 14155 1660 14391
rect 1896 14155 1983 14391
rect 2219 14155 2306 14391
rect 2542 14155 2629 14391
rect 2865 14155 2952 14391
rect 3188 14155 3275 14391
rect 3511 14155 3598 14391
rect 3834 14155 3921 14391
rect 4157 14155 4244 14391
rect 4480 14155 4567 14391
rect 4803 14155 4890 14391
rect 5126 14155 5213 14391
rect 5449 14155 5536 14391
rect 5772 14155 5859 14391
rect 6095 14155 6182 14391
rect 6418 14155 6505 14391
rect 6741 14155 6828 14391
rect 7064 14155 7150 14391
rect 7386 14155 7472 14391
rect 7708 14155 7794 14391
rect 8030 14155 8116 14391
rect 8352 14155 8438 14391
rect 8674 14155 8760 14391
rect 8996 14155 9082 14391
rect 9318 14155 9404 14391
rect 9640 14155 9726 14391
rect 9962 14155 10048 14391
rect 10284 14155 10370 14391
rect 10606 14155 10692 14391
rect 10928 14155 11014 14391
rect 11250 14155 11336 14391
rect 11572 14155 11658 14391
rect 11894 14155 11980 14391
rect 12216 14155 12302 14391
rect 12538 14155 12624 14391
rect 12860 14155 12946 14391
rect 13182 14155 13268 14391
rect 13504 14155 13590 14391
rect 13826 14155 13912 14391
rect 14148 14155 14234 14391
rect 14470 14155 14556 14391
rect 14792 14155 14878 14391
rect 15114 14155 15200 14391
rect 15436 14155 15522 14391
rect 15758 14155 15844 14391
rect 16080 14155 16166 14391
rect 16402 14155 16488 14391
rect 16724 14155 16810 14391
rect 17046 14155 17132 14391
rect 17368 14155 17454 14391
rect 17690 14155 17776 14391
rect 18012 14155 18098 14391
rect 18334 14155 18420 14391
rect 18656 14155 18742 14391
rect 18978 14155 19064 14391
rect 19300 14155 19386 14391
rect 19622 14155 19708 14391
rect 19944 14155 20030 14391
rect 20266 14155 20352 14391
rect 20588 14155 20674 14391
rect 20910 14155 20996 14391
rect 21232 14155 21318 14391
rect 21554 14155 21640 14391
rect 21876 14155 21962 14391
rect 22198 14155 22284 14391
rect 22520 14155 22606 14391
rect 22842 14155 22928 14391
rect 23164 14155 23250 14391
rect 23486 14155 23572 14391
rect 23808 14155 23894 14391
rect 24130 14155 24216 14391
rect 24452 14155 24640 14391
rect -3360 14055 24640 14155
rect -3360 13819 -3185 14055
rect -2949 13819 -2862 14055
rect -2626 13819 -2539 14055
rect -2303 13819 -2216 14055
rect -1980 13819 -1893 14055
rect -1657 13819 -1570 14055
rect -1334 13819 -1247 14055
rect -1011 13819 -924 14055
rect -688 13819 -601 14055
rect -365 13819 -278 14055
rect -42 13819 45 14055
rect 281 13819 368 14055
rect 604 13819 691 14055
rect 927 13819 1014 14055
rect 1250 13819 1337 14055
rect 1573 13819 1660 14055
rect 1896 13819 1983 14055
rect 2219 13819 2306 14055
rect 2542 13819 2629 14055
rect 2865 13819 2952 14055
rect 3188 13819 3275 14055
rect 3511 13819 3598 14055
rect 3834 13819 3921 14055
rect 4157 13819 4244 14055
rect 4480 13819 4567 14055
rect 4803 13819 4890 14055
rect 5126 13819 5213 14055
rect 5449 13819 5536 14055
rect 5772 13819 5859 14055
rect 6095 13819 6182 14055
rect 6418 13819 6505 14055
rect 6741 13819 6828 14055
rect 7064 13819 7150 14055
rect 7386 13819 7472 14055
rect 7708 13819 7794 14055
rect 8030 13819 8116 14055
rect 8352 13819 8438 14055
rect 8674 13819 8760 14055
rect 8996 13819 9082 14055
rect 9318 13819 9404 14055
rect 9640 13819 9726 14055
rect 9962 13819 10048 14055
rect 10284 13819 10370 14055
rect 10606 13819 10692 14055
rect 10928 13819 11014 14055
rect 11250 13819 11336 14055
rect 11572 13819 11658 14055
rect 11894 13819 11980 14055
rect 12216 13819 12302 14055
rect 12538 13819 12624 14055
rect 12860 13819 12946 14055
rect 13182 13819 13268 14055
rect 13504 13819 13590 14055
rect 13826 13819 13912 14055
rect 14148 13819 14234 14055
rect 14470 13819 14556 14055
rect 14792 13819 14878 14055
rect 15114 13819 15200 14055
rect 15436 13819 15522 14055
rect 15758 13819 15844 14055
rect 16080 13819 16166 14055
rect 16402 13819 16488 14055
rect 16724 13819 16810 14055
rect 17046 13819 17132 14055
rect 17368 13819 17454 14055
rect 17690 13819 17776 14055
rect 18012 13819 18098 14055
rect 18334 13819 18420 14055
rect 18656 13819 18742 14055
rect 18978 13819 19064 14055
rect 19300 13819 19386 14055
rect 19622 13819 19708 14055
rect 19944 13819 20030 14055
rect 20266 13819 20352 14055
rect 20588 13819 20674 14055
rect 20910 13819 20996 14055
rect 21232 13819 21318 14055
rect 21554 13819 21640 14055
rect 21876 13819 21962 14055
rect 22198 13819 22284 14055
rect 22520 13819 22606 14055
rect 22842 13819 22928 14055
rect 23164 13819 23250 14055
rect 23486 13819 23572 14055
rect 23808 13819 23894 14055
rect 24130 13819 24216 14055
rect 24452 13819 24640 14055
rect -3360 13719 24640 13819
rect -3360 13483 -3185 13719
rect -2949 13483 -2862 13719
rect -2626 13483 -2539 13719
rect -2303 13483 -2216 13719
rect -1980 13483 -1893 13719
rect -1657 13483 -1570 13719
rect -1334 13483 -1247 13719
rect -1011 13483 -924 13719
rect -688 13483 -601 13719
rect -365 13483 -278 13719
rect -42 13483 45 13719
rect 281 13483 368 13719
rect 604 13483 691 13719
rect 927 13483 1014 13719
rect 1250 13483 1337 13719
rect 1573 13483 1660 13719
rect 1896 13483 1983 13719
rect 2219 13483 2306 13719
rect 2542 13483 2629 13719
rect 2865 13483 2952 13719
rect 3188 13483 3275 13719
rect 3511 13483 3598 13719
rect 3834 13483 3921 13719
rect 4157 13483 4244 13719
rect 4480 13483 4567 13719
rect 4803 13483 4890 13719
rect 5126 13483 5213 13719
rect 5449 13483 5536 13719
rect 5772 13483 5859 13719
rect 6095 13483 6182 13719
rect 6418 13483 6505 13719
rect 6741 13483 6828 13719
rect 7064 13483 7150 13719
rect 7386 13483 7472 13719
rect 7708 13483 7794 13719
rect 8030 13483 8116 13719
rect 8352 13483 8438 13719
rect 8674 13483 8760 13719
rect 8996 13483 9082 13719
rect 9318 13483 9404 13719
rect 9640 13483 9726 13719
rect 9962 13483 10048 13719
rect 10284 13483 10370 13719
rect 10606 13483 10692 13719
rect 10928 13483 11014 13719
rect 11250 13483 11336 13719
rect 11572 13483 11658 13719
rect 11894 13483 11980 13719
rect 12216 13483 12302 13719
rect 12538 13483 12624 13719
rect 12860 13483 12946 13719
rect 13182 13483 13268 13719
rect 13504 13483 13590 13719
rect 13826 13483 13912 13719
rect 14148 13483 14234 13719
rect 14470 13483 14556 13719
rect 14792 13483 14878 13719
rect 15114 13483 15200 13719
rect 15436 13483 15522 13719
rect 15758 13483 15844 13719
rect 16080 13483 16166 13719
rect 16402 13483 16488 13719
rect 16724 13483 16810 13719
rect 17046 13483 17132 13719
rect 17368 13483 17454 13719
rect 17690 13483 17776 13719
rect 18012 13483 18098 13719
rect 18334 13483 18420 13719
rect 18656 13483 18742 13719
rect 18978 13483 19064 13719
rect 19300 13483 19386 13719
rect 19622 13483 19708 13719
rect 19944 13483 20030 13719
rect 20266 13483 20352 13719
rect 20588 13483 20674 13719
rect 20910 13483 20996 13719
rect 21232 13483 21318 13719
rect 21554 13483 21640 13719
rect 21876 13483 21962 13719
rect 22198 13483 22284 13719
rect 22520 13483 22606 13719
rect 22842 13483 22928 13719
rect 23164 13483 23250 13719
rect 23486 13483 23572 13719
rect 23808 13483 23894 13719
rect 24130 13483 24216 13719
rect 24452 13483 24640 13719
rect -3360 13458 24640 13483
rect -3360 13114 24640 13138
rect -3360 12878 -3185 13114
rect -2949 12878 -2862 13114
rect -2626 12878 -2539 13114
rect -2303 12878 -2216 13114
rect -1980 12878 -1893 13114
rect -1657 12878 -1570 13114
rect -1334 12878 -1247 13114
rect -1011 12878 -924 13114
rect -688 12878 -601 13114
rect -365 12878 -278 13114
rect -42 12878 45 13114
rect 281 12878 368 13114
rect 604 12878 691 13114
rect 927 12878 1014 13114
rect 1250 12878 1337 13114
rect 1573 12878 1660 13114
rect 1896 12878 1983 13114
rect 2219 12878 2306 13114
rect 2542 12878 2629 13114
rect 2865 12878 2952 13114
rect 3188 12878 3275 13114
rect 3511 12878 3598 13114
rect 3834 12878 3921 13114
rect 4157 12878 4244 13114
rect 4480 12878 4567 13114
rect 4803 12878 4890 13114
rect 5126 12878 5213 13114
rect 5449 12878 5536 13114
rect 5772 12878 5859 13114
rect 6095 12878 6182 13114
rect 6418 12878 6504 13114
rect 6740 12878 6826 13114
rect 7062 12878 7148 13114
rect 7384 12878 7470 13114
rect 7706 12878 7792 13114
rect 8028 12878 8114 13114
rect 8350 12878 8436 13114
rect 8672 12878 8758 13114
rect 8994 12878 9080 13114
rect 9316 12878 9402 13114
rect 9638 12878 9724 13114
rect 9960 12878 10046 13114
rect 10282 12878 10368 13114
rect 10604 12878 10690 13114
rect 10926 12878 11012 13114
rect 11248 12878 11334 13114
rect 11570 12878 11656 13114
rect 11892 12878 11978 13114
rect 12214 12878 12300 13114
rect 12536 12878 12622 13114
rect 12858 12878 12944 13114
rect 13180 12878 13266 13114
rect 13502 12878 13588 13114
rect 13824 12878 13910 13114
rect 14146 12878 14232 13114
rect 14468 12878 14554 13114
rect 14790 12878 14876 13114
rect 15112 12878 15198 13114
rect 15434 12878 15520 13114
rect 15756 12878 15842 13114
rect 16078 12878 16164 13114
rect 16400 12878 16486 13114
rect 16722 12878 16808 13114
rect 17044 12878 17130 13114
rect 17366 12878 17452 13114
rect 17688 12878 17774 13114
rect 18010 12878 18096 13114
rect 18332 12878 18418 13114
rect 18654 12878 18740 13114
rect 18976 12878 19062 13114
rect 19298 12878 19384 13114
rect 19620 12878 19706 13114
rect 19942 12878 20028 13114
rect 20264 12878 20350 13114
rect 20586 12878 20672 13114
rect 20908 12878 20994 13114
rect 21230 12878 21316 13114
rect 21552 12878 21638 13114
rect 21874 12878 21960 13114
rect 22196 12878 22282 13114
rect 22518 12878 22604 13114
rect 22840 12878 22926 13114
rect 23162 12878 23248 13114
rect 23484 12878 23570 13114
rect 23806 12878 23892 13114
rect 24128 12878 24214 13114
rect 24450 12878 24640 13114
rect -3360 12548 24640 12878
rect -3360 12312 -3185 12548
rect -2949 12312 -2862 12548
rect -2626 12312 -2539 12548
rect -2303 12312 -2216 12548
rect -1980 12312 -1893 12548
rect -1657 12312 -1570 12548
rect -1334 12312 -1247 12548
rect -1011 12312 -924 12548
rect -688 12312 -601 12548
rect -365 12312 -278 12548
rect -42 12312 45 12548
rect 281 12312 368 12548
rect 604 12312 691 12548
rect 927 12312 1014 12548
rect 1250 12312 1337 12548
rect 1573 12312 1660 12548
rect 1896 12312 1983 12548
rect 2219 12312 2306 12548
rect 2542 12312 2629 12548
rect 2865 12312 2952 12548
rect 3188 12312 3275 12548
rect 3511 12312 3598 12548
rect 3834 12312 3921 12548
rect 4157 12312 4244 12548
rect 4480 12312 4567 12548
rect 4803 12312 4890 12548
rect 5126 12312 5213 12548
rect 5449 12312 5536 12548
rect 5772 12312 5859 12548
rect 6095 12312 6182 12548
rect 6418 12312 6504 12548
rect 6740 12312 6826 12548
rect 7062 12312 7148 12548
rect 7384 12312 7470 12548
rect 7706 12312 7792 12548
rect 8028 12312 8114 12548
rect 8350 12312 8436 12548
rect 8672 12312 8758 12548
rect 8994 12312 9080 12548
rect 9316 12312 9402 12548
rect 9638 12312 9724 12548
rect 9960 12312 10046 12548
rect 10282 12312 10368 12548
rect 10604 12312 10690 12548
rect 10926 12312 11012 12548
rect 11248 12312 11334 12548
rect 11570 12312 11656 12548
rect 11892 12312 11978 12548
rect 12214 12312 12300 12548
rect 12536 12312 12622 12548
rect 12858 12312 12944 12548
rect 13180 12312 13266 12548
rect 13502 12312 13588 12548
rect 13824 12312 13910 12548
rect 14146 12312 14232 12548
rect 14468 12312 14554 12548
rect 14790 12312 14876 12548
rect 15112 12312 15198 12548
rect 15434 12312 15520 12548
rect 15756 12312 15842 12548
rect 16078 12312 16164 12548
rect 16400 12312 16486 12548
rect 16722 12312 16808 12548
rect 17044 12312 17130 12548
rect 17366 12312 17452 12548
rect 17688 12312 17774 12548
rect 18010 12312 18096 12548
rect 18332 12312 18418 12548
rect 18654 12312 18740 12548
rect 18976 12312 19062 12548
rect 19298 12312 19384 12548
rect 19620 12312 19706 12548
rect 19942 12312 20028 12548
rect 20264 12312 20350 12548
rect 20586 12312 20672 12548
rect 20908 12312 20994 12548
rect 21230 12312 21316 12548
rect 21552 12312 21638 12548
rect 21874 12312 21960 12548
rect 22196 12312 22282 12548
rect 22518 12312 22604 12548
rect 22840 12312 22926 12548
rect 23162 12312 23248 12548
rect 23484 12312 23570 12548
rect 23806 12312 23892 12548
rect 24128 12312 24214 12548
rect 24450 12312 24640 12548
rect -3360 12288 24640 12312
rect -3360 11944 24640 11968
rect -3360 11708 -3185 11944
rect -2949 11708 -2862 11944
rect -2626 11708 -2539 11944
rect -2303 11708 -2216 11944
rect -1980 11708 -1893 11944
rect -1657 11708 -1570 11944
rect -1334 11708 -1247 11944
rect -1011 11708 -924 11944
rect -688 11708 -601 11944
rect -365 11708 -278 11944
rect -42 11708 45 11944
rect 281 11708 368 11944
rect 604 11708 691 11944
rect 927 11708 1014 11944
rect 1250 11708 1337 11944
rect 1573 11708 1660 11944
rect 1896 11708 1983 11944
rect 2219 11708 2306 11944
rect 2542 11708 2629 11944
rect 2865 11708 2952 11944
rect 3188 11708 3275 11944
rect 3511 11708 3598 11944
rect 3834 11708 3921 11944
rect 4157 11708 4244 11944
rect 4480 11708 4567 11944
rect 4803 11708 4890 11944
rect 5126 11708 5213 11944
rect 5449 11708 5536 11944
rect 5772 11708 5859 11944
rect 6095 11708 6182 11944
rect 6418 11708 6504 11944
rect 6740 11708 6826 11944
rect 7062 11708 7148 11944
rect 7384 11708 7470 11944
rect 7706 11708 7792 11944
rect 8028 11708 8114 11944
rect 8350 11708 8436 11944
rect 8672 11708 8758 11944
rect 8994 11708 9080 11944
rect 9316 11708 9402 11944
rect 9638 11708 9724 11944
rect 9960 11708 10046 11944
rect 10282 11708 10368 11944
rect 10604 11708 10690 11944
rect 10926 11708 11012 11944
rect 11248 11708 11334 11944
rect 11570 11708 11656 11944
rect 11892 11708 11978 11944
rect 12214 11708 12300 11944
rect 12536 11708 12622 11944
rect 12858 11708 12944 11944
rect 13180 11708 13266 11944
rect 13502 11708 13588 11944
rect 13824 11708 13910 11944
rect 14146 11708 14232 11944
rect 14468 11708 14554 11944
rect 14790 11708 14876 11944
rect 15112 11708 15198 11944
rect 15434 11708 15520 11944
rect 15756 11708 15842 11944
rect 16078 11708 16164 11944
rect 16400 11708 16486 11944
rect 16722 11708 16808 11944
rect 17044 11708 17130 11944
rect 17366 11708 17452 11944
rect 17688 11708 17774 11944
rect 18010 11708 18096 11944
rect 18332 11708 18418 11944
rect 18654 11708 18740 11944
rect 18976 11708 19062 11944
rect 19298 11708 19384 11944
rect 19620 11708 19706 11944
rect 19942 11708 20028 11944
rect 20264 11708 20350 11944
rect 20586 11708 20672 11944
rect 20908 11708 20994 11944
rect 21230 11708 21316 11944
rect 21552 11708 21638 11944
rect 21874 11708 21960 11944
rect 22196 11708 22282 11944
rect 22518 11708 22604 11944
rect 22840 11708 22926 11944
rect 23162 11708 23248 11944
rect 23484 11708 23570 11944
rect 23806 11708 23892 11944
rect 24128 11708 24214 11944
rect 24450 11708 24640 11944
rect -3360 11378 24640 11708
rect -3360 11142 -3185 11378
rect -2949 11142 -2862 11378
rect -2626 11142 -2539 11378
rect -2303 11142 -2216 11378
rect -1980 11142 -1893 11378
rect -1657 11142 -1570 11378
rect -1334 11142 -1247 11378
rect -1011 11142 -924 11378
rect -688 11142 -601 11378
rect -365 11142 -278 11378
rect -42 11142 45 11378
rect 281 11142 368 11378
rect 604 11142 691 11378
rect 927 11142 1014 11378
rect 1250 11142 1337 11378
rect 1573 11142 1660 11378
rect 1896 11142 1983 11378
rect 2219 11142 2306 11378
rect 2542 11142 2629 11378
rect 2865 11142 2952 11378
rect 3188 11142 3275 11378
rect 3511 11142 3598 11378
rect 3834 11142 3921 11378
rect 4157 11142 4244 11378
rect 4480 11142 4567 11378
rect 4803 11142 4890 11378
rect 5126 11142 5213 11378
rect 5449 11142 5536 11378
rect 5772 11142 5859 11378
rect 6095 11142 6182 11378
rect 6418 11142 6504 11378
rect 6740 11142 6826 11378
rect 7062 11142 7148 11378
rect 7384 11142 7470 11378
rect 7706 11142 7792 11378
rect 8028 11142 8114 11378
rect 8350 11142 8436 11378
rect 8672 11142 8758 11378
rect 8994 11142 9080 11378
rect 9316 11142 9402 11378
rect 9638 11142 9724 11378
rect 9960 11142 10046 11378
rect 10282 11142 10368 11378
rect 10604 11142 10690 11378
rect 10926 11142 11012 11378
rect 11248 11142 11334 11378
rect 11570 11142 11656 11378
rect 11892 11142 11978 11378
rect 12214 11142 12300 11378
rect 12536 11142 12622 11378
rect 12858 11142 12944 11378
rect 13180 11142 13266 11378
rect 13502 11142 13588 11378
rect 13824 11142 13910 11378
rect 14146 11142 14232 11378
rect 14468 11142 14554 11378
rect 14790 11142 14876 11378
rect 15112 11142 15198 11378
rect 15434 11142 15520 11378
rect 15756 11142 15842 11378
rect 16078 11142 16164 11378
rect 16400 11142 16486 11378
rect 16722 11142 16808 11378
rect 17044 11142 17130 11378
rect 17366 11142 17452 11378
rect 17688 11142 17774 11378
rect 18010 11142 18096 11378
rect 18332 11142 18418 11378
rect 18654 11142 18740 11378
rect 18976 11142 19062 11378
rect 19298 11142 19384 11378
rect 19620 11142 19706 11378
rect 19942 11142 20028 11378
rect 20264 11142 20350 11378
rect 20586 11142 20672 11378
rect 20908 11142 20994 11378
rect 21230 11142 21316 11378
rect 21552 11142 21638 11378
rect 21874 11142 21960 11378
rect 22196 11142 22282 11378
rect 22518 11142 22604 11378
rect 22840 11142 22926 11378
rect 23162 11142 23248 11378
rect 23484 11142 23570 11378
rect 23806 11142 23892 11378
rect 24128 11142 24214 11378
rect 24450 11142 24640 11378
rect -3360 11118 24640 11142
rect -3360 8998 -2720 10798
rect 24000 8998 24640 10798
rect -3360 8654 24640 8678
rect -3360 8418 -3185 8654
rect -2949 8418 -2862 8654
rect -2626 8418 -2539 8654
rect -2303 8418 -2216 8654
rect -1980 8418 -1893 8654
rect -1657 8418 -1570 8654
rect -1334 8418 -1247 8654
rect -1011 8418 -924 8654
rect -688 8418 -601 8654
rect -365 8418 -278 8654
rect -42 8418 45 8654
rect 281 8418 368 8654
rect 604 8418 691 8654
rect 927 8418 1014 8654
rect 1250 8418 1337 8654
rect 1573 8418 1660 8654
rect 1896 8418 1983 8654
rect 2219 8418 2306 8654
rect 2542 8418 2629 8654
rect 2865 8418 2952 8654
rect 3188 8418 3275 8654
rect 3511 8418 3598 8654
rect 3834 8418 3921 8654
rect 4157 8418 4244 8654
rect 4480 8418 4567 8654
rect 4803 8418 4890 8654
rect 5126 8418 5213 8654
rect 5449 8418 5536 8654
rect 5772 8418 5859 8654
rect 6095 8418 6182 8654
rect 6418 8418 6505 8654
rect 6741 8418 6828 8654
rect 7064 8418 7150 8654
rect 7386 8418 7472 8654
rect 7708 8418 7794 8654
rect 8030 8418 8116 8654
rect 8352 8418 8438 8654
rect 8674 8418 8760 8654
rect 8996 8418 9082 8654
rect 9318 8418 9404 8654
rect 9640 8418 9726 8654
rect 9962 8418 10048 8654
rect 10284 8418 10370 8654
rect 10606 8418 10692 8654
rect 10928 8418 11014 8654
rect 11250 8418 11336 8654
rect 11572 8418 11658 8654
rect 11894 8418 11980 8654
rect 12216 8418 12302 8654
rect 12538 8418 12624 8654
rect 12860 8418 12946 8654
rect 13182 8418 13268 8654
rect 13504 8418 13590 8654
rect 13826 8418 13912 8654
rect 14148 8418 14234 8654
rect 14470 8418 14556 8654
rect 14792 8418 14878 8654
rect 15114 8418 15200 8654
rect 15436 8418 15522 8654
rect 15758 8418 15844 8654
rect 16080 8418 16166 8654
rect 16402 8418 16488 8654
rect 16724 8418 16810 8654
rect 17046 8418 17132 8654
rect 17368 8418 17454 8654
rect 17690 8418 17776 8654
rect 18012 8418 18098 8654
rect 18334 8418 18420 8654
rect 18656 8418 18742 8654
rect 18978 8418 19064 8654
rect 19300 8418 19386 8654
rect 19622 8418 19708 8654
rect 19944 8418 20030 8654
rect 20266 8418 20352 8654
rect 20588 8418 20674 8654
rect 20910 8418 20996 8654
rect 21232 8418 21318 8654
rect 21554 8418 21640 8654
rect 21876 8418 21962 8654
rect 22198 8418 22284 8654
rect 22520 8418 22606 8654
rect 22842 8418 22928 8654
rect 23164 8418 23250 8654
rect 23486 8418 23572 8654
rect 23808 8418 23894 8654
rect 24130 8418 24216 8654
rect 24452 8418 24640 8654
rect -3360 8048 24640 8418
rect -3360 7812 -3185 8048
rect -2949 7812 -2862 8048
rect -2626 7812 -2539 8048
rect -2303 7812 -2216 8048
rect -1980 7812 -1893 8048
rect -1657 7812 -1570 8048
rect -1334 7812 -1247 8048
rect -1011 7812 -924 8048
rect -688 7812 -601 8048
rect -365 7812 -278 8048
rect -42 7812 45 8048
rect 281 7812 368 8048
rect 604 7812 691 8048
rect 927 7812 1014 8048
rect 1250 7812 1337 8048
rect 1573 7812 1660 8048
rect 1896 7812 1983 8048
rect 2219 7812 2306 8048
rect 2542 7812 2629 8048
rect 2865 7812 2952 8048
rect 3188 7812 3275 8048
rect 3511 7812 3598 8048
rect 3834 7812 3921 8048
rect 4157 7812 4244 8048
rect 4480 7812 4567 8048
rect 4803 7812 4890 8048
rect 5126 7812 5213 8048
rect 5449 7812 5536 8048
rect 5772 7812 5859 8048
rect 6095 7812 6182 8048
rect 6418 7812 6505 8048
rect 6741 7812 6828 8048
rect 7064 7812 7150 8048
rect 7386 7812 7472 8048
rect 7708 7812 7794 8048
rect 8030 7812 8116 8048
rect 8352 7812 8438 8048
rect 8674 7812 8760 8048
rect 8996 7812 9082 8048
rect 9318 7812 9404 8048
rect 9640 7812 9726 8048
rect 9962 7812 10048 8048
rect 10284 7812 10370 8048
rect 10606 7812 10692 8048
rect 10928 7812 11014 8048
rect 11250 7812 11336 8048
rect 11572 7812 11658 8048
rect 11894 7812 11980 8048
rect 12216 7812 12302 8048
rect 12538 7812 12624 8048
rect 12860 7812 12946 8048
rect 13182 7812 13268 8048
rect 13504 7812 13590 8048
rect 13826 7812 13912 8048
rect 14148 7812 14234 8048
rect 14470 7812 14556 8048
rect 14792 7812 14878 8048
rect 15114 7812 15200 8048
rect 15436 7812 15522 8048
rect 15758 7812 15844 8048
rect 16080 7812 16166 8048
rect 16402 7812 16488 8048
rect 16724 7812 16810 8048
rect 17046 7812 17132 8048
rect 17368 7812 17454 8048
rect 17690 7812 17776 8048
rect 18012 7812 18098 8048
rect 18334 7812 18420 8048
rect 18656 7812 18742 8048
rect 18978 7812 19064 8048
rect 19300 7812 19386 8048
rect 19622 7812 19708 8048
rect 19944 7812 20030 8048
rect 20266 7812 20352 8048
rect 20588 7812 20674 8048
rect 20910 7812 20996 8048
rect 21232 7812 21318 8048
rect 21554 7812 21640 8048
rect 21876 7812 21962 8048
rect 22198 7812 22284 8048
rect 22520 7812 22606 8048
rect 22842 7812 22928 8048
rect 23164 7812 23250 8048
rect 23486 7812 23572 8048
rect 23808 7812 23894 8048
rect 24130 7812 24216 8048
rect 24452 7812 24640 8048
rect -3360 7788 24640 7812
rect -3360 7444 24640 7468
rect -3360 7208 -3185 7444
rect -2949 7208 -2862 7444
rect -2626 7208 -2539 7444
rect -2303 7208 -2216 7444
rect -1980 7208 -1893 7444
rect -1657 7208 -1570 7444
rect -1334 7208 -1247 7444
rect -1011 7208 -924 7444
rect -688 7208 -601 7444
rect -365 7208 -278 7444
rect -42 7208 45 7444
rect 281 7208 368 7444
rect 604 7208 691 7444
rect 927 7208 1014 7444
rect 1250 7208 1337 7444
rect 1573 7208 1660 7444
rect 1896 7208 1983 7444
rect 2219 7208 2306 7444
rect 2542 7208 2629 7444
rect 2865 7208 2952 7444
rect 3188 7208 3275 7444
rect 3511 7208 3598 7444
rect 3834 7208 3921 7444
rect 4157 7208 4244 7444
rect 4480 7208 4567 7444
rect 4803 7208 4890 7444
rect 5126 7208 5213 7444
rect 5449 7208 5536 7444
rect 5772 7208 5859 7444
rect 6095 7208 6182 7444
rect 6418 7208 6505 7444
rect 6741 7208 6828 7444
rect 7064 7208 7150 7444
rect 7386 7208 7472 7444
rect 7708 7208 7794 7444
rect 8030 7208 8116 7444
rect 8352 7208 8438 7444
rect 8674 7208 8760 7444
rect 8996 7208 9082 7444
rect 9318 7208 9404 7444
rect 9640 7208 9726 7444
rect 9962 7208 10048 7444
rect 10284 7208 10370 7444
rect 10606 7208 10692 7444
rect 10928 7208 11014 7444
rect 11250 7208 11336 7444
rect 11572 7208 11658 7444
rect 11894 7208 11980 7444
rect 12216 7208 12302 7444
rect 12538 7208 12624 7444
rect 12860 7208 12946 7444
rect 13182 7208 13268 7444
rect 13504 7208 13590 7444
rect 13826 7208 13912 7444
rect 14148 7208 14234 7444
rect 14470 7208 14556 7444
rect 14792 7208 14878 7444
rect 15114 7208 15200 7444
rect 15436 7208 15522 7444
rect 15758 7208 15844 7444
rect 16080 7208 16166 7444
rect 16402 7208 16488 7444
rect 16724 7208 16810 7444
rect 17046 7208 17132 7444
rect 17368 7208 17454 7444
rect 17690 7208 17776 7444
rect 18012 7208 18098 7444
rect 18334 7208 18420 7444
rect 18656 7208 18742 7444
rect 18978 7208 19064 7444
rect 19300 7208 19386 7444
rect 19622 7208 19708 7444
rect 19944 7208 20030 7444
rect 20266 7208 20352 7444
rect 20588 7208 20674 7444
rect 20910 7208 20996 7444
rect 21232 7208 21318 7444
rect 21554 7208 21640 7444
rect 21876 7208 21962 7444
rect 22198 7208 22284 7444
rect 22520 7208 22606 7444
rect 22842 7208 22928 7444
rect 23164 7208 23250 7444
rect 23486 7208 23572 7444
rect 23808 7208 23894 7444
rect 24130 7208 24216 7444
rect 24452 7208 24640 7444
rect -3360 7078 24640 7208
rect -3360 6842 -3185 7078
rect -2949 6842 -2862 7078
rect -2626 6842 -2539 7078
rect -2303 6842 -2216 7078
rect -1980 6842 -1893 7078
rect -1657 6842 -1570 7078
rect -1334 6842 -1247 7078
rect -1011 6842 -924 7078
rect -688 6842 -601 7078
rect -365 6842 -278 7078
rect -42 6842 45 7078
rect 281 6842 368 7078
rect 604 6842 691 7078
rect 927 6842 1014 7078
rect 1250 6842 1337 7078
rect 1573 6842 1660 7078
rect 1896 6842 1983 7078
rect 2219 6842 2306 7078
rect 2542 6842 2629 7078
rect 2865 6842 2952 7078
rect 3188 6842 3275 7078
rect 3511 6842 3598 7078
rect 3834 6842 3921 7078
rect 4157 6842 4244 7078
rect 4480 6842 4567 7078
rect 4803 6842 4890 7078
rect 5126 6842 5213 7078
rect 5449 6842 5536 7078
rect 5772 6842 5859 7078
rect 6095 6842 6182 7078
rect 6418 6842 6505 7078
rect 6741 6842 6828 7078
rect 7064 6842 7150 7078
rect 7386 6842 7472 7078
rect 7708 6842 7794 7078
rect 8030 6842 8116 7078
rect 8352 6842 8438 7078
rect 8674 6842 8760 7078
rect 8996 6842 9082 7078
rect 9318 6842 9404 7078
rect 9640 6842 9726 7078
rect 9962 6842 10048 7078
rect 10284 6842 10370 7078
rect 10606 6842 10692 7078
rect 10928 6842 11014 7078
rect 11250 6842 11336 7078
rect 11572 6842 11658 7078
rect 11894 6842 11980 7078
rect 12216 6842 12302 7078
rect 12538 6842 12624 7078
rect 12860 6842 12946 7078
rect 13182 6842 13268 7078
rect 13504 6842 13590 7078
rect 13826 6842 13912 7078
rect 14148 6842 14234 7078
rect 14470 6842 14556 7078
rect 14792 6842 14878 7078
rect 15114 6842 15200 7078
rect 15436 6842 15522 7078
rect 15758 6842 15844 7078
rect 16080 6842 16166 7078
rect 16402 6842 16488 7078
rect 16724 6842 16810 7078
rect 17046 6842 17132 7078
rect 17368 6842 17454 7078
rect 17690 6842 17776 7078
rect 18012 6842 18098 7078
rect 18334 6842 18420 7078
rect 18656 6842 18742 7078
rect 18978 6842 19064 7078
rect 19300 6842 19386 7078
rect 19622 6842 19708 7078
rect 19944 6842 20030 7078
rect 20266 6842 20352 7078
rect 20588 6842 20674 7078
rect 20910 6842 20996 7078
rect 21232 6842 21318 7078
rect 21554 6842 21640 7078
rect 21876 6842 21962 7078
rect 22198 6842 22284 7078
rect 22520 6842 22606 7078
rect 22842 6842 22928 7078
rect 23164 6842 23250 7078
rect 23486 6842 23572 7078
rect 23808 6842 23894 7078
rect 24130 6842 24216 7078
rect 24452 6842 24640 7078
rect -3360 6818 24640 6842
rect -3360 6474 24640 6498
rect -3360 6238 -3185 6474
rect -2949 6238 -2862 6474
rect -2626 6238 -2539 6474
rect -2303 6238 -2216 6474
rect -1980 6238 -1893 6474
rect -1657 6238 -1570 6474
rect -1334 6238 -1247 6474
rect -1011 6238 -924 6474
rect -688 6238 -601 6474
rect -365 6238 -278 6474
rect -42 6238 45 6474
rect 281 6238 368 6474
rect 604 6238 691 6474
rect 927 6238 1014 6474
rect 1250 6238 1337 6474
rect 1573 6238 1660 6474
rect 1896 6238 1983 6474
rect 2219 6238 2306 6474
rect 2542 6238 2629 6474
rect 2865 6238 2952 6474
rect 3188 6238 3275 6474
rect 3511 6238 3598 6474
rect 3834 6238 3921 6474
rect 4157 6238 4244 6474
rect 4480 6238 4567 6474
rect 4803 6238 4890 6474
rect 5126 6238 5213 6474
rect 5449 6238 5536 6474
rect 5772 6238 5859 6474
rect 6095 6238 6182 6474
rect 6418 6238 6505 6474
rect 6741 6238 6828 6474
rect 7064 6238 7150 6474
rect 7386 6238 7472 6474
rect 7708 6238 7794 6474
rect 8030 6238 8116 6474
rect 8352 6238 8438 6474
rect 8674 6238 8760 6474
rect 8996 6238 9082 6474
rect 9318 6238 9404 6474
rect 9640 6238 9726 6474
rect 9962 6238 10048 6474
rect 10284 6238 10370 6474
rect 10606 6238 10692 6474
rect 10928 6238 11014 6474
rect 11250 6238 11336 6474
rect 11572 6238 11658 6474
rect 11894 6238 11980 6474
rect 12216 6238 12302 6474
rect 12538 6238 12624 6474
rect 12860 6238 12946 6474
rect 13182 6238 13268 6474
rect 13504 6238 13590 6474
rect 13826 6238 13912 6474
rect 14148 6238 14234 6474
rect 14470 6238 14556 6474
rect 14792 6238 14878 6474
rect 15114 6238 15200 6474
rect 15436 6238 15522 6474
rect 15758 6238 15844 6474
rect 16080 6238 16166 6474
rect 16402 6238 16488 6474
rect 16724 6238 16810 6474
rect 17046 6238 17132 6474
rect 17368 6238 17454 6474
rect 17690 6238 17776 6474
rect 18012 6238 18098 6474
rect 18334 6238 18420 6474
rect 18656 6238 18742 6474
rect 18978 6238 19064 6474
rect 19300 6238 19386 6474
rect 19622 6238 19708 6474
rect 19944 6238 20030 6474
rect 20266 6238 20352 6474
rect 20588 6238 20674 6474
rect 20910 6238 20996 6474
rect 21232 6238 21318 6474
rect 21554 6238 21640 6474
rect 21876 6238 21962 6474
rect 22198 6238 22284 6474
rect 22520 6238 22606 6474
rect 22842 6238 22928 6474
rect 23164 6238 23250 6474
rect 23486 6238 23572 6474
rect 23808 6238 23894 6474
rect 24130 6238 24216 6474
rect 24452 6238 24640 6474
rect -3360 6108 24640 6238
rect -3360 5872 -3185 6108
rect -2949 5872 -2862 6108
rect -2626 5872 -2539 6108
rect -2303 5872 -2216 6108
rect -1980 5872 -1893 6108
rect -1657 5872 -1570 6108
rect -1334 5872 -1247 6108
rect -1011 5872 -924 6108
rect -688 5872 -601 6108
rect -365 5872 -278 6108
rect -42 5872 45 6108
rect 281 5872 368 6108
rect 604 5872 691 6108
rect 927 5872 1014 6108
rect 1250 5872 1337 6108
rect 1573 5872 1660 6108
rect 1896 5872 1983 6108
rect 2219 5872 2306 6108
rect 2542 5872 2629 6108
rect 2865 5872 2952 6108
rect 3188 5872 3275 6108
rect 3511 5872 3598 6108
rect 3834 5872 3921 6108
rect 4157 5872 4244 6108
rect 4480 5872 4567 6108
rect 4803 5872 4890 6108
rect 5126 5872 5213 6108
rect 5449 5872 5536 6108
rect 5772 5872 5859 6108
rect 6095 5872 6182 6108
rect 6418 5872 6505 6108
rect 6741 5872 6828 6108
rect 7064 5872 7150 6108
rect 7386 5872 7472 6108
rect 7708 5872 7794 6108
rect 8030 5872 8116 6108
rect 8352 5872 8438 6108
rect 8674 5872 8760 6108
rect 8996 5872 9082 6108
rect 9318 5872 9404 6108
rect 9640 5872 9726 6108
rect 9962 5872 10048 6108
rect 10284 5872 10370 6108
rect 10606 5872 10692 6108
rect 10928 5872 11014 6108
rect 11250 5872 11336 6108
rect 11572 5872 11658 6108
rect 11894 5872 11980 6108
rect 12216 5872 12302 6108
rect 12538 5872 12624 6108
rect 12860 5872 12946 6108
rect 13182 5872 13268 6108
rect 13504 5872 13590 6108
rect 13826 5872 13912 6108
rect 14148 5872 14234 6108
rect 14470 5872 14556 6108
rect 14792 5872 14878 6108
rect 15114 5872 15200 6108
rect 15436 5872 15522 6108
rect 15758 5872 15844 6108
rect 16080 5872 16166 6108
rect 16402 5872 16488 6108
rect 16724 5872 16810 6108
rect 17046 5872 17132 6108
rect 17368 5872 17454 6108
rect 17690 5872 17776 6108
rect 18012 5872 18098 6108
rect 18334 5872 18420 6108
rect 18656 5872 18742 6108
rect 18978 5872 19064 6108
rect 19300 5872 19386 6108
rect 19622 5872 19708 6108
rect 19944 5872 20030 6108
rect 20266 5872 20352 6108
rect 20588 5872 20674 6108
rect 20910 5872 20996 6108
rect 21232 5872 21318 6108
rect 21554 5872 21640 6108
rect 21876 5872 21962 6108
rect 22198 5872 22284 6108
rect 22520 5872 22606 6108
rect 22842 5872 22928 6108
rect 23164 5872 23250 6108
rect 23486 5872 23572 6108
rect 23808 5872 23894 6108
rect 24130 5872 24216 6108
rect 24452 5872 24640 6108
rect -3360 5848 24640 5872
rect -3360 5504 24640 5528
rect -3360 5268 -3185 5504
rect -2949 5268 -2862 5504
rect -2626 5268 -2539 5504
rect -2303 5268 -2216 5504
rect -1980 5268 -1893 5504
rect -1657 5268 -1570 5504
rect -1334 5268 -1247 5504
rect -1011 5268 -924 5504
rect -688 5268 -601 5504
rect -365 5268 -278 5504
rect -42 5268 45 5504
rect 281 5268 368 5504
rect 604 5268 691 5504
rect 927 5268 1014 5504
rect 1250 5268 1337 5504
rect 1573 5268 1660 5504
rect 1896 5268 1983 5504
rect 2219 5268 2306 5504
rect 2542 5268 2629 5504
rect 2865 5268 2952 5504
rect 3188 5268 3275 5504
rect 3511 5268 3598 5504
rect 3834 5268 3921 5504
rect 4157 5268 4244 5504
rect 4480 5268 4567 5504
rect 4803 5268 4890 5504
rect 5126 5268 5213 5504
rect 5449 5268 5536 5504
rect 5772 5268 5859 5504
rect 6095 5268 6182 5504
rect 6418 5268 6505 5504
rect 6741 5268 6828 5504
rect 7064 5268 7150 5504
rect 7386 5268 7472 5504
rect 7708 5268 7794 5504
rect 8030 5268 8116 5504
rect 8352 5268 8438 5504
rect 8674 5268 8760 5504
rect 8996 5268 9082 5504
rect 9318 5268 9404 5504
rect 9640 5268 9726 5504
rect 9962 5268 10048 5504
rect 10284 5268 10370 5504
rect 10606 5268 10692 5504
rect 10928 5268 11014 5504
rect 11250 5268 11336 5504
rect 11572 5268 11658 5504
rect 11894 5268 11980 5504
rect 12216 5268 12302 5504
rect 12538 5268 12624 5504
rect 12860 5268 12946 5504
rect 13182 5268 13268 5504
rect 13504 5268 13590 5504
rect 13826 5268 13912 5504
rect 14148 5268 14234 5504
rect 14470 5268 14556 5504
rect 14792 5268 14878 5504
rect 15114 5268 15200 5504
rect 15436 5268 15522 5504
rect 15758 5268 15844 5504
rect 16080 5268 16166 5504
rect 16402 5268 16488 5504
rect 16724 5268 16810 5504
rect 17046 5268 17132 5504
rect 17368 5268 17454 5504
rect 17690 5268 17776 5504
rect 18012 5268 18098 5504
rect 18334 5268 18420 5504
rect 18656 5268 18742 5504
rect 18978 5268 19064 5504
rect 19300 5268 19386 5504
rect 19622 5268 19708 5504
rect 19944 5268 20030 5504
rect 20266 5268 20352 5504
rect 20588 5268 20674 5504
rect 20910 5268 20996 5504
rect 21232 5268 21318 5504
rect 21554 5268 21640 5504
rect 21876 5268 21962 5504
rect 22198 5268 22284 5504
rect 22520 5268 22606 5504
rect 22842 5268 22928 5504
rect 23164 5268 23250 5504
rect 23486 5268 23572 5504
rect 23808 5268 23894 5504
rect 24130 5268 24216 5504
rect 24452 5268 24640 5504
rect -3360 4898 24640 5268
rect -3360 4662 -3185 4898
rect -2949 4662 -2862 4898
rect -2626 4662 -2539 4898
rect -2303 4662 -2216 4898
rect -1980 4662 -1893 4898
rect -1657 4662 -1570 4898
rect -1334 4662 -1247 4898
rect -1011 4662 -924 4898
rect -688 4662 -601 4898
rect -365 4662 -278 4898
rect -42 4662 45 4898
rect 281 4662 368 4898
rect 604 4662 691 4898
rect 927 4662 1014 4898
rect 1250 4662 1337 4898
rect 1573 4662 1660 4898
rect 1896 4662 1983 4898
rect 2219 4662 2306 4898
rect 2542 4662 2629 4898
rect 2865 4662 2952 4898
rect 3188 4662 3275 4898
rect 3511 4662 3598 4898
rect 3834 4662 3921 4898
rect 4157 4662 4244 4898
rect 4480 4662 4567 4898
rect 4803 4662 4890 4898
rect 5126 4662 5213 4898
rect 5449 4662 5536 4898
rect 5772 4662 5859 4898
rect 6095 4662 6182 4898
rect 6418 4662 6505 4898
rect 6741 4662 6828 4898
rect 7064 4662 7150 4898
rect 7386 4662 7472 4898
rect 7708 4662 7794 4898
rect 8030 4662 8116 4898
rect 8352 4662 8438 4898
rect 8674 4662 8760 4898
rect 8996 4662 9082 4898
rect 9318 4662 9404 4898
rect 9640 4662 9726 4898
rect 9962 4662 10048 4898
rect 10284 4662 10370 4898
rect 10606 4662 10692 4898
rect 10928 4662 11014 4898
rect 11250 4662 11336 4898
rect 11572 4662 11658 4898
rect 11894 4662 11980 4898
rect 12216 4662 12302 4898
rect 12538 4662 12624 4898
rect 12860 4662 12946 4898
rect 13182 4662 13268 4898
rect 13504 4662 13590 4898
rect 13826 4662 13912 4898
rect 14148 4662 14234 4898
rect 14470 4662 14556 4898
rect 14792 4662 14878 4898
rect 15114 4662 15200 4898
rect 15436 4662 15522 4898
rect 15758 4662 15844 4898
rect 16080 4662 16166 4898
rect 16402 4662 16488 4898
rect 16724 4662 16810 4898
rect 17046 4662 17132 4898
rect 17368 4662 17454 4898
rect 17690 4662 17776 4898
rect 18012 4662 18098 4898
rect 18334 4662 18420 4898
rect 18656 4662 18742 4898
rect 18978 4662 19064 4898
rect 19300 4662 19386 4898
rect 19622 4662 19708 4898
rect 19944 4662 20030 4898
rect 20266 4662 20352 4898
rect 20588 4662 20674 4898
rect 20910 4662 20996 4898
rect 21232 4662 21318 4898
rect 21554 4662 21640 4898
rect 21876 4662 21962 4898
rect 22198 4662 22284 4898
rect 22520 4662 22606 4898
rect 22842 4662 22928 4898
rect 23164 4662 23250 4898
rect 23486 4662 23572 4898
rect 23808 4662 23894 4898
rect 24130 4662 24216 4898
rect 24452 4662 24640 4898
rect -3360 4638 24640 4662
rect -3360 4294 24640 4318
rect -3360 4058 -3185 4294
rect -2949 4058 -2862 4294
rect -2626 4058 -2539 4294
rect -2303 4058 -2216 4294
rect -1980 4058 -1893 4294
rect -1657 4058 -1570 4294
rect -1334 4058 -1247 4294
rect -1011 4058 -924 4294
rect -688 4058 -601 4294
rect -365 4058 -278 4294
rect -42 4058 45 4294
rect 281 4058 368 4294
rect 604 4058 691 4294
rect 927 4058 1014 4294
rect 1250 4058 1337 4294
rect 1573 4058 1660 4294
rect 1896 4058 1983 4294
rect 2219 4058 2306 4294
rect 2542 4058 2629 4294
rect 2865 4058 2952 4294
rect 3188 4058 3275 4294
rect 3511 4058 3598 4294
rect 3834 4058 3921 4294
rect 4157 4058 4244 4294
rect 4480 4058 4567 4294
rect 4803 4058 4890 4294
rect 5126 4058 5213 4294
rect 5449 4058 5536 4294
rect 5772 4058 5859 4294
rect 6095 4058 6182 4294
rect 6418 4058 6505 4294
rect 6741 4058 6828 4294
rect 7064 4058 7150 4294
rect 7386 4058 7472 4294
rect 7708 4058 7794 4294
rect 8030 4058 8116 4294
rect 8352 4058 8438 4294
rect 8674 4058 8760 4294
rect 8996 4058 9082 4294
rect 9318 4058 9404 4294
rect 9640 4058 9726 4294
rect 9962 4058 10048 4294
rect 10284 4058 10370 4294
rect 10606 4058 10692 4294
rect 10928 4058 11014 4294
rect 11250 4058 11336 4294
rect 11572 4058 11658 4294
rect 11894 4058 11980 4294
rect 12216 4058 12302 4294
rect 12538 4058 12624 4294
rect 12860 4058 12946 4294
rect 13182 4058 13268 4294
rect 13504 4058 13590 4294
rect 13826 4058 13912 4294
rect 14148 4058 14234 4294
rect 14470 4058 14556 4294
rect 14792 4058 14878 4294
rect 15114 4058 15200 4294
rect 15436 4058 15522 4294
rect 15758 4058 15844 4294
rect 16080 4058 16166 4294
rect 16402 4058 16488 4294
rect 16724 4058 16810 4294
rect 17046 4058 17132 4294
rect 17368 4058 17454 4294
rect 17690 4058 17776 4294
rect 18012 4058 18098 4294
rect 18334 4058 18420 4294
rect 18656 4058 18742 4294
rect 18978 4058 19064 4294
rect 19300 4058 19386 4294
rect 19622 4058 19708 4294
rect 19944 4058 20030 4294
rect 20266 4058 20352 4294
rect 20588 4058 20674 4294
rect 20910 4058 20996 4294
rect 21232 4058 21318 4294
rect 21554 4058 21640 4294
rect 21876 4058 21962 4294
rect 22198 4058 22284 4294
rect 22520 4058 22606 4294
rect 22842 4058 22928 4294
rect 23164 4058 23250 4294
rect 23486 4058 23572 4294
rect 23808 4058 23894 4294
rect 24130 4058 24216 4294
rect 24452 4058 24640 4294
rect -3360 3688 24640 4058
rect -3360 3452 -3185 3688
rect -2949 3452 -2862 3688
rect -2626 3452 -2539 3688
rect -2303 3452 -2216 3688
rect -1980 3452 -1893 3688
rect -1657 3452 -1570 3688
rect -1334 3452 -1247 3688
rect -1011 3452 -924 3688
rect -688 3452 -601 3688
rect -365 3452 -278 3688
rect -42 3452 45 3688
rect 281 3452 368 3688
rect 604 3452 691 3688
rect 927 3452 1014 3688
rect 1250 3452 1337 3688
rect 1573 3452 1660 3688
rect 1896 3452 1983 3688
rect 2219 3452 2306 3688
rect 2542 3452 2629 3688
rect 2865 3452 2952 3688
rect 3188 3452 3275 3688
rect 3511 3452 3598 3688
rect 3834 3452 3921 3688
rect 4157 3452 4244 3688
rect 4480 3452 4567 3688
rect 4803 3452 4890 3688
rect 5126 3452 5213 3688
rect 5449 3452 5536 3688
rect 5772 3452 5859 3688
rect 6095 3452 6182 3688
rect 6418 3452 6505 3688
rect 6741 3452 6828 3688
rect 7064 3452 7150 3688
rect 7386 3452 7472 3688
rect 7708 3452 7794 3688
rect 8030 3452 8116 3688
rect 8352 3452 8438 3688
rect 8674 3452 8760 3688
rect 8996 3452 9082 3688
rect 9318 3452 9404 3688
rect 9640 3452 9726 3688
rect 9962 3452 10048 3688
rect 10284 3452 10370 3688
rect 10606 3452 10692 3688
rect 10928 3452 11014 3688
rect 11250 3452 11336 3688
rect 11572 3452 11658 3688
rect 11894 3452 11980 3688
rect 12216 3452 12302 3688
rect 12538 3452 12624 3688
rect 12860 3452 12946 3688
rect 13182 3452 13268 3688
rect 13504 3452 13590 3688
rect 13826 3452 13912 3688
rect 14148 3452 14234 3688
rect 14470 3452 14556 3688
rect 14792 3452 14878 3688
rect 15114 3452 15200 3688
rect 15436 3452 15522 3688
rect 15758 3452 15844 3688
rect 16080 3452 16166 3688
rect 16402 3452 16488 3688
rect 16724 3452 16810 3688
rect 17046 3452 17132 3688
rect 17368 3452 17454 3688
rect 17690 3452 17776 3688
rect 18012 3452 18098 3688
rect 18334 3452 18420 3688
rect 18656 3452 18742 3688
rect 18978 3452 19064 3688
rect 19300 3452 19386 3688
rect 19622 3452 19708 3688
rect 19944 3452 20030 3688
rect 20266 3452 20352 3688
rect 20588 3452 20674 3688
rect 20910 3452 20996 3688
rect 21232 3452 21318 3688
rect 21554 3452 21640 3688
rect 21876 3452 21962 3688
rect 22198 3452 22284 3688
rect 22520 3452 22606 3688
rect 22842 3452 22928 3688
rect 23164 3452 23250 3688
rect 23486 3452 23572 3688
rect 23808 3452 23894 3688
rect 24130 3452 24216 3688
rect 24452 3452 24640 3688
rect -3360 3428 24640 3452
rect -3360 3084 24640 3108
rect -3360 2848 -3185 3084
rect -2949 2848 -2862 3084
rect -2626 2848 -2539 3084
rect -2303 2848 -2216 3084
rect -1980 2848 -1893 3084
rect -1657 2848 -1570 3084
rect -1334 2848 -1247 3084
rect -1011 2848 -924 3084
rect -688 2848 -601 3084
rect -365 2848 -278 3084
rect -42 2848 45 3084
rect 281 2848 368 3084
rect 604 2848 691 3084
rect 927 2848 1014 3084
rect 1250 2848 1337 3084
rect 1573 2848 1660 3084
rect 1896 2848 1983 3084
rect 2219 2848 2306 3084
rect 2542 2848 2629 3084
rect 2865 2848 2952 3084
rect 3188 2848 3275 3084
rect 3511 2848 3598 3084
rect 3834 2848 3921 3084
rect 4157 2848 4244 3084
rect 4480 2848 4567 3084
rect 4803 2848 4890 3084
rect 5126 2848 5213 3084
rect 5449 2848 5536 3084
rect 5772 2848 5859 3084
rect 6095 2848 6182 3084
rect 6418 2848 6505 3084
rect 6741 2848 6828 3084
rect 7064 2848 7150 3084
rect 7386 2848 7472 3084
rect 7708 2848 7794 3084
rect 8030 2848 8116 3084
rect 8352 2848 8438 3084
rect 8674 2848 8760 3084
rect 8996 2848 9082 3084
rect 9318 2848 9404 3084
rect 9640 2848 9726 3084
rect 9962 2848 10048 3084
rect 10284 2848 10370 3084
rect 10606 2848 10692 3084
rect 10928 2848 11014 3084
rect 11250 2848 11336 3084
rect 11572 2848 11658 3084
rect 11894 2848 11980 3084
rect 12216 2848 12302 3084
rect 12538 2848 12624 3084
rect 12860 2848 12946 3084
rect 13182 2848 13268 3084
rect 13504 2848 13590 3084
rect 13826 2848 13912 3084
rect 14148 2848 14234 3084
rect 14470 2848 14556 3084
rect 14792 2848 14878 3084
rect 15114 2848 15200 3084
rect 15436 2848 15522 3084
rect 15758 2848 15844 3084
rect 16080 2848 16166 3084
rect 16402 2848 16488 3084
rect 16724 2848 16810 3084
rect 17046 2848 17132 3084
rect 17368 2848 17454 3084
rect 17690 2848 17776 3084
rect 18012 2848 18098 3084
rect 18334 2848 18420 3084
rect 18656 2848 18742 3084
rect 18978 2848 19064 3084
rect 19300 2848 19386 3084
rect 19622 2848 19708 3084
rect 19944 2848 20030 3084
rect 20266 2848 20352 3084
rect 20588 2848 20674 3084
rect 20910 2848 20996 3084
rect 21232 2848 21318 3084
rect 21554 2848 21640 3084
rect 21876 2848 21962 3084
rect 22198 2848 22284 3084
rect 22520 2848 22606 3084
rect 22842 2848 22928 3084
rect 23164 2848 23250 3084
rect 23486 2848 23572 3084
rect 23808 2848 23894 3084
rect 24130 2848 24216 3084
rect 24452 2848 24640 3084
rect -3360 2718 24640 2848
rect -3360 2482 -3185 2718
rect -2949 2482 -2862 2718
rect -2626 2482 -2539 2718
rect -2303 2482 -2216 2718
rect -1980 2482 -1893 2718
rect -1657 2482 -1570 2718
rect -1334 2482 -1247 2718
rect -1011 2482 -924 2718
rect -688 2482 -601 2718
rect -365 2482 -278 2718
rect -42 2482 45 2718
rect 281 2482 368 2718
rect 604 2482 691 2718
rect 927 2482 1014 2718
rect 1250 2482 1337 2718
rect 1573 2482 1660 2718
rect 1896 2482 1983 2718
rect 2219 2482 2306 2718
rect 2542 2482 2629 2718
rect 2865 2482 2952 2718
rect 3188 2482 3275 2718
rect 3511 2482 3598 2718
rect 3834 2482 3921 2718
rect 4157 2482 4244 2718
rect 4480 2482 4567 2718
rect 4803 2482 4890 2718
rect 5126 2482 5213 2718
rect 5449 2482 5536 2718
rect 5772 2482 5859 2718
rect 6095 2482 6182 2718
rect 6418 2482 6505 2718
rect 6741 2482 6828 2718
rect 7064 2482 7150 2718
rect 7386 2482 7472 2718
rect 7708 2482 7794 2718
rect 8030 2482 8116 2718
rect 8352 2482 8438 2718
rect 8674 2482 8760 2718
rect 8996 2482 9082 2718
rect 9318 2482 9404 2718
rect 9640 2482 9726 2718
rect 9962 2482 10048 2718
rect 10284 2482 10370 2718
rect 10606 2482 10692 2718
rect 10928 2482 11014 2718
rect 11250 2482 11336 2718
rect 11572 2482 11658 2718
rect 11894 2482 11980 2718
rect 12216 2482 12302 2718
rect 12538 2482 12624 2718
rect 12860 2482 12946 2718
rect 13182 2482 13268 2718
rect 13504 2482 13590 2718
rect 13826 2482 13912 2718
rect 14148 2482 14234 2718
rect 14470 2482 14556 2718
rect 14792 2482 14878 2718
rect 15114 2482 15200 2718
rect 15436 2482 15522 2718
rect 15758 2482 15844 2718
rect 16080 2482 16166 2718
rect 16402 2482 16488 2718
rect 16724 2482 16810 2718
rect 17046 2482 17132 2718
rect 17368 2482 17454 2718
rect 17690 2482 17776 2718
rect 18012 2482 18098 2718
rect 18334 2482 18420 2718
rect 18656 2482 18742 2718
rect 18978 2482 19064 2718
rect 19300 2482 19386 2718
rect 19622 2482 19708 2718
rect 19944 2482 20030 2718
rect 20266 2482 20352 2718
rect 20588 2482 20674 2718
rect 20910 2482 20996 2718
rect 21232 2482 21318 2718
rect 21554 2482 21640 2718
rect 21876 2482 21962 2718
rect 22198 2482 22284 2718
rect 22520 2482 22606 2718
rect 22842 2482 22928 2718
rect 23164 2482 23250 2718
rect 23486 2482 23572 2718
rect 23808 2482 23894 2718
rect 24130 2482 24216 2718
rect 24452 2482 24640 2718
rect -3360 2458 24640 2482
rect -3360 2114 24640 2138
rect -3360 1878 -3185 2114
rect -2949 1878 -2862 2114
rect -2626 1878 -2539 2114
rect -2303 1878 -2216 2114
rect -1980 1878 -1893 2114
rect -1657 1878 -1570 2114
rect -1334 1878 -1247 2114
rect -1011 1878 -924 2114
rect -688 1878 -601 2114
rect -365 1878 -278 2114
rect -42 1878 45 2114
rect 281 1878 368 2114
rect 604 1878 691 2114
rect 927 1878 1014 2114
rect 1250 1878 1337 2114
rect 1573 1878 1660 2114
rect 1896 1878 1983 2114
rect 2219 1878 2306 2114
rect 2542 1878 2629 2114
rect 2865 1878 2952 2114
rect 3188 1878 3275 2114
rect 3511 1878 3598 2114
rect 3834 1878 3921 2114
rect 4157 1878 4244 2114
rect 4480 1878 4567 2114
rect 4803 1878 4890 2114
rect 5126 1878 5213 2114
rect 5449 1878 5536 2114
rect 5772 1878 5859 2114
rect 6095 1878 6182 2114
rect 6418 1878 6505 2114
rect 6741 1878 6828 2114
rect 7064 1878 7150 2114
rect 7386 1878 7472 2114
rect 7708 1878 7794 2114
rect 8030 1878 8116 2114
rect 8352 1878 8438 2114
rect 8674 1878 8760 2114
rect 8996 1878 9082 2114
rect 9318 1878 9404 2114
rect 9640 1878 9726 2114
rect 9962 1878 10048 2114
rect 10284 1878 10370 2114
rect 10606 1878 10692 2114
rect 10928 1878 11014 2114
rect 11250 1878 11336 2114
rect 11572 1878 11658 2114
rect 11894 1878 11980 2114
rect 12216 1878 12302 2114
rect 12538 1878 12624 2114
rect 12860 1878 12946 2114
rect 13182 1878 13268 2114
rect 13504 1878 13590 2114
rect 13826 1878 13912 2114
rect 14148 1878 14234 2114
rect 14470 1878 14556 2114
rect 14792 1878 14878 2114
rect 15114 1878 15200 2114
rect 15436 1878 15522 2114
rect 15758 1878 15844 2114
rect 16080 1878 16166 2114
rect 16402 1878 16488 2114
rect 16724 1878 16810 2114
rect 17046 1878 17132 2114
rect 17368 1878 17454 2114
rect 17690 1878 17776 2114
rect 18012 1878 18098 2114
rect 18334 1878 18420 2114
rect 18656 1878 18742 2114
rect 18978 1878 19064 2114
rect 19300 1878 19386 2114
rect 19622 1878 19708 2114
rect 19944 1878 20030 2114
rect 20266 1878 20352 2114
rect 20588 1878 20674 2114
rect 20910 1878 20996 2114
rect 21232 1878 21318 2114
rect 21554 1878 21640 2114
rect 21876 1878 21962 2114
rect 22198 1878 22284 2114
rect 22520 1878 22606 2114
rect 22842 1878 22928 2114
rect 23164 1878 23250 2114
rect 23486 1878 23572 2114
rect 23808 1878 23894 2114
rect 24130 1878 24216 2114
rect 24452 1878 24640 2114
rect -3360 1508 24640 1878
rect -3360 1272 -3185 1508
rect -2949 1272 -2862 1508
rect -2626 1272 -2539 1508
rect -2303 1272 -2216 1508
rect -1980 1272 -1893 1508
rect -1657 1272 -1570 1508
rect -1334 1272 -1247 1508
rect -1011 1272 -924 1508
rect -688 1272 -601 1508
rect -365 1272 -278 1508
rect -42 1272 45 1508
rect 281 1272 368 1508
rect 604 1272 691 1508
rect 927 1272 1014 1508
rect 1250 1272 1337 1508
rect 1573 1272 1660 1508
rect 1896 1272 1983 1508
rect 2219 1272 2306 1508
rect 2542 1272 2629 1508
rect 2865 1272 2952 1508
rect 3188 1272 3275 1508
rect 3511 1272 3598 1508
rect 3834 1272 3921 1508
rect 4157 1272 4244 1508
rect 4480 1272 4567 1508
rect 4803 1272 4890 1508
rect 5126 1272 5213 1508
rect 5449 1272 5536 1508
rect 5772 1272 5859 1508
rect 6095 1272 6182 1508
rect 6418 1272 6505 1508
rect 6741 1272 6828 1508
rect 7064 1272 7150 1508
rect 7386 1272 7472 1508
rect 7708 1272 7794 1508
rect 8030 1272 8116 1508
rect 8352 1272 8438 1508
rect 8674 1272 8760 1508
rect 8996 1272 9082 1508
rect 9318 1272 9404 1508
rect 9640 1272 9726 1508
rect 9962 1272 10048 1508
rect 10284 1272 10370 1508
rect 10606 1272 10692 1508
rect 10928 1272 11014 1508
rect 11250 1272 11336 1508
rect 11572 1272 11658 1508
rect 11894 1272 11980 1508
rect 12216 1272 12302 1508
rect 12538 1272 12624 1508
rect 12860 1272 12946 1508
rect 13182 1272 13268 1508
rect 13504 1272 13590 1508
rect 13826 1272 13912 1508
rect 14148 1272 14234 1508
rect 14470 1272 14556 1508
rect 14792 1272 14878 1508
rect 15114 1272 15200 1508
rect 15436 1272 15522 1508
rect 15758 1272 15844 1508
rect 16080 1272 16166 1508
rect 16402 1272 16488 1508
rect 16724 1272 16810 1508
rect 17046 1272 17132 1508
rect 17368 1272 17454 1508
rect 17690 1272 17776 1508
rect 18012 1272 18098 1508
rect 18334 1272 18420 1508
rect 18656 1272 18742 1508
rect 18978 1272 19064 1508
rect 19300 1272 19386 1508
rect 19622 1272 19708 1508
rect 19944 1272 20030 1508
rect 20266 1272 20352 1508
rect 20588 1272 20674 1508
rect 20910 1272 20996 1508
rect 21232 1272 21318 1508
rect 21554 1272 21640 1508
rect 21876 1272 21962 1508
rect 22198 1272 22284 1508
rect 22520 1272 22606 1508
rect 22842 1272 22928 1508
rect 23164 1272 23250 1508
rect 23486 1272 23572 1508
rect 23808 1272 23894 1508
rect 24130 1272 24216 1508
rect 24452 1272 24640 1508
rect -3360 1248 24640 1272
rect -3360 903 24640 928
rect -3360 667 -3185 903
rect -2949 667 -2862 903
rect -2626 667 -2539 903
rect -2303 667 -2216 903
rect -1980 667 -1893 903
rect -1657 667 -1570 903
rect -1334 667 -1247 903
rect -1011 667 -924 903
rect -688 667 -601 903
rect -365 667 -278 903
rect -42 667 45 903
rect 281 667 368 903
rect 604 667 691 903
rect 927 667 1014 903
rect 1250 667 1337 903
rect 1573 667 1660 903
rect 1896 667 1983 903
rect 2219 667 2306 903
rect 2542 667 2629 903
rect 2865 667 2952 903
rect 3188 667 3275 903
rect 3511 667 3598 903
rect 3834 667 3921 903
rect 4157 667 4244 903
rect 4480 667 4567 903
rect 4803 667 4890 903
rect 5126 667 5213 903
rect 5449 667 5536 903
rect 5772 667 5859 903
rect 6095 667 6182 903
rect 6418 667 6505 903
rect 6741 667 6828 903
rect 7064 667 7150 903
rect 7386 667 7472 903
rect 7708 667 7794 903
rect 8030 667 8116 903
rect 8352 667 8438 903
rect 8674 667 8760 903
rect 8996 667 9082 903
rect 9318 667 9404 903
rect 9640 667 9726 903
rect 9962 667 10048 903
rect 10284 667 10370 903
rect 10606 667 10692 903
rect 10928 667 11014 903
rect 11250 667 11336 903
rect 11572 667 11658 903
rect 11894 667 11980 903
rect 12216 667 12302 903
rect 12538 667 12624 903
rect 12860 667 12946 903
rect 13182 667 13268 903
rect 13504 667 13590 903
rect 13826 667 13912 903
rect 14148 667 14234 903
rect 14470 667 14556 903
rect 14792 667 14878 903
rect 15114 667 15200 903
rect 15436 667 15522 903
rect 15758 667 15844 903
rect 16080 667 16166 903
rect 16402 667 16488 903
rect 16724 667 16810 903
rect 17046 667 17132 903
rect 17368 667 17454 903
rect 17690 667 17776 903
rect 18012 667 18098 903
rect 18334 667 18420 903
rect 18656 667 18742 903
rect 18978 667 19064 903
rect 19300 667 19386 903
rect 19622 667 19708 903
rect 19944 667 20030 903
rect 20266 667 20352 903
rect 20588 667 20674 903
rect 20910 667 20996 903
rect 21232 667 21318 903
rect 21554 667 21640 903
rect 21876 667 21962 903
rect 22198 667 22284 903
rect 22520 667 22606 903
rect 22842 667 22928 903
rect 23164 667 23250 903
rect 23486 667 23572 903
rect 23808 667 23894 903
rect 24130 667 24216 903
rect 24452 667 24640 903
rect -3360 521 24640 667
rect -3360 285 -3185 521
rect -2949 285 -2862 521
rect -2626 285 -2539 521
rect -2303 285 -2216 521
rect -1980 285 -1893 521
rect -1657 285 -1570 521
rect -1334 285 -1247 521
rect -1011 285 -924 521
rect -688 285 -601 521
rect -365 285 -278 521
rect -42 285 45 521
rect 281 285 368 521
rect 604 285 691 521
rect 927 285 1014 521
rect 1250 285 1337 521
rect 1573 285 1660 521
rect 1896 285 1983 521
rect 2219 285 2306 521
rect 2542 285 2629 521
rect 2865 285 2952 521
rect 3188 285 3275 521
rect 3511 285 3598 521
rect 3834 285 3921 521
rect 4157 285 4244 521
rect 4480 285 4567 521
rect 4803 285 4890 521
rect 5126 285 5213 521
rect 5449 285 5536 521
rect 5772 285 5859 521
rect 6095 285 6182 521
rect 6418 285 6505 521
rect 6741 285 6828 521
rect 7064 285 7150 521
rect 7386 285 7472 521
rect 7708 285 7794 521
rect 8030 285 8116 521
rect 8352 285 8438 521
rect 8674 285 8760 521
rect 8996 285 9082 521
rect 9318 285 9404 521
rect 9640 285 9726 521
rect 9962 285 10048 521
rect 10284 285 10370 521
rect 10606 285 10692 521
rect 10928 285 11014 521
rect 11250 285 11336 521
rect 11572 285 11658 521
rect 11894 285 11980 521
rect 12216 285 12302 521
rect 12538 285 12624 521
rect 12860 285 12946 521
rect 13182 285 13268 521
rect 13504 285 13590 521
rect 13826 285 13912 521
rect 14148 285 14234 521
rect 14470 285 14556 521
rect 14792 285 14878 521
rect 15114 285 15200 521
rect 15436 285 15522 521
rect 15758 285 15844 521
rect 16080 285 16166 521
rect 16402 285 16488 521
rect 16724 285 16810 521
rect 17046 285 17132 521
rect 17368 285 17454 521
rect 17690 285 17776 521
rect 18012 285 18098 521
rect 18334 285 18420 521
rect 18656 285 18742 521
rect 18978 285 19064 521
rect 19300 285 19386 521
rect 19622 285 19708 521
rect 19944 285 20030 521
rect 20266 285 20352 521
rect 20588 285 20674 521
rect 20910 285 20996 521
rect 21232 285 21318 521
rect 21554 285 21640 521
rect 21876 285 21962 521
rect 22198 285 22284 521
rect 22520 285 22606 521
rect 22842 285 22928 521
rect 23164 285 23250 521
rect 23486 285 23572 521
rect 23808 285 23894 521
rect 24130 285 24216 521
rect 24452 285 24640 521
rect -3360 139 24640 285
rect -3360 -97 -3185 139
rect -2949 -97 -2862 139
rect -2626 -97 -2539 139
rect -2303 -97 -2216 139
rect -1980 -97 -1893 139
rect -1657 -97 -1570 139
rect -1334 -97 -1247 139
rect -1011 -97 -924 139
rect -688 -97 -601 139
rect -365 -97 -278 139
rect -42 -97 45 139
rect 281 -97 368 139
rect 604 -97 691 139
rect 927 -97 1014 139
rect 1250 -97 1337 139
rect 1573 -97 1660 139
rect 1896 -97 1983 139
rect 2219 -97 2306 139
rect 2542 -97 2629 139
rect 2865 -97 2952 139
rect 3188 -97 3275 139
rect 3511 -97 3598 139
rect 3834 -97 3921 139
rect 4157 -97 4244 139
rect 4480 -97 4567 139
rect 4803 -97 4890 139
rect 5126 -97 5213 139
rect 5449 -97 5536 139
rect 5772 -97 5859 139
rect 6095 -97 6182 139
rect 6418 -97 6505 139
rect 6741 -97 6828 139
rect 7064 -97 7150 139
rect 7386 -97 7472 139
rect 7708 -97 7794 139
rect 8030 -97 8116 139
rect 8352 -97 8438 139
rect 8674 -97 8760 139
rect 8996 -97 9082 139
rect 9318 -97 9404 139
rect 9640 -97 9726 139
rect 9962 -97 10048 139
rect 10284 -97 10370 139
rect 10606 -97 10692 139
rect 10928 -97 11014 139
rect 11250 -97 11336 139
rect 11572 -97 11658 139
rect 11894 -97 11980 139
rect 12216 -97 12302 139
rect 12538 -97 12624 139
rect 12860 -97 12946 139
rect 13182 -97 13268 139
rect 13504 -97 13590 139
rect 13826 -97 13912 139
rect 14148 -97 14234 139
rect 14470 -97 14556 139
rect 14792 -97 14878 139
rect 15114 -97 15200 139
rect 15436 -97 15522 139
rect 15758 -97 15844 139
rect 16080 -97 16166 139
rect 16402 -97 16488 139
rect 16724 -97 16810 139
rect 17046 -97 17132 139
rect 17368 -97 17454 139
rect 17690 -97 17776 139
rect 18012 -97 18098 139
rect 18334 -97 18420 139
rect 18656 -97 18742 139
rect 18978 -97 19064 139
rect 19300 -97 19386 139
rect 19622 -97 19708 139
rect 19944 -97 20030 139
rect 20266 -97 20352 139
rect 20588 -97 20674 139
rect 20910 -97 20996 139
rect 21232 -97 21318 139
rect 21554 -97 21640 139
rect 21876 -97 21962 139
rect 22198 -97 22284 139
rect 22520 -97 22606 139
rect 22842 -97 22928 139
rect 23164 -97 23250 139
rect 23486 -97 23572 139
rect 23808 -97 23894 139
rect 24130 -97 24216 139
rect 24452 -97 24640 139
rect -3360 -122 24640 -97
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_0
timestamp 1666199351
transform 1 0 23000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_1
timestamp 1666199351
transform 1 0 22000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_2
timestamp 1666199351
transform 1 0 21000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_3
timestamp 1666199351
transform 1 0 20000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_4
timestamp 1666199351
transform 1 0 19000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_5
timestamp 1666199351
transform 1 0 18000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_6
timestamp 1666199351
transform 1 0 17000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_7
timestamp 1666199351
transform 1 0 16000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_8
timestamp 1666199351
transform 1 0 15000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_9
timestamp 1666199351
transform 1 0 -1000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_10
timestamp 1666199351
transform 1 0 -2000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_11
timestamp 1666199351
transform 1 0 -3000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_12
timestamp 1666199351
transform 1 0 0 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_13
timestamp 1666199351
transform 1 0 1000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_14
timestamp 1666199351
transform 1 0 2000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_15
timestamp 1666199351
transform 1 0 3000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_16
timestamp 1666199351
transform 1 0 4000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_17
timestamp 1666199351
transform 1 0 5000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_18
timestamp 1666199351
transform 1 0 6000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_19
timestamp 1666199351
transform 1 0 7000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_20
timestamp 1666199351
transform 1 0 8000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_21
timestamp 1666199351
transform 1 0 9000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_22
timestamp 1666199351
transform 1 0 14000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_23
timestamp 1666199351
transform 1 0 13000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_24
timestamp 1666199351
transform 1 0 12000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_25
timestamp 1666199351
transform 1 0 11000 0 1 -6457
box 0 6315 1000 45908
use sky130_fd_io__com_bus_slice  sky130_fd_io__com_bus_slice_26
timestamp 1666199351
transform 1 0 10000 0 1 -6457
box 0 6315 1000 45908
<< labels >>
flabel metal5 s 24386 34608 24640 39451 3 FreeSans 520 180 0 0 VSSIO
port 1 nsew
flabel metal5 s 24386 8998 24640 10798 3 FreeSans 520 180 0 0 VSSA
port 2 nsew
flabel metal5 s 24447 2458 24640 3108 3 FreeSans 520 180 0 0 VDDA
port 3 nsew
flabel metal5 s 24386 7788 24640 8678 3 FreeSans 520 180 0 0 VSSD
port 4 nsew
flabel metal5 s 24386 11118 24640 11968 3 FreeSans 520 180 0 0 VSSIO_Q
port 5 nsew
flabel metal5 s 24386 4638 24640 5528 3 FreeSans 520 180 0 0 VSSIO
port 1 nsew
flabel metal5 s 24386 5848 24640 6498 3 FreeSans 520 180 0 0 VSWITCH
port 6 nsew
flabel metal5 s 24386 6819 24640 7468 3 FreeSans 520 180 0 0 VSSA
port 2 nsew
flabel metal5 s 24386 1248 24640 2138 3 FreeSans 520 180 0 0 VCCD
port 7 nsew
flabel metal5 s 24386 12288 24640 13138 3 FreeSans 520 180 0 0 VDDIO_Q
port 8 nsew
flabel metal5 s 24386 13458 24640 18448 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew
flabel metal5 s 24386 -122 24640 928 3 FreeSans 520 180 0 0 VCCHIB
port 10 nsew
flabel metal5 s 24386 3428 24640 4318 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew
flabel metal5 s -3360 34608 -3106 39451 3 FreeSans 520 0 0 0 VSSIO
port 1 nsew
flabel metal5 s -3360 13458 -3106 18448 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew
flabel metal5 s -3360 7788 -3106 8678 3 FreeSans 520 0 0 0 VSSD
port 4 nsew
flabel metal5 s -3360 11118 -3106 11968 3 FreeSans 520 0 0 0 VSSIO_Q
port 5 nsew
flabel metal5 s -3360 5848 -3106 6498 3 FreeSans 520 0 0 0 VSWITCH
port 6 nsew
flabel metal5 s -3360 4638 -3106 5528 3 FreeSans 520 0 0 0 VSSIO
port 1 nsew
flabel metal5 s -3360 2458 -3167 3108 3 FreeSans 520 0 0 0 VDDA
port 3 nsew
flabel metal5 s -3360 3428 -3106 4318 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew
flabel metal5 s -3360 1248 -3106 2138 3 FreeSans 520 0 0 0 VCCD
port 7 nsew
flabel metal5 s -3360 12288 -3106 13138 3 FreeSans 520 0 0 0 VDDIO_Q
port 8 nsew
flabel metal5 s -3360 8998 -3106 10798 3 FreeSans 520 0 0 0 VSSA
port 2 nsew
flabel metal5 s -3360 6819 -3106 7468 3 FreeSans 520 0 0 0 VSSA
port 2 nsew
flabel metal5 s -3360 -122 -3106 928 3 FreeSans 520 0 0 0 VCCHIB
port 10 nsew
flabel metal4 s 24386 7768 24640 8698 3 FreeSans 520 180 0 0 VSSD
port 4 nsew
flabel metal4 s 24447 2438 24640 3128 3 FreeSans 520 180 0 0 VDDA
port 3 nsew
flabel metal4 s 24386 11098 24640 11988 3 FreeSans 520 180 0 0 VSSIO_Q
port 5 nsew
flabel metal4 s 24386 4618 24640 5548 3 FreeSans 520 180 0 0 VSSIO
port 1 nsew
flabel metal4 s 24386 5828 24640 6518 3 FreeSans 520 180 0 0 VSWITCH
port 6 nsew
flabel metal4 s 24386 9780 24640 10016 3 FreeSans 520 180 0 0 VSSA
port 2 nsew
flabel metal4 s 24386 10732 24640 10798 3 FreeSans 520 180 0 0 VSSA
port 2 nsew
flabel metal4 s 24386 -142 24640 948 3 FreeSans 520 180 0 0 VCCHIB
port 10 nsew
flabel metal4 s 24386 3408 24640 4338 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew
flabel metal4 s 24386 8998 24640 9064 3 FreeSans 520 180 0 0 VSSA
port 2 nsew
flabel metal4 s 24386 6798 24640 7488 3 FreeSans 520 180 0 0 VSSA
port 2 nsew
flabel metal4 s 24386 12268 24640 13158 3 FreeSans 520 180 0 0 VDDIO_Q
port 8 nsew
flabel metal4 s 24386 1228 24640 2158 3 FreeSans 520 180 0 0 VCCD
port 7 nsew
flabel metal4 s 24386 9124 24640 9720 3 FreeSans 520 180 0 0 AMUXBUS_B
port 11 nsew
flabel metal4 s 24386 34608 24640 39451 3 FreeSans 520 180 0 0 VSSIO
port 1 nsew
flabel metal4 s 24386 10076 24640 10672 3 FreeSans 520 180 0 0 AMUXBUS_A
port 12 nsew
flabel metal4 s 24386 13458 24640 18451 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew
flabel metal4 s -3360 34608 -3106 39451 3 FreeSans 520 0 0 0 VSSIO
port 1 nsew
flabel metal4 s -3360 3408 -3106 4338 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew
flabel metal4 s -3360 12268 -3106 13158 3 FreeSans 520 0 0 0 VDDIO_Q
port 8 nsew
flabel metal4 s -3360 13458 -3106 18451 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew
flabel metal4 s -3360 1228 -3106 2158 3 FreeSans 520 0 0 0 VCCD
port 7 nsew
flabel metal4 s -3360 8998 -3106 9064 3 FreeSans 520 0 0 0 VSSA
port 2 nsew
flabel metal4 s -3360 5828 -3106 6518 3 FreeSans 520 0 0 0 VSWITCH
port 6 nsew
flabel metal4 s -3360 -142 -3106 948 3 FreeSans 520 0 0 0 VCCHIB
port 10 nsew
flabel metal4 s -3360 9780 -3106 10016 3 FreeSans 520 0 0 0 VSSA
port 2 nsew
flabel metal4 s -3360 11098 -3106 11988 3 FreeSans 520 0 0 0 VSSIO_Q
port 5 nsew
flabel metal4 s -3360 4618 -3106 5548 3 FreeSans 520 0 0 0 VSSIO
port 1 nsew
flabel metal4 s -3360 2438 -3167 3128 3 FreeSans 520 0 0 0 VDDA
port 3 nsew
flabel metal4 s -3360 10076 -3106 10672 3 FreeSans 520 0 0 0 AMUXBUS_A
port 12 nsew
flabel metal4 s -3360 10732 -3106 10798 3 FreeSans 520 0 0 0 VSSA
port 2 nsew
flabel metal4 s -3360 6798 -3106 7488 3 FreeSans 520 0 0 0 VSSA
port 2 nsew
flabel metal4 s -3360 7768 -3106 8698 3 FreeSans 520 0 0 0 VSSD
port 4 nsew
flabel metal4 s -3360 9124 -3106 9720 3 FreeSans 520 0 0 0 AMUXBUS_B
port 11 nsew
<< properties >>
string GDS_END 31659838
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31363550
<< end >>
