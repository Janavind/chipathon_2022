magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 145 457 157
rect 741 145 1011 203
rect 1 21 1011 145
rect 29 -17 63 21
<< locali >>
rect 18 197 66 325
rect 350 153 425 219
rect 938 334 995 491
rect 961 149 995 334
rect 938 83 995 149
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 35 393 69 493
rect 103 427 169 527
rect 203 417 237 493
rect 291 451 370 527
rect 462 451 637 485
rect 203 393 569 417
rect 35 359 156 393
rect 122 292 156 359
rect 196 383 569 393
rect 196 365 237 383
rect 122 226 162 292
rect 122 161 156 226
rect 35 127 156 161
rect 196 182 230 365
rect 264 305 467 339
rect 264 248 298 305
rect 410 271 467 305
rect 501 315 569 383
rect 196 148 237 182
rect 501 207 535 315
rect 603 265 637 451
rect 671 427 705 527
rect 767 373 825 487
rect 684 307 825 373
rect 859 314 893 527
rect 603 233 756 265
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 237 148
rect 459 141 535 207
rect 574 199 756 233
rect 574 107 608 199
rect 790 149 825 307
rect 291 17 357 93
rect 476 73 608 107
rect 653 17 719 106
rect 767 83 825 149
rect 859 17 893 143
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 350 153 425 219 6 D
port 1 nsew signal input
rlabel locali s 18 197 66 325 6 SLEEP_B
port 2 nsew clock input
rlabel metal1 s 0 -48 1012 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 1011 145 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 741 145 1011 203 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 145 457 157 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1050 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 938 83 995 149 6 Q
port 7 nsew signal output
rlabel locali s 961 149 995 334 6 Q
port 7 nsew signal output
rlabel locali s 938 334 995 491 6 Q
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1012 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2376910
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2367978
<< end >>
