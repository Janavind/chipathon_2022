magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< pwell >>
rect 15 163 615 545
<< nmos >>
rect 171 189 201 519
rect 257 189 287 519
rect 343 189 373 519
rect 429 189 459 519
<< ndiff >>
rect 111 507 171 519
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 507 257 519
rect 201 473 212 507
rect 246 473 257 507
rect 201 439 257 473
rect 201 405 212 439
rect 246 405 257 439
rect 201 371 257 405
rect 201 337 212 371
rect 246 337 257 371
rect 201 303 257 337
rect 201 269 212 303
rect 246 269 257 303
rect 201 235 257 269
rect 201 201 212 235
rect 246 201 257 235
rect 201 189 257 201
rect 287 507 343 519
rect 287 473 298 507
rect 332 473 343 507
rect 287 439 343 473
rect 287 405 298 439
rect 332 405 343 439
rect 287 371 343 405
rect 287 337 298 371
rect 332 337 343 371
rect 287 303 343 337
rect 287 269 298 303
rect 332 269 343 303
rect 287 235 343 269
rect 287 201 298 235
rect 332 201 343 235
rect 287 189 343 201
rect 373 507 429 519
rect 373 473 384 507
rect 418 473 429 507
rect 373 439 429 473
rect 373 405 384 439
rect 418 405 429 439
rect 373 371 429 405
rect 373 337 384 371
rect 418 337 429 371
rect 373 303 429 337
rect 373 269 384 303
rect 418 269 429 303
rect 373 235 429 269
rect 373 201 384 235
rect 418 201 429 235
rect 373 189 429 201
rect 459 507 519 519
rect 459 473 470 507
rect 504 473 519 507
rect 459 439 519 473
rect 459 405 470 439
rect 504 405 519 439
rect 459 371 519 405
rect 459 337 470 371
rect 504 337 519 371
rect 459 303 519 337
rect 459 269 470 303
rect 504 269 519 303
rect 459 235 519 269
rect 459 201 470 235
rect 504 201 519 235
rect 459 189 519 201
<< ndiffc >>
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 473 246 507
rect 212 405 246 439
rect 212 337 246 371
rect 212 269 246 303
rect 212 201 246 235
rect 298 473 332 507
rect 298 405 332 439
rect 298 337 332 371
rect 298 269 332 303
rect 298 201 332 235
rect 384 473 418 507
rect 384 405 418 439
rect 384 337 418 371
rect 384 269 418 303
rect 384 201 418 235
rect 470 473 504 507
rect 470 405 504 439
rect 470 337 504 371
rect 470 269 504 303
rect 470 201 504 235
<< psubdiff >>
rect 41 507 111 519
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 519 507 589 519
rect 519 473 538 507
rect 572 473 589 507
rect 519 439 589 473
rect 519 405 538 439
rect 572 405 589 439
rect 519 371 589 405
rect 519 337 538 371
rect 572 337 589 371
rect 519 303 589 337
rect 519 269 538 303
rect 572 269 589 303
rect 519 235 589 269
rect 519 201 538 235
rect 572 201 589 235
rect 519 189 589 201
<< psubdiffcont >>
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 538 473 572 507
rect 538 405 572 439
rect 538 337 572 371
rect 538 269 572 303
rect 538 201 572 235
<< poly >>
rect 243 687 387 708
rect 120 595 201 611
rect 120 561 136 595
rect 170 561 201 595
rect 243 585 264 687
rect 366 585 387 687
rect 243 569 387 585
rect 429 595 510 611
rect 120 545 201 561
rect 171 519 201 545
rect 257 519 287 569
rect 343 519 373 569
rect 429 561 460 595
rect 494 561 510 595
rect 429 545 510 561
rect 429 519 459 545
rect 171 163 201 189
rect 120 147 201 163
rect 120 113 136 147
rect 170 113 201 147
rect 257 139 287 189
rect 343 139 373 189
rect 429 163 459 189
rect 429 147 510 163
rect 120 97 201 113
rect 243 123 387 139
rect 243 21 264 123
rect 366 21 387 123
rect 429 113 460 147
rect 494 113 510 147
rect 429 97 510 113
rect 243 0 387 21
<< polycont >>
rect 136 561 170 595
rect 264 585 366 687
rect 460 561 494 595
rect 136 113 170 147
rect 264 21 366 123
rect 460 113 494 147
<< locali >>
rect 248 689 382 708
rect 120 595 186 611
rect 120 561 136 595
rect 170 561 186 595
rect 248 583 262 689
rect 368 583 382 689
rect 248 569 382 583
rect 444 595 510 611
rect 120 545 186 561
rect 444 561 460 595
rect 494 561 510 595
rect 444 545 510 561
rect 120 523 160 545
rect 470 523 510 545
rect 41 507 160 523
rect 41 473 58 507
rect 92 479 126 507
rect 94 473 126 479
rect 41 445 60 473
rect 94 445 160 473
rect 41 439 160 445
rect 41 405 58 439
rect 92 407 126 439
rect 94 405 126 407
rect 41 373 60 405
rect 94 373 160 405
rect 41 371 160 373
rect 41 337 58 371
rect 92 337 126 371
rect 41 335 160 337
rect 41 303 60 335
rect 94 303 160 335
rect 41 269 58 303
rect 94 301 126 303
rect 92 269 126 301
rect 41 263 160 269
rect 41 235 60 263
rect 94 235 160 263
rect 41 201 58 235
rect 94 229 126 235
rect 92 201 126 229
rect 41 185 160 201
rect 212 507 246 523
rect 212 439 246 445
rect 212 371 246 373
rect 212 335 246 337
rect 212 263 246 269
rect 212 185 246 201
rect 298 507 332 523
rect 298 439 332 445
rect 298 371 332 373
rect 298 335 332 337
rect 298 263 332 269
rect 298 185 332 201
rect 384 507 418 523
rect 384 439 418 445
rect 384 371 418 373
rect 384 335 418 337
rect 384 263 418 269
rect 384 185 418 201
rect 470 507 589 523
rect 504 479 538 507
rect 504 473 536 479
rect 572 473 589 507
rect 470 445 536 473
rect 570 445 589 473
rect 470 439 589 445
rect 504 407 538 439
rect 504 405 536 407
rect 572 405 589 439
rect 470 373 536 405
rect 570 373 589 405
rect 470 371 589 373
rect 504 337 538 371
rect 572 337 589 371
rect 470 335 589 337
rect 470 303 536 335
rect 570 303 589 335
rect 504 301 536 303
rect 504 269 538 301
rect 572 269 589 303
rect 470 263 589 269
rect 470 235 536 263
rect 570 235 589 263
rect 504 229 536 235
rect 504 201 538 229
rect 572 201 589 235
rect 470 185 589 201
rect 120 163 160 185
rect 470 163 510 185
rect 120 147 186 163
rect 120 113 136 147
rect 170 113 186 147
rect 444 147 510 163
rect 120 97 186 113
rect 248 125 382 139
rect 248 19 262 125
rect 368 19 382 125
rect 444 113 460 147
rect 494 113 510 147
rect 444 97 510 113
rect 248 0 382 19
<< viali >>
rect 262 687 368 689
rect 262 585 264 687
rect 264 585 366 687
rect 366 585 368 687
rect 262 583 368 585
rect 60 473 92 479
rect 92 473 94 479
rect 60 445 94 473
rect 60 405 92 407
rect 92 405 94 407
rect 60 373 94 405
rect 60 303 94 335
rect 60 301 92 303
rect 92 301 94 303
rect 60 235 94 263
rect 60 229 92 235
rect 92 229 94 235
rect 212 473 246 479
rect 212 445 246 473
rect 212 405 246 407
rect 212 373 246 405
rect 212 303 246 335
rect 212 301 246 303
rect 212 235 246 263
rect 212 229 246 235
rect 298 473 332 479
rect 298 445 332 473
rect 298 405 332 407
rect 298 373 332 405
rect 298 303 332 335
rect 298 301 332 303
rect 298 235 332 263
rect 298 229 332 235
rect 384 473 418 479
rect 384 445 418 473
rect 384 405 418 407
rect 384 373 418 405
rect 384 303 418 335
rect 384 301 418 303
rect 384 235 418 263
rect 384 229 418 235
rect 536 473 538 479
rect 538 473 570 479
rect 536 445 570 473
rect 536 405 538 407
rect 538 405 570 407
rect 536 373 570 405
rect 536 303 570 335
rect 536 301 538 303
rect 538 301 570 303
rect 536 235 570 263
rect 536 229 538 235
rect 538 229 570 235
rect 262 123 368 125
rect 262 21 264 123
rect 264 21 366 123
rect 366 21 368 123
rect 262 19 368 21
<< metal1 >>
rect 250 689 380 708
rect 250 583 262 689
rect 368 583 380 689
rect 250 571 380 583
rect 41 479 100 507
rect 41 445 60 479
rect 94 445 100 479
rect 41 407 100 445
rect 41 373 60 407
rect 94 373 100 407
rect 41 335 100 373
rect 41 301 60 335
rect 94 301 100 335
rect 41 263 100 301
rect 41 229 60 263
rect 94 229 100 263
rect 41 201 100 229
rect 203 479 255 507
rect 203 445 212 479
rect 246 445 255 479
rect 203 407 255 445
rect 203 373 212 407
rect 246 373 255 407
rect 203 335 255 373
rect 203 323 212 335
rect 246 323 255 335
rect 203 263 255 271
rect 203 259 212 263
rect 246 259 255 263
rect 203 201 255 207
rect 289 501 341 507
rect 289 445 298 449
rect 332 445 341 449
rect 289 437 341 445
rect 289 373 298 385
rect 332 373 341 385
rect 289 335 341 373
rect 289 301 298 335
rect 332 301 341 335
rect 289 263 341 301
rect 289 229 298 263
rect 332 229 341 263
rect 289 201 341 229
rect 375 479 427 507
rect 375 445 384 479
rect 418 445 427 479
rect 375 407 427 445
rect 375 373 384 407
rect 418 373 427 407
rect 375 335 427 373
rect 375 323 384 335
rect 418 323 427 335
rect 375 263 427 271
rect 375 259 384 263
rect 418 259 427 263
rect 375 201 427 207
rect 530 479 589 507
rect 530 445 536 479
rect 570 445 589 479
rect 530 407 589 445
rect 530 373 536 407
rect 570 373 589 407
rect 530 335 589 373
rect 530 301 536 335
rect 570 301 589 335
rect 530 263 589 301
rect 530 229 536 263
rect 570 229 589 263
rect 530 201 589 229
rect 250 125 380 137
rect 250 19 262 125
rect 368 19 380 125
rect 250 0 380 19
<< via1 >>
rect 203 301 212 323
rect 212 301 246 323
rect 246 301 255 323
rect 203 271 255 301
rect 203 229 212 259
rect 212 229 246 259
rect 246 229 255 259
rect 203 207 255 229
rect 289 479 341 501
rect 289 449 298 479
rect 298 449 332 479
rect 332 449 341 479
rect 289 407 341 437
rect 289 385 298 407
rect 298 385 332 407
rect 332 385 341 407
rect 375 301 384 323
rect 384 301 418 323
rect 418 301 427 323
rect 375 271 427 301
rect 375 229 384 259
rect 384 229 418 259
rect 418 229 427 259
rect 375 207 427 229
<< metal2 >>
rect 14 501 616 507
rect 14 449 289 501
rect 341 449 616 501
rect 14 437 616 449
rect 14 385 289 437
rect 341 385 616 437
rect 14 379 616 385
rect 14 323 616 329
rect 14 271 203 323
rect 255 271 375 323
rect 427 271 616 323
rect 14 259 616 271
rect 14 207 203 259
rect 255 207 375 259
rect 427 207 616 259
rect 14 201 616 207
<< labels >>
flabel comment s 182 360 182 360 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 442 350 442 350 0 FreeSans 180 90 0 0 dummy_poly
flabel metal1 s 255 608 374 659 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 255 44 374 95 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 543 339 589 369 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 41 339 87 369 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal2 s 14 201 35 329 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 14 379 35 507 7 FreeSans 300 180 0 0 DRAIN
port 1 nsew
<< properties >>
string GDS_END 2907912
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 2896952
string device primitive
<< end >>
