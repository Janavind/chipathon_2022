magic
tech sky130A
timestamp 1666199351
<< properties >>
string GDS_END 238102
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 234194
<< end >>
