magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< dnwell >>
tri -500 6514 -414 6600 se
rect -414 6514 564 6600
tri 564 6514 650 6600 sw
rect -500 -514 650 6514
tri -500 -600 -414 -514 ne
rect -414 -600 564 -514
tri 564 -600 650 -514 nw
<< nwell >>
rect -10 0 160 6000
<< pwell >>
rect -1866 6874 2016 7008
rect -1866 6026 -1732 6874
rect 1882 6026 2016 6874
rect -1866 -26 -374 6026
rect 524 -26 2016 6026
rect -1866 -874 -1732 -26
rect 1882 -874 2016 -26
rect -1866 -1008 2016 -874
<< obsactive >>
rect -2044 -1182 2186 7182
<< locali >>
rect -1840 6900 1990 6982
rect -1840 -900 -1758 6900
rect -1662 5969 -1596 5991
rect -1662 5935 -1646 5969
rect -1612 5935 -1596 5969
rect -1662 5897 -1596 5935
rect -1662 5863 -1646 5897
rect -1612 5863 -1596 5897
rect -1662 5825 -1596 5863
rect -1662 5791 -1646 5825
rect -1612 5791 -1596 5825
rect -1662 5753 -1596 5791
rect -1662 5719 -1646 5753
rect -1612 5719 -1596 5753
rect -1662 5681 -1596 5719
rect -1662 5647 -1646 5681
rect -1612 5647 -1596 5681
rect -1662 5609 -1596 5647
rect -1662 5575 -1646 5609
rect -1612 5575 -1596 5609
rect -1662 5537 -1596 5575
rect -1662 5503 -1646 5537
rect -1612 5503 -1596 5537
rect -1662 5465 -1596 5503
rect -1662 5431 -1646 5465
rect -1612 5431 -1596 5465
rect -1662 5393 -1596 5431
rect -1662 5359 -1646 5393
rect -1612 5359 -1596 5393
rect -1662 5321 -1596 5359
rect -1662 5287 -1646 5321
rect -1612 5287 -1596 5321
rect -1662 5249 -1596 5287
rect -1662 5215 -1646 5249
rect -1612 5215 -1596 5249
rect -1662 5177 -1596 5215
rect -1662 5143 -1646 5177
rect -1612 5143 -1596 5177
rect -1662 5105 -1596 5143
rect -1662 5071 -1646 5105
rect -1612 5071 -1596 5105
rect -1662 5033 -1596 5071
rect -1662 4999 -1646 5033
rect -1612 4999 -1596 5033
rect -1662 4961 -1596 4999
rect -1662 4927 -1646 4961
rect -1612 4927 -1596 4961
rect -1662 4889 -1596 4927
rect -1662 4855 -1646 4889
rect -1612 4855 -1596 4889
rect -1662 4817 -1596 4855
rect -1662 4783 -1646 4817
rect -1612 4783 -1596 4817
rect -1662 4745 -1596 4783
rect -1662 4711 -1646 4745
rect -1612 4711 -1596 4745
rect -1662 4673 -1596 4711
rect -1662 4639 -1646 4673
rect -1612 4639 -1596 4673
rect -1662 4601 -1596 4639
rect -1662 4567 -1646 4601
rect -1612 4567 -1596 4601
rect -1662 4529 -1596 4567
rect -1662 4495 -1646 4529
rect -1612 4495 -1596 4529
rect -1662 4457 -1596 4495
rect -1662 4423 -1646 4457
rect -1612 4423 -1596 4457
rect -1662 4385 -1596 4423
rect -1662 4351 -1646 4385
rect -1612 4351 -1596 4385
rect -1662 4313 -1596 4351
rect -1662 4279 -1646 4313
rect -1612 4279 -1596 4313
rect -1662 4241 -1596 4279
rect -1662 4207 -1646 4241
rect -1612 4207 -1596 4241
rect -1662 4169 -1596 4207
rect -1662 4135 -1646 4169
rect -1612 4135 -1596 4169
rect -1662 4097 -1596 4135
rect -1662 4063 -1646 4097
rect -1612 4063 -1596 4097
rect -1662 4025 -1596 4063
rect -1662 3991 -1646 4025
rect -1612 3991 -1596 4025
rect -1662 3953 -1596 3991
rect -1662 3919 -1646 3953
rect -1612 3919 -1596 3953
rect -1662 3881 -1596 3919
rect -1662 3847 -1646 3881
rect -1612 3847 -1596 3881
rect -1662 3809 -1596 3847
rect -1662 3775 -1646 3809
rect -1612 3775 -1596 3809
rect -1662 3737 -1596 3775
rect -1662 3703 -1646 3737
rect -1612 3703 -1596 3737
rect -1662 3665 -1596 3703
rect -1662 3631 -1646 3665
rect -1612 3631 -1596 3665
rect -1662 3593 -1596 3631
rect -1662 3559 -1646 3593
rect -1612 3559 -1596 3593
rect -1662 3521 -1596 3559
rect -1662 3487 -1646 3521
rect -1612 3487 -1596 3521
rect -1662 3449 -1596 3487
rect -1662 3415 -1646 3449
rect -1612 3415 -1596 3449
rect -1662 3377 -1596 3415
rect -1662 3343 -1646 3377
rect -1612 3343 -1596 3377
rect -1662 3305 -1596 3343
rect -1662 3271 -1646 3305
rect -1612 3271 -1596 3305
rect -1662 3233 -1596 3271
rect -1662 3199 -1646 3233
rect -1612 3199 -1596 3233
rect -1662 3161 -1596 3199
rect -1662 3127 -1646 3161
rect -1612 3127 -1596 3161
rect -1662 3089 -1596 3127
rect -1662 3055 -1646 3089
rect -1612 3055 -1596 3089
rect -1662 3017 -1596 3055
rect -1662 2983 -1646 3017
rect -1612 2983 -1596 3017
rect -1662 2945 -1596 2983
rect -1662 2911 -1646 2945
rect -1612 2911 -1596 2945
rect -1662 2873 -1596 2911
rect -1662 2839 -1646 2873
rect -1612 2839 -1596 2873
rect -1662 2801 -1596 2839
rect -1662 2767 -1646 2801
rect -1612 2767 -1596 2801
rect -1662 2729 -1596 2767
rect -1662 2695 -1646 2729
rect -1612 2695 -1596 2729
rect -1662 2657 -1596 2695
rect -1662 2623 -1646 2657
rect -1612 2623 -1596 2657
rect -1662 2585 -1596 2623
rect -1662 2551 -1646 2585
rect -1612 2551 -1596 2585
rect -1662 2513 -1596 2551
rect -1662 2479 -1646 2513
rect -1612 2479 -1596 2513
rect -1662 2441 -1596 2479
rect -1662 2407 -1646 2441
rect -1612 2407 -1596 2441
rect -1662 2369 -1596 2407
rect -1662 2335 -1646 2369
rect -1612 2335 -1596 2369
rect -1662 2297 -1596 2335
rect -1662 2263 -1646 2297
rect -1612 2263 -1596 2297
rect -1662 2225 -1596 2263
rect -1662 2191 -1646 2225
rect -1612 2191 -1596 2225
rect -1662 2153 -1596 2191
rect -1662 2119 -1646 2153
rect -1612 2119 -1596 2153
rect -1662 2081 -1596 2119
rect -1662 2047 -1646 2081
rect -1612 2047 -1596 2081
rect -1662 2009 -1596 2047
rect -1662 1975 -1646 2009
rect -1612 1975 -1596 2009
rect -1662 1937 -1596 1975
rect -1662 1903 -1646 1937
rect -1612 1903 -1596 1937
rect -1662 1865 -1596 1903
rect -1662 1831 -1646 1865
rect -1612 1831 -1596 1865
rect -1662 1793 -1596 1831
rect -1662 1759 -1646 1793
rect -1612 1759 -1596 1793
rect -1662 1721 -1596 1759
rect -1662 1687 -1646 1721
rect -1612 1687 -1596 1721
rect -1662 1649 -1596 1687
rect -1662 1615 -1646 1649
rect -1612 1615 -1596 1649
rect -1662 1577 -1596 1615
rect -1662 1543 -1646 1577
rect -1612 1543 -1596 1577
rect -1662 1505 -1596 1543
rect -1662 1471 -1646 1505
rect -1612 1471 -1596 1505
rect -1662 1433 -1596 1471
rect -1662 1399 -1646 1433
rect -1612 1399 -1596 1433
rect -1662 1361 -1596 1399
rect -1662 1327 -1646 1361
rect -1612 1327 -1596 1361
rect -1662 1289 -1596 1327
rect -1662 1255 -1646 1289
rect -1612 1255 -1596 1289
rect -1662 1217 -1596 1255
rect -1662 1183 -1646 1217
rect -1612 1183 -1596 1217
rect -1662 1145 -1596 1183
rect -1662 1111 -1646 1145
rect -1612 1111 -1596 1145
rect -1662 1073 -1596 1111
rect -1662 1039 -1646 1073
rect -1612 1039 -1596 1073
rect -1662 1001 -1596 1039
rect -1662 967 -1646 1001
rect -1612 967 -1596 1001
rect -1662 929 -1596 967
rect -1662 895 -1646 929
rect -1612 895 -1596 929
rect -1662 857 -1596 895
rect -1662 823 -1646 857
rect -1612 823 -1596 857
rect -1662 785 -1596 823
rect -1662 751 -1646 785
rect -1612 751 -1596 785
rect -1662 713 -1596 751
rect -1662 679 -1646 713
rect -1612 679 -1596 713
rect -1662 641 -1596 679
rect -1662 607 -1646 641
rect -1612 607 -1596 641
rect -1662 569 -1596 607
rect -1662 535 -1646 569
rect -1612 535 -1596 569
rect -1662 497 -1596 535
rect -1662 463 -1646 497
rect -1612 463 -1596 497
rect -1662 425 -1596 463
rect -1662 391 -1646 425
rect -1612 391 -1596 425
rect -1662 353 -1596 391
rect -1662 319 -1646 353
rect -1612 319 -1596 353
rect -1662 281 -1596 319
rect -1662 247 -1646 281
rect -1612 247 -1596 281
rect -1662 209 -1596 247
rect -1662 175 -1646 209
rect -1612 175 -1596 209
rect -1662 137 -1596 175
rect -1662 103 -1646 137
rect -1612 103 -1596 137
rect -1662 65 -1596 103
rect -1662 31 -1646 65
rect -1612 31 -1596 65
rect -1662 9 -1596 31
rect -25 5969 175 6050
rect -25 31 22 5969
rect 128 31 175 5969
rect -25 -50 175 31
rect 1746 5969 1812 5991
rect 1746 5935 1762 5969
rect 1796 5935 1812 5969
rect 1746 5897 1812 5935
rect 1746 5863 1762 5897
rect 1796 5863 1812 5897
rect 1746 5825 1812 5863
rect 1746 5791 1762 5825
rect 1796 5791 1812 5825
rect 1746 5753 1812 5791
rect 1746 5719 1762 5753
rect 1796 5719 1812 5753
rect 1746 5681 1812 5719
rect 1746 5647 1762 5681
rect 1796 5647 1812 5681
rect 1746 5609 1812 5647
rect 1746 5575 1762 5609
rect 1796 5575 1812 5609
rect 1746 5537 1812 5575
rect 1746 5503 1762 5537
rect 1796 5503 1812 5537
rect 1746 5465 1812 5503
rect 1746 5431 1762 5465
rect 1796 5431 1812 5465
rect 1746 5393 1812 5431
rect 1746 5359 1762 5393
rect 1796 5359 1812 5393
rect 1746 5321 1812 5359
rect 1746 5287 1762 5321
rect 1796 5287 1812 5321
rect 1746 5249 1812 5287
rect 1746 5215 1762 5249
rect 1796 5215 1812 5249
rect 1746 5177 1812 5215
rect 1746 5143 1762 5177
rect 1796 5143 1812 5177
rect 1746 5105 1812 5143
rect 1746 5071 1762 5105
rect 1796 5071 1812 5105
rect 1746 5033 1812 5071
rect 1746 4999 1762 5033
rect 1796 4999 1812 5033
rect 1746 4961 1812 4999
rect 1746 4927 1762 4961
rect 1796 4927 1812 4961
rect 1746 4889 1812 4927
rect 1746 4855 1762 4889
rect 1796 4855 1812 4889
rect 1746 4817 1812 4855
rect 1746 4783 1762 4817
rect 1796 4783 1812 4817
rect 1746 4745 1812 4783
rect 1746 4711 1762 4745
rect 1796 4711 1812 4745
rect 1746 4673 1812 4711
rect 1746 4639 1762 4673
rect 1796 4639 1812 4673
rect 1746 4601 1812 4639
rect 1746 4567 1762 4601
rect 1796 4567 1812 4601
rect 1746 4529 1812 4567
rect 1746 4495 1762 4529
rect 1796 4495 1812 4529
rect 1746 4457 1812 4495
rect 1746 4423 1762 4457
rect 1796 4423 1812 4457
rect 1746 4385 1812 4423
rect 1746 4351 1762 4385
rect 1796 4351 1812 4385
rect 1746 4313 1812 4351
rect 1746 4279 1762 4313
rect 1796 4279 1812 4313
rect 1746 4241 1812 4279
rect 1746 4207 1762 4241
rect 1796 4207 1812 4241
rect 1746 4169 1812 4207
rect 1746 4135 1762 4169
rect 1796 4135 1812 4169
rect 1746 4097 1812 4135
rect 1746 4063 1762 4097
rect 1796 4063 1812 4097
rect 1746 4025 1812 4063
rect 1746 3991 1762 4025
rect 1796 3991 1812 4025
rect 1746 3953 1812 3991
rect 1746 3919 1762 3953
rect 1796 3919 1812 3953
rect 1746 3881 1812 3919
rect 1746 3847 1762 3881
rect 1796 3847 1812 3881
rect 1746 3809 1812 3847
rect 1746 3775 1762 3809
rect 1796 3775 1812 3809
rect 1746 3737 1812 3775
rect 1746 3703 1762 3737
rect 1796 3703 1812 3737
rect 1746 3665 1812 3703
rect 1746 3631 1762 3665
rect 1796 3631 1812 3665
rect 1746 3593 1812 3631
rect 1746 3559 1762 3593
rect 1796 3559 1812 3593
rect 1746 3521 1812 3559
rect 1746 3487 1762 3521
rect 1796 3487 1812 3521
rect 1746 3449 1812 3487
rect 1746 3415 1762 3449
rect 1796 3415 1812 3449
rect 1746 3377 1812 3415
rect 1746 3343 1762 3377
rect 1796 3343 1812 3377
rect 1746 3305 1812 3343
rect 1746 3271 1762 3305
rect 1796 3271 1812 3305
rect 1746 3233 1812 3271
rect 1746 3199 1762 3233
rect 1796 3199 1812 3233
rect 1746 3161 1812 3199
rect 1746 3127 1762 3161
rect 1796 3127 1812 3161
rect 1746 3089 1812 3127
rect 1746 3055 1762 3089
rect 1796 3055 1812 3089
rect 1746 3017 1812 3055
rect 1746 2983 1762 3017
rect 1796 2983 1812 3017
rect 1746 2945 1812 2983
rect 1746 2911 1762 2945
rect 1796 2911 1812 2945
rect 1746 2873 1812 2911
rect 1746 2839 1762 2873
rect 1796 2839 1812 2873
rect 1746 2801 1812 2839
rect 1746 2767 1762 2801
rect 1796 2767 1812 2801
rect 1746 2729 1812 2767
rect 1746 2695 1762 2729
rect 1796 2695 1812 2729
rect 1746 2657 1812 2695
rect 1746 2623 1762 2657
rect 1796 2623 1812 2657
rect 1746 2585 1812 2623
rect 1746 2551 1762 2585
rect 1796 2551 1812 2585
rect 1746 2513 1812 2551
rect 1746 2479 1762 2513
rect 1796 2479 1812 2513
rect 1746 2441 1812 2479
rect 1746 2407 1762 2441
rect 1796 2407 1812 2441
rect 1746 2369 1812 2407
rect 1746 2335 1762 2369
rect 1796 2335 1812 2369
rect 1746 2297 1812 2335
rect 1746 2263 1762 2297
rect 1796 2263 1812 2297
rect 1746 2225 1812 2263
rect 1746 2191 1762 2225
rect 1796 2191 1812 2225
rect 1746 2153 1812 2191
rect 1746 2119 1762 2153
rect 1796 2119 1812 2153
rect 1746 2081 1812 2119
rect 1746 2047 1762 2081
rect 1796 2047 1812 2081
rect 1746 2009 1812 2047
rect 1746 1975 1762 2009
rect 1796 1975 1812 2009
rect 1746 1937 1812 1975
rect 1746 1903 1762 1937
rect 1796 1903 1812 1937
rect 1746 1865 1812 1903
rect 1746 1831 1762 1865
rect 1796 1831 1812 1865
rect 1746 1793 1812 1831
rect 1746 1759 1762 1793
rect 1796 1759 1812 1793
rect 1746 1721 1812 1759
rect 1746 1687 1762 1721
rect 1796 1687 1812 1721
rect 1746 1649 1812 1687
rect 1746 1615 1762 1649
rect 1796 1615 1812 1649
rect 1746 1577 1812 1615
rect 1746 1543 1762 1577
rect 1796 1543 1812 1577
rect 1746 1505 1812 1543
rect 1746 1471 1762 1505
rect 1796 1471 1812 1505
rect 1746 1433 1812 1471
rect 1746 1399 1762 1433
rect 1796 1399 1812 1433
rect 1746 1361 1812 1399
rect 1746 1327 1762 1361
rect 1796 1327 1812 1361
rect 1746 1289 1812 1327
rect 1746 1255 1762 1289
rect 1796 1255 1812 1289
rect 1746 1217 1812 1255
rect 1746 1183 1762 1217
rect 1796 1183 1812 1217
rect 1746 1145 1812 1183
rect 1746 1111 1762 1145
rect 1796 1111 1812 1145
rect 1746 1073 1812 1111
rect 1746 1039 1762 1073
rect 1796 1039 1812 1073
rect 1746 1001 1812 1039
rect 1746 967 1762 1001
rect 1796 967 1812 1001
rect 1746 929 1812 967
rect 1746 895 1762 929
rect 1796 895 1812 929
rect 1746 857 1812 895
rect 1746 823 1762 857
rect 1796 823 1812 857
rect 1746 785 1812 823
rect 1746 751 1762 785
rect 1796 751 1812 785
rect 1746 713 1812 751
rect 1746 679 1762 713
rect 1796 679 1812 713
rect 1746 641 1812 679
rect 1746 607 1762 641
rect 1796 607 1812 641
rect 1746 569 1812 607
rect 1746 535 1762 569
rect 1796 535 1812 569
rect 1746 497 1812 535
rect 1746 463 1762 497
rect 1796 463 1812 497
rect 1746 425 1812 463
rect 1746 391 1762 425
rect 1796 391 1812 425
rect 1746 353 1812 391
rect 1746 319 1762 353
rect 1796 319 1812 353
rect 1746 281 1812 319
rect 1746 247 1762 281
rect 1796 247 1812 281
rect 1746 209 1812 247
rect 1746 175 1762 209
rect 1796 175 1812 209
rect 1746 137 1812 175
rect 1746 103 1762 137
rect 1796 103 1812 137
rect 1746 65 1812 103
rect 1746 31 1762 65
rect 1796 31 1812 65
rect 1746 9 1812 31
rect -296 -459 460 -443
rect -296 -493 -280 -459
rect -246 -493 -206 -459
rect -172 -493 -132 -459
rect -98 -493 -58 -459
rect -24 -493 16 -459
rect 50 -493 90 -459
rect 124 -493 164 -459
rect 198 -493 238 -459
rect 272 -493 312 -459
rect 346 -493 386 -459
rect 420 -493 460 -459
rect -296 -533 460 -493
rect -296 -567 -280 -533
rect -246 -567 -206 -533
rect -172 -567 -132 -533
rect -98 -567 -58 -533
rect -24 -567 16 -533
rect 50 -567 90 -533
rect 124 -567 164 -533
rect 198 -567 238 -533
rect 272 -567 312 -533
rect 346 -567 386 -533
rect 420 -567 460 -533
rect -296 -607 460 -567
rect -296 -641 -280 -607
rect -246 -641 -206 -607
rect -172 -641 -132 -607
rect -98 -641 -58 -607
rect -24 -641 16 -607
rect 50 -641 90 -607
rect 124 -641 164 -607
rect 198 -641 238 -607
rect 272 -641 312 -607
rect 346 -641 386 -607
rect 420 -641 460 -607
rect -296 -657 460 -641
rect 1908 -900 1990 6900
rect -1840 -982 1990 -900
<< viali >>
rect -1646 5935 -1612 5969
rect -1646 5863 -1612 5897
rect -1646 5791 -1612 5825
rect -1646 5719 -1612 5753
rect -1646 5647 -1612 5681
rect -1646 5575 -1612 5609
rect -1646 5503 -1612 5537
rect -1646 5431 -1612 5465
rect -1646 5359 -1612 5393
rect -1646 5287 -1612 5321
rect -1646 5215 -1612 5249
rect -1646 5143 -1612 5177
rect -1646 5071 -1612 5105
rect -1646 4999 -1612 5033
rect -1646 4927 -1612 4961
rect -1646 4855 -1612 4889
rect -1646 4783 -1612 4817
rect -1646 4711 -1612 4745
rect -1646 4639 -1612 4673
rect -1646 4567 -1612 4601
rect -1646 4495 -1612 4529
rect -1646 4423 -1612 4457
rect -1646 4351 -1612 4385
rect -1646 4279 -1612 4313
rect -1646 4207 -1612 4241
rect -1646 4135 -1612 4169
rect -1646 4063 -1612 4097
rect -1646 3991 -1612 4025
rect -1646 3919 -1612 3953
rect -1646 3847 -1612 3881
rect -1646 3775 -1612 3809
rect -1646 3703 -1612 3737
rect -1646 3631 -1612 3665
rect -1646 3559 -1612 3593
rect -1646 3487 -1612 3521
rect -1646 3415 -1612 3449
rect -1646 3343 -1612 3377
rect -1646 3271 -1612 3305
rect -1646 3199 -1612 3233
rect -1646 3127 -1612 3161
rect -1646 3055 -1612 3089
rect -1646 2983 -1612 3017
rect -1646 2911 -1612 2945
rect -1646 2839 -1612 2873
rect -1646 2767 -1612 2801
rect -1646 2695 -1612 2729
rect -1646 2623 -1612 2657
rect -1646 2551 -1612 2585
rect -1646 2479 -1612 2513
rect -1646 2407 -1612 2441
rect -1646 2335 -1612 2369
rect -1646 2263 -1612 2297
rect -1646 2191 -1612 2225
rect -1646 2119 -1612 2153
rect -1646 2047 -1612 2081
rect -1646 1975 -1612 2009
rect -1646 1903 -1612 1937
rect -1646 1831 -1612 1865
rect -1646 1759 -1612 1793
rect -1646 1687 -1612 1721
rect -1646 1615 -1612 1649
rect -1646 1543 -1612 1577
rect -1646 1471 -1612 1505
rect -1646 1399 -1612 1433
rect -1646 1327 -1612 1361
rect -1646 1255 -1612 1289
rect -1646 1183 -1612 1217
rect -1646 1111 -1612 1145
rect -1646 1039 -1612 1073
rect -1646 967 -1612 1001
rect -1646 895 -1612 929
rect -1646 823 -1612 857
rect -1646 751 -1612 785
rect -1646 679 -1612 713
rect -1646 607 -1612 641
rect -1646 535 -1612 569
rect -1646 463 -1612 497
rect -1646 391 -1612 425
rect -1646 319 -1612 353
rect -1646 247 -1612 281
rect -1646 175 -1612 209
rect -1646 103 -1612 137
rect -1646 31 -1612 65
rect 22 31 128 5969
rect 1762 5935 1796 5969
rect 1762 5863 1796 5897
rect 1762 5791 1796 5825
rect 1762 5719 1796 5753
rect 1762 5647 1796 5681
rect 1762 5575 1796 5609
rect 1762 5503 1796 5537
rect 1762 5431 1796 5465
rect 1762 5359 1796 5393
rect 1762 5287 1796 5321
rect 1762 5215 1796 5249
rect 1762 5143 1796 5177
rect 1762 5071 1796 5105
rect 1762 4999 1796 5033
rect 1762 4927 1796 4961
rect 1762 4855 1796 4889
rect 1762 4783 1796 4817
rect 1762 4711 1796 4745
rect 1762 4639 1796 4673
rect 1762 4567 1796 4601
rect 1762 4495 1796 4529
rect 1762 4423 1796 4457
rect 1762 4351 1796 4385
rect 1762 4279 1796 4313
rect 1762 4207 1796 4241
rect 1762 4135 1796 4169
rect 1762 4063 1796 4097
rect 1762 3991 1796 4025
rect 1762 3919 1796 3953
rect 1762 3847 1796 3881
rect 1762 3775 1796 3809
rect 1762 3703 1796 3737
rect 1762 3631 1796 3665
rect 1762 3559 1796 3593
rect 1762 3487 1796 3521
rect 1762 3415 1796 3449
rect 1762 3343 1796 3377
rect 1762 3271 1796 3305
rect 1762 3199 1796 3233
rect 1762 3127 1796 3161
rect 1762 3055 1796 3089
rect 1762 2983 1796 3017
rect 1762 2911 1796 2945
rect 1762 2839 1796 2873
rect 1762 2767 1796 2801
rect 1762 2695 1796 2729
rect 1762 2623 1796 2657
rect 1762 2551 1796 2585
rect 1762 2479 1796 2513
rect 1762 2407 1796 2441
rect 1762 2335 1796 2369
rect 1762 2263 1796 2297
rect 1762 2191 1796 2225
rect 1762 2119 1796 2153
rect 1762 2047 1796 2081
rect 1762 1975 1796 2009
rect 1762 1903 1796 1937
rect 1762 1831 1796 1865
rect 1762 1759 1796 1793
rect 1762 1687 1796 1721
rect 1762 1615 1796 1649
rect 1762 1543 1796 1577
rect 1762 1471 1796 1505
rect 1762 1399 1796 1433
rect 1762 1327 1796 1361
rect 1762 1255 1796 1289
rect 1762 1183 1796 1217
rect 1762 1111 1796 1145
rect 1762 1039 1796 1073
rect 1762 967 1796 1001
rect 1762 895 1796 929
rect 1762 823 1796 857
rect 1762 751 1796 785
rect 1762 679 1796 713
rect 1762 607 1796 641
rect 1762 535 1796 569
rect 1762 463 1796 497
rect 1762 391 1796 425
rect 1762 319 1796 353
rect 1762 247 1796 281
rect 1762 175 1796 209
rect 1762 103 1796 137
rect 1762 31 1796 65
rect -280 -493 -246 -459
rect -206 -493 -172 -459
rect -132 -493 -98 -459
rect -58 -493 -24 -459
rect 16 -493 50 -459
rect 90 -493 124 -459
rect 164 -493 198 -459
rect 238 -493 272 -459
rect 312 -493 346 -459
rect 386 -493 420 -459
rect -280 -567 -246 -533
rect -206 -567 -172 -533
rect -132 -567 -98 -533
rect -58 -567 -24 -533
rect 16 -567 50 -533
rect 90 -567 124 -533
rect 164 -567 198 -533
rect 238 -567 272 -533
rect 312 -567 346 -533
rect 386 -567 420 -533
rect -280 -641 -246 -607
rect -206 -641 -172 -607
rect -132 -641 -98 -607
rect -58 -641 -24 -607
rect 16 -641 50 -607
rect 90 -641 124 -607
rect 164 -641 198 -607
rect 238 -641 272 -607
rect 312 -641 346 -607
rect 386 -641 420 -607
<< metal1 >>
rect -1712 5969 -1112 6200
rect -1712 5935 -1646 5969
rect -1612 5935 -1112 5969
rect -1712 5897 -1112 5935
rect -1712 5863 -1646 5897
rect -1612 5863 -1112 5897
rect -1712 5825 -1112 5863
rect -1712 5791 -1646 5825
rect -1612 5791 -1112 5825
rect -1712 5753 -1112 5791
rect -1712 5719 -1646 5753
rect -1612 5719 -1112 5753
rect -1712 5681 -1112 5719
rect -1712 5647 -1646 5681
rect -1612 5647 -1112 5681
rect -1712 5609 -1112 5647
rect -1712 5575 -1646 5609
rect -1612 5575 -1112 5609
rect -1712 5537 -1112 5575
rect -1712 5503 -1646 5537
rect -1612 5503 -1112 5537
rect -1712 5465 -1112 5503
rect -1712 5431 -1646 5465
rect -1612 5431 -1112 5465
rect -1712 5393 -1112 5431
rect -1712 5359 -1646 5393
rect -1612 5359 -1112 5393
rect -1712 5321 -1112 5359
rect -1712 5287 -1646 5321
rect -1612 5287 -1112 5321
rect -1712 5249 -1112 5287
rect -1712 5215 -1646 5249
rect -1612 5215 -1112 5249
rect -1712 5177 -1112 5215
rect -1712 5143 -1646 5177
rect -1612 5143 -1112 5177
rect -1712 5105 -1112 5143
rect -1712 5071 -1646 5105
rect -1612 5071 -1112 5105
rect -1712 5033 -1112 5071
rect -1712 4999 -1646 5033
rect -1612 4999 -1112 5033
rect -1712 4961 -1112 4999
rect -1712 4927 -1646 4961
rect -1612 4927 -1112 4961
rect -1712 4889 -1112 4927
rect -1712 4855 -1646 4889
rect -1612 4855 -1112 4889
rect -1712 4817 -1112 4855
rect -1712 4783 -1646 4817
rect -1612 4783 -1112 4817
rect -1712 4745 -1112 4783
rect -1712 4711 -1646 4745
rect -1612 4711 -1112 4745
rect -1712 4673 -1112 4711
rect -1712 4639 -1646 4673
rect -1612 4639 -1112 4673
rect -1712 4601 -1112 4639
rect -1712 4567 -1646 4601
rect -1612 4567 -1112 4601
rect -1712 4529 -1112 4567
rect -1712 4495 -1646 4529
rect -1612 4495 -1112 4529
rect -1712 4457 -1112 4495
rect -1712 4423 -1646 4457
rect -1612 4423 -1112 4457
rect -1712 4385 -1112 4423
rect -1712 4351 -1646 4385
rect -1612 4351 -1112 4385
rect -1712 4313 -1112 4351
rect -1712 4279 -1646 4313
rect -1612 4279 -1112 4313
rect -1712 4241 -1112 4279
rect -1712 4207 -1646 4241
rect -1612 4207 -1112 4241
rect -1712 4169 -1112 4207
rect -1712 4135 -1646 4169
rect -1612 4135 -1112 4169
rect -1712 4097 -1112 4135
rect -1712 4063 -1646 4097
rect -1612 4063 -1112 4097
rect -1712 4025 -1112 4063
rect -1712 3991 -1646 4025
rect -1612 3991 -1112 4025
rect -1712 3953 -1112 3991
rect -1712 3919 -1646 3953
rect -1612 3919 -1112 3953
rect -1712 3881 -1112 3919
rect -1712 3847 -1646 3881
rect -1612 3847 -1112 3881
rect -1712 3809 -1112 3847
rect -1712 3775 -1646 3809
rect -1612 3775 -1112 3809
rect -1712 3737 -1112 3775
rect -1712 3703 -1646 3737
rect -1612 3703 -1112 3737
rect -1712 3665 -1112 3703
rect -1712 3631 -1646 3665
rect -1612 3631 -1112 3665
rect -1712 3593 -1112 3631
rect -1712 3559 -1646 3593
rect -1612 3559 -1112 3593
rect -1712 3521 -1112 3559
rect -1712 3487 -1646 3521
rect -1612 3487 -1112 3521
rect -1712 3449 -1112 3487
rect -1712 3415 -1646 3449
rect -1612 3415 -1112 3449
rect -1712 3377 -1112 3415
rect -1712 3343 -1646 3377
rect -1612 3343 -1112 3377
rect -1712 3305 -1112 3343
rect -1712 3271 -1646 3305
rect -1612 3271 -1112 3305
rect -1712 3233 -1112 3271
rect -1712 3199 -1646 3233
rect -1612 3199 -1112 3233
rect -1712 3161 -1112 3199
rect -1712 3127 -1646 3161
rect -1612 3127 -1112 3161
rect -1712 3089 -1112 3127
rect -1712 3055 -1646 3089
rect -1612 3055 -1112 3089
rect -1712 3017 -1112 3055
rect -1712 2983 -1646 3017
rect -1612 2983 -1112 3017
rect -1712 2945 -1112 2983
rect -1712 2911 -1646 2945
rect -1612 2911 -1112 2945
rect -1712 2873 -1112 2911
rect -1712 2839 -1646 2873
rect -1612 2839 -1112 2873
rect -1712 2801 -1112 2839
rect -1712 2767 -1646 2801
rect -1612 2767 -1112 2801
rect -1712 2729 -1112 2767
rect -1712 2695 -1646 2729
rect -1612 2695 -1112 2729
rect -1712 2657 -1112 2695
rect -1712 2623 -1646 2657
rect -1612 2623 -1112 2657
rect -1712 2585 -1112 2623
rect -1712 2551 -1646 2585
rect -1612 2551 -1112 2585
rect -1712 2513 -1112 2551
rect -1712 2479 -1646 2513
rect -1612 2479 -1112 2513
rect -1712 2441 -1112 2479
rect -1712 2407 -1646 2441
rect -1612 2407 -1112 2441
rect -1712 2369 -1112 2407
rect -1712 2335 -1646 2369
rect -1612 2335 -1112 2369
rect -1712 2297 -1112 2335
rect -1712 2263 -1646 2297
rect -1612 2263 -1112 2297
rect -1712 2225 -1112 2263
rect -1712 2191 -1646 2225
rect -1612 2191 -1112 2225
rect -1712 2153 -1112 2191
rect -1712 2119 -1646 2153
rect -1612 2119 -1112 2153
rect -1712 2081 -1112 2119
rect -1712 2047 -1646 2081
rect -1612 2047 -1112 2081
rect -1712 2009 -1112 2047
rect -1712 1975 -1646 2009
rect -1612 1975 -1112 2009
rect -1712 1937 -1112 1975
rect -1712 1903 -1646 1937
rect -1612 1903 -1112 1937
rect -1712 1865 -1112 1903
rect -1712 1831 -1646 1865
rect -1612 1831 -1112 1865
rect -1712 1793 -1112 1831
rect -1712 1759 -1646 1793
rect -1612 1759 -1112 1793
rect -1712 1721 -1112 1759
rect -1712 1687 -1646 1721
rect -1612 1687 -1112 1721
rect -1712 1649 -1112 1687
rect -1712 1615 -1646 1649
rect -1612 1615 -1112 1649
rect -1712 1577 -1112 1615
rect -1712 1543 -1646 1577
rect -1612 1543 -1112 1577
rect -1712 1505 -1112 1543
rect -1712 1471 -1646 1505
rect -1612 1471 -1112 1505
rect -1712 1433 -1112 1471
rect -1712 1399 -1646 1433
rect -1612 1399 -1112 1433
rect -1712 1361 -1112 1399
rect -1712 1327 -1646 1361
rect -1612 1327 -1112 1361
rect -1712 1289 -1112 1327
rect -1712 1255 -1646 1289
rect -1612 1255 -1112 1289
rect -1712 1217 -1112 1255
rect -1712 1183 -1646 1217
rect -1612 1183 -1112 1217
rect -1712 1145 -1112 1183
rect -1712 1111 -1646 1145
rect -1612 1111 -1112 1145
rect -1712 1073 -1112 1111
rect -1712 1039 -1646 1073
rect -1612 1039 -1112 1073
rect -1712 1001 -1112 1039
rect -1712 967 -1646 1001
rect -1612 967 -1112 1001
rect -1712 929 -1112 967
rect -1712 895 -1646 929
rect -1612 895 -1112 929
rect -1712 857 -1112 895
rect -1712 823 -1646 857
rect -1612 823 -1112 857
rect -1712 785 -1112 823
rect -1712 751 -1646 785
rect -1612 751 -1112 785
rect -1712 713 -1112 751
rect -1712 679 -1646 713
rect -1612 679 -1112 713
rect -1712 641 -1112 679
rect -1712 607 -1646 641
rect -1612 607 -1112 641
rect -1712 569 -1112 607
rect -1712 535 -1646 569
rect -1612 535 -1112 569
rect -1712 497 -1112 535
rect -1712 463 -1646 497
rect -1612 463 -1112 497
rect -1712 425 -1112 463
rect -1712 391 -1646 425
rect -1612 391 -1112 425
rect -1712 353 -1112 391
rect -1712 319 -1646 353
rect -1612 319 -1112 353
rect -1712 281 -1112 319
rect -1712 247 -1646 281
rect -1612 247 -1112 281
rect -1712 209 -1112 247
rect -1712 175 -1646 209
rect -1612 175 -1112 209
rect -1712 137 -1112 175
rect -1712 103 -1646 137
rect -1612 103 -1112 137
rect -1712 65 -1112 103
rect -1712 31 -1646 65
rect -1612 31 -1112 65
rect -1712 -200 -1112 31
rect -275 5969 425 6200
rect -275 31 22 5969
rect 128 31 425 5969
rect -275 -200 425 31
rect 1262 5969 1862 6200
rect 1262 5935 1762 5969
rect 1796 5935 1862 5969
rect 1262 5897 1862 5935
rect 1262 5863 1762 5897
rect 1796 5863 1862 5897
rect 1262 5825 1862 5863
rect 1262 5791 1762 5825
rect 1796 5791 1862 5825
rect 1262 5753 1862 5791
rect 1262 5719 1762 5753
rect 1796 5719 1862 5753
rect 1262 5681 1862 5719
rect 1262 5647 1762 5681
rect 1796 5647 1862 5681
rect 1262 5609 1862 5647
rect 1262 5575 1762 5609
rect 1796 5575 1862 5609
rect 1262 5537 1862 5575
rect 1262 5503 1762 5537
rect 1796 5503 1862 5537
rect 1262 5465 1862 5503
rect 1262 5431 1762 5465
rect 1796 5431 1862 5465
rect 1262 5393 1862 5431
rect 1262 5359 1762 5393
rect 1796 5359 1862 5393
rect 1262 5321 1862 5359
rect 1262 5287 1762 5321
rect 1796 5287 1862 5321
rect 1262 5249 1862 5287
rect 1262 5215 1762 5249
rect 1796 5215 1862 5249
rect 1262 5177 1862 5215
rect 1262 5143 1762 5177
rect 1796 5143 1862 5177
rect 1262 5105 1862 5143
rect 1262 5071 1762 5105
rect 1796 5071 1862 5105
rect 1262 5033 1862 5071
rect 1262 4999 1762 5033
rect 1796 4999 1862 5033
rect 1262 4961 1862 4999
rect 1262 4927 1762 4961
rect 1796 4927 1862 4961
rect 1262 4889 1862 4927
rect 1262 4855 1762 4889
rect 1796 4855 1862 4889
rect 1262 4817 1862 4855
rect 1262 4783 1762 4817
rect 1796 4783 1862 4817
rect 1262 4745 1862 4783
rect 1262 4711 1762 4745
rect 1796 4711 1862 4745
rect 1262 4673 1862 4711
rect 1262 4639 1762 4673
rect 1796 4639 1862 4673
rect 1262 4601 1862 4639
rect 1262 4567 1762 4601
rect 1796 4567 1862 4601
rect 1262 4529 1862 4567
rect 1262 4495 1762 4529
rect 1796 4495 1862 4529
rect 1262 4457 1862 4495
rect 1262 4423 1762 4457
rect 1796 4423 1862 4457
rect 1262 4385 1862 4423
rect 1262 4351 1762 4385
rect 1796 4351 1862 4385
rect 1262 4313 1862 4351
rect 1262 4279 1762 4313
rect 1796 4279 1862 4313
rect 1262 4241 1862 4279
rect 1262 4207 1762 4241
rect 1796 4207 1862 4241
rect 1262 4169 1862 4207
rect 1262 4135 1762 4169
rect 1796 4135 1862 4169
rect 1262 4097 1862 4135
rect 1262 4063 1762 4097
rect 1796 4063 1862 4097
rect 1262 4025 1862 4063
rect 1262 3991 1762 4025
rect 1796 3991 1862 4025
rect 1262 3953 1862 3991
rect 1262 3919 1762 3953
rect 1796 3919 1862 3953
rect 1262 3881 1862 3919
rect 1262 3847 1762 3881
rect 1796 3847 1862 3881
rect 1262 3809 1862 3847
rect 1262 3775 1762 3809
rect 1796 3775 1862 3809
rect 1262 3737 1862 3775
rect 1262 3703 1762 3737
rect 1796 3703 1862 3737
rect 1262 3665 1862 3703
rect 1262 3631 1762 3665
rect 1796 3631 1862 3665
rect 1262 3593 1862 3631
rect 1262 3559 1762 3593
rect 1796 3559 1862 3593
rect 1262 3521 1862 3559
rect 1262 3487 1762 3521
rect 1796 3487 1862 3521
rect 1262 3449 1862 3487
rect 1262 3415 1762 3449
rect 1796 3415 1862 3449
rect 1262 3377 1862 3415
rect 1262 3343 1762 3377
rect 1796 3343 1862 3377
rect 1262 3305 1862 3343
rect 1262 3271 1762 3305
rect 1796 3271 1862 3305
rect 1262 3233 1862 3271
rect 1262 3199 1762 3233
rect 1796 3199 1862 3233
rect 1262 3161 1862 3199
rect 1262 3127 1762 3161
rect 1796 3127 1862 3161
rect 1262 3089 1862 3127
rect 1262 3055 1762 3089
rect 1796 3055 1862 3089
rect 1262 3017 1862 3055
rect 1262 2983 1762 3017
rect 1796 2983 1862 3017
rect 1262 2945 1862 2983
rect 1262 2911 1762 2945
rect 1796 2911 1862 2945
rect 1262 2873 1862 2911
rect 1262 2839 1762 2873
rect 1796 2839 1862 2873
rect 1262 2801 1862 2839
rect 1262 2767 1762 2801
rect 1796 2767 1862 2801
rect 1262 2729 1862 2767
rect 1262 2695 1762 2729
rect 1796 2695 1862 2729
rect 1262 2657 1862 2695
rect 1262 2623 1762 2657
rect 1796 2623 1862 2657
rect 1262 2585 1862 2623
rect 1262 2551 1762 2585
rect 1796 2551 1862 2585
rect 1262 2513 1862 2551
rect 1262 2479 1762 2513
rect 1796 2479 1862 2513
rect 1262 2441 1862 2479
rect 1262 2407 1762 2441
rect 1796 2407 1862 2441
rect 1262 2369 1862 2407
rect 1262 2335 1762 2369
rect 1796 2335 1862 2369
rect 1262 2297 1862 2335
rect 1262 2263 1762 2297
rect 1796 2263 1862 2297
rect 1262 2225 1862 2263
rect 1262 2191 1762 2225
rect 1796 2191 1862 2225
rect 1262 2153 1862 2191
rect 1262 2119 1762 2153
rect 1796 2119 1862 2153
rect 1262 2081 1862 2119
rect 1262 2047 1762 2081
rect 1796 2047 1862 2081
rect 1262 2009 1862 2047
rect 1262 1975 1762 2009
rect 1796 1975 1862 2009
rect 1262 1937 1862 1975
rect 1262 1903 1762 1937
rect 1796 1903 1862 1937
rect 1262 1865 1862 1903
rect 1262 1831 1762 1865
rect 1796 1831 1862 1865
rect 1262 1793 1862 1831
rect 1262 1759 1762 1793
rect 1796 1759 1862 1793
rect 1262 1721 1862 1759
rect 1262 1687 1762 1721
rect 1796 1687 1862 1721
rect 1262 1649 1862 1687
rect 1262 1615 1762 1649
rect 1796 1615 1862 1649
rect 1262 1577 1862 1615
rect 1262 1543 1762 1577
rect 1796 1543 1862 1577
rect 1262 1505 1862 1543
rect 1262 1471 1762 1505
rect 1796 1471 1862 1505
rect 1262 1433 1862 1471
rect 1262 1399 1762 1433
rect 1796 1399 1862 1433
rect 1262 1361 1862 1399
rect 1262 1327 1762 1361
rect 1796 1327 1862 1361
rect 1262 1289 1862 1327
rect 1262 1255 1762 1289
rect 1796 1255 1862 1289
rect 1262 1217 1862 1255
rect 1262 1183 1762 1217
rect 1796 1183 1862 1217
rect 1262 1145 1862 1183
rect 1262 1111 1762 1145
rect 1796 1111 1862 1145
rect 1262 1073 1862 1111
rect 1262 1039 1762 1073
rect 1796 1039 1862 1073
rect 1262 1001 1862 1039
rect 1262 967 1762 1001
rect 1796 967 1862 1001
rect 1262 929 1862 967
rect 1262 895 1762 929
rect 1796 895 1862 929
rect 1262 857 1862 895
rect 1262 823 1762 857
rect 1796 823 1862 857
rect 1262 785 1862 823
rect 1262 751 1762 785
rect 1796 751 1862 785
rect 1262 713 1862 751
rect 1262 679 1762 713
rect 1796 679 1862 713
rect 1262 641 1862 679
rect 1262 607 1762 641
rect 1796 607 1862 641
rect 1262 569 1862 607
rect 1262 535 1762 569
rect 1796 535 1862 569
rect 1262 497 1862 535
rect 1262 463 1762 497
rect 1796 463 1862 497
rect 1262 425 1862 463
rect 1262 391 1762 425
rect 1796 391 1862 425
rect 1262 353 1862 391
rect 1262 319 1762 353
rect 1796 319 1862 353
rect 1262 281 1862 319
rect 1262 247 1762 281
rect 1796 247 1862 281
rect 1262 209 1862 247
rect 1262 175 1762 209
rect 1796 175 1862 209
rect 1262 137 1862 175
rect 1262 103 1762 137
rect 1796 103 1862 137
rect 1262 65 1862 103
rect 1262 31 1762 65
rect 1796 31 1862 65
rect 1262 -200 1862 31
rect -296 -450 460 -443
rect -296 -502 -289 -450
rect -237 -502 -215 -450
rect -163 -502 -141 -450
rect -89 -502 -67 -450
rect -15 -502 7 -450
rect 59 -502 81 -450
rect 133 -502 155 -450
rect 207 -502 229 -450
rect 281 -502 303 -450
rect 355 -502 377 -450
rect 429 -502 460 -450
rect -296 -524 460 -502
rect -296 -576 -289 -524
rect -237 -576 -215 -524
rect -163 -576 -141 -524
rect -89 -576 -67 -524
rect -15 -576 7 -524
rect 59 -576 81 -524
rect 133 -576 155 -524
rect 207 -576 229 -524
rect 281 -576 303 -524
rect 355 -576 377 -524
rect 429 -576 460 -524
rect -296 -598 460 -576
rect -296 -650 -289 -598
rect -237 -650 -215 -598
rect -163 -650 -141 -598
rect -89 -650 -67 -598
rect -15 -650 7 -598
rect 59 -650 81 -598
rect 133 -650 155 -598
rect 207 -650 229 -598
rect 281 -650 303 -598
rect 355 -650 377 -598
rect 429 -650 460 -598
rect -296 -657 460 -650
<< via1 >>
rect -289 -459 -237 -450
rect -289 -493 -280 -459
rect -280 -493 -246 -459
rect -246 -493 -237 -459
rect -289 -502 -237 -493
rect -215 -459 -163 -450
rect -215 -493 -206 -459
rect -206 -493 -172 -459
rect -172 -493 -163 -459
rect -215 -502 -163 -493
rect -141 -459 -89 -450
rect -141 -493 -132 -459
rect -132 -493 -98 -459
rect -98 -493 -89 -459
rect -141 -502 -89 -493
rect -67 -459 -15 -450
rect -67 -493 -58 -459
rect -58 -493 -24 -459
rect -24 -493 -15 -459
rect -67 -502 -15 -493
rect 7 -459 59 -450
rect 7 -493 16 -459
rect 16 -493 50 -459
rect 50 -493 59 -459
rect 7 -502 59 -493
rect 81 -459 133 -450
rect 81 -493 90 -459
rect 90 -493 124 -459
rect 124 -493 133 -459
rect 81 -502 133 -493
rect 155 -459 207 -450
rect 155 -493 164 -459
rect 164 -493 198 -459
rect 198 -493 207 -459
rect 155 -502 207 -493
rect 229 -459 281 -450
rect 229 -493 238 -459
rect 238 -493 272 -459
rect 272 -493 281 -459
rect 229 -502 281 -493
rect 303 -459 355 -450
rect 303 -493 312 -459
rect 312 -493 346 -459
rect 346 -493 355 -459
rect 303 -502 355 -493
rect 377 -459 429 -450
rect 377 -493 386 -459
rect 386 -493 420 -459
rect 420 -493 429 -459
rect 377 -502 429 -493
rect -289 -533 -237 -524
rect -289 -567 -280 -533
rect -280 -567 -246 -533
rect -246 -567 -237 -533
rect -289 -576 -237 -567
rect -215 -533 -163 -524
rect -215 -567 -206 -533
rect -206 -567 -172 -533
rect -172 -567 -163 -533
rect -215 -576 -163 -567
rect -141 -533 -89 -524
rect -141 -567 -132 -533
rect -132 -567 -98 -533
rect -98 -567 -89 -533
rect -141 -576 -89 -567
rect -67 -533 -15 -524
rect -67 -567 -58 -533
rect -58 -567 -24 -533
rect -24 -567 -15 -533
rect -67 -576 -15 -567
rect 7 -533 59 -524
rect 7 -567 16 -533
rect 16 -567 50 -533
rect 50 -567 59 -533
rect 7 -576 59 -567
rect 81 -533 133 -524
rect 81 -567 90 -533
rect 90 -567 124 -533
rect 124 -567 133 -533
rect 81 -576 133 -567
rect 155 -533 207 -524
rect 155 -567 164 -533
rect 164 -567 198 -533
rect 198 -567 207 -533
rect 155 -576 207 -567
rect 229 -533 281 -524
rect 229 -567 238 -533
rect 238 -567 272 -533
rect 272 -567 281 -533
rect 229 -576 281 -567
rect 303 -533 355 -524
rect 303 -567 312 -533
rect 312 -567 346 -533
rect 346 -567 355 -533
rect 303 -576 355 -567
rect 377 -533 429 -524
rect 377 -567 386 -533
rect 386 -567 420 -533
rect 420 -567 429 -533
rect 377 -576 429 -567
rect -289 -607 -237 -598
rect -289 -641 -280 -607
rect -280 -641 -246 -607
rect -246 -641 -237 -607
rect -289 -650 -237 -641
rect -215 -607 -163 -598
rect -215 -641 -206 -607
rect -206 -641 -172 -607
rect -172 -641 -163 -607
rect -215 -650 -163 -641
rect -141 -607 -89 -598
rect -141 -641 -132 -607
rect -132 -641 -98 -607
rect -98 -641 -89 -607
rect -141 -650 -89 -641
rect -67 -607 -15 -598
rect -67 -641 -58 -607
rect -58 -641 -24 -607
rect -24 -641 -15 -607
rect -67 -650 -15 -641
rect 7 -607 59 -598
rect 7 -641 16 -607
rect 16 -641 50 -607
rect 50 -641 59 -607
rect 7 -650 59 -641
rect 81 -607 133 -598
rect 81 -641 90 -607
rect 90 -641 124 -607
rect 124 -641 133 -607
rect 81 -650 133 -641
rect 155 -607 207 -598
rect 155 -641 164 -607
rect 164 -641 198 -607
rect 198 -641 207 -607
rect 155 -650 207 -641
rect 229 -607 281 -598
rect 229 -641 238 -607
rect 238 -641 272 -607
rect 272 -641 281 -607
rect 229 -650 281 -641
rect 303 -607 355 -598
rect 303 -641 312 -607
rect 312 -641 346 -607
rect 346 -641 355 -607
rect 303 -650 355 -641
rect 377 -607 429 -598
rect 377 -641 386 -607
rect 386 -641 420 -607
rect 420 -641 429 -607
rect 377 -650 429 -641
<< metal2 >>
rect -296 -450 460 -443
rect -296 -502 -289 -450
rect -237 -502 -215 -450
rect -163 -502 -141 -450
rect -89 -502 -67 -450
rect -15 -502 7 -450
rect 59 -502 81 -450
rect 133 -502 155 -450
rect 207 -502 229 -450
rect 281 -502 303 -450
rect 355 -502 377 -450
rect 429 -502 460 -450
rect -296 -524 460 -502
rect -296 -576 -289 -524
rect -237 -576 -215 -524
rect -163 -576 -141 -524
rect -89 -576 -67 -524
rect -15 -576 7 -524
rect 59 -576 81 -524
rect 133 -576 155 -524
rect 207 -576 229 -524
rect 281 -576 303 -524
rect 355 -576 377 -524
rect 429 -576 460 -524
rect -296 -598 460 -576
rect -296 -650 -289 -598
rect -237 -650 -215 -598
rect -163 -650 -141 -598
rect -89 -650 -67 -598
rect -15 -650 7 -598
rect 59 -650 81 -598
rect 133 -650 155 -598
rect 207 -650 229 -598
rect 281 -650 303 -598
rect 355 -650 377 -598
rect 429 -650 460 -598
rect -296 -657 460 -650
<< labels >>
flabel locali s 1835 6920 1990 6982 0 FreeSans 400 0 0 0 PSUB
port 1 nsew
flabel locali s 1779 28 1779 28 0 FreeSans 400 0 0 0 S
port 2 nsew
flabel locali s -1630 31 -1630 31 0 FreeSans 400 0 0 0 S
port 2 nsew
flabel locali s 8 43 142 47 0 FreeSans 400 0 0 0 D
port 3 nsew
flabel comment s 885 159 885 159 0 FreeSans 2000 0 0 0 S
flabel comment s -725 159 -725 159 0 FreeSans 2000 0 0 0 S
flabel comment s 67 159 67 159 0 FreeSans 2000 0 0 0 D
<< properties >>
string GDS_END 5673470
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5581804
<< end >>
