magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1471 203
rect 30 -17 64 21
<< locali >>
rect 103 333 169 493
rect 271 333 337 493
rect 439 333 505 493
rect 607 333 673 493
rect 775 333 841 493
rect 943 333 1009 493
rect 1111 333 1177 493
rect 1279 333 1345 493
rect 103 293 1345 333
rect 102 215 673 259
rect 728 215 824 293
rect 858 215 1261 255
rect 775 181 824 215
rect 1295 181 1345 293
rect 775 131 1345 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 18 299 69 527
rect 203 367 237 527
rect 371 367 405 527
rect 539 367 573 527
rect 707 367 741 527
rect 875 367 909 527
rect 1043 367 1077 527
rect 1211 367 1245 527
rect 1383 299 1454 527
rect 18 147 741 181
rect 18 51 85 147
rect 119 17 153 113
rect 187 51 253 147
rect 287 17 321 113
rect 355 51 421 147
rect 455 17 489 113
rect 523 51 589 147
rect 623 17 657 113
rect 691 97 741 147
rect 1379 97 1454 181
rect 691 51 1454 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel locali s 858 215 1261 255 6 A
port 1 nsew signal input
rlabel locali s 102 215 673 259 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 1472 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 1471 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1510 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 775 131 1345 181 6 Y
port 7 nsew signal output
rlabel locali s 1295 181 1345 293 6 Y
port 7 nsew signal output
rlabel locali s 775 181 824 215 6 Y
port 7 nsew signal output
rlabel locali s 728 215 824 293 6 Y
port 7 nsew signal output
rlabel locali s 103 293 1345 333 6 Y
port 7 nsew signal output
rlabel locali s 1279 333 1345 493 6 Y
port 7 nsew signal output
rlabel locali s 1111 333 1177 493 6 Y
port 7 nsew signal output
rlabel locali s 943 333 1009 493 6 Y
port 7 nsew signal output
rlabel locali s 775 333 841 493 6 Y
port 7 nsew signal output
rlabel locali s 607 333 673 493 6 Y
port 7 nsew signal output
rlabel locali s 439 333 505 493 6 Y
port 7 nsew signal output
rlabel locali s 271 333 337 493 6 Y
port 7 nsew signal output
rlabel locali s 103 333 169 493 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1472 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1729556
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1717264
<< end >>
