magic
tech sky130A
magscale 1 2
timestamp 1666199351
use sky130_fd_pr__dfm1sd2__example_5595914180836  sky130_fd_pr__dfm1sd2__example_5595914180836_0
timestamp 1666199351
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_5595914180835  sky130_fd_pr__hvdfm1sd__example_5595914180835_0
timestamp 1666199351
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_5595914180835  sky130_fd_pr__hvdfm1sd__example_5595914180835_1
timestamp 1666199351
transform 1 0 256 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 28882828
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 28881388
<< end >>
