magic
tech sky130A
magscale 1 2
timestamp 1666199351
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_0
timestamp 1666199351
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_1
timestamp 1666199351
transform 1 0 120 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 35318844
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35317922
<< end >>
