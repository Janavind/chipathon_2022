magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< obsli1 >>
rect 386 1816 424 1850
rect 458 1816 496 1850
rect 530 1816 568 1850
rect 602 1816 640 1850
rect 674 1816 712 1850
rect 746 1816 784 1850
rect 818 1816 856 1850
rect 890 1816 894 1850
rect 196 1663 230 1701
rect 196 1591 230 1629
rect 196 1519 230 1557
rect 196 1447 230 1485
rect 196 1375 230 1413
rect 196 1303 230 1341
rect 196 1231 230 1269
rect 196 1159 230 1197
rect 196 1087 230 1125
rect 196 1015 230 1053
rect 196 943 230 981
rect 196 871 230 909
rect 196 765 230 837
rect 307 741 341 1759
rect 391 741 497 1759
rect 545 741 651 1759
rect 699 741 805 1759
rect 855 741 889 1759
rect 969 1663 1003 1701
rect 969 1591 1003 1629
rect 969 1519 1003 1557
rect 969 1447 1003 1485
rect 969 1375 1003 1413
rect 969 1303 1003 1341
rect 969 1231 1003 1269
rect 969 1159 1003 1197
rect 969 1087 1003 1125
rect 969 1015 1003 1053
rect 969 943 1003 981
rect 969 871 1003 909
rect 969 765 1003 837
rect 386 650 424 684
rect 458 650 496 684
rect 530 650 568 684
rect 602 650 640 684
rect 674 650 712 684
rect 746 650 784 684
rect 818 650 856 684
rect 890 650 894 684
<< obsli1c >>
rect 352 1816 386 1850
rect 424 1816 458 1850
rect 496 1816 530 1850
rect 568 1816 602 1850
rect 640 1816 674 1850
rect 712 1816 746 1850
rect 784 1816 818 1850
rect 856 1816 890 1850
rect 196 1701 230 1735
rect 196 1629 230 1663
rect 196 1557 230 1591
rect 196 1485 230 1519
rect 196 1413 230 1447
rect 196 1341 230 1375
rect 196 1269 230 1303
rect 196 1197 230 1231
rect 196 1125 230 1159
rect 196 1053 230 1087
rect 196 981 230 1015
rect 196 909 230 943
rect 196 837 230 871
rect 969 1701 1003 1735
rect 969 1629 1003 1663
rect 969 1557 1003 1591
rect 969 1485 1003 1519
rect 969 1413 1003 1447
rect 969 1341 1003 1375
rect 969 1269 1003 1303
rect 969 1197 1003 1231
rect 969 1125 1003 1159
rect 969 1053 1003 1087
rect 969 981 1003 1015
rect 969 909 1003 943
rect 969 837 1003 871
rect 352 650 386 684
rect 424 650 458 684
rect 496 650 530 684
rect 568 650 602 684
rect 640 650 674 684
rect 712 650 746 684
rect 784 650 818 684
rect 856 650 890 684
<< metal1 >>
rect 340 1850 902 1862
rect 340 1816 352 1850
rect 386 1816 424 1850
rect 458 1816 496 1850
rect 530 1816 568 1850
rect 602 1816 640 1850
rect 674 1816 712 1850
rect 746 1816 784 1850
rect 818 1816 856 1850
rect 890 1816 902 1850
rect 340 1804 902 1816
rect 184 1735 242 1747
rect 184 1701 196 1735
rect 230 1701 242 1735
rect 184 1663 242 1701
rect 184 1629 196 1663
rect 230 1629 242 1663
rect 184 1591 242 1629
rect 184 1557 196 1591
rect 230 1557 242 1591
rect 184 1519 242 1557
rect 184 1485 196 1519
rect 230 1485 242 1519
rect 184 1447 242 1485
rect 184 1413 196 1447
rect 230 1413 242 1447
rect 184 1375 242 1413
rect 184 1341 196 1375
rect 230 1341 242 1375
rect 184 1303 242 1341
rect 184 1269 196 1303
rect 230 1269 242 1303
rect 184 1231 242 1269
rect 184 1197 196 1231
rect 230 1197 242 1231
rect 184 1159 242 1197
rect 184 1125 196 1159
rect 230 1125 242 1159
rect 184 1087 242 1125
rect 184 1053 196 1087
rect 230 1053 242 1087
rect 184 1015 242 1053
rect 184 981 196 1015
rect 230 981 242 1015
rect 184 943 242 981
rect 184 909 196 943
rect 230 909 242 943
rect 184 871 242 909
rect 184 837 196 871
rect 230 837 242 871
rect 184 753 242 837
rect 957 1735 1015 1747
rect 957 1701 969 1735
rect 1003 1701 1015 1735
rect 957 1663 1015 1701
rect 957 1629 969 1663
rect 1003 1629 1015 1663
rect 957 1591 1015 1629
rect 957 1557 969 1591
rect 1003 1557 1015 1591
rect 957 1519 1015 1557
rect 957 1485 969 1519
rect 1003 1485 1015 1519
rect 957 1447 1015 1485
rect 957 1413 969 1447
rect 1003 1413 1015 1447
rect 957 1375 1015 1413
rect 957 1341 969 1375
rect 1003 1341 1015 1375
rect 957 1303 1015 1341
rect 957 1269 969 1303
rect 1003 1269 1015 1303
rect 957 1231 1015 1269
rect 957 1197 969 1231
rect 1003 1197 1015 1231
rect 957 1159 1015 1197
rect 957 1125 969 1159
rect 1003 1125 1015 1159
rect 957 1087 1015 1125
rect 957 1053 969 1087
rect 1003 1053 1015 1087
rect 957 1015 1015 1053
rect 957 981 969 1015
rect 1003 981 1015 1015
rect 957 943 1015 981
rect 957 909 969 943
rect 1003 909 1015 943
rect 957 871 1015 909
rect 957 837 969 871
rect 1003 837 1015 871
rect 957 753 1015 837
rect 340 684 902 696
rect 340 650 352 684
rect 386 650 424 684
rect 458 650 496 684
rect 530 650 568 684
rect 602 650 640 684
rect 674 650 712 684
rect 746 650 784 684
rect 818 650 856 684
rect 890 650 902 684
rect 340 638 902 650
<< obsm1 >>
rect 298 1747 350 1776
rect 540 1747 656 1776
rect 846 1747 898 1776
rect 298 753 353 1747
rect 381 753 507 1747
rect 535 753 661 1747
rect 689 753 815 1747
rect 843 753 901 1747
rect 298 724 350 753
rect 540 724 656 753
rect 846 724 898 753
<< obsm2 >>
rect 158 1626 1042 2428
rect 158 1456 350 1626
rect 158 1044 214 1456
rect 386 1428 502 1570
rect 540 1456 656 1626
rect 694 1428 810 1570
rect 846 1456 1042 1626
rect 386 1072 810 1428
rect 158 874 350 1044
rect 386 930 502 1072
rect 540 874 656 1044
rect 694 930 810 1072
rect 986 1044 1042 1456
rect 846 874 1042 1044
rect 158 72 1042 874
<< metal3 >>
rect 0 2000 1200 2500
rect 0 1000 1200 1500
rect 0 0 1200 500
<< labels >>
rlabel metal1 s 957 753 1015 1747 6 BULK
port 1 nsew
rlabel metal1 s 184 753 242 1747 6 BULK
port 1 nsew
rlabel metal3 s 0 1000 1200 1500 6 DRAIN
port 2 nsew
rlabel metal1 s 340 1804 902 1862 6 GATE
port 3 nsew
rlabel metal1 s 340 638 902 696 6 GATE
port 3 nsew
rlabel metal3 s 0 2000 1200 2500 6 SOURCE
port 4 nsew
rlabel metal3 s 0 0 1200 500 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1200 2500
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9881838
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9849760
<< end >>
