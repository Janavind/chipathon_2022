magic
tech sky130A
magscale 1 2
timestamp 1666199351
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1666199351
transform 1 0 -50 0 1 8
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1666199351
transform 1 0 -46 0 1 -1242
box 0 0 1 1
<< properties >>
string GDS_END 32655954
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 32654146
<< end >>
