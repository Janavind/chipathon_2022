magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< poly >>
rect 1671 435 1701 648
rect 2295 559 2325 648
rect 2277 543 2343 559
rect 2277 509 2293 543
rect 2327 509 2343 543
rect 2277 493 2343 509
rect 2919 435 2949 648
rect 3543 559 3573 648
rect 3525 543 3591 559
rect 3525 509 3541 543
rect 3575 509 3591 543
rect 3525 493 3591 509
rect 4167 435 4197 648
rect 4791 559 4821 648
rect 4773 543 4839 559
rect 4773 509 4789 543
rect 4823 509 4839 543
rect 4773 493 4839 509
rect 5415 435 5445 648
rect 6039 559 6069 648
rect 6021 543 6087 559
rect 6021 509 6037 543
rect 6071 509 6087 543
rect 6021 493 6087 509
rect 6663 435 6693 648
rect 7287 559 7317 648
rect 7269 543 7335 559
rect 7269 509 7285 543
rect 7319 509 7335 543
rect 7269 493 7335 509
rect 7911 435 7941 648
rect 8535 559 8565 648
rect 8517 543 8583 559
rect 8517 509 8533 543
rect 8567 509 8583 543
rect 8517 493 8583 509
rect 9159 435 9189 648
rect 9783 559 9813 648
rect 9765 543 9831 559
rect 9765 509 9781 543
rect 9815 509 9831 543
rect 9765 493 9831 509
rect 10407 435 10437 648
rect 11031 559 11061 648
rect 11013 543 11079 559
rect 11013 509 11029 543
rect 11063 509 11079 543
rect 11013 493 11079 509
rect 11655 435 11685 648
rect 12279 559 12309 648
rect 12261 543 12327 559
rect 12261 509 12277 543
rect 12311 509 12327 543
rect 12261 493 12327 509
rect 12903 435 12933 648
rect 13527 559 13557 648
rect 13509 543 13575 559
rect 13509 509 13525 543
rect 13559 509 13575 543
rect 13509 493 13575 509
rect 14151 435 14181 648
rect 14775 559 14805 648
rect 14757 543 14823 559
rect 14757 509 14773 543
rect 14807 509 14823 543
rect 14757 493 14823 509
rect 15399 435 15429 648
rect 16023 559 16053 648
rect 16005 543 16071 559
rect 16005 509 16021 543
rect 16055 509 16071 543
rect 16005 493 16071 509
rect 16647 435 16677 648
rect 17271 559 17301 648
rect 17253 543 17319 559
rect 17253 509 17269 543
rect 17303 509 17319 543
rect 17253 493 17319 509
rect 17895 435 17925 648
rect 18519 559 18549 648
rect 18501 543 18567 559
rect 18501 509 18517 543
rect 18551 509 18567 543
rect 18501 493 18567 509
rect 19143 435 19173 648
rect 19767 559 19797 648
rect 19749 543 19815 559
rect 19749 509 19765 543
rect 19799 509 19815 543
rect 19749 493 19815 509
rect 20391 435 20421 648
rect 21015 559 21045 648
rect 20997 543 21063 559
rect 20997 509 21013 543
rect 21047 509 21063 543
rect 20997 493 21063 509
rect 21639 435 21669 648
rect 22263 559 22293 648
rect 22245 543 22311 559
rect 22245 509 22261 543
rect 22295 509 22311 543
rect 22245 493 22311 509
rect 22887 435 22917 648
rect 23511 559 23541 648
rect 23493 543 23559 559
rect 23493 509 23509 543
rect 23543 509 23559 543
rect 23493 493 23559 509
rect 24135 435 24165 648
rect 24759 559 24789 648
rect 24741 543 24807 559
rect 24741 509 24757 543
rect 24791 509 24807 543
rect 24741 493 24807 509
rect 25383 435 25413 648
rect 26007 559 26037 648
rect 25989 543 26055 559
rect 25989 509 26005 543
rect 26039 509 26055 543
rect 25989 493 26055 509
rect 26631 435 26661 648
rect 27255 559 27285 648
rect 27237 543 27303 559
rect 27237 509 27253 543
rect 27287 509 27303 543
rect 27237 493 27303 509
rect 27879 435 27909 648
rect 28503 559 28533 648
rect 28485 543 28551 559
rect 28485 509 28501 543
rect 28535 509 28551 543
rect 28485 493 28551 509
rect 29127 435 29157 648
rect 29751 559 29781 648
rect 29733 543 29799 559
rect 29733 509 29749 543
rect 29783 509 29799 543
rect 29733 493 29799 509
rect 30375 435 30405 648
rect 30999 559 31029 648
rect 30981 543 31047 559
rect 30981 509 30997 543
rect 31031 509 31047 543
rect 30981 493 31047 509
rect 31623 435 31653 648
rect 32247 559 32277 648
rect 32229 543 32295 559
rect 32229 509 32245 543
rect 32279 509 32295 543
rect 32229 493 32295 509
rect 32871 435 32901 648
rect 33495 559 33525 648
rect 33477 543 33543 559
rect 33477 509 33493 543
rect 33527 509 33543 543
rect 33477 493 33543 509
rect 34119 435 34149 648
rect 34743 559 34773 648
rect 34725 543 34791 559
rect 34725 509 34741 543
rect 34775 509 34791 543
rect 34725 493 34791 509
rect 35367 435 35397 648
rect 35991 559 36021 648
rect 35973 543 36039 559
rect 35973 509 35989 543
rect 36023 509 36039 543
rect 35973 493 36039 509
rect 36615 435 36645 648
rect 37239 559 37269 648
rect 37221 543 37287 559
rect 37221 509 37237 543
rect 37271 509 37287 543
rect 37221 493 37287 509
rect 37863 435 37893 648
rect 38487 559 38517 648
rect 38469 543 38535 559
rect 38469 509 38485 543
rect 38519 509 38535 543
rect 38469 493 38535 509
rect 39111 435 39141 648
rect 39735 559 39765 648
rect 39717 543 39783 559
rect 39717 509 39733 543
rect 39767 509 39783 543
rect 39717 493 39783 509
rect 40359 435 40389 648
rect 40983 559 41013 648
rect 40965 543 41031 559
rect 40965 509 40981 543
rect 41015 509 41031 543
rect 40965 493 41031 509
rect 1653 419 1719 435
rect 1653 385 1669 419
rect 1703 385 1719 419
rect 1653 369 1719 385
rect 2901 419 2967 435
rect 2901 385 2917 419
rect 2951 385 2967 419
rect 2901 369 2967 385
rect 4149 419 4215 435
rect 4149 385 4165 419
rect 4199 385 4215 419
rect 4149 369 4215 385
rect 5397 419 5463 435
rect 5397 385 5413 419
rect 5447 385 5463 419
rect 5397 369 5463 385
rect 6645 419 6711 435
rect 6645 385 6661 419
rect 6695 385 6711 419
rect 6645 369 6711 385
rect 7893 419 7959 435
rect 7893 385 7909 419
rect 7943 385 7959 419
rect 7893 369 7959 385
rect 9141 419 9207 435
rect 9141 385 9157 419
rect 9191 385 9207 419
rect 9141 369 9207 385
rect 10389 419 10455 435
rect 10389 385 10405 419
rect 10439 385 10455 419
rect 10389 369 10455 385
rect 11637 419 11703 435
rect 11637 385 11653 419
rect 11687 385 11703 419
rect 11637 369 11703 385
rect 12885 419 12951 435
rect 12885 385 12901 419
rect 12935 385 12951 419
rect 12885 369 12951 385
rect 14133 419 14199 435
rect 14133 385 14149 419
rect 14183 385 14199 419
rect 14133 369 14199 385
rect 15381 419 15447 435
rect 15381 385 15397 419
rect 15431 385 15447 419
rect 15381 369 15447 385
rect 16629 419 16695 435
rect 16629 385 16645 419
rect 16679 385 16695 419
rect 16629 369 16695 385
rect 17877 419 17943 435
rect 17877 385 17893 419
rect 17927 385 17943 419
rect 17877 369 17943 385
rect 19125 419 19191 435
rect 19125 385 19141 419
rect 19175 385 19191 419
rect 19125 369 19191 385
rect 20373 419 20439 435
rect 20373 385 20389 419
rect 20423 385 20439 419
rect 20373 369 20439 385
rect 21621 419 21687 435
rect 21621 385 21637 419
rect 21671 385 21687 419
rect 21621 369 21687 385
rect 22869 419 22935 435
rect 22869 385 22885 419
rect 22919 385 22935 419
rect 22869 369 22935 385
rect 24117 419 24183 435
rect 24117 385 24133 419
rect 24167 385 24183 419
rect 24117 369 24183 385
rect 25365 419 25431 435
rect 25365 385 25381 419
rect 25415 385 25431 419
rect 25365 369 25431 385
rect 26613 419 26679 435
rect 26613 385 26629 419
rect 26663 385 26679 419
rect 26613 369 26679 385
rect 27861 419 27927 435
rect 27861 385 27877 419
rect 27911 385 27927 419
rect 27861 369 27927 385
rect 29109 419 29175 435
rect 29109 385 29125 419
rect 29159 385 29175 419
rect 29109 369 29175 385
rect 30357 419 30423 435
rect 30357 385 30373 419
rect 30407 385 30423 419
rect 30357 369 30423 385
rect 31605 419 31671 435
rect 31605 385 31621 419
rect 31655 385 31671 419
rect 31605 369 31671 385
rect 32853 419 32919 435
rect 32853 385 32869 419
rect 32903 385 32919 419
rect 32853 369 32919 385
rect 34101 419 34167 435
rect 34101 385 34117 419
rect 34151 385 34167 419
rect 34101 369 34167 385
rect 35349 419 35415 435
rect 35349 385 35365 419
rect 35399 385 35415 419
rect 35349 369 35415 385
rect 36597 419 36663 435
rect 36597 385 36613 419
rect 36647 385 36663 419
rect 36597 369 36663 385
rect 37845 419 37911 435
rect 37845 385 37861 419
rect 37895 385 37911 419
rect 37845 369 37911 385
rect 39093 419 39159 435
rect 39093 385 39109 419
rect 39143 385 39159 419
rect 39093 369 39159 385
rect 40341 419 40407 435
rect 40341 385 40357 419
rect 40391 385 40407 419
rect 40341 369 40407 385
<< polycont >>
rect 2293 509 2327 543
rect 3541 509 3575 543
rect 4789 509 4823 543
rect 6037 509 6071 543
rect 7285 509 7319 543
rect 8533 509 8567 543
rect 9781 509 9815 543
rect 11029 509 11063 543
rect 12277 509 12311 543
rect 13525 509 13559 543
rect 14773 509 14807 543
rect 16021 509 16055 543
rect 17269 509 17303 543
rect 18517 509 18551 543
rect 19765 509 19799 543
rect 21013 509 21047 543
rect 22261 509 22295 543
rect 23509 509 23543 543
rect 24757 509 24791 543
rect 26005 509 26039 543
rect 27253 509 27287 543
rect 28501 509 28535 543
rect 29749 509 29783 543
rect 30997 509 31031 543
rect 32245 509 32279 543
rect 33493 509 33527 543
rect 34741 509 34775 543
rect 35989 509 36023 543
rect 37237 509 37271 543
rect 38485 509 38519 543
rect 39733 509 39767 543
rect 40981 509 41015 543
rect 1669 385 1703 419
rect 2917 385 2951 419
rect 4165 385 4199 419
rect 5413 385 5447 419
rect 6661 385 6695 419
rect 7909 385 7943 419
rect 9157 385 9191 419
rect 10405 385 10439 419
rect 11653 385 11687 419
rect 12901 385 12935 419
rect 14149 385 14183 419
rect 15397 385 15431 419
rect 16645 385 16679 419
rect 17893 385 17927 419
rect 19141 385 19175 419
rect 20389 385 20423 419
rect 21637 385 21671 419
rect 22885 385 22919 419
rect 24133 385 24167 419
rect 25381 385 25415 419
rect 26629 385 26663 419
rect 27877 385 27911 419
rect 29125 385 29159 419
rect 30373 385 30407 419
rect 31621 385 31655 419
rect 32869 385 32903 419
rect 34117 385 34151 419
rect 35365 385 35399 419
rect 36613 385 36647 419
rect 37861 385 37895 419
rect 39109 385 39143 419
rect 40357 385 40391 419
<< locali >>
rect 2293 543 2327 559
rect 2293 493 2327 509
rect 3541 543 3575 559
rect 3541 493 3575 509
rect 4789 543 4823 559
rect 4789 493 4823 509
rect 6037 543 6071 559
rect 6037 493 6071 509
rect 7285 543 7319 559
rect 7285 493 7319 509
rect 8533 543 8567 559
rect 8533 493 8567 509
rect 9781 543 9815 559
rect 9781 493 9815 509
rect 11029 543 11063 559
rect 11029 493 11063 509
rect 12277 543 12311 559
rect 12277 493 12311 509
rect 13525 543 13559 559
rect 13525 493 13559 509
rect 14773 543 14807 559
rect 14773 493 14807 509
rect 16021 543 16055 559
rect 16021 493 16055 509
rect 17269 543 17303 559
rect 17269 493 17303 509
rect 18517 543 18551 559
rect 18517 493 18551 509
rect 19765 543 19799 559
rect 19765 493 19799 509
rect 21013 543 21047 559
rect 21013 493 21047 509
rect 22261 543 22295 559
rect 22261 493 22295 509
rect 23509 543 23543 559
rect 23509 493 23543 509
rect 24757 543 24791 559
rect 24757 493 24791 509
rect 26005 543 26039 559
rect 26005 493 26039 509
rect 27253 543 27287 559
rect 27253 493 27287 509
rect 28501 543 28535 559
rect 28501 493 28535 509
rect 29749 543 29783 559
rect 29749 493 29783 509
rect 30997 543 31031 559
rect 30997 493 31031 509
rect 32245 543 32279 559
rect 32245 493 32279 509
rect 33493 543 33527 559
rect 33493 493 33527 509
rect 34741 543 34775 559
rect 34741 493 34775 509
rect 35989 543 36023 559
rect 35989 493 36023 509
rect 37237 543 37271 559
rect 37237 493 37271 509
rect 38485 543 38519 559
rect 38485 493 38519 509
rect 39733 543 39767 559
rect 39733 493 39767 509
rect 40981 543 41015 559
rect 40981 493 41015 509
rect 1669 419 1703 435
rect 1669 369 1703 385
rect 2917 419 2951 435
rect 2917 369 2951 385
rect 4165 419 4199 435
rect 4165 369 4199 385
rect 5413 419 5447 435
rect 5413 369 5447 385
rect 6661 419 6695 435
rect 6661 369 6695 385
rect 7909 419 7943 435
rect 7909 369 7943 385
rect 9157 419 9191 435
rect 9157 369 9191 385
rect 10405 419 10439 435
rect 10405 369 10439 385
rect 11653 419 11687 435
rect 11653 369 11687 385
rect 12901 419 12935 435
rect 12901 369 12935 385
rect 14149 419 14183 435
rect 14149 369 14183 385
rect 15397 419 15431 435
rect 15397 369 15431 385
rect 16645 419 16679 435
rect 16645 369 16679 385
rect 17893 419 17927 435
rect 17893 369 17927 385
rect 19141 419 19175 435
rect 19141 369 19175 385
rect 20389 419 20423 435
rect 20389 369 20423 385
rect 21637 419 21671 435
rect 21637 369 21671 385
rect 22885 419 22919 435
rect 22885 369 22919 385
rect 24133 419 24167 435
rect 24133 369 24167 385
rect 25381 419 25415 435
rect 25381 369 25415 385
rect 26629 419 26663 435
rect 26629 369 26663 385
rect 27877 419 27911 435
rect 27877 369 27911 385
rect 29125 419 29159 435
rect 29125 369 29159 385
rect 30373 419 30407 435
rect 30373 369 30407 385
rect 31621 419 31655 435
rect 31621 369 31655 385
rect 32869 419 32903 435
rect 32869 369 32903 385
rect 34117 419 34151 435
rect 34117 369 34151 385
rect 35365 419 35399 435
rect 35365 369 35399 385
rect 36613 419 36647 435
rect 36613 369 36647 385
rect 37861 419 37895 435
rect 37861 369 37895 385
rect 39109 419 39143 435
rect 39109 369 39143 385
rect 40357 419 40391 435
rect 40357 369 40391 385
<< viali >>
rect 2293 509 2327 543
rect 3541 509 3575 543
rect 4789 509 4823 543
rect 6037 509 6071 543
rect 7285 509 7319 543
rect 8533 509 8567 543
rect 9781 509 9815 543
rect 11029 509 11063 543
rect 12277 509 12311 543
rect 13525 509 13559 543
rect 14773 509 14807 543
rect 16021 509 16055 543
rect 17269 509 17303 543
rect 18517 509 18551 543
rect 19765 509 19799 543
rect 21013 509 21047 543
rect 22261 509 22295 543
rect 23509 509 23543 543
rect 24757 509 24791 543
rect 26005 509 26039 543
rect 27253 509 27287 543
rect 28501 509 28535 543
rect 29749 509 29783 543
rect 30997 509 31031 543
rect 32245 509 32279 543
rect 33493 509 33527 543
rect 34741 509 34775 543
rect 35989 509 36023 543
rect 37237 509 37271 543
rect 38485 509 38519 543
rect 39733 509 39767 543
rect 40981 509 41015 543
rect 1669 385 1703 419
rect 2917 385 2951 419
rect 4165 385 4199 419
rect 5413 385 5447 419
rect 6661 385 6695 419
rect 7909 385 7943 419
rect 9157 385 9191 419
rect 10405 385 10439 419
rect 11653 385 11687 419
rect 12901 385 12935 419
rect 14149 385 14183 419
rect 15397 385 15431 419
rect 16645 385 16679 419
rect 17893 385 17927 419
rect 19141 385 19175 419
rect 20389 385 20423 419
rect 21637 385 21671 419
rect 22885 385 22919 419
rect 24133 385 24167 419
rect 25381 385 25415 419
rect 26629 385 26663 419
rect 27877 385 27911 419
rect 29125 385 29159 419
rect 30373 385 30407 419
rect 31621 385 31655 419
rect 32869 385 32903 419
rect 34117 385 34151 419
rect 35365 385 35399 419
rect 36613 385 36647 419
rect 37861 385 37895 419
rect 39109 385 39143 419
rect 40357 385 40391 419
<< metal1 >>
rect 1454 1880 1482 1936
rect 1918 1880 1946 1936
rect 2050 1880 2078 1936
rect 2514 1880 2542 1936
rect 2702 1880 2730 1936
rect 3166 1880 3194 1936
rect 3298 1880 3326 1936
rect 3762 1880 3790 1936
rect 3950 1880 3978 1936
rect 4414 1880 4442 1936
rect 4546 1880 4574 1936
rect 5010 1880 5038 1936
rect 5198 1880 5226 1936
rect 5662 1880 5690 1936
rect 5794 1880 5822 1936
rect 6258 1880 6286 1936
rect 6446 1880 6474 1936
rect 6910 1880 6938 1936
rect 7042 1880 7070 1936
rect 7506 1880 7534 1936
rect 7694 1880 7722 1936
rect 8158 1880 8186 1936
rect 8290 1880 8318 1936
rect 8754 1880 8782 1936
rect 8942 1880 8970 1936
rect 9406 1880 9434 1936
rect 9538 1880 9566 1936
rect 10002 1880 10030 1936
rect 10190 1880 10218 1936
rect 10654 1880 10682 1936
rect 10786 1880 10814 1936
rect 11250 1880 11278 1936
rect 11438 1880 11466 1936
rect 11902 1880 11930 1936
rect 12034 1880 12062 1936
rect 12498 1880 12526 1936
rect 12686 1880 12714 1936
rect 13150 1880 13178 1936
rect 13282 1880 13310 1936
rect 13746 1880 13774 1936
rect 13934 1880 13962 1936
rect 14398 1880 14426 1936
rect 14530 1880 14558 1936
rect 14994 1880 15022 1936
rect 15182 1880 15210 1936
rect 15646 1880 15674 1936
rect 15778 1880 15806 1936
rect 16242 1880 16270 1936
rect 16430 1880 16458 1936
rect 16894 1880 16922 1936
rect 17026 1880 17054 1936
rect 17490 1880 17518 1936
rect 17678 1880 17706 1936
rect 18142 1880 18170 1936
rect 18274 1880 18302 1936
rect 18738 1880 18766 1936
rect 18926 1880 18954 1936
rect 19390 1880 19418 1936
rect 19522 1880 19550 1936
rect 19986 1880 20014 1936
rect 20174 1880 20202 1936
rect 20638 1880 20666 1936
rect 20770 1880 20798 1936
rect 21234 1880 21262 1936
rect 21422 1880 21450 1936
rect 21886 1880 21914 1936
rect 22018 1880 22046 1936
rect 22482 1880 22510 1936
rect 22670 1880 22698 1936
rect 23134 1880 23162 1936
rect 23266 1880 23294 1936
rect 23730 1880 23758 1936
rect 23918 1880 23946 1936
rect 24382 1880 24410 1936
rect 24514 1880 24542 1936
rect 24978 1880 25006 1936
rect 25166 1880 25194 1936
rect 25630 1880 25658 1936
rect 25762 1880 25790 1936
rect 26226 1880 26254 1936
rect 26414 1880 26442 1936
rect 26878 1880 26906 1936
rect 27010 1880 27038 1936
rect 27474 1880 27502 1936
rect 27662 1880 27690 1936
rect 28126 1880 28154 1936
rect 28258 1880 28286 1936
rect 28722 1880 28750 1936
rect 28910 1880 28938 1936
rect 29374 1880 29402 1936
rect 29506 1880 29534 1936
rect 29970 1880 29998 1936
rect 30158 1880 30186 1936
rect 30622 1880 30650 1936
rect 30754 1880 30782 1936
rect 31218 1880 31246 1936
rect 31406 1880 31434 1936
rect 31870 1880 31898 1936
rect 32002 1880 32030 1936
rect 32466 1880 32494 1936
rect 32654 1880 32682 1936
rect 33118 1880 33146 1936
rect 33250 1880 33278 1936
rect 33714 1880 33742 1936
rect 33902 1880 33930 1936
rect 34366 1880 34394 1936
rect 34498 1880 34526 1936
rect 34962 1880 34990 1936
rect 35150 1880 35178 1936
rect 35614 1880 35642 1936
rect 35746 1880 35774 1936
rect 36210 1880 36238 1936
rect 36398 1880 36426 1936
rect 36862 1880 36890 1936
rect 36994 1880 37022 1936
rect 37458 1880 37486 1936
rect 37646 1880 37674 1936
rect 38110 1880 38138 1936
rect 38242 1880 38270 1936
rect 38706 1880 38734 1936
rect 38894 1880 38922 1936
rect 39358 1880 39386 1936
rect 39490 1880 39518 1936
rect 39954 1880 39982 1936
rect 40142 1880 40170 1936
rect 40606 1880 40634 1936
rect 40738 1880 40766 1936
rect 41202 1880 41230 1936
rect 1454 274 1482 620
rect 1654 376 1660 428
rect 1712 376 1718 428
rect 1436 222 1442 274
rect 1494 222 1500 274
rect 1918 150 1946 620
rect 2050 150 2078 620
rect 2278 500 2284 552
rect 2336 500 2342 552
rect 2514 274 2542 620
rect 2702 274 2730 620
rect 2902 376 2908 428
rect 2960 376 2966 428
rect 2496 222 2502 274
rect 2554 222 2560 274
rect 2684 222 2690 274
rect 2742 222 2748 274
rect 3166 150 3194 620
rect 3298 150 3326 620
rect 3526 500 3532 552
rect 3584 500 3590 552
rect 3762 274 3790 620
rect 3950 274 3978 620
rect 4150 376 4156 428
rect 4208 376 4214 428
rect 3744 222 3750 274
rect 3802 222 3808 274
rect 3932 222 3938 274
rect 3990 222 3996 274
rect 4414 150 4442 620
rect 4546 150 4574 620
rect 4774 500 4780 552
rect 4832 500 4838 552
rect 5010 274 5038 620
rect 5198 274 5226 620
rect 5398 376 5404 428
rect 5456 376 5462 428
rect 4992 222 4998 274
rect 5050 222 5056 274
rect 5180 222 5186 274
rect 5238 222 5244 274
rect 5662 150 5690 620
rect 5794 150 5822 620
rect 6022 500 6028 552
rect 6080 500 6086 552
rect 6258 274 6286 620
rect 6446 274 6474 620
rect 6646 376 6652 428
rect 6704 376 6710 428
rect 6240 222 6246 274
rect 6298 222 6304 274
rect 6428 222 6434 274
rect 6486 222 6492 274
rect 6910 150 6938 620
rect 7042 150 7070 620
rect 7270 500 7276 552
rect 7328 500 7334 552
rect 7506 274 7534 620
rect 7694 274 7722 620
rect 7894 376 7900 428
rect 7952 376 7958 428
rect 7488 222 7494 274
rect 7546 222 7552 274
rect 7676 222 7682 274
rect 7734 222 7740 274
rect 8158 150 8186 620
rect 8290 150 8318 620
rect 8518 500 8524 552
rect 8576 500 8582 552
rect 8754 274 8782 620
rect 8942 274 8970 620
rect 9142 376 9148 428
rect 9200 376 9206 428
rect 8736 222 8742 274
rect 8794 222 8800 274
rect 8924 222 8930 274
rect 8982 222 8988 274
rect 9406 150 9434 620
rect 9538 150 9566 620
rect 9766 500 9772 552
rect 9824 500 9830 552
rect 10002 274 10030 620
rect 10190 274 10218 620
rect 10390 376 10396 428
rect 10448 376 10454 428
rect 9984 222 9990 274
rect 10042 222 10048 274
rect 10172 222 10178 274
rect 10230 222 10236 274
rect 10654 150 10682 620
rect 10786 150 10814 620
rect 11014 500 11020 552
rect 11072 500 11078 552
rect 11250 274 11278 620
rect 11438 274 11466 620
rect 11638 376 11644 428
rect 11696 376 11702 428
rect 11232 222 11238 274
rect 11290 222 11296 274
rect 11420 222 11426 274
rect 11478 222 11484 274
rect 11902 150 11930 620
rect 12034 150 12062 620
rect 12262 500 12268 552
rect 12320 500 12326 552
rect 12498 274 12526 620
rect 12686 274 12714 620
rect 12886 376 12892 428
rect 12944 376 12950 428
rect 12480 222 12486 274
rect 12538 222 12544 274
rect 12668 222 12674 274
rect 12726 222 12732 274
rect 13150 150 13178 620
rect 13282 150 13310 620
rect 13510 500 13516 552
rect 13568 500 13574 552
rect 13746 274 13774 620
rect 13934 274 13962 620
rect 14134 376 14140 428
rect 14192 376 14198 428
rect 13728 222 13734 274
rect 13786 222 13792 274
rect 13916 222 13922 274
rect 13974 222 13980 274
rect 14398 150 14426 620
rect 14530 150 14558 620
rect 14758 500 14764 552
rect 14816 500 14822 552
rect 14994 274 15022 620
rect 15182 274 15210 620
rect 15382 376 15388 428
rect 15440 376 15446 428
rect 14976 222 14982 274
rect 15034 222 15040 274
rect 15164 222 15170 274
rect 15222 222 15228 274
rect 15646 150 15674 620
rect 15778 150 15806 620
rect 16006 500 16012 552
rect 16064 500 16070 552
rect 16242 274 16270 620
rect 16430 274 16458 620
rect 16630 376 16636 428
rect 16688 376 16694 428
rect 16224 222 16230 274
rect 16282 222 16288 274
rect 16412 222 16418 274
rect 16470 222 16476 274
rect 16894 150 16922 620
rect 17026 150 17054 620
rect 17254 500 17260 552
rect 17312 500 17318 552
rect 17490 274 17518 620
rect 17678 274 17706 620
rect 17878 376 17884 428
rect 17936 376 17942 428
rect 17472 222 17478 274
rect 17530 222 17536 274
rect 17660 222 17666 274
rect 17718 222 17724 274
rect 18142 150 18170 620
rect 18274 150 18302 620
rect 18502 500 18508 552
rect 18560 500 18566 552
rect 18738 274 18766 620
rect 18926 274 18954 620
rect 19126 376 19132 428
rect 19184 376 19190 428
rect 18720 222 18726 274
rect 18778 222 18784 274
rect 18908 222 18914 274
rect 18966 222 18972 274
rect 19390 150 19418 620
rect 19522 150 19550 620
rect 19750 500 19756 552
rect 19808 500 19814 552
rect 19986 274 20014 620
rect 20174 274 20202 620
rect 20374 376 20380 428
rect 20432 376 20438 428
rect 19968 222 19974 274
rect 20026 222 20032 274
rect 20156 222 20162 274
rect 20214 222 20220 274
rect 20638 150 20666 620
rect 20770 150 20798 620
rect 20998 500 21004 552
rect 21056 500 21062 552
rect 21234 274 21262 620
rect 21422 274 21450 620
rect 21622 376 21628 428
rect 21680 376 21686 428
rect 21216 222 21222 274
rect 21274 222 21280 274
rect 21404 222 21410 274
rect 21462 222 21468 274
rect 21886 150 21914 620
rect 22018 150 22046 620
rect 22246 500 22252 552
rect 22304 500 22310 552
rect 22482 274 22510 620
rect 22670 274 22698 620
rect 22870 376 22876 428
rect 22928 376 22934 428
rect 22464 222 22470 274
rect 22522 222 22528 274
rect 22652 222 22658 274
rect 22710 222 22716 274
rect 23134 150 23162 620
rect 23266 150 23294 620
rect 23494 500 23500 552
rect 23552 500 23558 552
rect 23730 274 23758 620
rect 23918 274 23946 620
rect 24118 376 24124 428
rect 24176 376 24182 428
rect 23712 222 23718 274
rect 23770 222 23776 274
rect 23900 222 23906 274
rect 23958 222 23964 274
rect 24382 150 24410 620
rect 24514 150 24542 620
rect 24742 500 24748 552
rect 24800 500 24806 552
rect 24978 274 25006 620
rect 25166 274 25194 620
rect 25366 376 25372 428
rect 25424 376 25430 428
rect 24960 222 24966 274
rect 25018 222 25024 274
rect 25148 222 25154 274
rect 25206 222 25212 274
rect 25630 150 25658 620
rect 25762 150 25790 620
rect 25990 500 25996 552
rect 26048 500 26054 552
rect 26226 274 26254 620
rect 26414 274 26442 620
rect 26614 376 26620 428
rect 26672 376 26678 428
rect 26208 222 26214 274
rect 26266 222 26272 274
rect 26396 222 26402 274
rect 26454 222 26460 274
rect 26878 150 26906 620
rect 27010 150 27038 620
rect 27238 500 27244 552
rect 27296 500 27302 552
rect 27474 274 27502 620
rect 27662 274 27690 620
rect 27862 376 27868 428
rect 27920 376 27926 428
rect 27456 222 27462 274
rect 27514 222 27520 274
rect 27644 222 27650 274
rect 27702 222 27708 274
rect 28126 150 28154 620
rect 28258 150 28286 620
rect 28486 500 28492 552
rect 28544 500 28550 552
rect 28722 274 28750 620
rect 28910 274 28938 620
rect 29110 376 29116 428
rect 29168 376 29174 428
rect 28704 222 28710 274
rect 28762 222 28768 274
rect 28892 222 28898 274
rect 28950 222 28956 274
rect 29374 150 29402 620
rect 29506 150 29534 620
rect 29734 500 29740 552
rect 29792 500 29798 552
rect 29970 274 29998 620
rect 30158 274 30186 620
rect 30358 376 30364 428
rect 30416 376 30422 428
rect 29952 222 29958 274
rect 30010 222 30016 274
rect 30140 222 30146 274
rect 30198 222 30204 274
rect 30622 150 30650 620
rect 30754 150 30782 620
rect 30982 500 30988 552
rect 31040 500 31046 552
rect 31218 274 31246 620
rect 31406 274 31434 620
rect 31606 376 31612 428
rect 31664 376 31670 428
rect 31200 222 31206 274
rect 31258 222 31264 274
rect 31388 222 31394 274
rect 31446 222 31452 274
rect 31870 150 31898 620
rect 32002 150 32030 620
rect 32230 500 32236 552
rect 32288 500 32294 552
rect 32466 274 32494 620
rect 32654 274 32682 620
rect 32854 376 32860 428
rect 32912 376 32918 428
rect 32448 222 32454 274
rect 32506 222 32512 274
rect 32636 222 32642 274
rect 32694 222 32700 274
rect 33118 150 33146 620
rect 33250 150 33278 620
rect 33478 500 33484 552
rect 33536 500 33542 552
rect 33714 274 33742 620
rect 33902 274 33930 620
rect 34102 376 34108 428
rect 34160 376 34166 428
rect 33696 222 33702 274
rect 33754 222 33760 274
rect 33884 222 33890 274
rect 33942 222 33948 274
rect 34366 150 34394 620
rect 34498 150 34526 620
rect 34726 500 34732 552
rect 34784 500 34790 552
rect 34962 274 34990 620
rect 35150 274 35178 620
rect 35350 376 35356 428
rect 35408 376 35414 428
rect 34944 222 34950 274
rect 35002 222 35008 274
rect 35132 222 35138 274
rect 35190 222 35196 274
rect 35614 150 35642 620
rect 35746 150 35774 620
rect 35974 500 35980 552
rect 36032 500 36038 552
rect 36210 274 36238 620
rect 36398 274 36426 620
rect 36598 376 36604 428
rect 36656 376 36662 428
rect 36192 222 36198 274
rect 36250 222 36256 274
rect 36380 222 36386 274
rect 36438 222 36444 274
rect 36862 150 36890 620
rect 36994 150 37022 620
rect 37222 500 37228 552
rect 37280 500 37286 552
rect 37458 274 37486 620
rect 37646 274 37674 620
rect 37846 376 37852 428
rect 37904 376 37910 428
rect 37440 222 37446 274
rect 37498 222 37504 274
rect 37628 222 37634 274
rect 37686 222 37692 274
rect 38110 150 38138 620
rect 38242 150 38270 620
rect 38470 500 38476 552
rect 38528 500 38534 552
rect 38706 274 38734 620
rect 38894 274 38922 620
rect 39094 376 39100 428
rect 39152 376 39158 428
rect 38688 222 38694 274
rect 38746 222 38752 274
rect 38876 222 38882 274
rect 38934 222 38940 274
rect 39358 150 39386 620
rect 39490 150 39518 620
rect 39718 500 39724 552
rect 39776 500 39782 552
rect 39954 274 39982 620
rect 40142 274 40170 620
rect 40342 376 40348 428
rect 40400 376 40406 428
rect 39936 222 39942 274
rect 39994 222 40000 274
rect 40124 222 40130 274
rect 40182 222 40188 274
rect 40606 150 40634 620
rect 40738 150 40766 620
rect 40966 500 40972 552
rect 41024 500 41030 552
rect 41202 274 41230 620
rect 41184 222 41190 274
rect 41242 222 41248 274
rect 1900 98 1906 150
rect 1958 98 1964 150
rect 2032 98 2038 150
rect 2090 98 2096 150
rect 3148 98 3154 150
rect 3206 98 3212 150
rect 3280 98 3286 150
rect 3338 98 3344 150
rect 4396 98 4402 150
rect 4454 98 4460 150
rect 4528 98 4534 150
rect 4586 98 4592 150
rect 5644 98 5650 150
rect 5702 98 5708 150
rect 5776 98 5782 150
rect 5834 98 5840 150
rect 6892 98 6898 150
rect 6950 98 6956 150
rect 7024 98 7030 150
rect 7082 98 7088 150
rect 8140 98 8146 150
rect 8198 98 8204 150
rect 8272 98 8278 150
rect 8330 98 8336 150
rect 9388 98 9394 150
rect 9446 98 9452 150
rect 9520 98 9526 150
rect 9578 98 9584 150
rect 10636 98 10642 150
rect 10694 98 10700 150
rect 10768 98 10774 150
rect 10826 98 10832 150
rect 11884 98 11890 150
rect 11942 98 11948 150
rect 12016 98 12022 150
rect 12074 98 12080 150
rect 13132 98 13138 150
rect 13190 98 13196 150
rect 13264 98 13270 150
rect 13322 98 13328 150
rect 14380 98 14386 150
rect 14438 98 14444 150
rect 14512 98 14518 150
rect 14570 98 14576 150
rect 15628 98 15634 150
rect 15686 98 15692 150
rect 15760 98 15766 150
rect 15818 98 15824 150
rect 16876 98 16882 150
rect 16934 98 16940 150
rect 17008 98 17014 150
rect 17066 98 17072 150
rect 18124 98 18130 150
rect 18182 98 18188 150
rect 18256 98 18262 150
rect 18314 98 18320 150
rect 19372 98 19378 150
rect 19430 98 19436 150
rect 19504 98 19510 150
rect 19562 98 19568 150
rect 20620 98 20626 150
rect 20678 98 20684 150
rect 20752 98 20758 150
rect 20810 98 20816 150
rect 21868 98 21874 150
rect 21926 98 21932 150
rect 22000 98 22006 150
rect 22058 98 22064 150
rect 23116 98 23122 150
rect 23174 98 23180 150
rect 23248 98 23254 150
rect 23306 98 23312 150
rect 24364 98 24370 150
rect 24422 98 24428 150
rect 24496 98 24502 150
rect 24554 98 24560 150
rect 25612 98 25618 150
rect 25670 98 25676 150
rect 25744 98 25750 150
rect 25802 98 25808 150
rect 26860 98 26866 150
rect 26918 98 26924 150
rect 26992 98 26998 150
rect 27050 98 27056 150
rect 28108 98 28114 150
rect 28166 98 28172 150
rect 28240 98 28246 150
rect 28298 98 28304 150
rect 29356 98 29362 150
rect 29414 98 29420 150
rect 29488 98 29494 150
rect 29546 98 29552 150
rect 30604 98 30610 150
rect 30662 98 30668 150
rect 30736 98 30742 150
rect 30794 98 30800 150
rect 31852 98 31858 150
rect 31910 98 31916 150
rect 31984 98 31990 150
rect 32042 98 32048 150
rect 33100 98 33106 150
rect 33158 98 33164 150
rect 33232 98 33238 150
rect 33290 98 33296 150
rect 34348 98 34354 150
rect 34406 98 34412 150
rect 34480 98 34486 150
rect 34538 98 34544 150
rect 35596 98 35602 150
rect 35654 98 35660 150
rect 35728 98 35734 150
rect 35786 98 35792 150
rect 36844 98 36850 150
rect 36902 98 36908 150
rect 36976 98 36982 150
rect 37034 98 37040 150
rect 38092 98 38098 150
rect 38150 98 38156 150
rect 38224 98 38230 150
rect 38282 98 38288 150
rect 39340 98 39346 150
rect 39398 98 39404 150
rect 39472 98 39478 150
rect 39530 98 39536 150
rect 40588 98 40594 150
rect 40646 98 40652 150
rect 40720 98 40726 150
rect 40778 98 40784 150
<< via1 >>
rect 1660 419 1712 428
rect 1660 385 1669 419
rect 1669 385 1703 419
rect 1703 385 1712 419
rect 1660 376 1712 385
rect 1442 222 1494 274
rect 2284 543 2336 552
rect 2284 509 2293 543
rect 2293 509 2327 543
rect 2327 509 2336 543
rect 2284 500 2336 509
rect 2908 419 2960 428
rect 2908 385 2917 419
rect 2917 385 2951 419
rect 2951 385 2960 419
rect 2908 376 2960 385
rect 2502 222 2554 274
rect 2690 222 2742 274
rect 3532 543 3584 552
rect 3532 509 3541 543
rect 3541 509 3575 543
rect 3575 509 3584 543
rect 3532 500 3584 509
rect 4156 419 4208 428
rect 4156 385 4165 419
rect 4165 385 4199 419
rect 4199 385 4208 419
rect 4156 376 4208 385
rect 3750 222 3802 274
rect 3938 222 3990 274
rect 4780 543 4832 552
rect 4780 509 4789 543
rect 4789 509 4823 543
rect 4823 509 4832 543
rect 4780 500 4832 509
rect 5404 419 5456 428
rect 5404 385 5413 419
rect 5413 385 5447 419
rect 5447 385 5456 419
rect 5404 376 5456 385
rect 4998 222 5050 274
rect 5186 222 5238 274
rect 6028 543 6080 552
rect 6028 509 6037 543
rect 6037 509 6071 543
rect 6071 509 6080 543
rect 6028 500 6080 509
rect 6652 419 6704 428
rect 6652 385 6661 419
rect 6661 385 6695 419
rect 6695 385 6704 419
rect 6652 376 6704 385
rect 6246 222 6298 274
rect 6434 222 6486 274
rect 7276 543 7328 552
rect 7276 509 7285 543
rect 7285 509 7319 543
rect 7319 509 7328 543
rect 7276 500 7328 509
rect 7900 419 7952 428
rect 7900 385 7909 419
rect 7909 385 7943 419
rect 7943 385 7952 419
rect 7900 376 7952 385
rect 7494 222 7546 274
rect 7682 222 7734 274
rect 8524 543 8576 552
rect 8524 509 8533 543
rect 8533 509 8567 543
rect 8567 509 8576 543
rect 8524 500 8576 509
rect 9148 419 9200 428
rect 9148 385 9157 419
rect 9157 385 9191 419
rect 9191 385 9200 419
rect 9148 376 9200 385
rect 8742 222 8794 274
rect 8930 222 8982 274
rect 9772 543 9824 552
rect 9772 509 9781 543
rect 9781 509 9815 543
rect 9815 509 9824 543
rect 9772 500 9824 509
rect 10396 419 10448 428
rect 10396 385 10405 419
rect 10405 385 10439 419
rect 10439 385 10448 419
rect 10396 376 10448 385
rect 9990 222 10042 274
rect 10178 222 10230 274
rect 11020 543 11072 552
rect 11020 509 11029 543
rect 11029 509 11063 543
rect 11063 509 11072 543
rect 11020 500 11072 509
rect 11644 419 11696 428
rect 11644 385 11653 419
rect 11653 385 11687 419
rect 11687 385 11696 419
rect 11644 376 11696 385
rect 11238 222 11290 274
rect 11426 222 11478 274
rect 12268 543 12320 552
rect 12268 509 12277 543
rect 12277 509 12311 543
rect 12311 509 12320 543
rect 12268 500 12320 509
rect 12892 419 12944 428
rect 12892 385 12901 419
rect 12901 385 12935 419
rect 12935 385 12944 419
rect 12892 376 12944 385
rect 12486 222 12538 274
rect 12674 222 12726 274
rect 13516 543 13568 552
rect 13516 509 13525 543
rect 13525 509 13559 543
rect 13559 509 13568 543
rect 13516 500 13568 509
rect 14140 419 14192 428
rect 14140 385 14149 419
rect 14149 385 14183 419
rect 14183 385 14192 419
rect 14140 376 14192 385
rect 13734 222 13786 274
rect 13922 222 13974 274
rect 14764 543 14816 552
rect 14764 509 14773 543
rect 14773 509 14807 543
rect 14807 509 14816 543
rect 14764 500 14816 509
rect 15388 419 15440 428
rect 15388 385 15397 419
rect 15397 385 15431 419
rect 15431 385 15440 419
rect 15388 376 15440 385
rect 14982 222 15034 274
rect 15170 222 15222 274
rect 16012 543 16064 552
rect 16012 509 16021 543
rect 16021 509 16055 543
rect 16055 509 16064 543
rect 16012 500 16064 509
rect 16636 419 16688 428
rect 16636 385 16645 419
rect 16645 385 16679 419
rect 16679 385 16688 419
rect 16636 376 16688 385
rect 16230 222 16282 274
rect 16418 222 16470 274
rect 17260 543 17312 552
rect 17260 509 17269 543
rect 17269 509 17303 543
rect 17303 509 17312 543
rect 17260 500 17312 509
rect 17884 419 17936 428
rect 17884 385 17893 419
rect 17893 385 17927 419
rect 17927 385 17936 419
rect 17884 376 17936 385
rect 17478 222 17530 274
rect 17666 222 17718 274
rect 18508 543 18560 552
rect 18508 509 18517 543
rect 18517 509 18551 543
rect 18551 509 18560 543
rect 18508 500 18560 509
rect 19132 419 19184 428
rect 19132 385 19141 419
rect 19141 385 19175 419
rect 19175 385 19184 419
rect 19132 376 19184 385
rect 18726 222 18778 274
rect 18914 222 18966 274
rect 19756 543 19808 552
rect 19756 509 19765 543
rect 19765 509 19799 543
rect 19799 509 19808 543
rect 19756 500 19808 509
rect 20380 419 20432 428
rect 20380 385 20389 419
rect 20389 385 20423 419
rect 20423 385 20432 419
rect 20380 376 20432 385
rect 19974 222 20026 274
rect 20162 222 20214 274
rect 21004 543 21056 552
rect 21004 509 21013 543
rect 21013 509 21047 543
rect 21047 509 21056 543
rect 21004 500 21056 509
rect 21628 419 21680 428
rect 21628 385 21637 419
rect 21637 385 21671 419
rect 21671 385 21680 419
rect 21628 376 21680 385
rect 21222 222 21274 274
rect 21410 222 21462 274
rect 22252 543 22304 552
rect 22252 509 22261 543
rect 22261 509 22295 543
rect 22295 509 22304 543
rect 22252 500 22304 509
rect 22876 419 22928 428
rect 22876 385 22885 419
rect 22885 385 22919 419
rect 22919 385 22928 419
rect 22876 376 22928 385
rect 22470 222 22522 274
rect 22658 222 22710 274
rect 23500 543 23552 552
rect 23500 509 23509 543
rect 23509 509 23543 543
rect 23543 509 23552 543
rect 23500 500 23552 509
rect 24124 419 24176 428
rect 24124 385 24133 419
rect 24133 385 24167 419
rect 24167 385 24176 419
rect 24124 376 24176 385
rect 23718 222 23770 274
rect 23906 222 23958 274
rect 24748 543 24800 552
rect 24748 509 24757 543
rect 24757 509 24791 543
rect 24791 509 24800 543
rect 24748 500 24800 509
rect 25372 419 25424 428
rect 25372 385 25381 419
rect 25381 385 25415 419
rect 25415 385 25424 419
rect 25372 376 25424 385
rect 24966 222 25018 274
rect 25154 222 25206 274
rect 25996 543 26048 552
rect 25996 509 26005 543
rect 26005 509 26039 543
rect 26039 509 26048 543
rect 25996 500 26048 509
rect 26620 419 26672 428
rect 26620 385 26629 419
rect 26629 385 26663 419
rect 26663 385 26672 419
rect 26620 376 26672 385
rect 26214 222 26266 274
rect 26402 222 26454 274
rect 27244 543 27296 552
rect 27244 509 27253 543
rect 27253 509 27287 543
rect 27287 509 27296 543
rect 27244 500 27296 509
rect 27868 419 27920 428
rect 27868 385 27877 419
rect 27877 385 27911 419
rect 27911 385 27920 419
rect 27868 376 27920 385
rect 27462 222 27514 274
rect 27650 222 27702 274
rect 28492 543 28544 552
rect 28492 509 28501 543
rect 28501 509 28535 543
rect 28535 509 28544 543
rect 28492 500 28544 509
rect 29116 419 29168 428
rect 29116 385 29125 419
rect 29125 385 29159 419
rect 29159 385 29168 419
rect 29116 376 29168 385
rect 28710 222 28762 274
rect 28898 222 28950 274
rect 29740 543 29792 552
rect 29740 509 29749 543
rect 29749 509 29783 543
rect 29783 509 29792 543
rect 29740 500 29792 509
rect 30364 419 30416 428
rect 30364 385 30373 419
rect 30373 385 30407 419
rect 30407 385 30416 419
rect 30364 376 30416 385
rect 29958 222 30010 274
rect 30146 222 30198 274
rect 30988 543 31040 552
rect 30988 509 30997 543
rect 30997 509 31031 543
rect 31031 509 31040 543
rect 30988 500 31040 509
rect 31612 419 31664 428
rect 31612 385 31621 419
rect 31621 385 31655 419
rect 31655 385 31664 419
rect 31612 376 31664 385
rect 31206 222 31258 274
rect 31394 222 31446 274
rect 32236 543 32288 552
rect 32236 509 32245 543
rect 32245 509 32279 543
rect 32279 509 32288 543
rect 32236 500 32288 509
rect 32860 419 32912 428
rect 32860 385 32869 419
rect 32869 385 32903 419
rect 32903 385 32912 419
rect 32860 376 32912 385
rect 32454 222 32506 274
rect 32642 222 32694 274
rect 33484 543 33536 552
rect 33484 509 33493 543
rect 33493 509 33527 543
rect 33527 509 33536 543
rect 33484 500 33536 509
rect 34108 419 34160 428
rect 34108 385 34117 419
rect 34117 385 34151 419
rect 34151 385 34160 419
rect 34108 376 34160 385
rect 33702 222 33754 274
rect 33890 222 33942 274
rect 34732 543 34784 552
rect 34732 509 34741 543
rect 34741 509 34775 543
rect 34775 509 34784 543
rect 34732 500 34784 509
rect 35356 419 35408 428
rect 35356 385 35365 419
rect 35365 385 35399 419
rect 35399 385 35408 419
rect 35356 376 35408 385
rect 34950 222 35002 274
rect 35138 222 35190 274
rect 35980 543 36032 552
rect 35980 509 35989 543
rect 35989 509 36023 543
rect 36023 509 36032 543
rect 35980 500 36032 509
rect 36604 419 36656 428
rect 36604 385 36613 419
rect 36613 385 36647 419
rect 36647 385 36656 419
rect 36604 376 36656 385
rect 36198 222 36250 274
rect 36386 222 36438 274
rect 37228 543 37280 552
rect 37228 509 37237 543
rect 37237 509 37271 543
rect 37271 509 37280 543
rect 37228 500 37280 509
rect 37852 419 37904 428
rect 37852 385 37861 419
rect 37861 385 37895 419
rect 37895 385 37904 419
rect 37852 376 37904 385
rect 37446 222 37498 274
rect 37634 222 37686 274
rect 38476 543 38528 552
rect 38476 509 38485 543
rect 38485 509 38519 543
rect 38519 509 38528 543
rect 38476 500 38528 509
rect 39100 419 39152 428
rect 39100 385 39109 419
rect 39109 385 39143 419
rect 39143 385 39152 419
rect 39100 376 39152 385
rect 38694 222 38746 274
rect 38882 222 38934 274
rect 39724 543 39776 552
rect 39724 509 39733 543
rect 39733 509 39767 543
rect 39767 509 39776 543
rect 39724 500 39776 509
rect 40348 419 40400 428
rect 40348 385 40357 419
rect 40357 385 40391 419
rect 40391 385 40400 419
rect 40348 376 40400 385
rect 39942 222 39994 274
rect 40130 222 40182 274
rect 40972 543 41024 552
rect 40972 509 40981 543
rect 40981 509 41015 543
rect 41015 509 41024 543
rect 40972 500 41024 509
rect 41190 222 41242 274
rect 1906 98 1958 150
rect 2038 98 2090 150
rect 3154 98 3206 150
rect 3286 98 3338 150
rect 4402 98 4454 150
rect 4534 98 4586 150
rect 5650 98 5702 150
rect 5782 98 5834 150
rect 6898 98 6950 150
rect 7030 98 7082 150
rect 8146 98 8198 150
rect 8278 98 8330 150
rect 9394 98 9446 150
rect 9526 98 9578 150
rect 10642 98 10694 150
rect 10774 98 10826 150
rect 11890 98 11942 150
rect 12022 98 12074 150
rect 13138 98 13190 150
rect 13270 98 13322 150
rect 14386 98 14438 150
rect 14518 98 14570 150
rect 15634 98 15686 150
rect 15766 98 15818 150
rect 16882 98 16934 150
rect 17014 98 17066 150
rect 18130 98 18182 150
rect 18262 98 18314 150
rect 19378 98 19430 150
rect 19510 98 19562 150
rect 20626 98 20678 150
rect 20758 98 20810 150
rect 21874 98 21926 150
rect 22006 98 22058 150
rect 23122 98 23174 150
rect 23254 98 23306 150
rect 24370 98 24422 150
rect 24502 98 24554 150
rect 25618 98 25670 150
rect 25750 98 25802 150
rect 26866 98 26918 150
rect 26998 98 27050 150
rect 28114 98 28166 150
rect 28246 98 28298 150
rect 29362 98 29414 150
rect 29494 98 29546 150
rect 30610 98 30662 150
rect 30742 98 30794 150
rect 31858 98 31910 150
rect 31990 98 32042 150
rect 33106 98 33158 150
rect 33238 98 33290 150
rect 34354 98 34406 150
rect 34486 98 34538 150
rect 35602 98 35654 150
rect 35734 98 35786 150
rect 36850 98 36902 150
rect 36982 98 37034 150
rect 38098 98 38150 150
rect 38230 98 38282 150
rect 39346 98 39398 150
rect 39478 98 39530 150
rect 40594 98 40646 150
rect 40726 98 40778 150
<< metal2 >>
rect 2282 554 2338 563
rect 2282 489 2338 498
rect 3530 554 3586 563
rect 3530 489 3586 498
rect 4778 554 4834 563
rect 4778 489 4834 498
rect 6026 554 6082 563
rect 6026 489 6082 498
rect 7274 554 7330 563
rect 7274 489 7330 498
rect 8522 554 8578 563
rect 8522 489 8578 498
rect 9770 554 9826 563
rect 9770 489 9826 498
rect 11018 554 11074 563
rect 11018 489 11074 498
rect 12266 554 12322 563
rect 12266 489 12322 498
rect 13514 554 13570 563
rect 13514 489 13570 498
rect 14762 554 14818 563
rect 14762 489 14818 498
rect 16010 554 16066 563
rect 16010 489 16066 498
rect 17258 554 17314 563
rect 17258 489 17314 498
rect 18506 554 18562 563
rect 18506 489 18562 498
rect 19754 554 19810 563
rect 19754 489 19810 498
rect 21002 554 21058 563
rect 21002 489 21058 498
rect 22250 554 22306 563
rect 22250 489 22306 498
rect 23498 554 23554 563
rect 23498 489 23554 498
rect 24746 554 24802 563
rect 24746 489 24802 498
rect 25994 554 26050 563
rect 25994 489 26050 498
rect 27242 554 27298 563
rect 27242 489 27298 498
rect 28490 554 28546 563
rect 28490 489 28546 498
rect 29738 554 29794 563
rect 29738 489 29794 498
rect 30986 554 31042 563
rect 30986 489 31042 498
rect 32234 554 32290 563
rect 32234 489 32290 498
rect 33482 554 33538 563
rect 33482 489 33538 498
rect 34730 554 34786 563
rect 34730 489 34786 498
rect 35978 554 36034 563
rect 35978 489 36034 498
rect 37226 554 37282 563
rect 37226 489 37282 498
rect 38474 554 38530 563
rect 38474 489 38530 498
rect 39722 554 39778 563
rect 39722 489 39778 498
rect 40970 554 41026 563
rect 40970 489 41026 498
rect 1658 430 1714 439
rect 1658 365 1714 374
rect 2906 430 2962 439
rect 2906 365 2962 374
rect 4154 430 4210 439
rect 4154 365 4210 374
rect 5402 430 5458 439
rect 5402 365 5458 374
rect 6650 430 6706 439
rect 6650 365 6706 374
rect 7898 430 7954 439
rect 7898 365 7954 374
rect 9146 430 9202 439
rect 9146 365 9202 374
rect 10394 430 10450 439
rect 10394 365 10450 374
rect 11642 430 11698 439
rect 11642 365 11698 374
rect 12890 430 12946 439
rect 12890 365 12946 374
rect 14138 430 14194 439
rect 14138 365 14194 374
rect 15386 430 15442 439
rect 15386 365 15442 374
rect 16634 430 16690 439
rect 16634 365 16690 374
rect 17882 430 17938 439
rect 17882 365 17938 374
rect 19130 430 19186 439
rect 19130 365 19186 374
rect 20378 430 20434 439
rect 20378 365 20434 374
rect 21626 430 21682 439
rect 21626 365 21682 374
rect 22874 430 22930 439
rect 22874 365 22930 374
rect 24122 430 24178 439
rect 24122 365 24178 374
rect 25370 430 25426 439
rect 25370 365 25426 374
rect 26618 430 26674 439
rect 26618 365 26674 374
rect 27866 430 27922 439
rect 27866 365 27922 374
rect 29114 430 29170 439
rect 29114 365 29170 374
rect 30362 430 30418 439
rect 30362 365 30418 374
rect 31610 430 31666 439
rect 31610 365 31666 374
rect 32858 430 32914 439
rect 32858 365 32914 374
rect 34106 430 34162 439
rect 34106 365 34162 374
rect 35354 430 35410 439
rect 35354 365 35410 374
rect 36602 430 36658 439
rect 36602 365 36658 374
rect 37850 430 37906 439
rect 37850 365 37906 374
rect 39098 430 39154 439
rect 39098 365 39154 374
rect 40346 430 40402 439
rect 40346 365 40402 374
rect 1440 276 1496 285
rect 1440 211 1496 220
rect 2500 276 2556 285
rect 2500 211 2556 220
rect 2688 276 2744 285
rect 2688 211 2744 220
rect 3748 276 3804 285
rect 3748 211 3804 220
rect 3936 276 3992 285
rect 3936 211 3992 220
rect 4996 276 5052 285
rect 4996 211 5052 220
rect 5184 276 5240 285
rect 5184 211 5240 220
rect 6244 276 6300 285
rect 6244 211 6300 220
rect 6432 276 6488 285
rect 6432 211 6488 220
rect 7492 276 7548 285
rect 7492 211 7548 220
rect 7680 276 7736 285
rect 7680 211 7736 220
rect 8740 276 8796 285
rect 8740 211 8796 220
rect 8928 276 8984 285
rect 8928 211 8984 220
rect 9988 276 10044 285
rect 9988 211 10044 220
rect 10176 276 10232 285
rect 10176 211 10232 220
rect 11236 276 11292 285
rect 11236 211 11292 220
rect 11424 276 11480 285
rect 11424 211 11480 220
rect 12484 276 12540 285
rect 12484 211 12540 220
rect 12672 276 12728 285
rect 12672 211 12728 220
rect 13732 276 13788 285
rect 13732 211 13788 220
rect 13920 276 13976 285
rect 13920 211 13976 220
rect 14980 276 15036 285
rect 14980 211 15036 220
rect 15168 276 15224 285
rect 15168 211 15224 220
rect 16228 276 16284 285
rect 16228 211 16284 220
rect 16416 276 16472 285
rect 16416 211 16472 220
rect 17476 276 17532 285
rect 17476 211 17532 220
rect 17664 276 17720 285
rect 17664 211 17720 220
rect 18724 276 18780 285
rect 18724 211 18780 220
rect 18912 276 18968 285
rect 18912 211 18968 220
rect 19972 276 20028 285
rect 19972 211 20028 220
rect 20160 276 20216 285
rect 20160 211 20216 220
rect 21220 276 21276 285
rect 21220 211 21276 220
rect 21408 276 21464 285
rect 21408 211 21464 220
rect 22468 276 22524 285
rect 22468 211 22524 220
rect 22656 276 22712 285
rect 22656 211 22712 220
rect 23716 276 23772 285
rect 23716 211 23772 220
rect 23904 276 23960 285
rect 23904 211 23960 220
rect 24964 276 25020 285
rect 24964 211 25020 220
rect 25152 276 25208 285
rect 25152 211 25208 220
rect 26212 276 26268 285
rect 26212 211 26268 220
rect 26400 276 26456 285
rect 26400 211 26456 220
rect 27460 276 27516 285
rect 27460 211 27516 220
rect 27648 276 27704 285
rect 27648 211 27704 220
rect 28708 276 28764 285
rect 28708 211 28764 220
rect 28896 276 28952 285
rect 28896 211 28952 220
rect 29956 276 30012 285
rect 29956 211 30012 220
rect 30144 276 30200 285
rect 30144 211 30200 220
rect 31204 276 31260 285
rect 31204 211 31260 220
rect 31392 276 31448 285
rect 31392 211 31448 220
rect 32452 276 32508 285
rect 32452 211 32508 220
rect 32640 276 32696 285
rect 32640 211 32696 220
rect 33700 276 33756 285
rect 33700 211 33756 220
rect 33888 276 33944 285
rect 33888 211 33944 220
rect 34948 276 35004 285
rect 34948 211 35004 220
rect 35136 276 35192 285
rect 35136 211 35192 220
rect 36196 276 36252 285
rect 36196 211 36252 220
rect 36384 276 36440 285
rect 36384 211 36440 220
rect 37444 276 37500 285
rect 37444 211 37500 220
rect 37632 276 37688 285
rect 37632 211 37688 220
rect 38692 276 38748 285
rect 38692 211 38748 220
rect 38880 276 38936 285
rect 38880 211 38936 220
rect 39940 276 39996 285
rect 39940 211 39996 220
rect 40128 276 40184 285
rect 40128 211 40184 220
rect 41188 276 41244 285
rect 41188 211 41244 220
rect 1904 152 1960 161
rect 1904 87 1960 96
rect 2036 152 2092 161
rect 2036 87 2092 96
rect 3152 152 3208 161
rect 3152 87 3208 96
rect 3284 152 3340 161
rect 3284 87 3340 96
rect 4400 152 4456 161
rect 4400 87 4456 96
rect 4532 152 4588 161
rect 4532 87 4588 96
rect 5648 152 5704 161
rect 5648 87 5704 96
rect 5780 152 5836 161
rect 5780 87 5836 96
rect 6896 152 6952 161
rect 6896 87 6952 96
rect 7028 152 7084 161
rect 7028 87 7084 96
rect 8144 152 8200 161
rect 8144 87 8200 96
rect 8276 152 8332 161
rect 8276 87 8332 96
rect 9392 152 9448 161
rect 9392 87 9448 96
rect 9524 152 9580 161
rect 9524 87 9580 96
rect 10640 152 10696 161
rect 10640 87 10696 96
rect 10772 152 10828 161
rect 10772 87 10828 96
rect 11888 152 11944 161
rect 11888 87 11944 96
rect 12020 152 12076 161
rect 12020 87 12076 96
rect 13136 152 13192 161
rect 13136 87 13192 96
rect 13268 152 13324 161
rect 13268 87 13324 96
rect 14384 152 14440 161
rect 14384 87 14440 96
rect 14516 152 14572 161
rect 14516 87 14572 96
rect 15632 152 15688 161
rect 15632 87 15688 96
rect 15764 152 15820 161
rect 15764 87 15820 96
rect 16880 152 16936 161
rect 16880 87 16936 96
rect 17012 152 17068 161
rect 17012 87 17068 96
rect 18128 152 18184 161
rect 18128 87 18184 96
rect 18260 152 18316 161
rect 18260 87 18316 96
rect 19376 152 19432 161
rect 19376 87 19432 96
rect 19508 152 19564 161
rect 19508 87 19564 96
rect 20624 152 20680 161
rect 20624 87 20680 96
rect 20756 152 20812 161
rect 20756 87 20812 96
rect 21872 152 21928 161
rect 21872 87 21928 96
rect 22004 152 22060 161
rect 22004 87 22060 96
rect 23120 152 23176 161
rect 23120 87 23176 96
rect 23252 152 23308 161
rect 23252 87 23308 96
rect 24368 152 24424 161
rect 24368 87 24424 96
rect 24500 152 24556 161
rect 24500 87 24556 96
rect 25616 152 25672 161
rect 25616 87 25672 96
rect 25748 152 25804 161
rect 25748 87 25804 96
rect 26864 152 26920 161
rect 26864 87 26920 96
rect 26996 152 27052 161
rect 26996 87 27052 96
rect 28112 152 28168 161
rect 28112 87 28168 96
rect 28244 152 28300 161
rect 28244 87 28300 96
rect 29360 152 29416 161
rect 29360 87 29416 96
rect 29492 152 29548 161
rect 29492 87 29548 96
rect 30608 152 30664 161
rect 30608 87 30664 96
rect 30740 152 30796 161
rect 30740 87 30796 96
rect 31856 152 31912 161
rect 31856 87 31912 96
rect 31988 152 32044 161
rect 31988 87 32044 96
rect 33104 152 33160 161
rect 33104 87 33160 96
rect 33236 152 33292 161
rect 33236 87 33292 96
rect 34352 152 34408 161
rect 34352 87 34408 96
rect 34484 152 34540 161
rect 34484 87 34540 96
rect 35600 152 35656 161
rect 35600 87 35656 96
rect 35732 152 35788 161
rect 35732 87 35788 96
rect 36848 152 36904 161
rect 36848 87 36904 96
rect 36980 152 37036 161
rect 36980 87 37036 96
rect 38096 152 38152 161
rect 38096 87 38152 96
rect 38228 152 38284 161
rect 38228 87 38284 96
rect 39344 152 39400 161
rect 39344 87 39400 96
rect 39476 152 39532 161
rect 39476 87 39532 96
rect 40592 152 40648 161
rect 40592 87 40648 96
rect 40724 152 40780 161
rect 40724 87 40780 96
<< via2 >>
rect 2282 552 2338 554
rect 2282 500 2284 552
rect 2284 500 2336 552
rect 2336 500 2338 552
rect 2282 498 2338 500
rect 3530 552 3586 554
rect 3530 500 3532 552
rect 3532 500 3584 552
rect 3584 500 3586 552
rect 3530 498 3586 500
rect 4778 552 4834 554
rect 4778 500 4780 552
rect 4780 500 4832 552
rect 4832 500 4834 552
rect 4778 498 4834 500
rect 6026 552 6082 554
rect 6026 500 6028 552
rect 6028 500 6080 552
rect 6080 500 6082 552
rect 6026 498 6082 500
rect 7274 552 7330 554
rect 7274 500 7276 552
rect 7276 500 7328 552
rect 7328 500 7330 552
rect 7274 498 7330 500
rect 8522 552 8578 554
rect 8522 500 8524 552
rect 8524 500 8576 552
rect 8576 500 8578 552
rect 8522 498 8578 500
rect 9770 552 9826 554
rect 9770 500 9772 552
rect 9772 500 9824 552
rect 9824 500 9826 552
rect 9770 498 9826 500
rect 11018 552 11074 554
rect 11018 500 11020 552
rect 11020 500 11072 552
rect 11072 500 11074 552
rect 11018 498 11074 500
rect 12266 552 12322 554
rect 12266 500 12268 552
rect 12268 500 12320 552
rect 12320 500 12322 552
rect 12266 498 12322 500
rect 13514 552 13570 554
rect 13514 500 13516 552
rect 13516 500 13568 552
rect 13568 500 13570 552
rect 13514 498 13570 500
rect 14762 552 14818 554
rect 14762 500 14764 552
rect 14764 500 14816 552
rect 14816 500 14818 552
rect 14762 498 14818 500
rect 16010 552 16066 554
rect 16010 500 16012 552
rect 16012 500 16064 552
rect 16064 500 16066 552
rect 16010 498 16066 500
rect 17258 552 17314 554
rect 17258 500 17260 552
rect 17260 500 17312 552
rect 17312 500 17314 552
rect 17258 498 17314 500
rect 18506 552 18562 554
rect 18506 500 18508 552
rect 18508 500 18560 552
rect 18560 500 18562 552
rect 18506 498 18562 500
rect 19754 552 19810 554
rect 19754 500 19756 552
rect 19756 500 19808 552
rect 19808 500 19810 552
rect 19754 498 19810 500
rect 21002 552 21058 554
rect 21002 500 21004 552
rect 21004 500 21056 552
rect 21056 500 21058 552
rect 21002 498 21058 500
rect 22250 552 22306 554
rect 22250 500 22252 552
rect 22252 500 22304 552
rect 22304 500 22306 552
rect 22250 498 22306 500
rect 23498 552 23554 554
rect 23498 500 23500 552
rect 23500 500 23552 552
rect 23552 500 23554 552
rect 23498 498 23554 500
rect 24746 552 24802 554
rect 24746 500 24748 552
rect 24748 500 24800 552
rect 24800 500 24802 552
rect 24746 498 24802 500
rect 25994 552 26050 554
rect 25994 500 25996 552
rect 25996 500 26048 552
rect 26048 500 26050 552
rect 25994 498 26050 500
rect 27242 552 27298 554
rect 27242 500 27244 552
rect 27244 500 27296 552
rect 27296 500 27298 552
rect 27242 498 27298 500
rect 28490 552 28546 554
rect 28490 500 28492 552
rect 28492 500 28544 552
rect 28544 500 28546 552
rect 28490 498 28546 500
rect 29738 552 29794 554
rect 29738 500 29740 552
rect 29740 500 29792 552
rect 29792 500 29794 552
rect 29738 498 29794 500
rect 30986 552 31042 554
rect 30986 500 30988 552
rect 30988 500 31040 552
rect 31040 500 31042 552
rect 30986 498 31042 500
rect 32234 552 32290 554
rect 32234 500 32236 552
rect 32236 500 32288 552
rect 32288 500 32290 552
rect 32234 498 32290 500
rect 33482 552 33538 554
rect 33482 500 33484 552
rect 33484 500 33536 552
rect 33536 500 33538 552
rect 33482 498 33538 500
rect 34730 552 34786 554
rect 34730 500 34732 552
rect 34732 500 34784 552
rect 34784 500 34786 552
rect 34730 498 34786 500
rect 35978 552 36034 554
rect 35978 500 35980 552
rect 35980 500 36032 552
rect 36032 500 36034 552
rect 35978 498 36034 500
rect 37226 552 37282 554
rect 37226 500 37228 552
rect 37228 500 37280 552
rect 37280 500 37282 552
rect 37226 498 37282 500
rect 38474 552 38530 554
rect 38474 500 38476 552
rect 38476 500 38528 552
rect 38528 500 38530 552
rect 38474 498 38530 500
rect 39722 552 39778 554
rect 39722 500 39724 552
rect 39724 500 39776 552
rect 39776 500 39778 552
rect 39722 498 39778 500
rect 40970 552 41026 554
rect 40970 500 40972 552
rect 40972 500 41024 552
rect 41024 500 41026 552
rect 40970 498 41026 500
rect 1658 428 1714 430
rect 1658 376 1660 428
rect 1660 376 1712 428
rect 1712 376 1714 428
rect 1658 374 1714 376
rect 2906 428 2962 430
rect 2906 376 2908 428
rect 2908 376 2960 428
rect 2960 376 2962 428
rect 2906 374 2962 376
rect 4154 428 4210 430
rect 4154 376 4156 428
rect 4156 376 4208 428
rect 4208 376 4210 428
rect 4154 374 4210 376
rect 5402 428 5458 430
rect 5402 376 5404 428
rect 5404 376 5456 428
rect 5456 376 5458 428
rect 5402 374 5458 376
rect 6650 428 6706 430
rect 6650 376 6652 428
rect 6652 376 6704 428
rect 6704 376 6706 428
rect 6650 374 6706 376
rect 7898 428 7954 430
rect 7898 376 7900 428
rect 7900 376 7952 428
rect 7952 376 7954 428
rect 7898 374 7954 376
rect 9146 428 9202 430
rect 9146 376 9148 428
rect 9148 376 9200 428
rect 9200 376 9202 428
rect 9146 374 9202 376
rect 10394 428 10450 430
rect 10394 376 10396 428
rect 10396 376 10448 428
rect 10448 376 10450 428
rect 10394 374 10450 376
rect 11642 428 11698 430
rect 11642 376 11644 428
rect 11644 376 11696 428
rect 11696 376 11698 428
rect 11642 374 11698 376
rect 12890 428 12946 430
rect 12890 376 12892 428
rect 12892 376 12944 428
rect 12944 376 12946 428
rect 12890 374 12946 376
rect 14138 428 14194 430
rect 14138 376 14140 428
rect 14140 376 14192 428
rect 14192 376 14194 428
rect 14138 374 14194 376
rect 15386 428 15442 430
rect 15386 376 15388 428
rect 15388 376 15440 428
rect 15440 376 15442 428
rect 15386 374 15442 376
rect 16634 428 16690 430
rect 16634 376 16636 428
rect 16636 376 16688 428
rect 16688 376 16690 428
rect 16634 374 16690 376
rect 17882 428 17938 430
rect 17882 376 17884 428
rect 17884 376 17936 428
rect 17936 376 17938 428
rect 17882 374 17938 376
rect 19130 428 19186 430
rect 19130 376 19132 428
rect 19132 376 19184 428
rect 19184 376 19186 428
rect 19130 374 19186 376
rect 20378 428 20434 430
rect 20378 376 20380 428
rect 20380 376 20432 428
rect 20432 376 20434 428
rect 20378 374 20434 376
rect 21626 428 21682 430
rect 21626 376 21628 428
rect 21628 376 21680 428
rect 21680 376 21682 428
rect 21626 374 21682 376
rect 22874 428 22930 430
rect 22874 376 22876 428
rect 22876 376 22928 428
rect 22928 376 22930 428
rect 22874 374 22930 376
rect 24122 428 24178 430
rect 24122 376 24124 428
rect 24124 376 24176 428
rect 24176 376 24178 428
rect 24122 374 24178 376
rect 25370 428 25426 430
rect 25370 376 25372 428
rect 25372 376 25424 428
rect 25424 376 25426 428
rect 25370 374 25426 376
rect 26618 428 26674 430
rect 26618 376 26620 428
rect 26620 376 26672 428
rect 26672 376 26674 428
rect 26618 374 26674 376
rect 27866 428 27922 430
rect 27866 376 27868 428
rect 27868 376 27920 428
rect 27920 376 27922 428
rect 27866 374 27922 376
rect 29114 428 29170 430
rect 29114 376 29116 428
rect 29116 376 29168 428
rect 29168 376 29170 428
rect 29114 374 29170 376
rect 30362 428 30418 430
rect 30362 376 30364 428
rect 30364 376 30416 428
rect 30416 376 30418 428
rect 30362 374 30418 376
rect 31610 428 31666 430
rect 31610 376 31612 428
rect 31612 376 31664 428
rect 31664 376 31666 428
rect 31610 374 31666 376
rect 32858 428 32914 430
rect 32858 376 32860 428
rect 32860 376 32912 428
rect 32912 376 32914 428
rect 32858 374 32914 376
rect 34106 428 34162 430
rect 34106 376 34108 428
rect 34108 376 34160 428
rect 34160 376 34162 428
rect 34106 374 34162 376
rect 35354 428 35410 430
rect 35354 376 35356 428
rect 35356 376 35408 428
rect 35408 376 35410 428
rect 35354 374 35410 376
rect 36602 428 36658 430
rect 36602 376 36604 428
rect 36604 376 36656 428
rect 36656 376 36658 428
rect 36602 374 36658 376
rect 37850 428 37906 430
rect 37850 376 37852 428
rect 37852 376 37904 428
rect 37904 376 37906 428
rect 37850 374 37906 376
rect 39098 428 39154 430
rect 39098 376 39100 428
rect 39100 376 39152 428
rect 39152 376 39154 428
rect 39098 374 39154 376
rect 40346 428 40402 430
rect 40346 376 40348 428
rect 40348 376 40400 428
rect 40400 376 40402 428
rect 40346 374 40402 376
rect 1440 274 1496 276
rect 1440 222 1442 274
rect 1442 222 1494 274
rect 1494 222 1496 274
rect 1440 220 1496 222
rect 2500 274 2556 276
rect 2500 222 2502 274
rect 2502 222 2554 274
rect 2554 222 2556 274
rect 2500 220 2556 222
rect 2688 274 2744 276
rect 2688 222 2690 274
rect 2690 222 2742 274
rect 2742 222 2744 274
rect 2688 220 2744 222
rect 3748 274 3804 276
rect 3748 222 3750 274
rect 3750 222 3802 274
rect 3802 222 3804 274
rect 3748 220 3804 222
rect 3936 274 3992 276
rect 3936 222 3938 274
rect 3938 222 3990 274
rect 3990 222 3992 274
rect 3936 220 3992 222
rect 4996 274 5052 276
rect 4996 222 4998 274
rect 4998 222 5050 274
rect 5050 222 5052 274
rect 4996 220 5052 222
rect 5184 274 5240 276
rect 5184 222 5186 274
rect 5186 222 5238 274
rect 5238 222 5240 274
rect 5184 220 5240 222
rect 6244 274 6300 276
rect 6244 222 6246 274
rect 6246 222 6298 274
rect 6298 222 6300 274
rect 6244 220 6300 222
rect 6432 274 6488 276
rect 6432 222 6434 274
rect 6434 222 6486 274
rect 6486 222 6488 274
rect 6432 220 6488 222
rect 7492 274 7548 276
rect 7492 222 7494 274
rect 7494 222 7546 274
rect 7546 222 7548 274
rect 7492 220 7548 222
rect 7680 274 7736 276
rect 7680 222 7682 274
rect 7682 222 7734 274
rect 7734 222 7736 274
rect 7680 220 7736 222
rect 8740 274 8796 276
rect 8740 222 8742 274
rect 8742 222 8794 274
rect 8794 222 8796 274
rect 8740 220 8796 222
rect 8928 274 8984 276
rect 8928 222 8930 274
rect 8930 222 8982 274
rect 8982 222 8984 274
rect 8928 220 8984 222
rect 9988 274 10044 276
rect 9988 222 9990 274
rect 9990 222 10042 274
rect 10042 222 10044 274
rect 9988 220 10044 222
rect 10176 274 10232 276
rect 10176 222 10178 274
rect 10178 222 10230 274
rect 10230 222 10232 274
rect 10176 220 10232 222
rect 11236 274 11292 276
rect 11236 222 11238 274
rect 11238 222 11290 274
rect 11290 222 11292 274
rect 11236 220 11292 222
rect 11424 274 11480 276
rect 11424 222 11426 274
rect 11426 222 11478 274
rect 11478 222 11480 274
rect 11424 220 11480 222
rect 12484 274 12540 276
rect 12484 222 12486 274
rect 12486 222 12538 274
rect 12538 222 12540 274
rect 12484 220 12540 222
rect 12672 274 12728 276
rect 12672 222 12674 274
rect 12674 222 12726 274
rect 12726 222 12728 274
rect 12672 220 12728 222
rect 13732 274 13788 276
rect 13732 222 13734 274
rect 13734 222 13786 274
rect 13786 222 13788 274
rect 13732 220 13788 222
rect 13920 274 13976 276
rect 13920 222 13922 274
rect 13922 222 13974 274
rect 13974 222 13976 274
rect 13920 220 13976 222
rect 14980 274 15036 276
rect 14980 222 14982 274
rect 14982 222 15034 274
rect 15034 222 15036 274
rect 14980 220 15036 222
rect 15168 274 15224 276
rect 15168 222 15170 274
rect 15170 222 15222 274
rect 15222 222 15224 274
rect 15168 220 15224 222
rect 16228 274 16284 276
rect 16228 222 16230 274
rect 16230 222 16282 274
rect 16282 222 16284 274
rect 16228 220 16284 222
rect 16416 274 16472 276
rect 16416 222 16418 274
rect 16418 222 16470 274
rect 16470 222 16472 274
rect 16416 220 16472 222
rect 17476 274 17532 276
rect 17476 222 17478 274
rect 17478 222 17530 274
rect 17530 222 17532 274
rect 17476 220 17532 222
rect 17664 274 17720 276
rect 17664 222 17666 274
rect 17666 222 17718 274
rect 17718 222 17720 274
rect 17664 220 17720 222
rect 18724 274 18780 276
rect 18724 222 18726 274
rect 18726 222 18778 274
rect 18778 222 18780 274
rect 18724 220 18780 222
rect 18912 274 18968 276
rect 18912 222 18914 274
rect 18914 222 18966 274
rect 18966 222 18968 274
rect 18912 220 18968 222
rect 19972 274 20028 276
rect 19972 222 19974 274
rect 19974 222 20026 274
rect 20026 222 20028 274
rect 19972 220 20028 222
rect 20160 274 20216 276
rect 20160 222 20162 274
rect 20162 222 20214 274
rect 20214 222 20216 274
rect 20160 220 20216 222
rect 21220 274 21276 276
rect 21220 222 21222 274
rect 21222 222 21274 274
rect 21274 222 21276 274
rect 21220 220 21276 222
rect 21408 274 21464 276
rect 21408 222 21410 274
rect 21410 222 21462 274
rect 21462 222 21464 274
rect 21408 220 21464 222
rect 22468 274 22524 276
rect 22468 222 22470 274
rect 22470 222 22522 274
rect 22522 222 22524 274
rect 22468 220 22524 222
rect 22656 274 22712 276
rect 22656 222 22658 274
rect 22658 222 22710 274
rect 22710 222 22712 274
rect 22656 220 22712 222
rect 23716 274 23772 276
rect 23716 222 23718 274
rect 23718 222 23770 274
rect 23770 222 23772 274
rect 23716 220 23772 222
rect 23904 274 23960 276
rect 23904 222 23906 274
rect 23906 222 23958 274
rect 23958 222 23960 274
rect 23904 220 23960 222
rect 24964 274 25020 276
rect 24964 222 24966 274
rect 24966 222 25018 274
rect 25018 222 25020 274
rect 24964 220 25020 222
rect 25152 274 25208 276
rect 25152 222 25154 274
rect 25154 222 25206 274
rect 25206 222 25208 274
rect 25152 220 25208 222
rect 26212 274 26268 276
rect 26212 222 26214 274
rect 26214 222 26266 274
rect 26266 222 26268 274
rect 26212 220 26268 222
rect 26400 274 26456 276
rect 26400 222 26402 274
rect 26402 222 26454 274
rect 26454 222 26456 274
rect 26400 220 26456 222
rect 27460 274 27516 276
rect 27460 222 27462 274
rect 27462 222 27514 274
rect 27514 222 27516 274
rect 27460 220 27516 222
rect 27648 274 27704 276
rect 27648 222 27650 274
rect 27650 222 27702 274
rect 27702 222 27704 274
rect 27648 220 27704 222
rect 28708 274 28764 276
rect 28708 222 28710 274
rect 28710 222 28762 274
rect 28762 222 28764 274
rect 28708 220 28764 222
rect 28896 274 28952 276
rect 28896 222 28898 274
rect 28898 222 28950 274
rect 28950 222 28952 274
rect 28896 220 28952 222
rect 29956 274 30012 276
rect 29956 222 29958 274
rect 29958 222 30010 274
rect 30010 222 30012 274
rect 29956 220 30012 222
rect 30144 274 30200 276
rect 30144 222 30146 274
rect 30146 222 30198 274
rect 30198 222 30200 274
rect 30144 220 30200 222
rect 31204 274 31260 276
rect 31204 222 31206 274
rect 31206 222 31258 274
rect 31258 222 31260 274
rect 31204 220 31260 222
rect 31392 274 31448 276
rect 31392 222 31394 274
rect 31394 222 31446 274
rect 31446 222 31448 274
rect 31392 220 31448 222
rect 32452 274 32508 276
rect 32452 222 32454 274
rect 32454 222 32506 274
rect 32506 222 32508 274
rect 32452 220 32508 222
rect 32640 274 32696 276
rect 32640 222 32642 274
rect 32642 222 32694 274
rect 32694 222 32696 274
rect 32640 220 32696 222
rect 33700 274 33756 276
rect 33700 222 33702 274
rect 33702 222 33754 274
rect 33754 222 33756 274
rect 33700 220 33756 222
rect 33888 274 33944 276
rect 33888 222 33890 274
rect 33890 222 33942 274
rect 33942 222 33944 274
rect 33888 220 33944 222
rect 34948 274 35004 276
rect 34948 222 34950 274
rect 34950 222 35002 274
rect 35002 222 35004 274
rect 34948 220 35004 222
rect 35136 274 35192 276
rect 35136 222 35138 274
rect 35138 222 35190 274
rect 35190 222 35192 274
rect 35136 220 35192 222
rect 36196 274 36252 276
rect 36196 222 36198 274
rect 36198 222 36250 274
rect 36250 222 36252 274
rect 36196 220 36252 222
rect 36384 274 36440 276
rect 36384 222 36386 274
rect 36386 222 36438 274
rect 36438 222 36440 274
rect 36384 220 36440 222
rect 37444 274 37500 276
rect 37444 222 37446 274
rect 37446 222 37498 274
rect 37498 222 37500 274
rect 37444 220 37500 222
rect 37632 274 37688 276
rect 37632 222 37634 274
rect 37634 222 37686 274
rect 37686 222 37688 274
rect 37632 220 37688 222
rect 38692 274 38748 276
rect 38692 222 38694 274
rect 38694 222 38746 274
rect 38746 222 38748 274
rect 38692 220 38748 222
rect 38880 274 38936 276
rect 38880 222 38882 274
rect 38882 222 38934 274
rect 38934 222 38936 274
rect 38880 220 38936 222
rect 39940 274 39996 276
rect 39940 222 39942 274
rect 39942 222 39994 274
rect 39994 222 39996 274
rect 39940 220 39996 222
rect 40128 274 40184 276
rect 40128 222 40130 274
rect 40130 222 40182 274
rect 40182 222 40184 274
rect 40128 220 40184 222
rect 41188 274 41244 276
rect 41188 222 41190 274
rect 41190 222 41242 274
rect 41242 222 41244 274
rect 41188 220 41244 222
rect 1904 150 1960 152
rect 1904 98 1906 150
rect 1906 98 1958 150
rect 1958 98 1960 150
rect 1904 96 1960 98
rect 2036 150 2092 152
rect 2036 98 2038 150
rect 2038 98 2090 150
rect 2090 98 2092 150
rect 2036 96 2092 98
rect 3152 150 3208 152
rect 3152 98 3154 150
rect 3154 98 3206 150
rect 3206 98 3208 150
rect 3152 96 3208 98
rect 3284 150 3340 152
rect 3284 98 3286 150
rect 3286 98 3338 150
rect 3338 98 3340 150
rect 3284 96 3340 98
rect 4400 150 4456 152
rect 4400 98 4402 150
rect 4402 98 4454 150
rect 4454 98 4456 150
rect 4400 96 4456 98
rect 4532 150 4588 152
rect 4532 98 4534 150
rect 4534 98 4586 150
rect 4586 98 4588 150
rect 4532 96 4588 98
rect 5648 150 5704 152
rect 5648 98 5650 150
rect 5650 98 5702 150
rect 5702 98 5704 150
rect 5648 96 5704 98
rect 5780 150 5836 152
rect 5780 98 5782 150
rect 5782 98 5834 150
rect 5834 98 5836 150
rect 5780 96 5836 98
rect 6896 150 6952 152
rect 6896 98 6898 150
rect 6898 98 6950 150
rect 6950 98 6952 150
rect 6896 96 6952 98
rect 7028 150 7084 152
rect 7028 98 7030 150
rect 7030 98 7082 150
rect 7082 98 7084 150
rect 7028 96 7084 98
rect 8144 150 8200 152
rect 8144 98 8146 150
rect 8146 98 8198 150
rect 8198 98 8200 150
rect 8144 96 8200 98
rect 8276 150 8332 152
rect 8276 98 8278 150
rect 8278 98 8330 150
rect 8330 98 8332 150
rect 8276 96 8332 98
rect 9392 150 9448 152
rect 9392 98 9394 150
rect 9394 98 9446 150
rect 9446 98 9448 150
rect 9392 96 9448 98
rect 9524 150 9580 152
rect 9524 98 9526 150
rect 9526 98 9578 150
rect 9578 98 9580 150
rect 9524 96 9580 98
rect 10640 150 10696 152
rect 10640 98 10642 150
rect 10642 98 10694 150
rect 10694 98 10696 150
rect 10640 96 10696 98
rect 10772 150 10828 152
rect 10772 98 10774 150
rect 10774 98 10826 150
rect 10826 98 10828 150
rect 10772 96 10828 98
rect 11888 150 11944 152
rect 11888 98 11890 150
rect 11890 98 11942 150
rect 11942 98 11944 150
rect 11888 96 11944 98
rect 12020 150 12076 152
rect 12020 98 12022 150
rect 12022 98 12074 150
rect 12074 98 12076 150
rect 12020 96 12076 98
rect 13136 150 13192 152
rect 13136 98 13138 150
rect 13138 98 13190 150
rect 13190 98 13192 150
rect 13136 96 13192 98
rect 13268 150 13324 152
rect 13268 98 13270 150
rect 13270 98 13322 150
rect 13322 98 13324 150
rect 13268 96 13324 98
rect 14384 150 14440 152
rect 14384 98 14386 150
rect 14386 98 14438 150
rect 14438 98 14440 150
rect 14384 96 14440 98
rect 14516 150 14572 152
rect 14516 98 14518 150
rect 14518 98 14570 150
rect 14570 98 14572 150
rect 14516 96 14572 98
rect 15632 150 15688 152
rect 15632 98 15634 150
rect 15634 98 15686 150
rect 15686 98 15688 150
rect 15632 96 15688 98
rect 15764 150 15820 152
rect 15764 98 15766 150
rect 15766 98 15818 150
rect 15818 98 15820 150
rect 15764 96 15820 98
rect 16880 150 16936 152
rect 16880 98 16882 150
rect 16882 98 16934 150
rect 16934 98 16936 150
rect 16880 96 16936 98
rect 17012 150 17068 152
rect 17012 98 17014 150
rect 17014 98 17066 150
rect 17066 98 17068 150
rect 17012 96 17068 98
rect 18128 150 18184 152
rect 18128 98 18130 150
rect 18130 98 18182 150
rect 18182 98 18184 150
rect 18128 96 18184 98
rect 18260 150 18316 152
rect 18260 98 18262 150
rect 18262 98 18314 150
rect 18314 98 18316 150
rect 18260 96 18316 98
rect 19376 150 19432 152
rect 19376 98 19378 150
rect 19378 98 19430 150
rect 19430 98 19432 150
rect 19376 96 19432 98
rect 19508 150 19564 152
rect 19508 98 19510 150
rect 19510 98 19562 150
rect 19562 98 19564 150
rect 19508 96 19564 98
rect 20624 150 20680 152
rect 20624 98 20626 150
rect 20626 98 20678 150
rect 20678 98 20680 150
rect 20624 96 20680 98
rect 20756 150 20812 152
rect 20756 98 20758 150
rect 20758 98 20810 150
rect 20810 98 20812 150
rect 20756 96 20812 98
rect 21872 150 21928 152
rect 21872 98 21874 150
rect 21874 98 21926 150
rect 21926 98 21928 150
rect 21872 96 21928 98
rect 22004 150 22060 152
rect 22004 98 22006 150
rect 22006 98 22058 150
rect 22058 98 22060 150
rect 22004 96 22060 98
rect 23120 150 23176 152
rect 23120 98 23122 150
rect 23122 98 23174 150
rect 23174 98 23176 150
rect 23120 96 23176 98
rect 23252 150 23308 152
rect 23252 98 23254 150
rect 23254 98 23306 150
rect 23306 98 23308 150
rect 23252 96 23308 98
rect 24368 150 24424 152
rect 24368 98 24370 150
rect 24370 98 24422 150
rect 24422 98 24424 150
rect 24368 96 24424 98
rect 24500 150 24556 152
rect 24500 98 24502 150
rect 24502 98 24554 150
rect 24554 98 24556 150
rect 24500 96 24556 98
rect 25616 150 25672 152
rect 25616 98 25618 150
rect 25618 98 25670 150
rect 25670 98 25672 150
rect 25616 96 25672 98
rect 25748 150 25804 152
rect 25748 98 25750 150
rect 25750 98 25802 150
rect 25802 98 25804 150
rect 25748 96 25804 98
rect 26864 150 26920 152
rect 26864 98 26866 150
rect 26866 98 26918 150
rect 26918 98 26920 150
rect 26864 96 26920 98
rect 26996 150 27052 152
rect 26996 98 26998 150
rect 26998 98 27050 150
rect 27050 98 27052 150
rect 26996 96 27052 98
rect 28112 150 28168 152
rect 28112 98 28114 150
rect 28114 98 28166 150
rect 28166 98 28168 150
rect 28112 96 28168 98
rect 28244 150 28300 152
rect 28244 98 28246 150
rect 28246 98 28298 150
rect 28298 98 28300 150
rect 28244 96 28300 98
rect 29360 150 29416 152
rect 29360 98 29362 150
rect 29362 98 29414 150
rect 29414 98 29416 150
rect 29360 96 29416 98
rect 29492 150 29548 152
rect 29492 98 29494 150
rect 29494 98 29546 150
rect 29546 98 29548 150
rect 29492 96 29548 98
rect 30608 150 30664 152
rect 30608 98 30610 150
rect 30610 98 30662 150
rect 30662 98 30664 150
rect 30608 96 30664 98
rect 30740 150 30796 152
rect 30740 98 30742 150
rect 30742 98 30794 150
rect 30794 98 30796 150
rect 30740 96 30796 98
rect 31856 150 31912 152
rect 31856 98 31858 150
rect 31858 98 31910 150
rect 31910 98 31912 150
rect 31856 96 31912 98
rect 31988 150 32044 152
rect 31988 98 31990 150
rect 31990 98 32042 150
rect 32042 98 32044 150
rect 31988 96 32044 98
rect 33104 150 33160 152
rect 33104 98 33106 150
rect 33106 98 33158 150
rect 33158 98 33160 150
rect 33104 96 33160 98
rect 33236 150 33292 152
rect 33236 98 33238 150
rect 33238 98 33290 150
rect 33290 98 33292 150
rect 33236 96 33292 98
rect 34352 150 34408 152
rect 34352 98 34354 150
rect 34354 98 34406 150
rect 34406 98 34408 150
rect 34352 96 34408 98
rect 34484 150 34540 152
rect 34484 98 34486 150
rect 34486 98 34538 150
rect 34538 98 34540 150
rect 34484 96 34540 98
rect 35600 150 35656 152
rect 35600 98 35602 150
rect 35602 98 35654 150
rect 35654 98 35656 150
rect 35600 96 35656 98
rect 35732 150 35788 152
rect 35732 98 35734 150
rect 35734 98 35786 150
rect 35786 98 35788 150
rect 35732 96 35788 98
rect 36848 150 36904 152
rect 36848 98 36850 150
rect 36850 98 36902 150
rect 36902 98 36904 150
rect 36848 96 36904 98
rect 36980 150 37036 152
rect 36980 98 36982 150
rect 36982 98 37034 150
rect 37034 98 37036 150
rect 36980 96 37036 98
rect 38096 150 38152 152
rect 38096 98 38098 150
rect 38098 98 38150 150
rect 38150 98 38152 150
rect 38096 96 38152 98
rect 38228 150 38284 152
rect 38228 98 38230 150
rect 38230 98 38282 150
rect 38282 98 38284 150
rect 38228 96 38284 98
rect 39344 150 39400 152
rect 39344 98 39346 150
rect 39346 98 39398 150
rect 39398 98 39400 150
rect 39344 96 39400 98
rect 39476 150 39532 152
rect 39476 98 39478 150
rect 39478 98 39530 150
rect 39530 98 39532 150
rect 39476 96 39532 98
rect 40592 150 40648 152
rect 40592 98 40594 150
rect 40594 98 40646 150
rect 40646 98 40648 150
rect 40592 96 40648 98
rect 40724 150 40780 152
rect 40724 98 40726 150
rect 40726 98 40778 150
rect 40778 98 40780 150
rect 40724 96 40780 98
<< metal3 >>
rect 1949 1234 2047 1332
rect 3197 1234 3295 1332
rect 4445 1234 4543 1332
rect 5693 1234 5791 1332
rect 6941 1234 7039 1332
rect 8189 1234 8287 1332
rect 9437 1234 9535 1332
rect 10685 1234 10783 1332
rect 11933 1234 12031 1332
rect 13181 1234 13279 1332
rect 14429 1234 14527 1332
rect 15677 1234 15775 1332
rect 16925 1234 17023 1332
rect 18173 1234 18271 1332
rect 19421 1234 19519 1332
rect 20669 1234 20767 1332
rect 21917 1234 22015 1332
rect 23165 1234 23263 1332
rect 24413 1234 24511 1332
rect 25661 1234 25759 1332
rect 26909 1234 27007 1332
rect 28157 1234 28255 1332
rect 29405 1234 29503 1332
rect 30653 1234 30751 1332
rect 31901 1234 31999 1332
rect 33149 1234 33247 1332
rect 34397 1234 34495 1332
rect 35645 1234 35743 1332
rect 36893 1234 36991 1332
rect 38141 1234 38239 1332
rect 39389 1234 39487 1332
rect 40637 1234 40735 1332
rect 2277 556 2343 559
rect 3525 556 3591 559
rect 4773 556 4839 559
rect 6021 556 6087 559
rect 7269 556 7335 559
rect 8517 556 8583 559
rect 9765 556 9831 559
rect 11013 556 11079 559
rect 12261 556 12327 559
rect 13509 556 13575 559
rect 14757 556 14823 559
rect 16005 556 16071 559
rect 17253 556 17319 559
rect 18501 556 18567 559
rect 19749 556 19815 559
rect 20997 556 21063 559
rect 22245 556 22311 559
rect 23493 556 23559 559
rect 24741 556 24807 559
rect 25989 556 26055 559
rect 27237 556 27303 559
rect 28485 556 28551 559
rect 29733 556 29799 559
rect 30981 556 31047 559
rect 32229 556 32295 559
rect 33477 556 33543 559
rect 34725 556 34791 559
rect 35973 556 36039 559
rect 37221 556 37287 559
rect 38469 556 38535 559
rect 39717 556 39783 559
rect 40965 556 41031 559
rect 0 554 41310 556
rect 0 498 2282 554
rect 2338 498 3530 554
rect 3586 498 4778 554
rect 4834 498 6026 554
rect 6082 498 7274 554
rect 7330 498 8522 554
rect 8578 498 9770 554
rect 9826 498 11018 554
rect 11074 498 12266 554
rect 12322 498 13514 554
rect 13570 498 14762 554
rect 14818 498 16010 554
rect 16066 498 17258 554
rect 17314 498 18506 554
rect 18562 498 19754 554
rect 19810 498 21002 554
rect 21058 498 22250 554
rect 22306 498 23498 554
rect 23554 498 24746 554
rect 24802 498 25994 554
rect 26050 498 27242 554
rect 27298 498 28490 554
rect 28546 498 29738 554
rect 29794 498 30986 554
rect 31042 498 32234 554
rect 32290 498 33482 554
rect 33538 498 34730 554
rect 34786 498 35978 554
rect 36034 498 37226 554
rect 37282 498 38474 554
rect 38530 498 39722 554
rect 39778 498 40970 554
rect 41026 498 41310 554
rect 0 496 41310 498
rect 2277 493 2343 496
rect 3525 493 3591 496
rect 4773 493 4839 496
rect 6021 493 6087 496
rect 7269 493 7335 496
rect 8517 493 8583 496
rect 9765 493 9831 496
rect 11013 493 11079 496
rect 12261 493 12327 496
rect 13509 493 13575 496
rect 14757 493 14823 496
rect 16005 493 16071 496
rect 17253 493 17319 496
rect 18501 493 18567 496
rect 19749 493 19815 496
rect 20997 493 21063 496
rect 22245 493 22311 496
rect 23493 493 23559 496
rect 24741 493 24807 496
rect 25989 493 26055 496
rect 27237 493 27303 496
rect 28485 493 28551 496
rect 29733 493 29799 496
rect 30981 493 31047 496
rect 32229 493 32295 496
rect 33477 493 33543 496
rect 34725 493 34791 496
rect 35973 493 36039 496
rect 37221 493 37287 496
rect 38469 493 38535 496
rect 39717 493 39783 496
rect 40965 493 41031 496
rect 1653 432 1719 435
rect 2901 432 2967 435
rect 4149 432 4215 435
rect 5397 432 5463 435
rect 6645 432 6711 435
rect 7893 432 7959 435
rect 9141 432 9207 435
rect 10389 432 10455 435
rect 11637 432 11703 435
rect 12885 432 12951 435
rect 14133 432 14199 435
rect 15381 432 15447 435
rect 16629 432 16695 435
rect 17877 432 17943 435
rect 19125 432 19191 435
rect 20373 432 20439 435
rect 21621 432 21687 435
rect 22869 432 22935 435
rect 24117 432 24183 435
rect 25365 432 25431 435
rect 26613 432 26679 435
rect 27861 432 27927 435
rect 29109 432 29175 435
rect 30357 432 30423 435
rect 31605 432 31671 435
rect 32853 432 32919 435
rect 34101 432 34167 435
rect 35349 432 35415 435
rect 36597 432 36663 435
rect 37845 432 37911 435
rect 39093 432 39159 435
rect 40341 432 40407 435
rect 0 430 41310 432
rect 0 374 1658 430
rect 1714 374 2906 430
rect 2962 374 4154 430
rect 4210 374 5402 430
rect 5458 374 6650 430
rect 6706 374 7898 430
rect 7954 374 9146 430
rect 9202 374 10394 430
rect 10450 374 11642 430
rect 11698 374 12890 430
rect 12946 374 14138 430
rect 14194 374 15386 430
rect 15442 374 16634 430
rect 16690 374 17882 430
rect 17938 374 19130 430
rect 19186 374 20378 430
rect 20434 374 21626 430
rect 21682 374 22874 430
rect 22930 374 24122 430
rect 24178 374 25370 430
rect 25426 374 26618 430
rect 26674 374 27866 430
rect 27922 374 29114 430
rect 29170 374 30362 430
rect 30418 374 31610 430
rect 31666 374 32858 430
rect 32914 374 34106 430
rect 34162 374 35354 430
rect 35410 374 36602 430
rect 36658 374 37850 430
rect 37906 374 39098 430
rect 39154 374 40346 430
rect 40402 374 41310 430
rect 0 372 41310 374
rect 1653 369 1719 372
rect 2901 369 2967 372
rect 4149 369 4215 372
rect 5397 369 5463 372
rect 6645 369 6711 372
rect 7893 369 7959 372
rect 9141 369 9207 372
rect 10389 369 10455 372
rect 11637 369 11703 372
rect 12885 369 12951 372
rect 14133 369 14199 372
rect 15381 369 15447 372
rect 16629 369 16695 372
rect 17877 369 17943 372
rect 19125 369 19191 372
rect 20373 369 20439 372
rect 21621 369 21687 372
rect 22869 369 22935 372
rect 24117 369 24183 372
rect 25365 369 25431 372
rect 26613 369 26679 372
rect 27861 369 27927 372
rect 29109 369 29175 372
rect 30357 369 30423 372
rect 31605 369 31671 372
rect 32853 369 32919 372
rect 34101 369 34167 372
rect 35349 369 35415 372
rect 36597 369 36663 372
rect 37845 369 37911 372
rect 39093 369 39159 372
rect 40341 369 40407 372
rect 1435 278 1501 281
rect 2495 278 2561 281
rect 1435 276 2561 278
rect 1435 220 1440 276
rect 1496 220 2500 276
rect 2556 220 2561 276
rect 1435 218 2561 220
rect 1435 215 1501 218
rect 2495 215 2561 218
rect 2683 278 2749 281
rect 3743 278 3809 281
rect 2683 276 3809 278
rect 2683 220 2688 276
rect 2744 220 3748 276
rect 3804 220 3809 276
rect 2683 218 3809 220
rect 2683 215 2749 218
rect 3743 215 3809 218
rect 3931 278 3997 281
rect 4991 278 5057 281
rect 3931 276 5057 278
rect 3931 220 3936 276
rect 3992 220 4996 276
rect 5052 220 5057 276
rect 3931 218 5057 220
rect 3931 215 3997 218
rect 4991 215 5057 218
rect 5179 278 5245 281
rect 6239 278 6305 281
rect 5179 276 6305 278
rect 5179 220 5184 276
rect 5240 220 6244 276
rect 6300 220 6305 276
rect 5179 218 6305 220
rect 5179 215 5245 218
rect 6239 215 6305 218
rect 6427 278 6493 281
rect 7487 278 7553 281
rect 6427 276 7553 278
rect 6427 220 6432 276
rect 6488 220 7492 276
rect 7548 220 7553 276
rect 6427 218 7553 220
rect 6427 215 6493 218
rect 7487 215 7553 218
rect 7675 278 7741 281
rect 8735 278 8801 281
rect 7675 276 8801 278
rect 7675 220 7680 276
rect 7736 220 8740 276
rect 8796 220 8801 276
rect 7675 218 8801 220
rect 7675 215 7741 218
rect 8735 215 8801 218
rect 8923 278 8989 281
rect 9983 278 10049 281
rect 8923 276 10049 278
rect 8923 220 8928 276
rect 8984 220 9988 276
rect 10044 220 10049 276
rect 8923 218 10049 220
rect 8923 215 8989 218
rect 9983 215 10049 218
rect 10171 278 10237 281
rect 11231 278 11297 281
rect 10171 276 11297 278
rect 10171 220 10176 276
rect 10232 220 11236 276
rect 11292 220 11297 276
rect 10171 218 11297 220
rect 10171 215 10237 218
rect 11231 215 11297 218
rect 11419 278 11485 281
rect 12479 278 12545 281
rect 11419 276 12545 278
rect 11419 220 11424 276
rect 11480 220 12484 276
rect 12540 220 12545 276
rect 11419 218 12545 220
rect 11419 215 11485 218
rect 12479 215 12545 218
rect 12667 278 12733 281
rect 13727 278 13793 281
rect 12667 276 13793 278
rect 12667 220 12672 276
rect 12728 220 13732 276
rect 13788 220 13793 276
rect 12667 218 13793 220
rect 12667 215 12733 218
rect 13727 215 13793 218
rect 13915 278 13981 281
rect 14975 278 15041 281
rect 13915 276 15041 278
rect 13915 220 13920 276
rect 13976 220 14980 276
rect 15036 220 15041 276
rect 13915 218 15041 220
rect 13915 215 13981 218
rect 14975 215 15041 218
rect 15163 278 15229 281
rect 16223 278 16289 281
rect 15163 276 16289 278
rect 15163 220 15168 276
rect 15224 220 16228 276
rect 16284 220 16289 276
rect 15163 218 16289 220
rect 15163 215 15229 218
rect 16223 215 16289 218
rect 16411 278 16477 281
rect 17471 278 17537 281
rect 16411 276 17537 278
rect 16411 220 16416 276
rect 16472 220 17476 276
rect 17532 220 17537 276
rect 16411 218 17537 220
rect 16411 215 16477 218
rect 17471 215 17537 218
rect 17659 278 17725 281
rect 18719 278 18785 281
rect 17659 276 18785 278
rect 17659 220 17664 276
rect 17720 220 18724 276
rect 18780 220 18785 276
rect 17659 218 18785 220
rect 17659 215 17725 218
rect 18719 215 18785 218
rect 18907 278 18973 281
rect 19967 278 20033 281
rect 18907 276 20033 278
rect 18907 220 18912 276
rect 18968 220 19972 276
rect 20028 220 20033 276
rect 18907 218 20033 220
rect 18907 215 18973 218
rect 19967 215 20033 218
rect 20155 278 20221 281
rect 21215 278 21281 281
rect 20155 276 21281 278
rect 20155 220 20160 276
rect 20216 220 21220 276
rect 21276 220 21281 276
rect 20155 218 21281 220
rect 20155 215 20221 218
rect 21215 215 21281 218
rect 21403 278 21469 281
rect 22463 278 22529 281
rect 21403 276 22529 278
rect 21403 220 21408 276
rect 21464 220 22468 276
rect 22524 220 22529 276
rect 21403 218 22529 220
rect 21403 215 21469 218
rect 22463 215 22529 218
rect 22651 278 22717 281
rect 23711 278 23777 281
rect 22651 276 23777 278
rect 22651 220 22656 276
rect 22712 220 23716 276
rect 23772 220 23777 276
rect 22651 218 23777 220
rect 22651 215 22717 218
rect 23711 215 23777 218
rect 23899 278 23965 281
rect 24959 278 25025 281
rect 23899 276 25025 278
rect 23899 220 23904 276
rect 23960 220 24964 276
rect 25020 220 25025 276
rect 23899 218 25025 220
rect 23899 215 23965 218
rect 24959 215 25025 218
rect 25147 278 25213 281
rect 26207 278 26273 281
rect 25147 276 26273 278
rect 25147 220 25152 276
rect 25208 220 26212 276
rect 26268 220 26273 276
rect 25147 218 26273 220
rect 25147 215 25213 218
rect 26207 215 26273 218
rect 26395 278 26461 281
rect 27455 278 27521 281
rect 26395 276 27521 278
rect 26395 220 26400 276
rect 26456 220 27460 276
rect 27516 220 27521 276
rect 26395 218 27521 220
rect 26395 215 26461 218
rect 27455 215 27521 218
rect 27643 278 27709 281
rect 28703 278 28769 281
rect 27643 276 28769 278
rect 27643 220 27648 276
rect 27704 220 28708 276
rect 28764 220 28769 276
rect 27643 218 28769 220
rect 27643 215 27709 218
rect 28703 215 28769 218
rect 28891 278 28957 281
rect 29951 278 30017 281
rect 28891 276 30017 278
rect 28891 220 28896 276
rect 28952 220 29956 276
rect 30012 220 30017 276
rect 28891 218 30017 220
rect 28891 215 28957 218
rect 29951 215 30017 218
rect 30139 278 30205 281
rect 31199 278 31265 281
rect 30139 276 31265 278
rect 30139 220 30144 276
rect 30200 220 31204 276
rect 31260 220 31265 276
rect 30139 218 31265 220
rect 30139 215 30205 218
rect 31199 215 31265 218
rect 31387 278 31453 281
rect 32447 278 32513 281
rect 31387 276 32513 278
rect 31387 220 31392 276
rect 31448 220 32452 276
rect 32508 220 32513 276
rect 31387 218 32513 220
rect 31387 215 31453 218
rect 32447 215 32513 218
rect 32635 278 32701 281
rect 33695 278 33761 281
rect 32635 276 33761 278
rect 32635 220 32640 276
rect 32696 220 33700 276
rect 33756 220 33761 276
rect 32635 218 33761 220
rect 32635 215 32701 218
rect 33695 215 33761 218
rect 33883 278 33949 281
rect 34943 278 35009 281
rect 33883 276 35009 278
rect 33883 220 33888 276
rect 33944 220 34948 276
rect 35004 220 35009 276
rect 33883 218 35009 220
rect 33883 215 33949 218
rect 34943 215 35009 218
rect 35131 278 35197 281
rect 36191 278 36257 281
rect 35131 276 36257 278
rect 35131 220 35136 276
rect 35192 220 36196 276
rect 36252 220 36257 276
rect 35131 218 36257 220
rect 35131 215 35197 218
rect 36191 215 36257 218
rect 36379 278 36445 281
rect 37439 278 37505 281
rect 36379 276 37505 278
rect 36379 220 36384 276
rect 36440 220 37444 276
rect 37500 220 37505 276
rect 36379 218 37505 220
rect 36379 215 36445 218
rect 37439 215 37505 218
rect 37627 278 37693 281
rect 38687 278 38753 281
rect 37627 276 38753 278
rect 37627 220 37632 276
rect 37688 220 38692 276
rect 38748 220 38753 276
rect 37627 218 38753 220
rect 37627 215 37693 218
rect 38687 215 38753 218
rect 38875 278 38941 281
rect 39935 278 40001 281
rect 38875 276 40001 278
rect 38875 220 38880 276
rect 38936 220 39940 276
rect 39996 220 40001 276
rect 38875 218 40001 220
rect 38875 215 38941 218
rect 39935 215 40001 218
rect 40123 278 40189 281
rect 41183 278 41249 281
rect 40123 276 41249 278
rect 40123 220 40128 276
rect 40184 220 41188 276
rect 41244 220 41249 276
rect 40123 218 41249 220
rect 40123 215 40189 218
rect 41183 215 41249 218
rect 1899 154 1965 157
rect 2031 154 2097 157
rect 1899 152 2097 154
rect 1899 96 1904 152
rect 1960 96 2036 152
rect 2092 96 2097 152
rect 1899 94 2097 96
rect 1899 91 1965 94
rect 2031 91 2097 94
rect 3147 154 3213 157
rect 3279 154 3345 157
rect 3147 152 3345 154
rect 3147 96 3152 152
rect 3208 96 3284 152
rect 3340 96 3345 152
rect 3147 94 3345 96
rect 3147 91 3213 94
rect 3279 91 3345 94
rect 4395 154 4461 157
rect 4527 154 4593 157
rect 4395 152 4593 154
rect 4395 96 4400 152
rect 4456 96 4532 152
rect 4588 96 4593 152
rect 4395 94 4593 96
rect 4395 91 4461 94
rect 4527 91 4593 94
rect 5643 154 5709 157
rect 5775 154 5841 157
rect 5643 152 5841 154
rect 5643 96 5648 152
rect 5704 96 5780 152
rect 5836 96 5841 152
rect 5643 94 5841 96
rect 5643 91 5709 94
rect 5775 91 5841 94
rect 6891 154 6957 157
rect 7023 154 7089 157
rect 6891 152 7089 154
rect 6891 96 6896 152
rect 6952 96 7028 152
rect 7084 96 7089 152
rect 6891 94 7089 96
rect 6891 91 6957 94
rect 7023 91 7089 94
rect 8139 154 8205 157
rect 8271 154 8337 157
rect 8139 152 8337 154
rect 8139 96 8144 152
rect 8200 96 8276 152
rect 8332 96 8337 152
rect 8139 94 8337 96
rect 8139 91 8205 94
rect 8271 91 8337 94
rect 9387 154 9453 157
rect 9519 154 9585 157
rect 9387 152 9585 154
rect 9387 96 9392 152
rect 9448 96 9524 152
rect 9580 96 9585 152
rect 9387 94 9585 96
rect 9387 91 9453 94
rect 9519 91 9585 94
rect 10635 154 10701 157
rect 10767 154 10833 157
rect 10635 152 10833 154
rect 10635 96 10640 152
rect 10696 96 10772 152
rect 10828 96 10833 152
rect 10635 94 10833 96
rect 10635 91 10701 94
rect 10767 91 10833 94
rect 11883 154 11949 157
rect 12015 154 12081 157
rect 11883 152 12081 154
rect 11883 96 11888 152
rect 11944 96 12020 152
rect 12076 96 12081 152
rect 11883 94 12081 96
rect 11883 91 11949 94
rect 12015 91 12081 94
rect 13131 154 13197 157
rect 13263 154 13329 157
rect 13131 152 13329 154
rect 13131 96 13136 152
rect 13192 96 13268 152
rect 13324 96 13329 152
rect 13131 94 13329 96
rect 13131 91 13197 94
rect 13263 91 13329 94
rect 14379 154 14445 157
rect 14511 154 14577 157
rect 14379 152 14577 154
rect 14379 96 14384 152
rect 14440 96 14516 152
rect 14572 96 14577 152
rect 14379 94 14577 96
rect 14379 91 14445 94
rect 14511 91 14577 94
rect 15627 154 15693 157
rect 15759 154 15825 157
rect 15627 152 15825 154
rect 15627 96 15632 152
rect 15688 96 15764 152
rect 15820 96 15825 152
rect 15627 94 15825 96
rect 15627 91 15693 94
rect 15759 91 15825 94
rect 16875 154 16941 157
rect 17007 154 17073 157
rect 16875 152 17073 154
rect 16875 96 16880 152
rect 16936 96 17012 152
rect 17068 96 17073 152
rect 16875 94 17073 96
rect 16875 91 16941 94
rect 17007 91 17073 94
rect 18123 154 18189 157
rect 18255 154 18321 157
rect 18123 152 18321 154
rect 18123 96 18128 152
rect 18184 96 18260 152
rect 18316 96 18321 152
rect 18123 94 18321 96
rect 18123 91 18189 94
rect 18255 91 18321 94
rect 19371 154 19437 157
rect 19503 154 19569 157
rect 19371 152 19569 154
rect 19371 96 19376 152
rect 19432 96 19508 152
rect 19564 96 19569 152
rect 19371 94 19569 96
rect 19371 91 19437 94
rect 19503 91 19569 94
rect 20619 154 20685 157
rect 20751 154 20817 157
rect 20619 152 20817 154
rect 20619 96 20624 152
rect 20680 96 20756 152
rect 20812 96 20817 152
rect 20619 94 20817 96
rect 20619 91 20685 94
rect 20751 91 20817 94
rect 21867 154 21933 157
rect 21999 154 22065 157
rect 21867 152 22065 154
rect 21867 96 21872 152
rect 21928 96 22004 152
rect 22060 96 22065 152
rect 21867 94 22065 96
rect 21867 91 21933 94
rect 21999 91 22065 94
rect 23115 154 23181 157
rect 23247 154 23313 157
rect 23115 152 23313 154
rect 23115 96 23120 152
rect 23176 96 23252 152
rect 23308 96 23313 152
rect 23115 94 23313 96
rect 23115 91 23181 94
rect 23247 91 23313 94
rect 24363 154 24429 157
rect 24495 154 24561 157
rect 24363 152 24561 154
rect 24363 96 24368 152
rect 24424 96 24500 152
rect 24556 96 24561 152
rect 24363 94 24561 96
rect 24363 91 24429 94
rect 24495 91 24561 94
rect 25611 154 25677 157
rect 25743 154 25809 157
rect 25611 152 25809 154
rect 25611 96 25616 152
rect 25672 96 25748 152
rect 25804 96 25809 152
rect 25611 94 25809 96
rect 25611 91 25677 94
rect 25743 91 25809 94
rect 26859 154 26925 157
rect 26991 154 27057 157
rect 26859 152 27057 154
rect 26859 96 26864 152
rect 26920 96 26996 152
rect 27052 96 27057 152
rect 26859 94 27057 96
rect 26859 91 26925 94
rect 26991 91 27057 94
rect 28107 154 28173 157
rect 28239 154 28305 157
rect 28107 152 28305 154
rect 28107 96 28112 152
rect 28168 96 28244 152
rect 28300 96 28305 152
rect 28107 94 28305 96
rect 28107 91 28173 94
rect 28239 91 28305 94
rect 29355 154 29421 157
rect 29487 154 29553 157
rect 29355 152 29553 154
rect 29355 96 29360 152
rect 29416 96 29492 152
rect 29548 96 29553 152
rect 29355 94 29553 96
rect 29355 91 29421 94
rect 29487 91 29553 94
rect 30603 154 30669 157
rect 30735 154 30801 157
rect 30603 152 30801 154
rect 30603 96 30608 152
rect 30664 96 30740 152
rect 30796 96 30801 152
rect 30603 94 30801 96
rect 30603 91 30669 94
rect 30735 91 30801 94
rect 31851 154 31917 157
rect 31983 154 32049 157
rect 31851 152 32049 154
rect 31851 96 31856 152
rect 31912 96 31988 152
rect 32044 96 32049 152
rect 31851 94 32049 96
rect 31851 91 31917 94
rect 31983 91 32049 94
rect 33099 154 33165 157
rect 33231 154 33297 157
rect 33099 152 33297 154
rect 33099 96 33104 152
rect 33160 96 33236 152
rect 33292 96 33297 152
rect 33099 94 33297 96
rect 33099 91 33165 94
rect 33231 91 33297 94
rect 34347 154 34413 157
rect 34479 154 34545 157
rect 34347 152 34545 154
rect 34347 96 34352 152
rect 34408 96 34484 152
rect 34540 96 34545 152
rect 34347 94 34545 96
rect 34347 91 34413 94
rect 34479 91 34545 94
rect 35595 154 35661 157
rect 35727 154 35793 157
rect 35595 152 35793 154
rect 35595 96 35600 152
rect 35656 96 35732 152
rect 35788 96 35793 152
rect 35595 94 35793 96
rect 35595 91 35661 94
rect 35727 91 35793 94
rect 36843 154 36909 157
rect 36975 154 37041 157
rect 36843 152 37041 154
rect 36843 96 36848 152
rect 36904 96 36980 152
rect 37036 96 37041 152
rect 36843 94 37041 96
rect 36843 91 36909 94
rect 36975 91 37041 94
rect 38091 154 38157 157
rect 38223 154 38289 157
rect 38091 152 38289 154
rect 38091 96 38096 152
rect 38152 96 38228 152
rect 38284 96 38289 152
rect 38091 94 38289 96
rect 38091 91 38157 94
rect 38223 91 38289 94
rect 39339 154 39405 157
rect 39471 154 39537 157
rect 39339 152 39537 154
rect 39339 96 39344 152
rect 39400 96 39476 152
rect 39532 96 39537 152
rect 39339 94 39537 96
rect 39339 91 39405 94
rect 39471 91 39537 94
rect 40587 154 40653 157
rect 40719 154 40785 157
rect 40587 152 40785 154
rect 40587 96 40592 152
rect 40648 96 40724 152
rect 40780 96 40785 152
rect 40587 94 40785 96
rect 40587 91 40653 94
rect 40719 91 40785 94
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_0
timestamp 1666199351
transform -1 0 6366 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_1
timestamp 1666199351
transform 1 0 5118 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_2
timestamp 1666199351
transform -1 0 5118 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_3
timestamp 1666199351
transform 1 0 3870 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_4
timestamp 1666199351
transform -1 0 3870 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_5
timestamp 1666199351
transform 1 0 2622 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_6
timestamp 1666199351
transform -1 0 2622 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_7
timestamp 1666199351
transform 1 0 1374 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_8
timestamp 1666199351
transform -1 0 11358 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_9
timestamp 1666199351
transform 1 0 10110 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_10
timestamp 1666199351
transform -1 0 10110 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_11
timestamp 1666199351
transform 1 0 8862 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_12
timestamp 1666199351
transform -1 0 8862 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_13
timestamp 1666199351
transform 1 0 7614 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_14
timestamp 1666199351
transform -1 0 7614 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_15
timestamp 1666199351
transform 1 0 6366 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_16
timestamp 1666199351
transform -1 0 16350 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_17
timestamp 1666199351
transform 1 0 15102 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_18
timestamp 1666199351
transform -1 0 15102 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_19
timestamp 1666199351
transform 1 0 13854 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_20
timestamp 1666199351
transform -1 0 13854 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_21
timestamp 1666199351
transform 1 0 12606 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_22
timestamp 1666199351
transform -1 0 12606 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_23
timestamp 1666199351
transform 1 0 11358 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_24
timestamp 1666199351
transform -1 0 21342 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_25
timestamp 1666199351
transform 1 0 20094 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_26
timestamp 1666199351
transform -1 0 20094 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_27
timestamp 1666199351
transform 1 0 18846 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_28
timestamp 1666199351
transform -1 0 18846 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_29
timestamp 1666199351
transform 1 0 17598 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_30
timestamp 1666199351
transform -1 0 17598 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_31
timestamp 1666199351
transform 1 0 16350 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_32
timestamp 1666199351
transform -1 0 26334 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_33
timestamp 1666199351
transform 1 0 25086 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_34
timestamp 1666199351
transform -1 0 25086 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_35
timestamp 1666199351
transform 1 0 23838 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_36
timestamp 1666199351
transform -1 0 23838 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_37
timestamp 1666199351
transform 1 0 22590 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_38
timestamp 1666199351
transform -1 0 22590 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_39
timestamp 1666199351
transform 1 0 21342 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_40
timestamp 1666199351
transform -1 0 31326 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_41
timestamp 1666199351
transform 1 0 30078 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_42
timestamp 1666199351
transform -1 0 30078 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_43
timestamp 1666199351
transform 1 0 28830 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_44
timestamp 1666199351
transform -1 0 28830 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_45
timestamp 1666199351
transform 1 0 27582 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_46
timestamp 1666199351
transform -1 0 27582 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_47
timestamp 1666199351
transform 1 0 26334 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_48
timestamp 1666199351
transform -1 0 36318 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_49
timestamp 1666199351
transform 1 0 35070 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_50
timestamp 1666199351
transform -1 0 35070 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_51
timestamp 1666199351
transform 1 0 33822 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_52
timestamp 1666199351
transform -1 0 33822 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_53
timestamp 1666199351
transform 1 0 32574 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_54
timestamp 1666199351
transform -1 0 32574 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_55
timestamp 1666199351
transform 1 0 31326 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_56
timestamp 1666199351
transform -1 0 41310 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_57
timestamp 1666199351
transform 1 0 40062 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_58
timestamp 1666199351
transform -1 0 40062 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_59
timestamp 1666199351
transform 1 0 38814 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_60
timestamp 1666199351
transform -1 0 38814 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_61
timestamp 1666199351
transform 1 0 37566 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_62
timestamp 1666199351
transform -1 0 37566 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_63
timestamp 1666199351
transform 1 0 36318 0 1 620
box 65 0 675 1316
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_0
timestamp 1666199351
transform 1 0 6021 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_1
timestamp 1666199351
transform 1 0 5397 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_2
timestamp 1666199351
transform 1 0 4773 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_3
timestamp 1666199351
transform 1 0 4149 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_4
timestamp 1666199351
transform 1 0 3525 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_5
timestamp 1666199351
transform 1 0 2901 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_6
timestamp 1666199351
transform 1 0 2277 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_7
timestamp 1666199351
transform 1 0 1653 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_8
timestamp 1666199351
transform 1 0 11013 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_9
timestamp 1666199351
transform 1 0 10389 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_10
timestamp 1666199351
transform 1 0 9765 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_11
timestamp 1666199351
transform 1 0 9141 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_12
timestamp 1666199351
transform 1 0 8517 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_13
timestamp 1666199351
transform 1 0 7893 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_14
timestamp 1666199351
transform 1 0 7269 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_15
timestamp 1666199351
transform 1 0 6645 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_16
timestamp 1666199351
transform 1 0 12261 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_17
timestamp 1666199351
transform 1 0 11637 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_18
timestamp 1666199351
transform 1 0 16005 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_19
timestamp 1666199351
transform 1 0 15381 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_20
timestamp 1666199351
transform 1 0 14757 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_21
timestamp 1666199351
transform 1 0 14133 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_22
timestamp 1666199351
transform 1 0 13509 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_23
timestamp 1666199351
transform 1 0 12885 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_24
timestamp 1666199351
transform 1 0 20997 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_25
timestamp 1666199351
transform 1 0 20373 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_26
timestamp 1666199351
transform 1 0 19749 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_27
timestamp 1666199351
transform 1 0 19125 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_28
timestamp 1666199351
transform 1 0 18501 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_29
timestamp 1666199351
transform 1 0 17877 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_30
timestamp 1666199351
transform 1 0 17253 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_31
timestamp 1666199351
transform 1 0 16629 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_32
timestamp 1666199351
transform 1 0 25989 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_33
timestamp 1666199351
transform 1 0 25365 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_34
timestamp 1666199351
transform 1 0 24741 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_35
timestamp 1666199351
transform 1 0 24117 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_36
timestamp 1666199351
transform 1 0 23493 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_37
timestamp 1666199351
transform 1 0 22869 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_38
timestamp 1666199351
transform 1 0 22245 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_39
timestamp 1666199351
transform 1 0 21621 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_40
timestamp 1666199351
transform 1 0 30981 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_41
timestamp 1666199351
transform 1 0 30357 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_42
timestamp 1666199351
transform 1 0 29733 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_43
timestamp 1666199351
transform 1 0 29109 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_44
timestamp 1666199351
transform 1 0 28485 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_45
timestamp 1666199351
transform 1 0 27861 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_46
timestamp 1666199351
transform 1 0 27237 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_47
timestamp 1666199351
transform 1 0 26613 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_48
timestamp 1666199351
transform 1 0 33477 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_49
timestamp 1666199351
transform 1 0 32853 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_50
timestamp 1666199351
transform 1 0 32229 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_51
timestamp 1666199351
transform 1 0 31605 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_52
timestamp 1666199351
transform 1 0 35973 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_53
timestamp 1666199351
transform 1 0 35349 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_54
timestamp 1666199351
transform 1 0 34725 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_55
timestamp 1666199351
transform 1 0 34101 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_56
timestamp 1666199351
transform 1 0 40965 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_57
timestamp 1666199351
transform 1 0 40341 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_58
timestamp 1666199351
transform 1 0 39717 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_59
timestamp 1666199351
transform 1 0 39093 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_60
timestamp 1666199351
transform 1 0 38469 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_61
timestamp 1666199351
transform 1 0 37845 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_62
timestamp 1666199351
transform 1 0 37221 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_24  sky130_sram_1kbyte_1rw1r_32x256_8_contact_24_63
timestamp 1666199351
transform 1 0 36597 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_0
timestamp 1666199351
transform 1 0 6025 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_1
timestamp 1666199351
transform 1 0 5401 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_2
timestamp 1666199351
transform 1 0 4777 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_3
timestamp 1666199351
transform 1 0 4153 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_4
timestamp 1666199351
transform 1 0 3529 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_5
timestamp 1666199351
transform 1 0 2905 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_6
timestamp 1666199351
transform 1 0 2281 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_7
timestamp 1666199351
transform 1 0 1657 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_8
timestamp 1666199351
transform 1 0 11017 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_9
timestamp 1666199351
transform 1 0 10393 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_10
timestamp 1666199351
transform 1 0 9769 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_11
timestamp 1666199351
transform 1 0 9145 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_12
timestamp 1666199351
transform 1 0 8521 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_13
timestamp 1666199351
transform 1 0 7897 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_14
timestamp 1666199351
transform 1 0 7273 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_15
timestamp 1666199351
transform 1 0 6649 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_16
timestamp 1666199351
transform 1 0 12265 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_17
timestamp 1666199351
transform 1 0 11641 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_18
timestamp 1666199351
transform 1 0 16009 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_19
timestamp 1666199351
transform 1 0 15385 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_20
timestamp 1666199351
transform 1 0 14761 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_21
timestamp 1666199351
transform 1 0 14137 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_22
timestamp 1666199351
transform 1 0 13513 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_23
timestamp 1666199351
transform 1 0 12889 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_24
timestamp 1666199351
transform 1 0 21001 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_25
timestamp 1666199351
transform 1 0 20377 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_26
timestamp 1666199351
transform 1 0 19753 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_27
timestamp 1666199351
transform 1 0 19129 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_28
timestamp 1666199351
transform 1 0 18505 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_29
timestamp 1666199351
transform 1 0 17881 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_30
timestamp 1666199351
transform 1 0 17257 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_31
timestamp 1666199351
transform 1 0 16633 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_32
timestamp 1666199351
transform 1 0 25993 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_33
timestamp 1666199351
transform 1 0 25369 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_34
timestamp 1666199351
transform 1 0 24745 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_35
timestamp 1666199351
transform 1 0 24121 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_36
timestamp 1666199351
transform 1 0 23497 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_37
timestamp 1666199351
transform 1 0 22873 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_38
timestamp 1666199351
transform 1 0 22249 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_39
timestamp 1666199351
transform 1 0 21625 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_40
timestamp 1666199351
transform 1 0 30985 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_41
timestamp 1666199351
transform 1 0 30361 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_42
timestamp 1666199351
transform 1 0 29737 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_43
timestamp 1666199351
transform 1 0 29113 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_44
timestamp 1666199351
transform 1 0 28489 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_45
timestamp 1666199351
transform 1 0 27865 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_46
timestamp 1666199351
transform 1 0 27241 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_47
timestamp 1666199351
transform 1 0 26617 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_48
timestamp 1666199351
transform 1 0 33481 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_49
timestamp 1666199351
transform 1 0 32857 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_50
timestamp 1666199351
transform 1 0 32233 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_51
timestamp 1666199351
transform 1 0 31609 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_52
timestamp 1666199351
transform 1 0 35977 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_53
timestamp 1666199351
transform 1 0 35353 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_54
timestamp 1666199351
transform 1 0 34729 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_55
timestamp 1666199351
transform 1 0 34105 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_56
timestamp 1666199351
transform 1 0 40969 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_57
timestamp 1666199351
transform 1 0 40345 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_58
timestamp 1666199351
transform 1 0 39721 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_59
timestamp 1666199351
transform 1 0 39097 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_60
timestamp 1666199351
transform 1 0 38473 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_61
timestamp 1666199351
transform 1 0 37849 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_62
timestamp 1666199351
transform 1 0 37225 0 1 493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_25  sky130_sram_1kbyte_1rw1r_32x256_8_contact_25_63
timestamp 1666199351
transform 1 0 36601 0 1 369
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_0
timestamp 1666199351
transform 1 0 3280 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_1
timestamp 1666199351
transform 1 0 3744 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_2
timestamp 1666199351
transform 1 0 3148 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_3
timestamp 1666199351
transform 1 0 2684 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_4
timestamp 1666199351
transform 1 0 2032 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_5
timestamp 1666199351
transform 1 0 2496 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_6
timestamp 1666199351
transform 1 0 1900 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_7
timestamp 1666199351
transform 1 0 1436 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_8
timestamp 1666199351
transform 1 0 5776 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_9
timestamp 1666199351
transform 1 0 6240 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_10
timestamp 1666199351
transform 1 0 5644 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_11
timestamp 1666199351
transform 1 0 5180 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_12
timestamp 1666199351
transform 1 0 6022 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_13
timestamp 1666199351
transform 1 0 5398 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_14
timestamp 1666199351
transform 1 0 4774 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_15
timestamp 1666199351
transform 1 0 4150 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_16
timestamp 1666199351
transform 1 0 3526 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_17
timestamp 1666199351
transform 1 0 2902 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_18
timestamp 1666199351
transform 1 0 2278 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_19
timestamp 1666199351
transform 1 0 1654 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_20
timestamp 1666199351
transform 1 0 4528 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_21
timestamp 1666199351
transform 1 0 4992 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_22
timestamp 1666199351
transform 1 0 4396 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_23
timestamp 1666199351
transform 1 0 3932 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_24
timestamp 1666199351
transform 1 0 11014 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_25
timestamp 1666199351
transform 1 0 10390 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_26
timestamp 1666199351
transform 1 0 9766 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_27
timestamp 1666199351
transform 1 0 9142 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_28
timestamp 1666199351
transform 1 0 8518 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_29
timestamp 1666199351
transform 1 0 7894 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_30
timestamp 1666199351
transform 1 0 7270 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_31
timestamp 1666199351
transform 1 0 6646 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_32
timestamp 1666199351
transform 1 0 8272 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_33
timestamp 1666199351
transform 1 0 8736 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_34
timestamp 1666199351
transform 1 0 8140 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_35
timestamp 1666199351
transform 1 0 7676 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_36
timestamp 1666199351
transform 1 0 7024 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_37
timestamp 1666199351
transform 1 0 7488 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_38
timestamp 1666199351
transform 1 0 6892 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_39
timestamp 1666199351
transform 1 0 6428 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_40
timestamp 1666199351
transform 1 0 10768 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_41
timestamp 1666199351
transform 1 0 11232 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_42
timestamp 1666199351
transform 1 0 10636 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_43
timestamp 1666199351
transform 1 0 10172 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_44
timestamp 1666199351
transform 1 0 9520 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_45
timestamp 1666199351
transform 1 0 9984 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_46
timestamp 1666199351
transform 1 0 9388 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_47
timestamp 1666199351
transform 1 0 8924 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_48
timestamp 1666199351
transform 1 0 12262 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_49
timestamp 1666199351
transform 1 0 11638 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_50
timestamp 1666199351
transform 1 0 15760 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_51
timestamp 1666199351
transform 1 0 16224 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_52
timestamp 1666199351
transform 1 0 15628 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_53
timestamp 1666199351
transform 1 0 15164 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_54
timestamp 1666199351
transform 1 0 14512 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_55
timestamp 1666199351
transform 1 0 14976 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_56
timestamp 1666199351
transform 1 0 14380 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_57
timestamp 1666199351
transform 1 0 13916 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_58
timestamp 1666199351
transform 1 0 13264 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_59
timestamp 1666199351
transform 1 0 13728 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_60
timestamp 1666199351
transform 1 0 13132 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_61
timestamp 1666199351
transform 1 0 12668 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_62
timestamp 1666199351
transform 1 0 12016 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_63
timestamp 1666199351
transform 1 0 12480 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_64
timestamp 1666199351
transform 1 0 11884 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_65
timestamp 1666199351
transform 1 0 11420 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_66
timestamp 1666199351
transform 1 0 16006 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_67
timestamp 1666199351
transform 1 0 15382 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_68
timestamp 1666199351
transform 1 0 14758 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_69
timestamp 1666199351
transform 1 0 14134 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_70
timestamp 1666199351
transform 1 0 13510 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_71
timestamp 1666199351
transform 1 0 12886 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_72
timestamp 1666199351
transform 1 0 20998 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_73
timestamp 1666199351
transform 1 0 20374 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_74
timestamp 1666199351
transform 1 0 19750 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_75
timestamp 1666199351
transform 1 0 19126 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_76
timestamp 1666199351
transform 1 0 18502 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_77
timestamp 1666199351
transform 1 0 17878 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_78
timestamp 1666199351
transform 1 0 17254 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_79
timestamp 1666199351
transform 1 0 16630 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_80
timestamp 1666199351
transform 1 0 20752 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_81
timestamp 1666199351
transform 1 0 21216 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_82
timestamp 1666199351
transform 1 0 20620 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_83
timestamp 1666199351
transform 1 0 20156 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_84
timestamp 1666199351
transform 1 0 19504 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_85
timestamp 1666199351
transform 1 0 19968 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_86
timestamp 1666199351
transform 1 0 19372 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_87
timestamp 1666199351
transform 1 0 18908 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_88
timestamp 1666199351
transform 1 0 18256 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_89
timestamp 1666199351
transform 1 0 18720 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_90
timestamp 1666199351
transform 1 0 18124 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_91
timestamp 1666199351
transform 1 0 17660 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_92
timestamp 1666199351
transform 1 0 17008 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_93
timestamp 1666199351
transform 1 0 17472 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_94
timestamp 1666199351
transform 1 0 16876 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_95
timestamp 1666199351
transform 1 0 16412 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_96
timestamp 1666199351
transform 1 0 25990 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_97
timestamp 1666199351
transform 1 0 25366 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_98
timestamp 1666199351
transform 1 0 24742 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_99
timestamp 1666199351
transform 1 0 24118 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_100
timestamp 1666199351
transform 1 0 23494 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_101
timestamp 1666199351
transform 1 0 22870 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_102
timestamp 1666199351
transform 1 0 22246 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_103
timestamp 1666199351
transform 1 0 21622 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_104
timestamp 1666199351
transform 1 0 24496 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_105
timestamp 1666199351
transform 1 0 24960 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_106
timestamp 1666199351
transform 1 0 24364 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_107
timestamp 1666199351
transform 1 0 23900 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_108
timestamp 1666199351
transform 1 0 23248 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_109
timestamp 1666199351
transform 1 0 23712 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_110
timestamp 1666199351
transform 1 0 23116 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_111
timestamp 1666199351
transform 1 0 22652 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_112
timestamp 1666199351
transform 1 0 22000 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_113
timestamp 1666199351
transform 1 0 22464 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_114
timestamp 1666199351
transform 1 0 21868 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_115
timestamp 1666199351
transform 1 0 21404 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_116
timestamp 1666199351
transform 1 0 25744 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_117
timestamp 1666199351
transform 1 0 26208 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_118
timestamp 1666199351
transform 1 0 25612 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_119
timestamp 1666199351
transform 1 0 25148 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_120
timestamp 1666199351
transform 1 0 30982 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_121
timestamp 1666199351
transform 1 0 30358 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_122
timestamp 1666199351
transform 1 0 29734 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_123
timestamp 1666199351
transform 1 0 29110 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_124
timestamp 1666199351
transform 1 0 30736 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_125
timestamp 1666199351
transform 1 0 31200 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_126
timestamp 1666199351
transform 1 0 30604 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_127
timestamp 1666199351
transform 1 0 30140 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_128
timestamp 1666199351
transform 1 0 29488 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_129
timestamp 1666199351
transform 1 0 29952 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_130
timestamp 1666199351
transform 1 0 29356 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_131
timestamp 1666199351
transform 1 0 28892 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_132
timestamp 1666199351
transform 1 0 28240 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_133
timestamp 1666199351
transform 1 0 28704 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_134
timestamp 1666199351
transform 1 0 28108 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_135
timestamp 1666199351
transform 1 0 27644 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_136
timestamp 1666199351
transform 1 0 26992 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_137
timestamp 1666199351
transform 1 0 27456 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_138
timestamp 1666199351
transform 1 0 26860 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_139
timestamp 1666199351
transform 1 0 26396 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_140
timestamp 1666199351
transform 1 0 28486 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_141
timestamp 1666199351
transform 1 0 27862 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_142
timestamp 1666199351
transform 1 0 27238 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_143
timestamp 1666199351
transform 1 0 26614 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_144
timestamp 1666199351
transform 1 0 33478 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_145
timestamp 1666199351
transform 1 0 32854 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_146
timestamp 1666199351
transform 1 0 32230 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_147
timestamp 1666199351
transform 1 0 31606 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_148
timestamp 1666199351
transform 1 0 35974 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_149
timestamp 1666199351
transform 1 0 35350 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_150
timestamp 1666199351
transform 1 0 35728 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_151
timestamp 1666199351
transform 1 0 36192 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_152
timestamp 1666199351
transform 1 0 35596 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_153
timestamp 1666199351
transform 1 0 35132 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_154
timestamp 1666199351
transform 1 0 34480 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_155
timestamp 1666199351
transform 1 0 34944 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_156
timestamp 1666199351
transform 1 0 34348 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_157
timestamp 1666199351
transform 1 0 33884 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_158
timestamp 1666199351
transform 1 0 33232 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_159
timestamp 1666199351
transform 1 0 33696 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_160
timestamp 1666199351
transform 1 0 33100 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_161
timestamp 1666199351
transform 1 0 32636 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_162
timestamp 1666199351
transform 1 0 31984 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_163
timestamp 1666199351
transform 1 0 32448 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_164
timestamp 1666199351
transform 1 0 31852 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_165
timestamp 1666199351
transform 1 0 31388 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_166
timestamp 1666199351
transform 1 0 34726 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_167
timestamp 1666199351
transform 1 0 34102 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_168
timestamp 1666199351
transform 1 0 40720 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_169
timestamp 1666199351
transform 1 0 41184 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_170
timestamp 1666199351
transform 1 0 40588 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_171
timestamp 1666199351
transform 1 0 40124 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_172
timestamp 1666199351
transform 1 0 39472 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_173
timestamp 1666199351
transform 1 0 39936 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_174
timestamp 1666199351
transform 1 0 39340 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_175
timestamp 1666199351
transform 1 0 38876 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_176
timestamp 1666199351
transform 1 0 38224 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_177
timestamp 1666199351
transform 1 0 38688 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_178
timestamp 1666199351
transform 1 0 38092 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_179
timestamp 1666199351
transform 1 0 37628 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_180
timestamp 1666199351
transform 1 0 36976 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_181
timestamp 1666199351
transform 1 0 37440 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_182
timestamp 1666199351
transform 1 0 36844 0 1 92
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_183
timestamp 1666199351
transform 1 0 36380 0 1 216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_184
timestamp 1666199351
transform 1 0 40966 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_185
timestamp 1666199351
transform 1 0 40342 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_186
timestamp 1666199351
transform 1 0 39718 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_187
timestamp 1666199351
transform 1 0 39094 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_188
timestamp 1666199351
transform 1 0 38470 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_189
timestamp 1666199351
transform 1 0 37846 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_190
timestamp 1666199351
transform 1 0 37222 0 1 494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_26  sky130_sram_1kbyte_1rw1r_32x256_8_contact_26_191
timestamp 1666199351
transform 1 0 36598 0 1 370
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_0
timestamp 1666199351
transform 1 0 3279 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_1
timestamp 1666199351
transform 1 0 3743 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_2
timestamp 1666199351
transform 1 0 3147 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_3
timestamp 1666199351
transform 1 0 2683 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_4
timestamp 1666199351
transform 1 0 2031 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_5
timestamp 1666199351
transform 1 0 2495 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_6
timestamp 1666199351
transform 1 0 1899 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_7
timestamp 1666199351
transform 1 0 1435 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_8
timestamp 1666199351
transform 1 0 5775 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_9
timestamp 1666199351
transform 1 0 6239 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_10
timestamp 1666199351
transform 1 0 5643 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_11
timestamp 1666199351
transform 1 0 5179 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_12
timestamp 1666199351
transform 1 0 6021 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_13
timestamp 1666199351
transform 1 0 5397 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_14
timestamp 1666199351
transform 1 0 4773 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_15
timestamp 1666199351
transform 1 0 4149 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_16
timestamp 1666199351
transform 1 0 3525 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_17
timestamp 1666199351
transform 1 0 2901 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_18
timestamp 1666199351
transform 1 0 2277 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_19
timestamp 1666199351
transform 1 0 1653 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_20
timestamp 1666199351
transform 1 0 4527 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_21
timestamp 1666199351
transform 1 0 4991 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_22
timestamp 1666199351
transform 1 0 4395 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_23
timestamp 1666199351
transform 1 0 3931 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_24
timestamp 1666199351
transform 1 0 11013 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_25
timestamp 1666199351
transform 1 0 10389 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_26
timestamp 1666199351
transform 1 0 9765 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_27
timestamp 1666199351
transform 1 0 9141 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_28
timestamp 1666199351
transform 1 0 8517 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_29
timestamp 1666199351
transform 1 0 7893 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_30
timestamp 1666199351
transform 1 0 7269 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_31
timestamp 1666199351
transform 1 0 6645 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_32
timestamp 1666199351
transform 1 0 8271 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_33
timestamp 1666199351
transform 1 0 8735 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_34
timestamp 1666199351
transform 1 0 8139 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_35
timestamp 1666199351
transform 1 0 7675 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_36
timestamp 1666199351
transform 1 0 7023 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_37
timestamp 1666199351
transform 1 0 7487 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_38
timestamp 1666199351
transform 1 0 6891 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_39
timestamp 1666199351
transform 1 0 6427 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_40
timestamp 1666199351
transform 1 0 10767 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_41
timestamp 1666199351
transform 1 0 11231 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_42
timestamp 1666199351
transform 1 0 10635 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_43
timestamp 1666199351
transform 1 0 10171 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_44
timestamp 1666199351
transform 1 0 9519 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_45
timestamp 1666199351
transform 1 0 9983 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_46
timestamp 1666199351
transform 1 0 9387 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_47
timestamp 1666199351
transform 1 0 8923 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_48
timestamp 1666199351
transform 1 0 12261 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_49
timestamp 1666199351
transform 1 0 11637 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_50
timestamp 1666199351
transform 1 0 15759 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_51
timestamp 1666199351
transform 1 0 16223 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_52
timestamp 1666199351
transform 1 0 15627 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_53
timestamp 1666199351
transform 1 0 15163 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_54
timestamp 1666199351
transform 1 0 14511 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_55
timestamp 1666199351
transform 1 0 14975 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_56
timestamp 1666199351
transform 1 0 14379 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_57
timestamp 1666199351
transform 1 0 13915 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_58
timestamp 1666199351
transform 1 0 13263 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_59
timestamp 1666199351
transform 1 0 13727 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_60
timestamp 1666199351
transform 1 0 13131 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_61
timestamp 1666199351
transform 1 0 12667 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_62
timestamp 1666199351
transform 1 0 12015 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_63
timestamp 1666199351
transform 1 0 12479 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_64
timestamp 1666199351
transform 1 0 11883 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_65
timestamp 1666199351
transform 1 0 11419 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_66
timestamp 1666199351
transform 1 0 16005 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_67
timestamp 1666199351
transform 1 0 15381 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_68
timestamp 1666199351
transform 1 0 14757 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_69
timestamp 1666199351
transform 1 0 14133 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_70
timestamp 1666199351
transform 1 0 13509 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_71
timestamp 1666199351
transform 1 0 12885 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_72
timestamp 1666199351
transform 1 0 20997 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_73
timestamp 1666199351
transform 1 0 20373 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_74
timestamp 1666199351
transform 1 0 19749 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_75
timestamp 1666199351
transform 1 0 19125 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_76
timestamp 1666199351
transform 1 0 18501 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_77
timestamp 1666199351
transform 1 0 17877 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_78
timestamp 1666199351
transform 1 0 17253 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_79
timestamp 1666199351
transform 1 0 16629 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_80
timestamp 1666199351
transform 1 0 20751 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_81
timestamp 1666199351
transform 1 0 21215 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_82
timestamp 1666199351
transform 1 0 20619 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_83
timestamp 1666199351
transform 1 0 20155 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_84
timestamp 1666199351
transform 1 0 19503 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_85
timestamp 1666199351
transform 1 0 19967 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_86
timestamp 1666199351
transform 1 0 19371 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_87
timestamp 1666199351
transform 1 0 18907 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_88
timestamp 1666199351
transform 1 0 18255 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_89
timestamp 1666199351
transform 1 0 18719 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_90
timestamp 1666199351
transform 1 0 18123 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_91
timestamp 1666199351
transform 1 0 17659 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_92
timestamp 1666199351
transform 1 0 17007 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_93
timestamp 1666199351
transform 1 0 17471 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_94
timestamp 1666199351
transform 1 0 16875 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_95
timestamp 1666199351
transform 1 0 16411 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_96
timestamp 1666199351
transform 1 0 25989 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_97
timestamp 1666199351
transform 1 0 25365 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_98
timestamp 1666199351
transform 1 0 24741 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_99
timestamp 1666199351
transform 1 0 24117 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_100
timestamp 1666199351
transform 1 0 23493 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_101
timestamp 1666199351
transform 1 0 22869 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_102
timestamp 1666199351
transform 1 0 22245 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_103
timestamp 1666199351
transform 1 0 21621 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_104
timestamp 1666199351
transform 1 0 24495 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_105
timestamp 1666199351
transform 1 0 24959 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_106
timestamp 1666199351
transform 1 0 24363 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_107
timestamp 1666199351
transform 1 0 23899 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_108
timestamp 1666199351
transform 1 0 23247 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_109
timestamp 1666199351
transform 1 0 23711 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_110
timestamp 1666199351
transform 1 0 23115 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_111
timestamp 1666199351
transform 1 0 22651 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_112
timestamp 1666199351
transform 1 0 21999 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_113
timestamp 1666199351
transform 1 0 22463 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_114
timestamp 1666199351
transform 1 0 21867 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_115
timestamp 1666199351
transform 1 0 21403 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_116
timestamp 1666199351
transform 1 0 25743 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_117
timestamp 1666199351
transform 1 0 26207 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_118
timestamp 1666199351
transform 1 0 25611 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_119
timestamp 1666199351
transform 1 0 25147 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_120
timestamp 1666199351
transform 1 0 30981 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_121
timestamp 1666199351
transform 1 0 30357 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_122
timestamp 1666199351
transform 1 0 29733 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_123
timestamp 1666199351
transform 1 0 29109 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_124
timestamp 1666199351
transform 1 0 30735 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_125
timestamp 1666199351
transform 1 0 31199 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_126
timestamp 1666199351
transform 1 0 30603 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_127
timestamp 1666199351
transform 1 0 30139 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_128
timestamp 1666199351
transform 1 0 29487 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_129
timestamp 1666199351
transform 1 0 29951 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_130
timestamp 1666199351
transform 1 0 29355 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_131
timestamp 1666199351
transform 1 0 28891 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_132
timestamp 1666199351
transform 1 0 28239 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_133
timestamp 1666199351
transform 1 0 28703 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_134
timestamp 1666199351
transform 1 0 28107 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_135
timestamp 1666199351
transform 1 0 27643 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_136
timestamp 1666199351
transform 1 0 26991 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_137
timestamp 1666199351
transform 1 0 27455 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_138
timestamp 1666199351
transform 1 0 26859 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_139
timestamp 1666199351
transform 1 0 26395 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_140
timestamp 1666199351
transform 1 0 28485 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_141
timestamp 1666199351
transform 1 0 27861 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_142
timestamp 1666199351
transform 1 0 27237 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_143
timestamp 1666199351
transform 1 0 26613 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_144
timestamp 1666199351
transform 1 0 33477 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_145
timestamp 1666199351
transform 1 0 32853 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_146
timestamp 1666199351
transform 1 0 32229 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_147
timestamp 1666199351
transform 1 0 31605 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_148
timestamp 1666199351
transform 1 0 35973 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_149
timestamp 1666199351
transform 1 0 35349 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_150
timestamp 1666199351
transform 1 0 35727 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_151
timestamp 1666199351
transform 1 0 36191 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_152
timestamp 1666199351
transform 1 0 35595 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_153
timestamp 1666199351
transform 1 0 35131 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_154
timestamp 1666199351
transform 1 0 34479 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_155
timestamp 1666199351
transform 1 0 34943 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_156
timestamp 1666199351
transform 1 0 34347 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_157
timestamp 1666199351
transform 1 0 33883 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_158
timestamp 1666199351
transform 1 0 33231 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_159
timestamp 1666199351
transform 1 0 33695 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_160
timestamp 1666199351
transform 1 0 33099 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_161
timestamp 1666199351
transform 1 0 32635 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_162
timestamp 1666199351
transform 1 0 31983 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_163
timestamp 1666199351
transform 1 0 32447 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_164
timestamp 1666199351
transform 1 0 31851 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_165
timestamp 1666199351
transform 1 0 31387 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_166
timestamp 1666199351
transform 1 0 34725 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_167
timestamp 1666199351
transform 1 0 34101 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_168
timestamp 1666199351
transform 1 0 40719 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_169
timestamp 1666199351
transform 1 0 41183 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_170
timestamp 1666199351
transform 1 0 40587 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_171
timestamp 1666199351
transform 1 0 40123 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_172
timestamp 1666199351
transform 1 0 39471 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_173
timestamp 1666199351
transform 1 0 39935 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_174
timestamp 1666199351
transform 1 0 39339 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_175
timestamp 1666199351
transform 1 0 38875 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_176
timestamp 1666199351
transform 1 0 38223 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_177
timestamp 1666199351
transform 1 0 38687 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_178
timestamp 1666199351
transform 1 0 38091 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_179
timestamp 1666199351
transform 1 0 37627 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_180
timestamp 1666199351
transform 1 0 36975 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_181
timestamp 1666199351
transform 1 0 37439 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_182
timestamp 1666199351
transform 1 0 36843 0 1 87
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_183
timestamp 1666199351
transform 1 0 36379 0 1 211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_184
timestamp 1666199351
transform 1 0 40965 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_185
timestamp 1666199351
transform 1 0 40341 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_186
timestamp 1666199351
transform 1 0 39717 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_187
timestamp 1666199351
transform 1 0 39093 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_188
timestamp 1666199351
transform 1 0 38469 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_189
timestamp 1666199351
transform 1 0 37845 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_190
timestamp 1666199351
transform 1 0 37221 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_27  sky130_sram_1kbyte_1rw1r_32x256_8_contact_27_191
timestamp 1666199351
transform 1 0 36597 0 1 365
box 0 0 1 1
<< labels >>
rlabel metal3 s 0 372 41310 432 4 sel_0
port 1 nsew
rlabel metal3 s 0 496 41310 556 4 sel_1
port 2 nsew
rlabel metal3 s 18173 1234 18271 1332 4 gnd
port 3 nsew
rlabel metal3 s 18222 1283 18222 1283 4 gnd
port 3 nsew
rlabel metal3 s 36893 1234 36991 1332 4 gnd
port 3 nsew
rlabel metal3 s 14429 1234 14527 1332 4 gnd
port 3 nsew
rlabel metal3 s 14478 1283 14478 1283 4 gnd
port 3 nsew
rlabel metal3 s 9437 1234 9535 1332 4 gnd
port 3 nsew
rlabel metal3 s 19421 1234 19519 1332 4 gnd
port 3 nsew
rlabel metal3 s 8189 1234 8287 1332 4 gnd
port 3 nsew
rlabel metal3 s 23165 1234 23263 1332 4 gnd
port 3 nsew
rlabel metal3 s 33149 1234 33247 1332 4 gnd
port 3 nsew
rlabel metal3 s 16925 1234 17023 1332 4 gnd
port 3 nsew
rlabel metal3 s 13181 1234 13279 1332 4 gnd
port 3 nsew
rlabel metal3 s 25661 1234 25759 1332 4 gnd
port 3 nsew
rlabel metal3 s 11933 1234 12031 1332 4 gnd
port 3 nsew
rlabel metal3 s 38141 1234 38239 1332 4 gnd
port 3 nsew
rlabel metal3 s 38190 1283 38190 1283 4 gnd
port 3 nsew
rlabel metal3 s 20669 1234 20767 1332 4 gnd
port 3 nsew
rlabel metal3 s 20718 1283 20718 1283 4 gnd
port 3 nsew
rlabel metal3 s 21917 1234 22015 1332 4 gnd
port 3 nsew
rlabel metal3 s 15677 1234 15775 1332 4 gnd
port 3 nsew
rlabel metal3 s 10685 1234 10783 1332 4 gnd
port 3 nsew
rlabel metal3 s 10734 1283 10734 1283 4 gnd
port 3 nsew
rlabel metal3 s 30653 1234 30751 1332 4 gnd
port 3 nsew
rlabel metal3 s 30702 1283 30702 1283 4 gnd
port 3 nsew
rlabel metal3 s 1949 1234 2047 1332 4 gnd
port 3 nsew
rlabel metal3 s 1998 1283 1998 1283 4 gnd
port 3 nsew
rlabel metal3 s 29405 1234 29503 1332 4 gnd
port 3 nsew
rlabel metal3 s 26909 1234 27007 1332 4 gnd
port 3 nsew
rlabel metal3 s 26958 1283 26958 1283 4 gnd
port 3 nsew
rlabel metal3 s 6941 1234 7039 1332 4 gnd
port 3 nsew
rlabel metal3 s 5693 1234 5791 1332 4 gnd
port 3 nsew
rlabel metal3 s 5742 1283 5742 1283 4 gnd
port 3 nsew
rlabel metal3 s 3197 1234 3295 1332 4 gnd
port 3 nsew
rlabel metal3 s 3246 1283 3246 1283 4 gnd
port 3 nsew
rlabel metal3 s 35645 1234 35743 1332 4 gnd
port 3 nsew
rlabel metal3 s 24413 1234 24511 1332 4 gnd
port 3 nsew
rlabel metal3 s 24462 1283 24462 1283 4 gnd
port 3 nsew
rlabel metal3 s 31901 1234 31999 1332 4 gnd
port 3 nsew
rlabel metal3 s 34397 1234 34495 1332 4 gnd
port 3 nsew
rlabel metal3 s 34446 1283 34446 1283 4 gnd
port 3 nsew
rlabel metal3 s 39389 1234 39487 1332 4 gnd
port 3 nsew
rlabel metal3 s 40637 1234 40735 1332 4 gnd
port 3 nsew
rlabel metal3 s 4445 1234 4543 1332 4 gnd
port 3 nsew
rlabel metal3 s 4494 1283 4494 1283 4 gnd
port 3 nsew
rlabel metal3 s 28157 1234 28255 1332 4 gnd
port 3 nsew
rlabel metal1 s 21422 248 21450 620 4 bl_out_16
port 4 nsew
rlabel metal1 s 22670 248 22698 620 4 bl_out_17
port 5 nsew
rlabel metal1 s 23918 248 23946 620 4 bl_out_18
port 6 nsew
rlabel metal1 s 25166 248 25194 620 4 bl_out_19
port 7 nsew
rlabel metal1 s 26414 248 26442 620 4 bl_out_20
port 8 nsew
rlabel metal1 s 27662 248 27690 620 4 bl_out_21
port 9 nsew
rlabel metal1 s 28910 248 28938 620 4 bl_out_22
port 10 nsew
rlabel metal1 s 30158 248 30186 620 4 bl_out_23
port 11 nsew
rlabel metal1 s 31406 248 31434 620 4 bl_out_24
port 12 nsew
rlabel metal1 s 32654 248 32682 620 4 bl_out_25
port 13 nsew
rlabel metal1 s 33902 248 33930 620 4 bl_out_26
port 14 nsew
rlabel metal1 s 35150 248 35178 620 4 bl_out_27
port 15 nsew
rlabel metal1 s 36398 248 36426 620 4 bl_out_28
port 16 nsew
rlabel metal1 s 37646 248 37674 620 4 bl_out_29
port 17 nsew
rlabel metal1 s 38894 248 38922 620 4 bl_out_30
port 18 nsew
rlabel metal1 s 40142 248 40170 620 4 bl_out_31
port 19 nsew
rlabel metal1 s 21422 1880 21450 1936 4 bl_32
port 20 nsew
rlabel metal1 s 21886 1880 21914 1936 4 br_32
port 21 nsew
rlabel metal1 s 22482 1880 22510 1936 4 bl_33
port 22 nsew
rlabel metal1 s 22018 1880 22046 1936 4 br_33
port 23 nsew
rlabel metal1 s 22670 1880 22698 1936 4 bl_34
port 24 nsew
rlabel metal1 s 23134 1880 23162 1936 4 br_34
port 25 nsew
rlabel metal1 s 23730 1880 23758 1936 4 bl_35
port 26 nsew
rlabel metal1 s 23266 1880 23294 1936 4 br_35
port 27 nsew
rlabel metal1 s 23918 1880 23946 1936 4 bl_36
port 28 nsew
rlabel metal1 s 24382 1880 24410 1936 4 br_36
port 29 nsew
rlabel metal1 s 24978 1880 25006 1936 4 bl_37
port 30 nsew
rlabel metal1 s 24514 1880 24542 1936 4 br_37
port 31 nsew
rlabel metal1 s 25166 1880 25194 1936 4 bl_38
port 32 nsew
rlabel metal1 s 25630 1880 25658 1936 4 br_38
port 33 nsew
rlabel metal1 s 26226 1880 26254 1936 4 bl_39
port 34 nsew
rlabel metal1 s 25762 1880 25790 1936 4 br_39
port 35 nsew
rlabel metal1 s 26414 1880 26442 1936 4 bl_40
port 36 nsew
rlabel metal1 s 26878 1880 26906 1936 4 br_40
port 37 nsew
rlabel metal1 s 27474 1880 27502 1936 4 bl_41
port 38 nsew
rlabel metal1 s 27010 1880 27038 1936 4 br_41
port 39 nsew
rlabel metal1 s 27662 1880 27690 1936 4 bl_42
port 40 nsew
rlabel metal1 s 28126 1880 28154 1936 4 br_42
port 41 nsew
rlabel metal1 s 28722 1880 28750 1936 4 bl_43
port 42 nsew
rlabel metal1 s 28258 1880 28286 1936 4 br_43
port 43 nsew
rlabel metal1 s 28910 1880 28938 1936 4 bl_44
port 44 nsew
rlabel metal1 s 29374 1880 29402 1936 4 br_44
port 45 nsew
rlabel metal1 s 29970 1880 29998 1936 4 bl_45
port 46 nsew
rlabel metal1 s 29506 1880 29534 1936 4 br_45
port 47 nsew
rlabel metal1 s 30158 1880 30186 1936 4 bl_46
port 48 nsew
rlabel metal1 s 30622 1880 30650 1936 4 br_46
port 49 nsew
rlabel metal1 s 31218 1880 31246 1936 4 bl_47
port 50 nsew
rlabel metal1 s 30754 1880 30782 1936 4 br_47
port 51 nsew
rlabel metal1 s 31406 1880 31434 1936 4 bl_48
port 52 nsew
rlabel metal1 s 31870 1880 31898 1936 4 br_48
port 53 nsew
rlabel metal1 s 32466 1880 32494 1936 4 bl_49
port 54 nsew
rlabel metal1 s 32002 1880 32030 1936 4 br_49
port 55 nsew
rlabel metal1 s 32654 1880 32682 1936 4 bl_50
port 56 nsew
rlabel metal1 s 33118 1880 33146 1936 4 br_50
port 57 nsew
rlabel metal1 s 33714 1880 33742 1936 4 bl_51
port 58 nsew
rlabel metal1 s 33250 1880 33278 1936 4 br_51
port 59 nsew
rlabel metal1 s 33902 1880 33930 1936 4 bl_52
port 60 nsew
rlabel metal1 s 34366 1880 34394 1936 4 br_52
port 61 nsew
rlabel metal1 s 34962 1880 34990 1936 4 bl_53
port 62 nsew
rlabel metal1 s 34498 1880 34526 1936 4 br_53
port 63 nsew
rlabel metal1 s 35150 1880 35178 1936 4 bl_54
port 64 nsew
rlabel metal1 s 35614 1880 35642 1936 4 br_54
port 65 nsew
rlabel metal1 s 36210 1880 36238 1936 4 bl_55
port 66 nsew
rlabel metal1 s 35746 1880 35774 1936 4 br_55
port 67 nsew
rlabel metal1 s 36398 1880 36426 1936 4 bl_56
port 68 nsew
rlabel metal1 s 36862 1880 36890 1936 4 br_56
port 69 nsew
rlabel metal1 s 37458 1880 37486 1936 4 bl_57
port 70 nsew
rlabel metal1 s 36994 1880 37022 1936 4 br_57
port 71 nsew
rlabel metal1 s 37646 1880 37674 1936 4 bl_58
port 72 nsew
rlabel metal1 s 38110 1880 38138 1936 4 br_58
port 73 nsew
rlabel metal1 s 38706 1880 38734 1936 4 bl_59
port 74 nsew
rlabel metal1 s 38242 1880 38270 1936 4 br_59
port 75 nsew
rlabel metal1 s 38894 1880 38922 1936 4 bl_60
port 76 nsew
rlabel metal1 s 39358 1880 39386 1936 4 br_60
port 77 nsew
rlabel metal1 s 39954 1880 39982 1936 4 bl_61
port 78 nsew
rlabel metal1 s 39490 1880 39518 1936 4 br_61
port 79 nsew
rlabel metal1 s 40142 1880 40170 1936 4 bl_62
port 80 nsew
rlabel metal1 s 40606 1880 40634 1936 4 br_62
port 81 nsew
rlabel metal1 s 41202 1880 41230 1936 4 bl_63
port 82 nsew
rlabel metal1 s 40738 1880 40766 1936 4 br_63
port 83 nsew
rlabel metal1 s 16430 1880 16458 1936 4 bl_24
port 84 nsew
rlabel metal1 s 16894 1880 16922 1936 4 br_24
port 85 nsew
rlabel metal1 s 17490 1880 17518 1936 4 bl_25
port 86 nsew
rlabel metal1 s 17026 1880 17054 1936 4 br_25
port 87 nsew
rlabel metal1 s 17678 1880 17706 1936 4 bl_26
port 88 nsew
rlabel metal1 s 18142 1880 18170 1936 4 br_26
port 89 nsew
rlabel metal1 s 18738 1880 18766 1936 4 bl_27
port 90 nsew
rlabel metal1 s 18274 1880 18302 1936 4 br_27
port 91 nsew
rlabel metal1 s 18926 1880 18954 1936 4 bl_28
port 92 nsew
rlabel metal1 s 19390 1880 19418 1936 4 br_28
port 93 nsew
rlabel metal1 s 19986 1880 20014 1936 4 bl_29
port 94 nsew
rlabel metal1 s 19522 1880 19550 1936 4 br_29
port 95 nsew
rlabel metal1 s 20174 1880 20202 1936 4 bl_30
port 96 nsew
rlabel metal1 s 20638 1880 20666 1936 4 br_30
port 97 nsew
rlabel metal1 s 21234 1880 21262 1936 4 bl_31
port 98 nsew
rlabel metal1 s 20770 1880 20798 1936 4 br_31
port 99 nsew
rlabel metal1 s 1454 248 1482 620 4 bl_out_0
port 100 nsew
rlabel metal1 s 2702 248 2730 620 4 bl_out_1
port 101 nsew
rlabel metal1 s 3950 248 3978 620 4 bl_out_2
port 102 nsew
rlabel metal1 s 5198 248 5226 620 4 bl_out_3
port 103 nsew
rlabel metal1 s 6446 248 6474 620 4 bl_out_4
port 104 nsew
rlabel metal1 s 7694 248 7722 620 4 bl_out_5
port 105 nsew
rlabel metal1 s 8942 248 8970 620 4 bl_out_6
port 106 nsew
rlabel metal1 s 10190 248 10218 620 4 bl_out_7
port 107 nsew
rlabel metal1 s 11438 248 11466 620 4 bl_out_8
port 108 nsew
rlabel metal1 s 12686 248 12714 620 4 bl_out_9
port 109 nsew
rlabel metal1 s 13934 248 13962 620 4 bl_out_10
port 110 nsew
rlabel metal1 s 15182 248 15210 620 4 bl_out_11
port 111 nsew
rlabel metal1 s 16430 248 16458 620 4 bl_out_12
port 112 nsew
rlabel metal1 s 17678 248 17706 620 4 bl_out_13
port 113 nsew
rlabel metal1 s 18926 248 18954 620 4 bl_out_14
port 114 nsew
rlabel metal1 s 20174 248 20202 620 4 bl_out_15
port 115 nsew
rlabel metal1 s 1454 1880 1482 1936 4 bl_0
port 116 nsew
rlabel metal1 s 1918 1880 1946 1936 4 br_0
port 117 nsew
rlabel metal1 s 2514 1880 2542 1936 4 bl_1
port 118 nsew
rlabel metal1 s 2050 1880 2078 1936 4 br_1
port 119 nsew
rlabel metal1 s 2702 1880 2730 1936 4 bl_2
port 120 nsew
rlabel metal1 s 3166 1880 3194 1936 4 br_2
port 121 nsew
rlabel metal1 s 3762 1880 3790 1936 4 bl_3
port 122 nsew
rlabel metal1 s 3298 1880 3326 1936 4 br_3
port 123 nsew
rlabel metal1 s 3950 1880 3978 1936 4 bl_4
port 124 nsew
rlabel metal1 s 4414 1880 4442 1936 4 br_4
port 125 nsew
rlabel metal1 s 5010 1880 5038 1936 4 bl_5
port 126 nsew
rlabel metal1 s 4546 1880 4574 1936 4 br_5
port 127 nsew
rlabel metal1 s 5198 1880 5226 1936 4 bl_6
port 128 nsew
rlabel metal1 s 5662 1880 5690 1936 4 br_6
port 129 nsew
rlabel metal1 s 6258 1880 6286 1936 4 bl_7
port 130 nsew
rlabel metal1 s 5794 1880 5822 1936 4 br_7
port 131 nsew
rlabel metal1 s 6446 1880 6474 1936 4 bl_8
port 132 nsew
rlabel metal1 s 6910 1880 6938 1936 4 br_8
port 133 nsew
rlabel metal1 s 7506 1880 7534 1936 4 bl_9
port 134 nsew
rlabel metal1 s 7042 1880 7070 1936 4 br_9
port 135 nsew
rlabel metal1 s 7694 1880 7722 1936 4 bl_10
port 136 nsew
rlabel metal1 s 8158 1880 8186 1936 4 br_10
port 137 nsew
rlabel metal1 s 8754 1880 8782 1936 4 bl_11
port 138 nsew
rlabel metal1 s 8290 1880 8318 1936 4 br_11
port 139 nsew
rlabel metal1 s 8942 1880 8970 1936 4 bl_12
port 140 nsew
rlabel metal1 s 9406 1880 9434 1936 4 br_12
port 141 nsew
rlabel metal1 s 10002 1880 10030 1936 4 bl_13
port 142 nsew
rlabel metal1 s 9538 1880 9566 1936 4 br_13
port 143 nsew
rlabel metal1 s 10190 1880 10218 1936 4 bl_14
port 144 nsew
rlabel metal1 s 10654 1880 10682 1936 4 br_14
port 145 nsew
rlabel metal1 s 11250 1880 11278 1936 4 bl_15
port 146 nsew
rlabel metal1 s 10786 1880 10814 1936 4 br_15
port 147 nsew
rlabel metal1 s 11438 1880 11466 1936 4 bl_16
port 148 nsew
rlabel metal1 s 11902 1880 11930 1936 4 br_16
port 149 nsew
rlabel metal1 s 12498 1880 12526 1936 4 bl_17
port 150 nsew
rlabel metal1 s 12034 1880 12062 1936 4 br_17
port 151 nsew
rlabel metal1 s 12686 1880 12714 1936 4 bl_18
port 152 nsew
rlabel metal1 s 13150 1880 13178 1936 4 br_18
port 153 nsew
rlabel metal1 s 13746 1880 13774 1936 4 bl_19
port 154 nsew
rlabel metal1 s 13282 1880 13310 1936 4 br_19
port 155 nsew
rlabel metal1 s 13934 1880 13962 1936 4 bl_20
port 156 nsew
rlabel metal1 s 14398 1880 14426 1936 4 br_20
port 157 nsew
rlabel metal1 s 14994 1880 15022 1936 4 bl_21
port 158 nsew
rlabel metal1 s 14530 1880 14558 1936 4 br_21
port 159 nsew
rlabel metal1 s 15182 1880 15210 1936 4 bl_22
port 160 nsew
rlabel metal1 s 15646 1880 15674 1936 4 br_22
port 161 nsew
rlabel metal1 s 16242 1880 16270 1936 4 bl_23
port 162 nsew
rlabel metal1 s 15778 1880 15806 1936 4 br_23
port 163 nsew
rlabel metal1 s 1918 124 1946 620 4 br_out_0
port 164 nsew
rlabel metal1 s 11902 124 11930 620 4 br_out_8
port 165 nsew
rlabel metal1 s 6910 124 6938 620 4 br_out_4
port 166 nsew
rlabel metal1 s 13150 124 13178 620 4 br_out_9
port 167 nsew
rlabel metal1 s 4414 124 4442 620 4 br_out_2
port 168 nsew
rlabel metal1 s 14398 124 14426 620 4 br_out_10
port 169 nsew
rlabel metal1 s 8158 124 8186 620 4 br_out_5
port 170 nsew
rlabel metal1 s 15646 124 15674 620 4 br_out_11
port 171 nsew
rlabel metal1 s 3166 124 3194 620 4 br_out_1
port 172 nsew
rlabel metal1 s 16894 124 16922 620 4 br_out_12
port 173 nsew
rlabel metal1 s 9406 124 9434 620 4 br_out_6
port 174 nsew
rlabel metal1 s 18142 124 18170 620 4 br_out_13
port 175 nsew
rlabel metal1 s 5662 124 5690 620 4 br_out_3
port 176 nsew
rlabel metal1 s 19390 124 19418 620 4 br_out_14
port 177 nsew
rlabel metal1 s 10654 124 10682 620 4 br_out_7
port 178 nsew
rlabel metal1 s 20638 124 20666 620 4 br_out_15
port 179 nsew
rlabel metal1 s 21886 124 21914 620 4 br_out_16
port 180 nsew
rlabel metal1 s 31870 124 31898 620 4 br_out_24
port 181 nsew
rlabel metal1 s 26878 124 26906 620 4 br_out_20
port 182 nsew
rlabel metal1 s 33118 124 33146 620 4 br_out_25
port 183 nsew
rlabel metal1 s 24382 124 24410 620 4 br_out_18
port 184 nsew
rlabel metal1 s 34366 124 34394 620 4 br_out_26
port 185 nsew
rlabel metal1 s 28126 124 28154 620 4 br_out_21
port 186 nsew
rlabel metal1 s 35614 124 35642 620 4 br_out_27
port 187 nsew
rlabel metal1 s 23134 124 23162 620 4 br_out_17
port 188 nsew
rlabel metal1 s 36862 124 36890 620 4 br_out_28
port 189 nsew
rlabel metal1 s 29374 124 29402 620 4 br_out_22
port 190 nsew
rlabel metal1 s 38110 124 38138 620 4 br_out_29
port 191 nsew
rlabel metal1 s 25630 124 25658 620 4 br_out_19
port 192 nsew
rlabel metal1 s 39358 124 39386 620 4 br_out_30
port 193 nsew
rlabel metal1 s 30622 124 30650 620 4 br_out_23
port 194 nsew
rlabel metal1 s 40606 124 40634 620 4 br_out_31
port 195 nsew
<< properties >>
string FIXED_BBOX 40719 87 40785 161
string GDS_END 947598
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 833508
<< end >>
