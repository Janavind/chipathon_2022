magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 163 187 203
rect 453 163 643 203
rect 1 67 643 163
rect 30 27 643 67
rect 30 -17 64 27
rect 456 21 643 27
<< locali >>
rect 17 215 85 391
rect 358 425 453 493
rect 572 353 627 493
rect 397 145 479 249
rect 593 147 627 353
rect 397 61 437 145
rect 575 51 627 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 425 69 527
rect 119 249 153 493
rect 201 426 324 527
rect 201 319 251 392
rect 285 391 324 426
rect 487 418 530 527
rect 285 353 351 391
rect 395 319 538 378
rect 201 285 559 319
rect 119 199 278 249
rect 119 181 169 199
rect 17 17 69 181
rect 103 97 169 181
rect 312 114 363 285
rect 205 61 363 114
rect 513 199 559 285
rect 475 17 541 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 17 215 85 391 6 A_N
port 1 nsew signal input
rlabel locali s 358 425 453 493 6 B
port 2 nsew signal input
rlabel locali s 397 61 437 145 6 C
port 3 nsew signal input
rlabel locali s 397 145 479 249 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 456 21 643 27 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 30 -17 64 27 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 30 27 643 67 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 67 643 163 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 453 163 643 203 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 163 187 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 575 51 627 147 6 X
port 8 nsew signal output
rlabel locali s 593 147 627 353 6 X
port 8 nsew signal output
rlabel locali s 572 353 627 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3877840
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3871498
<< end >>
