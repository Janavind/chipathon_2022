magic
tech sky130B
magscale 1 2
timestamp 1666464484
use sky130_fd_pr__dfm1sd__example_55959141808169  sky130_fd_pr__dfm1sd__example_55959141808169_0
timestamp 1666464484
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfm1sd__example_55959141808169  sky130_fd_pr__dfm1sd__example_55959141808169_1
timestamp 1666464484
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808170  sky130_fd_pr__hvdfm1sd2__example_55959141808170_0
timestamp 1666464484
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808170  sky130_fd_pr__hvdfm1sd2__example_55959141808170_1
timestamp 1666464484
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808170  sky130_fd_pr__hvdfm1sd2__example_55959141808170_2
timestamp 1666464484
transform 1 0 412 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 35448958
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35446354
<< end >>
