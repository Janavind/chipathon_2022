magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 182 157 456 203
rect 1 21 456 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 264 47 294 177
rect 348 47 378 177
<< scpmoshvt >>
rect 91 297 121 381
rect 163 297 193 381
rect 264 297 294 497
rect 348 297 378 497
<< ndiff >>
rect 208 131 264 177
rect 27 103 79 131
rect 27 69 35 103
rect 69 69 79 103
rect 27 47 79 69
rect 109 103 163 131
rect 109 69 119 103
rect 153 69 163 103
rect 109 47 163 69
rect 193 103 264 131
rect 193 69 219 103
rect 253 69 264 103
rect 193 47 264 69
rect 294 130 348 177
rect 294 96 304 130
rect 338 96 348 130
rect 294 47 348 96
rect 378 95 430 177
rect 378 61 388 95
rect 422 61 430 95
rect 378 47 430 61
<< pdiff >>
rect 208 487 264 497
rect 208 453 220 487
rect 254 453 264 487
rect 208 419 264 453
rect 208 385 220 419
rect 254 385 264 419
rect 208 381 264 385
rect 39 349 91 381
rect 39 315 47 349
rect 81 315 91 349
rect 39 297 91 315
rect 121 297 163 381
rect 193 297 264 381
rect 294 485 348 497
rect 294 451 304 485
rect 338 451 348 485
rect 294 417 348 451
rect 294 383 304 417
rect 338 383 348 417
rect 294 297 348 383
rect 378 485 430 497
rect 378 451 388 485
rect 422 451 430 485
rect 378 297 430 451
<< ndiffc >>
rect 35 69 69 103
rect 119 69 153 103
rect 219 69 253 103
rect 304 96 338 130
rect 388 61 422 95
<< pdiffc >>
rect 220 453 254 487
rect 220 385 254 419
rect 47 315 81 349
rect 304 451 338 485
rect 304 383 338 417
rect 388 451 422 485
<< poly >>
rect 264 497 294 523
rect 348 497 378 523
rect 91 381 121 407
rect 163 381 193 407
rect 91 265 121 297
rect 25 249 121 265
rect 25 215 35 249
rect 69 215 121 249
rect 25 199 121 215
rect 163 265 193 297
rect 264 265 294 297
rect 348 265 378 297
rect 163 249 217 265
rect 163 215 173 249
rect 207 215 217 249
rect 163 199 217 215
rect 264 249 378 265
rect 264 215 289 249
rect 323 215 378 249
rect 264 199 378 215
rect 79 131 109 199
rect 163 131 193 199
rect 264 177 294 199
rect 348 177 378 199
rect 79 21 109 47
rect 163 21 193 47
rect 264 21 294 47
rect 348 21 378 47
<< polycont >>
rect 35 215 69 249
rect 173 215 207 249
rect 289 215 323 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 220 487 254 527
rect 220 419 254 453
rect 31 349 103 368
rect 220 367 254 385
rect 288 485 354 493
rect 288 451 304 485
rect 338 451 354 485
rect 288 417 354 451
rect 388 485 422 527
rect 388 435 422 451
rect 288 383 304 417
rect 338 401 354 417
rect 338 383 443 401
rect 288 367 443 383
rect 31 315 47 349
rect 81 333 103 349
rect 81 315 323 333
rect 31 299 323 315
rect 30 249 69 265
rect 30 215 35 249
rect 30 153 69 215
rect 103 119 139 299
rect 173 249 255 265
rect 207 215 255 249
rect 173 153 255 215
rect 289 249 323 299
rect 289 199 323 215
rect 357 165 443 367
rect 304 131 443 165
rect 304 130 338 131
rect 21 103 69 119
rect 21 69 35 103
rect 21 17 69 69
rect 103 103 161 119
rect 103 69 119 103
rect 153 69 161 103
rect 103 51 161 69
rect 207 103 270 119
rect 207 69 219 103
rect 253 69 270 103
rect 304 77 338 96
rect 372 95 438 97
rect 207 17 270 69
rect 372 61 388 95
rect 422 61 438 95
rect 372 17 438 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 398 357 432 391 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 or2_2
rlabel metal1 s 0 -48 460 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 988668
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 984310
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 2.720 2.300 2.720 
<< end >>
