magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1099 203
rect 30 -17 64 21
<< scnmos >>
rect 80 47 110 177
rect 166 47 196 177
rect 252 47 282 177
rect 338 47 368 177
rect 528 47 558 177
rect 614 47 644 177
rect 716 47 746 177
rect 818 47 848 177
rect 904 47 934 177
rect 990 47 1020 177
<< scpmoshvt >>
rect 144 297 174 497
rect 230 297 260 497
rect 316 297 346 497
rect 402 297 432 497
rect 492 297 522 497
rect 578 297 608 497
rect 732 297 762 497
rect 818 297 848 497
rect 904 297 934 497
rect 990 297 1020 497
<< ndiff >>
rect 27 93 80 177
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 161 166 177
rect 110 127 121 161
rect 155 127 166 161
rect 110 47 166 127
rect 196 89 252 177
rect 196 55 207 89
rect 241 55 252 89
rect 196 47 252 55
rect 282 159 338 177
rect 282 125 293 159
rect 327 125 338 159
rect 282 47 338 125
rect 368 93 421 177
rect 368 59 379 93
rect 413 59 421 93
rect 368 47 421 59
rect 475 93 528 177
rect 475 59 483 93
rect 517 59 528 93
rect 475 47 528 59
rect 558 169 614 177
rect 558 135 569 169
rect 603 135 614 169
rect 558 47 614 135
rect 644 157 716 177
rect 644 123 671 157
rect 705 123 716 157
rect 644 89 716 123
rect 644 55 671 89
rect 705 55 716 89
rect 644 47 716 55
rect 746 89 818 177
rect 746 55 771 89
rect 805 55 818 89
rect 746 47 818 55
rect 848 157 904 177
rect 848 123 859 157
rect 893 123 904 157
rect 848 47 904 123
rect 934 89 990 177
rect 934 55 945 89
rect 979 55 990 89
rect 934 47 990 55
rect 1020 157 1073 177
rect 1020 123 1031 157
rect 1065 123 1073 157
rect 1020 47 1073 123
<< pdiff >>
rect 91 485 144 497
rect 91 451 99 485
rect 133 451 144 485
rect 91 408 144 451
rect 91 374 99 408
rect 133 374 144 408
rect 91 297 144 374
rect 174 477 230 497
rect 174 443 185 477
rect 219 443 230 477
rect 174 385 230 443
rect 174 351 185 385
rect 219 351 230 385
rect 174 297 230 351
rect 260 485 316 497
rect 260 451 271 485
rect 305 451 316 485
rect 260 408 316 451
rect 260 374 271 408
rect 305 374 316 408
rect 260 297 316 374
rect 346 477 402 497
rect 346 443 357 477
rect 391 443 402 477
rect 346 385 402 443
rect 346 351 357 385
rect 391 351 402 385
rect 346 297 402 351
rect 432 485 492 497
rect 432 451 447 485
rect 481 451 492 485
rect 432 297 492 451
rect 522 477 578 497
rect 522 443 533 477
rect 567 443 578 477
rect 522 409 578 443
rect 522 375 533 409
rect 567 375 578 409
rect 522 297 578 375
rect 608 489 732 497
rect 608 455 619 489
rect 653 455 687 489
rect 721 455 732 489
rect 608 297 732 455
rect 762 297 818 497
rect 848 489 904 497
rect 848 455 859 489
rect 893 455 904 489
rect 848 421 904 455
rect 848 387 859 421
rect 893 387 904 421
rect 848 297 904 387
rect 934 297 990 497
rect 1020 489 1077 497
rect 1020 455 1031 489
rect 1065 455 1077 489
rect 1020 421 1077 455
rect 1020 387 1031 421
rect 1065 387 1077 421
rect 1020 297 1077 387
<< ndiffc >>
rect 35 59 69 93
rect 121 127 155 161
rect 207 55 241 89
rect 293 125 327 159
rect 379 59 413 93
rect 483 59 517 93
rect 569 135 603 169
rect 671 123 705 157
rect 671 55 705 89
rect 771 55 805 89
rect 859 123 893 157
rect 945 55 979 89
rect 1031 123 1065 157
<< pdiffc >>
rect 99 451 133 485
rect 99 374 133 408
rect 185 443 219 477
rect 185 351 219 385
rect 271 451 305 485
rect 271 374 305 408
rect 357 443 391 477
rect 357 351 391 385
rect 447 451 481 485
rect 533 443 567 477
rect 533 375 567 409
rect 619 455 653 489
rect 687 455 721 489
rect 859 455 893 489
rect 859 387 893 421
rect 1031 455 1065 489
rect 1031 387 1065 421
<< poly >>
rect 144 497 174 523
rect 230 497 260 523
rect 316 497 346 523
rect 402 497 432 523
rect 492 497 522 523
rect 578 497 608 523
rect 732 497 762 523
rect 818 497 848 523
rect 904 497 934 523
rect 990 497 1020 523
rect 144 265 174 297
rect 230 265 260 297
rect 316 265 346 297
rect 402 265 432 297
rect 80 249 432 265
rect 80 215 110 249
rect 144 215 178 249
rect 212 215 246 249
rect 280 215 314 249
rect 348 215 382 249
rect 416 215 432 249
rect 80 199 432 215
rect 492 265 522 297
rect 578 265 608 297
rect 732 265 762 297
rect 492 249 644 265
rect 492 215 513 249
rect 547 215 581 249
rect 615 215 644 249
rect 492 199 644 215
rect 687 249 762 265
rect 687 215 703 249
rect 737 215 762 249
rect 687 199 762 215
rect 818 265 848 297
rect 904 265 934 297
rect 990 265 1020 297
rect 818 249 948 265
rect 818 215 828 249
rect 862 215 904 249
rect 938 215 948 249
rect 818 199 948 215
rect 990 249 1056 265
rect 990 215 1006 249
rect 1040 215 1056 249
rect 990 199 1056 215
rect 80 177 110 199
rect 166 177 196 199
rect 252 177 282 199
rect 338 177 368 199
rect 528 177 558 199
rect 614 177 644 199
rect 716 177 746 199
rect 818 177 848 199
rect 904 177 934 199
rect 990 177 1020 199
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 338 21 368 47
rect 528 21 558 47
rect 614 21 644 47
rect 716 21 746 47
rect 818 21 848 47
rect 904 21 934 47
rect 990 21 1020 47
<< polycont >>
rect 110 215 144 249
rect 178 215 212 249
rect 246 215 280 249
rect 314 215 348 249
rect 382 215 416 249
rect 513 215 547 249
rect 581 215 615 249
rect 703 215 737 249
rect 828 215 862 249
rect 904 215 938 249
rect 1006 215 1040 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 83 485 149 527
rect 83 451 99 485
rect 133 451 149 485
rect 83 408 149 451
rect 83 374 99 408
rect 133 374 149 408
rect 183 477 221 493
rect 183 443 185 477
rect 219 443 221 477
rect 183 385 221 443
rect 183 351 185 385
rect 219 351 221 385
rect 255 485 321 527
rect 255 451 271 485
rect 305 451 321 485
rect 255 408 321 451
rect 255 374 271 408
rect 305 374 321 408
rect 355 477 391 493
rect 355 443 357 477
rect 427 485 497 527
rect 427 451 447 485
rect 481 451 497 485
rect 531 477 569 493
rect 355 385 391 443
rect 531 443 533 477
rect 567 443 569 477
rect 603 489 737 527
rect 1015 489 1087 527
rect 603 455 619 489
rect 653 455 687 489
rect 721 455 737 489
rect 843 455 859 489
rect 893 455 909 489
rect 531 421 569 443
rect 843 421 909 455
rect 531 417 859 421
rect 183 340 221 351
rect 355 351 357 385
rect 355 340 391 351
rect 18 306 391 340
rect 425 409 859 417
rect 425 375 533 409
rect 567 387 859 409
rect 893 387 909 421
rect 1015 455 1031 489
rect 1065 455 1087 489
rect 1015 421 1087 455
rect 1015 387 1031 421
rect 1065 387 1087 421
rect 567 375 909 387
rect 425 366 569 375
rect 18 161 64 306
rect 425 267 463 366
rect 98 249 463 267
rect 98 215 110 249
rect 144 215 178 249
rect 212 215 246 249
rect 280 215 314 249
rect 348 215 382 249
rect 416 215 463 249
rect 497 249 631 323
rect 497 215 513 249
rect 547 215 581 249
rect 615 215 631 249
rect 696 299 1080 341
rect 696 249 757 299
rect 696 215 703 249
rect 737 215 757 249
rect 98 199 463 215
rect 423 174 463 199
rect 696 198 757 215
rect 828 249 938 265
rect 862 215 904 249
rect 828 199 938 215
rect 1006 249 1080 299
rect 1040 215 1080 249
rect 1006 199 1080 215
rect 423 169 619 174
rect 18 127 121 161
rect 155 159 343 161
rect 155 127 293 159
rect 119 125 293 127
rect 327 125 343 159
rect 423 135 569 169
rect 603 135 619 169
rect 423 131 619 135
rect 119 123 343 125
rect 655 123 671 157
rect 705 123 859 157
rect 893 123 1031 157
rect 1065 123 1081 157
rect 655 97 721 123
rect 467 93 721 97
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 191 55 207 89
rect 241 55 257 89
rect 191 17 257 55
rect 363 59 379 93
rect 413 59 429 93
rect 363 17 429 59
rect 467 59 483 93
rect 517 89 721 93
rect 517 59 671 89
rect 467 55 671 59
rect 705 55 721 89
rect 467 51 721 55
rect 755 55 771 89
rect 805 55 823 89
rect 755 17 823 55
rect 929 55 945 89
rect 979 55 995 89
rect 929 17 995 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 1046 289 1080 323 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 862 221 896 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 586 289 620 323 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 30 153 64 187 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 o21a_4
rlabel metal1 s 0 -48 1104 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_END 1287542
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1279618
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 5.520 0.000 
<< end >>
