magic
tech sky130A
magscale 1 2
timestamp 1666464484
use sky130_fd_pr__hvdfm1sd2__example_5595914180827  sky130_fd_pr__hvdfm1sd2__example_5595914180827_0
timestamp 1666464484
transform 1 0 160 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808233  sky130_fd_pr__hvdfm1sd__example_55959141808233_0
timestamp 1666464484
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808233  sky130_fd_pr__hvdfm1sd__example_55959141808233_1
timestamp 1666464484
transform 1 0 376 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 240694
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 239252
<< end >>
