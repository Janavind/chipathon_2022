magic
tech sky130A
magscale 1 2
timestamp 1666464484
use sky130_fd_pr__dfl1sd__example_55959141808504  sky130_fd_pr__dfl1sd__example_55959141808504_0
timestamp 1666464484
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808462  sky130_fd_pr__hvdfl1sd2__example_55959141808462_0
timestamp 1666464484
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808278  sky130_fd_pr__hvdfl1sd__example_55959141808278_0
timestamp 1666464484
transform -1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 29612212
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 29610770
<< end >>
