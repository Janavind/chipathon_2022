magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect 1167 10569 1701 10901
<< pwell >>
rect 1260 11244 1646 11436
rect 1560 11232 1646 11244
<< mvnmos >>
rect 1339 11270 1459 11410
<< mvpmos >>
rect 1286 10635 1406 10835
rect 1462 10635 1582 10835
<< mvndiff >>
rect 1286 11398 1339 11410
rect 1286 11364 1294 11398
rect 1328 11364 1339 11398
rect 1286 11330 1339 11364
rect 1286 11296 1294 11330
rect 1328 11296 1339 11330
rect 1286 11270 1339 11296
rect 1459 11398 1512 11410
rect 1459 11364 1470 11398
rect 1504 11364 1512 11398
rect 1459 11330 1512 11364
rect 1459 11296 1470 11330
rect 1504 11296 1512 11330
rect 1459 11270 1512 11296
<< mvpdiff >>
rect 1233 10823 1286 10835
rect 1233 10789 1241 10823
rect 1275 10789 1286 10823
rect 1233 10755 1286 10789
rect 1233 10721 1241 10755
rect 1275 10721 1286 10755
rect 1233 10687 1286 10721
rect 1233 10653 1241 10687
rect 1275 10653 1286 10687
rect 1233 10635 1286 10653
rect 1406 10823 1462 10835
rect 1406 10789 1417 10823
rect 1451 10789 1462 10823
rect 1406 10755 1462 10789
rect 1406 10721 1417 10755
rect 1451 10721 1462 10755
rect 1406 10687 1462 10721
rect 1406 10653 1417 10687
rect 1451 10653 1462 10687
rect 1406 10635 1462 10653
rect 1582 10823 1635 10835
rect 1582 10789 1593 10823
rect 1627 10789 1635 10823
rect 1582 10755 1635 10789
rect 1582 10721 1593 10755
rect 1627 10721 1635 10755
rect 1582 10687 1635 10721
rect 1582 10653 1593 10687
rect 1627 10653 1635 10687
rect 1582 10635 1635 10653
<< mvndiffc >>
rect 1294 11364 1328 11398
rect 1294 11296 1328 11330
rect 1470 11364 1504 11398
rect 1470 11296 1504 11330
<< mvpdiffc >>
rect 1241 10789 1275 10823
rect 1241 10721 1275 10755
rect 1241 10653 1275 10687
rect 1417 10789 1451 10823
rect 1417 10721 1451 10755
rect 1417 10653 1451 10687
rect 1593 10789 1627 10823
rect 1593 10721 1627 10755
rect 1593 10653 1627 10687
<< psubdiff >>
rect 1586 11386 1620 11410
rect 1586 11316 1620 11352
rect 1586 11258 1620 11282
<< psubdiffcont >>
rect 1586 11352 1620 11386
rect 1586 11282 1620 11316
<< poly >>
rect 1339 11410 1459 11436
rect 1339 11244 1459 11270
rect 1343 11228 1477 11244
rect 1343 11194 1359 11228
rect 1393 11194 1427 11228
rect 1461 11194 1477 11228
rect 1343 11178 1477 11194
rect 1286 10835 1406 10861
rect 1462 10835 1582 10861
rect 1286 10602 1406 10635
rect 1462 10602 1582 10635
rect 1285 10586 1582 10602
rect 1285 10552 1301 10586
rect 1335 10552 1378 10586
rect 1412 10552 1455 10586
rect 1489 10552 1532 10586
rect 1566 10552 1582 10586
rect 1285 10536 1582 10552
<< polycont >>
rect 1359 11194 1393 11228
rect 1427 11194 1461 11228
rect 1301 10552 1335 10586
rect 1378 10552 1412 10586
rect 1455 10552 1489 10586
rect 1532 10552 1566 10586
<< locali >>
rect 1176 15232 1210 15270
rect 1294 11402 1328 11414
rect 1294 11330 1328 11364
rect 1294 11280 1328 11296
rect 1470 11398 1485 11414
rect 1519 11380 1586 11414
rect 1504 11364 1586 11380
rect 1470 11352 1586 11364
rect 1470 11342 1620 11352
rect 1470 11330 1485 11342
rect 1519 11308 1586 11342
rect 1504 11296 1586 11308
rect 1470 11282 1586 11296
rect 1470 11280 1620 11282
rect 1586 11258 1620 11280
rect 1343 11194 1344 11228
rect 1393 11194 1416 11228
rect 1461 11194 1477 11228
rect 1241 10823 1275 10837
rect 1241 10755 1275 10765
rect 1241 10687 1275 10721
rect 1417 10823 1451 10839
rect 1417 10755 1451 10789
rect 1417 10714 1451 10721
rect 1593 10823 1627 10837
rect 1593 10755 1627 10765
rect 1425 10687 1463 10714
rect 1451 10680 1463 10687
rect 1593 10687 1627 10721
rect 1241 10637 1275 10653
rect 1417 10637 1451 10653
rect 1593 10637 1627 10653
rect 1286 10586 1336 10593
rect 1286 10559 1301 10586
rect 1285 10552 1301 10559
rect 1335 10559 1336 10586
rect 1370 10586 1420 10593
rect 1370 10559 1378 10586
rect 1335 10552 1378 10559
rect 1412 10559 1420 10586
rect 1454 10586 1503 10593
rect 1454 10559 1455 10586
rect 1412 10552 1455 10559
rect 1489 10559 1503 10586
rect 1489 10552 1532 10559
rect 1566 10552 1582 10586
rect 14597 1107 14657 1143
rect 14706 801 14740 839
rect 14937 838 15009 850
rect 14937 800 15043 838
rect 15171 810 15209 844
rect 14937 766 15009 800
rect 14937 754 15013 766
rect 14597 511 14657 547
<< viali >>
rect 1176 15270 1210 15304
rect 1176 15198 1210 15232
rect 1294 11398 1328 11402
rect 1294 11368 1328 11398
rect 1294 11296 1328 11330
rect 1485 11398 1519 11414
rect 1485 11380 1504 11398
rect 1504 11380 1519 11398
rect 1586 11386 1620 11414
rect 1586 11380 1620 11386
rect 1485 11330 1519 11342
rect 1485 11308 1504 11330
rect 1504 11308 1519 11330
rect 1586 11316 1620 11342
rect 1586 11308 1620 11316
rect 1344 11194 1359 11228
rect 1359 11194 1378 11228
rect 1416 11194 1427 11228
rect 1427 11194 1450 11228
rect 1241 10837 1275 10871
rect 1241 10789 1275 10799
rect 1241 10765 1275 10789
rect 1593 10837 1627 10871
rect 1593 10789 1627 10799
rect 1593 10765 1627 10789
rect 1391 10687 1425 10714
rect 1391 10680 1417 10687
rect 1417 10680 1425 10687
rect 1463 10680 1497 10714
rect 1252 10559 1286 10593
rect 1336 10559 1370 10593
rect 1420 10559 1454 10593
rect 1503 10586 1537 10593
rect 1503 10559 1532 10586
rect 1532 10559 1537 10586
rect 14706 839 14740 873
rect 14706 767 14740 801
rect 15009 838 15043 872
rect 15137 810 15171 844
rect 15209 810 15243 844
rect 15009 766 15043 800
<< metal1 >>
rect 1689 16916 1717 16944
rect 1243 16169 1295 16175
rect 1243 16105 1295 16117
rect 1243 16047 1295 16053
rect 1818 16169 1870 16175
rect 1818 16105 1870 16117
tri 1870 16083 1896 16109 sw
rect 1870 16075 1896 16083
tri 1896 16075 1904 16083 sw
tri 2723 16075 2731 16083 se
rect 2731 16077 2783 16083
rect 1870 16053 2731 16075
rect 1818 16047 2731 16053
tri 2697 16013 2731 16047 ne
rect 2731 16013 2783 16025
rect 1327 15997 1379 16003
rect 1327 15933 1379 15945
rect 1327 15875 1379 15881
rect 1818 15997 2701 16003
rect 1870 15975 2649 15997
rect 1818 15933 1870 15945
tri 1870 15923 1922 15975 nw
tri 2615 15941 2649 15975 ne
rect 2731 15955 2783 15961
rect 2649 15933 2701 15945
rect 1818 15875 1870 15881
rect 2649 15875 2701 15881
rect 1170 15304 1216 15316
rect 1170 15270 1176 15304
rect 1210 15270 1216 15304
rect 1772 15295 1800 15323
rect 1170 15232 1216 15270
rect 1170 15198 1176 15232
rect 1210 15198 1216 15232
rect 1460 15212 1488 15240
rect 1170 15186 1216 15198
rect 1716 15162 1744 15190
rect 2043 15038 2579 15090
rect 2631 15038 2643 15090
rect 2695 15038 2701 15090
rect 2731 15055 2783 15061
tri 2699 14976 2731 15008 se
rect 2731 14991 2783 15003
rect 1226 14924 1232 14976
rect 1284 14924 1296 14976
rect 1348 14924 1354 14976
rect 2156 14970 2208 14976
tri 2697 14974 2699 14976 se
rect 2699 14974 2731 14976
rect 2088 14941 2116 14969
tri 2122 14924 2128 14930 ne
rect 2128 14924 2156 14930
tri 2128 14896 2156 14924 ne
rect 2406 14966 2731 14974
rect 2378 14939 2731 14966
rect 2783 14939 2788 14974
rect 2378 14938 2788 14939
rect 2406 14928 2788 14938
rect 2156 14906 2208 14918
rect 2156 14848 2208 14854
rect 2414 14295 2442 14323
rect 2265 11538 2293 11566
rect 3884 11473 3912 11501
rect 1479 11420 1835 11426
rect 1479 11414 1717 11420
rect 1288 11402 1421 11414
rect 1288 11368 1294 11402
rect 1328 11368 1421 11402
rect 1288 11330 1299 11368
rect 1288 11296 1294 11330
rect 1351 11316 1363 11368
rect 1415 11316 1421 11368
rect 1328 11296 1421 11316
rect 1479 11380 1485 11414
rect 1519 11380 1586 11414
rect 1620 11380 1717 11414
rect 1479 11368 1717 11380
rect 1769 11368 1783 11420
rect 3072 11397 3100 11425
rect 1479 11354 1835 11368
rect 1479 11342 1717 11354
rect 1479 11308 1485 11342
rect 1519 11308 1586 11342
rect 1620 11308 1717 11342
rect 1479 11302 1717 11308
rect 1769 11302 1783 11354
rect 1479 11296 1835 11302
rect 1288 11284 1421 11296
rect 1240 11248 1292 11254
tri 1292 11234 1312 11254 sw
rect 3420 11239 3448 11267
rect 1292 11228 1462 11234
rect 1292 11196 1344 11228
rect 1240 11194 1344 11196
rect 1378 11194 1416 11228
rect 1450 11194 1462 11228
rect 1240 11188 1462 11194
rect 1240 11184 1292 11188
tri 1292 11154 1326 11188 nw
rect 3614 11164 3654 11200
rect 1240 11126 1292 11132
tri 1240 11116 1250 11126 ne
rect 1250 11062 1282 11126
tri 1282 11116 1292 11126 nw
rect 1320 11078 1326 11130
rect 1378 11078 1390 11130
rect 1442 11127 1448 11130
tri 1448 11127 1451 11130 sw
rect 1442 11106 1451 11127
tri 1451 11106 1472 11127 sw
rect 3614 11106 3642 11164
rect 1442 11078 3642 11106
tri 3745 11089 3783 11127 se
rect 3783 11099 4126 11127
rect 3783 11089 3791 11099
tri 3791 11089 3801 11099 nw
tri 3737 11081 3745 11089 se
rect 3745 11081 3783 11089
tri 3783 11081 3791 11089 nw
rect 4332 11086 4338 11138
rect 4390 11086 4402 11138
rect 4454 11086 4460 11138
rect 4808 11089 4814 11141
rect 4866 11089 4878 11141
rect 4930 11089 4936 11141
tri 3734 11078 3737 11081 se
rect 3737 11078 3752 11081
tri 3732 11076 3734 11078 se
rect 3734 11076 3752 11078
tri 1250 11050 1262 11062 ne
rect 1262 11050 1282 11062
tri 1282 11050 1308 11076 sw
tri 3706 11050 3732 11076 se
rect 3732 11050 3752 11076
tri 3752 11050 3783 11081 nw
tri 1262 11030 1282 11050 ne
rect 1282 11030 3732 11050
tri 3732 11030 3752 11050 nw
tri 1282 11022 1290 11030 ne
rect 1290 11022 3724 11030
tri 3724 11022 3732 11030 nw
tri 1085 10871 1117 10903 ne
rect 1117 10871 1633 10903
tri 1117 10837 1151 10871 ne
rect 1151 10837 1241 10871
rect 1275 10837 1593 10871
rect 1627 10837 1633 10871
tri 1151 10799 1189 10837 ne
rect 1189 10799 1633 10837
tri 1189 10795 1193 10799 ne
rect 1193 10795 1241 10799
tri 1193 10767 1221 10795 ne
rect 1221 10767 1241 10795
tri 1221 10765 1223 10767 ne
rect 1223 10765 1241 10767
rect 1275 10765 1593 10799
rect 1627 10765 1633 10799
rect 1740 10767 1746 10819
rect 1798 10767 1810 10819
rect 1862 10795 1868 10819
rect 4801 10795 4807 10798
rect 1862 10767 4807 10795
tri 1223 10753 1235 10765 ne
rect 1235 10753 1633 10765
rect 4801 10746 4807 10767
rect 4859 10746 4871 10798
rect 4923 10746 4929 10798
rect 1315 10669 1321 10721
rect 1373 10669 1385 10721
rect 1437 10720 1443 10721
rect 1437 10714 1509 10720
rect 1437 10680 1463 10714
rect 1497 10680 1509 10714
rect 1437 10674 1509 10680
rect 1437 10669 1443 10674
rect 2903 10660 2909 10674
tri 1969 10636 1993 10660 se
rect 1993 10636 2909 10660
tri 1963 10630 1969 10636 se
rect 1969 10632 2909 10636
rect 1969 10630 1993 10632
rect 1240 10624 1292 10630
tri 1962 10629 1963 10630 se
rect 1963 10629 1993 10630
tri 1292 10616 1305 10629 sw
tri 1949 10616 1962 10629 se
rect 1962 10616 1993 10629
tri 1993 10616 2009 10632 nw
rect 2903 10622 2909 10632
rect 2961 10622 2973 10674
rect 3025 10636 4346 10674
rect 3025 10622 3031 10636
rect 4340 10622 4346 10636
rect 4398 10622 4410 10674
rect 4462 10622 4468 10674
rect 1292 10599 1305 10616
tri 1305 10599 1322 10616 sw
tri 1932 10599 1949 10616 se
rect 1292 10593 1549 10599
rect 1148 10567 1200 10573
rect 1148 10503 1200 10515
rect 1292 10572 1336 10593
rect 1240 10560 1252 10572
rect 1286 10560 1336 10572
rect 1292 10559 1336 10560
rect 1370 10559 1420 10593
rect 1454 10559 1503 10593
rect 1537 10559 1549 10593
tri 1905 10572 1932 10599 se
rect 1932 10572 1949 10599
tri 1949 10572 1993 10616 nw
rect 1292 10553 1549 10559
tri 1886 10553 1905 10572 se
rect 1292 10528 1301 10553
tri 1301 10528 1326 10553 nw
tri 1861 10528 1886 10553 se
rect 1886 10528 1905 10553
tri 1905 10528 1949 10572 nw
tri 1292 10519 1301 10528 nw
tri 1852 10519 1861 10528 se
rect 1240 10502 1292 10508
tri 1835 10502 1852 10519 se
rect 1852 10502 1861 10519
tri 1834 10501 1835 10502 se
rect 1835 10501 1861 10502
tri 1200 10484 1217 10501 sw
tri 1817 10484 1834 10501 se
rect 1834 10484 1861 10501
tri 1861 10484 1905 10528 nw
rect 1200 10473 1217 10484
tri 1217 10473 1228 10484 sw
tri 1806 10473 1817 10484 se
rect 1817 10473 1850 10484
tri 1850 10473 1861 10484 nw
rect 1200 10451 1822 10473
rect 1148 10445 1822 10451
tri 1822 10445 1850 10473 nw
rect 15305 2718 15311 2770
rect 15363 2718 15378 2770
rect 15430 2718 15444 2770
rect 15496 2718 15502 2770
rect 15305 2698 15502 2718
rect 15305 2646 15311 2698
rect 15363 2646 15378 2698
rect 15430 2646 15444 2698
rect 15496 2646 15502 2698
rect 15305 2626 15502 2646
rect 15305 2574 15311 2626
rect 15363 2574 15378 2626
rect 15430 2574 15444 2626
rect 15496 2574 15502 2626
rect 16316 2358 16344 2386
tri 16397 2339 16403 2345 ne
rect 16403 2339 16409 2391
rect 16461 2339 16473 2391
rect 16525 2339 16531 2391
tri 16531 2339 16537 2345 nw
rect 15008 1867 15014 1919
rect 15066 1867 15078 1919
rect 15130 1867 15136 1919
tri 15300 1873 15301 1874 se
tri 15136 1867 15142 1873 nw
tri 15294 1867 15300 1873 se
rect 15300 1867 15348 1873
tri 15252 1825 15294 1867 se
rect 15294 1825 15348 1867
rect 15134 1773 15140 1825
rect 15192 1773 15204 1825
rect 15256 1773 15348 1825
tri 15348 1773 15448 1873 nw
rect 16373 1799 16401 1827
rect 15578 1751 15606 1779
rect 16158 1723 16210 1729
rect 16158 1657 16210 1671
rect 16158 1599 16210 1605
rect 15661 1459 15689 1487
tri 15265 1227 15379 1341 se
rect 15379 1335 16531 1341
rect 15379 1283 16479 1335
rect 15379 1271 16531 1283
rect 15379 1227 16479 1271
tri 14775 1213 14789 1227 se
rect 14789 1213 14795 1227
tri 14771 1209 14775 1213 se
rect 14775 1209 14795 1213
rect 14789 1175 14795 1209
rect 14847 1175 14860 1227
rect 14789 1163 14860 1175
tri 14230 1111 14236 1117 sw
rect 14789 1111 14795 1163
rect 14847 1111 14860 1163
rect 14976 1213 14982 1227
tri 14982 1213 14996 1227 sw
tri 15251 1213 15265 1227 se
rect 15265 1219 16479 1227
rect 15265 1213 16531 1219
rect 14976 1209 14996 1213
tri 14996 1209 15000 1213 sw
tri 15247 1209 15251 1213 se
rect 15251 1209 15391 1213
tri 15391 1209 15395 1213 nw
rect 14976 1183 14982 1209
rect 15293 1183 15365 1209
tri 15365 1183 15391 1209 nw
rect 14976 1155 14983 1183
rect 15293 1155 15337 1183
tri 15337 1155 15365 1183 nw
rect 14976 1111 14982 1155
tri 15293 1111 15337 1155 nw
rect 14230 1079 14236 1111
tri 14236 1079 14268 1111 sw
rect 14230 1027 15312 1079
rect 15364 1027 15378 1079
rect 15430 1027 15444 1079
rect 15496 1027 15502 1079
rect 14230 967 15502 1027
rect 14230 915 15312 967
rect 15364 915 15378 967
rect 15430 915 15444 967
rect 15496 915 15502 967
rect 14696 875 14908 885
rect 14696 873 14856 875
rect 14696 839 14706 873
rect 14740 839 14856 873
rect 14696 823 14856 839
rect 14696 811 14908 823
rect 14696 801 14856 811
rect 14696 767 14706 801
rect 14740 767 14856 801
rect 14696 759 14856 767
rect 14696 753 14908 759
rect 15000 878 15052 884
rect 15000 814 15052 826
rect 15125 844 15255 850
rect 15125 810 15137 844
rect 15171 810 15209 844
rect 15243 810 15255 844
rect 15125 804 15255 810
rect 15000 754 15052 762
rect 14816 486 14844 514
rect 15293 445 16206 543
tri 16710 -367 16766 -311 se
rect 15995 -369 16766 -367
rect 15995 -421 16001 -369
rect 16053 -421 16065 -369
rect 16117 -421 16766 -369
rect 15995 -423 16766 -421
<< via1 >>
rect 1243 16117 1295 16169
rect 1243 16053 1295 16105
rect 1818 16117 1870 16169
rect 1818 16053 1870 16105
rect 2731 16025 2783 16077
rect 1327 15945 1379 15997
rect 1327 15881 1379 15933
rect 1818 15945 1870 15997
rect 1818 15881 1870 15933
rect 2649 15945 2701 15997
rect 2731 15961 2783 16013
rect 2649 15881 2701 15933
rect 2579 15038 2631 15090
rect 2643 15038 2695 15090
rect 2731 15003 2783 15055
rect 1232 14924 1284 14976
rect 1296 14924 1348 14976
rect 2156 14918 2208 14970
rect 2731 14939 2783 14991
rect 2156 14854 2208 14906
rect 1299 11330 1351 11368
rect 1299 11316 1328 11330
rect 1328 11316 1351 11330
rect 1363 11316 1415 11368
rect 1717 11368 1769 11420
rect 1783 11368 1835 11420
rect 1717 11302 1769 11354
rect 1783 11302 1835 11354
rect 1240 11196 1292 11248
rect 1240 11132 1292 11184
rect 1326 11078 1378 11130
rect 1390 11078 1442 11130
rect 4338 11086 4390 11138
rect 4402 11086 4454 11138
rect 4814 11089 4866 11141
rect 4878 11089 4930 11141
rect 1746 10767 1798 10819
rect 1810 10767 1862 10819
rect 4807 10746 4859 10798
rect 4871 10746 4923 10798
rect 1321 10669 1373 10721
rect 1385 10714 1437 10721
rect 1385 10680 1391 10714
rect 1391 10680 1425 10714
rect 1425 10680 1437 10714
rect 1385 10669 1437 10680
rect 1240 10593 1292 10624
rect 2909 10622 2961 10674
rect 2973 10622 3025 10674
rect 4346 10622 4398 10674
rect 4410 10622 4462 10674
rect 1148 10515 1200 10567
rect 1148 10451 1200 10503
rect 1240 10572 1252 10593
rect 1252 10572 1286 10593
rect 1286 10572 1292 10593
rect 1240 10559 1252 10560
rect 1252 10559 1286 10560
rect 1286 10559 1292 10560
rect 1240 10508 1292 10559
rect 15311 2718 15363 2770
rect 15378 2718 15430 2770
rect 15444 2718 15496 2770
rect 15311 2646 15363 2698
rect 15378 2646 15430 2698
rect 15444 2646 15496 2698
rect 15311 2574 15363 2626
rect 15378 2574 15430 2626
rect 15444 2574 15496 2626
rect 16409 2339 16461 2391
rect 16473 2339 16525 2391
rect 15014 1867 15066 1919
rect 15078 1867 15130 1919
rect 15140 1773 15192 1825
rect 15204 1773 15256 1825
rect 16158 1671 16210 1723
rect 16158 1605 16210 1657
rect 16479 1283 16531 1335
rect 14795 1175 14847 1227
rect 14795 1111 14847 1163
rect 14860 1111 14976 1227
rect 16479 1219 16531 1271
rect 15312 1027 15364 1079
rect 15378 1027 15430 1079
rect 15444 1027 15496 1079
rect 15312 915 15364 967
rect 15378 915 15430 967
rect 15444 915 15496 967
rect 14856 823 14908 875
rect 14856 759 14908 811
rect 15000 872 15052 878
rect 15000 838 15009 872
rect 15009 838 15043 872
rect 15043 838 15052 872
rect 15000 826 15052 838
rect 15000 800 15052 814
rect 15000 766 15009 800
rect 15009 766 15043 800
rect 15043 766 15052 800
rect 15000 762 15052 766
rect 16001 -421 16053 -369
rect 16065 -421 16117 -369
<< metal2 >>
rect 1243 16169 1295 16175
rect 1818 16169 1870 16175
tri 1804 16134 1818 16148 se
tri 1295 16117 1312 16134 sw
tri 1787 16117 1804 16134 se
rect 1804 16117 1818 16134
rect 1243 16105 1312 16117
tri 1312 16105 1324 16117 sw
tri 1775 16105 1787 16117 se
rect 1787 16105 1870 16117
rect 1295 16084 1324 16105
tri 1324 16084 1345 16105 sw
tri 1754 16084 1775 16105 se
rect 1775 16084 1818 16105
rect 1295 16053 1818 16084
rect 1243 16047 1870 16053
rect 2731 16077 2783 16083
rect 2731 16013 2783 16025
rect 1327 15997 1870 16003
rect 1379 15975 1818 15997
rect 1379 15945 1405 15975
tri 1405 15945 1435 15975 nw
tri 1763 15945 1793 15975 ne
rect 1793 15945 1818 15975
rect 1327 15933 1393 15945
tri 1393 15933 1405 15945 nw
tri 1793 15933 1805 15945 ne
rect 1805 15933 1870 15945
tri 1379 15919 1393 15933 nw
tri 1805 15920 1818 15933 ne
rect 1327 15875 1379 15881
rect 1818 15875 1870 15881
rect 2649 15997 2701 16003
rect 2649 15933 2701 15945
tri 2615 15090 2649 15124 se
rect 2649 15090 2701 15881
rect 2573 15038 2579 15090
rect 2631 15038 2643 15090
rect 2695 15038 2701 15090
rect 2731 15055 2783 15961
rect 2731 14991 2783 15003
rect 2156 14981 2212 14990
rect 1160 14924 1232 14976
rect 1284 14924 1296 14976
rect 1348 14924 1354 14976
rect 2731 14933 2783 14939
rect 1160 10573 1200 14924
rect 2208 14918 2212 14925
rect 2156 14906 2212 14918
rect 2208 14901 2212 14906
rect 2156 14836 2212 14845
tri 1717 11774 1719 11776 ne
rect 1719 11774 1868 11776
tri 1868 11774 1870 11776 nw
rect 1719 11426 1835 11774
tri 1835 11741 1868 11774 nw
rect 1717 11420 1835 11426
rect 1769 11368 1783 11420
rect 1293 11316 1299 11368
rect 1351 11316 1363 11368
rect 1415 11316 1421 11368
rect 1148 10567 1200 10573
rect 1148 10503 1200 10515
rect 1240 11248 1292 11254
rect 1240 11184 1292 11196
rect 1240 11126 1292 11132
rect 1381 11130 1421 11316
rect 1717 11354 1835 11368
rect 1769 11302 1783 11354
rect 1717 11296 1835 11302
rect 1240 10630 1286 11126
rect 1320 11078 1326 11130
rect 1378 11078 1390 11130
rect 1442 11078 1448 11130
rect 4332 11086 4338 11138
rect 4390 11086 4402 11138
rect 4454 11086 4460 11138
rect 4808 11089 4814 11141
rect 4866 11089 4878 11141
rect 4930 11089 4936 11141
rect 1381 10721 1421 11078
rect 1778 10912 1834 10921
tri 1744 10819 1778 10853 se
rect 1778 10832 1834 10856
tri 1834 10819 1868 10853 sw
rect 1740 10767 1746 10819
rect 1798 10767 1810 10776
rect 1862 10767 1868 10819
rect 1315 10669 1321 10721
rect 1373 10669 1385 10721
rect 1437 10669 1443 10721
rect 2903 10674 2912 10676
rect 2968 10674 2992 10676
rect 1240 10624 1292 10630
rect 2903 10622 2909 10674
rect 2968 10622 2973 10674
rect 2903 10620 2912 10622
rect 2968 10620 2992 10622
rect 3048 10620 3057 10676
rect 4342 10674 4380 11086
rect 4831 10798 4859 11089
rect 4801 10746 4807 10798
rect 4859 10746 4871 10798
rect 4923 10746 4929 10798
rect 4340 10622 4346 10674
rect 4398 10622 4410 10674
rect 4462 10622 4468 10674
rect 1240 10560 1292 10572
rect 1240 10502 1292 10508
rect 1148 10445 1200 10451
rect 16390 7730 16446 7739
rect 16095 7674 16390 7707
rect 16095 7661 16446 7674
rect 16095 5106 16141 7661
rect 16390 7650 16446 7661
rect 16390 7585 16446 7594
tri 16141 5106 16161 5126 sw
tri 16095 5040 16161 5106 ne
tri 16161 5040 16227 5106 sw
tri 16161 4974 16227 5040 ne
tri 16227 4980 16287 5040 sw
rect 16227 4974 16287 4980
tri 16287 4974 16293 4980 sw
tri 16227 4914 16287 4974 ne
rect 16287 4934 16293 4974
tri 16293 4934 16333 4974 sw
tri 16221 2975 16287 3041 se
rect 16287 3021 16333 4934
tri 16287 2975 16333 3021 nw
tri 16164 2918 16221 2975 se
rect 16221 2918 16230 2975
tri 16230 2918 16287 2975 nw
rect 15305 2718 15311 2770
rect 15363 2718 15378 2770
rect 15430 2718 15444 2770
rect 15496 2718 15502 2770
rect 15305 2698 15502 2718
rect 15305 2646 15311 2698
rect 15363 2646 15378 2698
rect 15430 2646 15444 2698
rect 15496 2646 15502 2698
rect 15305 2626 15502 2646
rect 15305 2574 15311 2626
rect 15363 2574 15378 2626
rect 15430 2574 15444 2626
rect 15496 2574 15502 2626
rect 15008 1867 15014 1919
rect 15066 1867 15078 1919
rect 15130 1867 15136 1919
tri 15008 1850 15025 1867 ne
rect 15025 1850 15119 1867
tri 15119 1850 15136 1867 nw
rect 15025 1825 15094 1850
tri 15094 1825 15119 1850 nw
rect 14789 1377 14983 1386
rect 14845 1321 14927 1377
rect 14789 1277 14983 1321
rect 14845 1227 14927 1277
rect 14789 1176 14795 1221
rect 14847 1175 14860 1227
rect 14976 1176 14983 1221
rect 14845 1163 14860 1175
rect 14789 1111 14795 1120
rect 14847 1111 14860 1163
rect 14976 1111 14983 1120
tri 15017 1027 15025 1035 se
rect 15025 1027 15077 1825
tri 15077 1808 15094 1825 nw
rect 15134 1773 15140 1825
rect 15192 1773 15204 1825
rect 15256 1773 15262 1825
tri 15134 1723 15184 1773 ne
rect 15184 1723 15237 1773
tri 15237 1748 15262 1773 nw
tri 15184 1722 15185 1723 ne
tri 15161 1027 15185 1051 se
rect 15185 1029 15237 1723
rect 15185 1027 15235 1029
tri 15235 1027 15237 1029 nw
rect 15305 1079 15502 2574
tri 16158 1729 16164 1735 se
rect 16164 1729 16210 2918
tri 16210 2898 16230 2918 nw
rect 16403 2339 16409 2391
rect 16461 2339 16473 2391
rect 16525 2339 16531 2391
tri 16445 2305 16479 2339 ne
rect 16158 1723 16210 1729
rect 16158 1657 16210 1671
rect 16158 1599 16210 1605
rect 16479 1335 16531 2339
rect 16479 1271 16531 1283
rect 16479 1213 16531 1219
rect 15305 1027 15312 1079
rect 15364 1027 15378 1079
rect 15430 1027 15444 1079
rect 15496 1027 15502 1079
tri 14967 977 15017 1027 se
rect 15017 1013 15077 1027
rect 15017 977 15041 1013
tri 15041 977 15077 1013 nw
tri 15111 977 15161 1027 se
rect 15161 977 15185 1027
tri 15185 977 15235 1027 nw
tri 14957 967 14967 977 se
rect 14967 967 15031 977
tri 15031 967 15041 977 nw
tri 15101 967 15111 977 se
rect 15111 967 15175 977
tri 15175 967 15185 977 nw
rect 15305 967 15502 1027
tri 14951 961 14957 967 se
rect 14957 961 15025 967
tri 15025 961 15031 967 nw
tri 15095 961 15101 967 se
rect 15101 961 15123 967
tri 14905 915 14951 961 se
rect 14951 915 14979 961
tri 14979 915 15025 961 nw
tri 15049 915 15095 961 se
rect 15095 915 15123 961
tri 15123 915 15175 967 nw
rect 15305 915 15312 967
rect 15364 915 15378 967
rect 15430 915 15444 967
rect 15496 915 15502 967
tri 14893 903 14905 915 se
rect 14905 903 14967 915
tri 14967 903 14979 915 nw
tri 15037 903 15049 915 se
rect 15049 903 15111 915
tri 15111 903 15123 915 nw
tri 14877 887 14893 903 se
rect 14893 891 14955 903
tri 14955 891 14967 903 nw
tri 15025 891 15037 903 se
rect 15037 891 15092 903
rect 14893 887 14951 891
tri 14951 887 14955 891 nw
tri 15021 887 15025 891 se
rect 15025 887 15092 891
tri 14874 884 14877 887 se
rect 14877 884 14948 887
tri 14948 884 14951 887 nw
tri 15018 884 15021 887 se
rect 15021 884 15092 887
tri 15092 884 15111 903 nw
tri 14871 881 14874 884 se
rect 14874 881 14945 884
tri 14945 881 14948 884 nw
rect 14856 878 14942 881
tri 14942 878 14945 881 nw
rect 15000 878 15052 884
rect 14856 875 14908 878
tri 14908 844 14942 878 nw
rect 14856 811 14908 823
rect 14856 753 14908 759
tri 15052 844 15092 884 nw
rect 15000 814 15052 826
rect 15000 756 15052 762
rect 15969 -423 15978 -367
rect 16034 -369 16058 -367
rect 16114 -369 16123 -367
rect 16053 -421 16058 -369
rect 16117 -421 16123 -369
rect 16034 -423 16058 -421
rect 16114 -423 16123 -421
<< via2 >>
rect 2156 14970 2212 14981
rect 2156 14925 2208 14970
rect 2208 14925 2212 14970
rect 2156 14854 2208 14901
rect 2208 14854 2212 14901
rect 2156 14845 2212 14854
rect 1778 10856 1834 10912
rect 1778 10819 1834 10832
rect 1778 10776 1798 10819
rect 1798 10776 1810 10819
rect 1810 10776 1834 10819
rect 2912 10674 2968 10676
rect 2992 10674 3048 10676
rect 2912 10622 2961 10674
rect 2961 10622 2968 10674
rect 2992 10622 3025 10674
rect 3025 10622 3048 10674
rect 2912 10620 2968 10622
rect 2992 10620 3048 10622
rect 16390 7674 16446 7730
rect 16390 7594 16446 7650
rect 14789 1321 14845 1377
rect 14927 1321 14983 1377
rect 14789 1227 14845 1277
rect 14927 1227 14983 1277
rect 14789 1221 14795 1227
rect 14795 1221 14845 1227
rect 14789 1175 14795 1176
rect 14795 1175 14845 1176
rect 14927 1221 14976 1227
rect 14976 1221 14983 1227
rect 14789 1163 14845 1175
rect 14789 1120 14795 1163
rect 14795 1120 14845 1163
rect 14927 1120 14976 1176
rect 14976 1120 14983 1176
rect 15978 -369 16034 -367
rect 16058 -369 16114 -367
rect 15978 -421 16001 -369
rect 16001 -421 16034 -369
rect 16058 -421 16065 -369
rect 16065 -421 16114 -369
rect 15978 -423 16034 -421
rect 16058 -423 16114 -421
<< metal3 >>
rect 2151 14981 2217 14990
rect 2151 14925 2156 14981
rect 2212 14925 2217 14981
rect 2151 14901 2217 14925
rect 2151 14845 2156 14901
rect 2212 14845 2217 14901
tri 2123 14801 2151 14829 se
rect 2151 14801 2217 14845
tri 2121 14799 2123 14801 se
rect 2123 14799 2215 14801
tri 2215 14799 2217 14801 nw
tri 2027 14705 2121 14799 se
tri 2121 14705 2215 14799 nw
tri 1933 14611 2027 14705 se
tri 2027 14611 2121 14705 nw
tri 1839 14517 1933 14611 se
tri 1933 14517 2027 14611 nw
tri 1773 14451 1839 14517 se
rect 1773 10912 1839 14451
tri 1839 14423 1933 14517 nw
rect 1773 10856 1778 10912
rect 1834 10856 1839 10912
rect 1773 10832 1839 10856
rect 1773 10776 1778 10832
rect 1834 10776 1839 10832
rect 1773 7114 1839 10776
rect 2907 10676 3053 10681
rect 2907 10620 2912 10676
rect 2968 10620 2992 10676
rect 3048 10620 3053 10676
rect 2907 10615 3053 10620
tri 2907 10600 2922 10615 ne
rect 2922 10600 3038 10615
tri 3038 10600 3053 10615 nw
tri 2892 7735 2922 7765 se
rect 2922 7735 2988 10600
tri 2988 10550 3038 10600 nw
tri 2887 7730 2892 7735 se
rect 2892 7730 2988 7735
tri 2851 7694 2887 7730 se
rect 2887 7694 2988 7730
rect 16385 7730 16541 7735
tri 2988 7694 3007 7713 sw
rect 2851 7630 2857 7694
rect 2921 7630 2937 7694
rect 3001 7630 3007 7694
rect 16385 7674 16390 7730
rect 16446 7694 16541 7730
rect 16385 7650 16391 7674
rect 16385 7594 16390 7650
rect 16455 7630 16471 7694
rect 16535 7630 16541 7694
rect 16446 7594 16541 7630
rect 16385 7589 16541 7594
tri 1773 7103 1784 7114 ne
rect 1784 7103 1839 7114
tri 1839 7103 1878 7142 sw
tri 1784 7048 1839 7103 ne
rect 1839 7048 1878 7103
tri 1839 7009 1878 7048 ne
tri 1878 7009 1972 7103 sw
tri 1878 6915 1972 7009 ne
tri 1972 6915 2066 7009 sw
tri 1972 6821 2066 6915 ne
tri 2066 6821 2160 6915 sw
tri 2066 6727 2160 6821 ne
tri 2160 6727 2254 6821 sw
tri 2160 6633 2254 6727 ne
tri 2254 6633 2348 6727 sw
tri 2254 6605 2282 6633 ne
tri 2270 1277 2282 1289 se
rect 2282 1277 2348 6633
tri 2220 1227 2270 1277 se
rect 2270 1261 2348 1277
rect 2270 1227 2314 1261
tri 2314 1227 2348 1261 nw
rect 14510 2356 14996 2491
tri 14996 2356 15131 2491 sw
rect 14510 1377 15131 2356
rect 14510 1321 14789 1377
rect 14845 1321 14927 1377
rect 14983 1321 15131 1377
rect 14510 1277 15131 1321
tri 1787 1221 1793 1227 se
rect 1793 1221 2308 1227
tri 2308 1221 2314 1227 nw
rect 14510 1221 14789 1277
rect 14845 1221 14927 1277
rect 14983 1221 15131 1277
tri 1742 1176 1787 1221 se
rect 1787 1176 2263 1221
tri 2263 1176 2308 1221 nw
rect 14510 1176 15131 1221
tri 1699 1133 1742 1176 se
rect 1742 1161 2248 1176
tri 2248 1161 2263 1176 nw
rect 1742 1133 1793 1161
tri 1793 1133 1821 1161 nw
tri 1686 1120 1699 1133 se
rect 1699 1120 1780 1133
tri 1780 1120 1793 1133 nw
rect 14510 1120 14789 1176
rect 14845 1120 14927 1176
rect 14983 1120 15131 1176
tri 1680 1114 1686 1120 se
rect 1686 1114 1774 1120
tri 1774 1114 1780 1120 nw
tri 1670 -363 1680 -353 se
rect 1680 -363 1746 1114
tri 1746 1086 1774 1114 nw
rect 14510 1111 15131 1120
tri 1746 -363 1826 -283 sw
rect 1670 -427 1676 -363
rect 1740 -427 1756 -363
rect 1820 -427 1826 -363
rect 15973 -363 16119 -362
rect 15973 -367 15979 -363
rect 16043 -367 16059 -363
rect 15973 -423 15978 -367
rect 16043 -423 16058 -367
rect 15973 -427 15979 -423
rect 16043 -427 16059 -423
rect 16123 -427 16129 -363
rect 15973 -428 16119 -427
<< via3 >>
rect 2857 7630 2921 7694
rect 2937 7630 3001 7694
rect 16391 7674 16446 7694
rect 16446 7674 16455 7694
rect 16391 7650 16455 7674
rect 16391 7630 16446 7650
rect 16446 7630 16455 7650
rect 16471 7630 16535 7694
rect 1676 -427 1740 -363
rect 1756 -427 1820 -363
rect 15979 -367 16043 -363
rect 16059 -367 16123 -363
rect 15979 -423 16034 -367
rect 16034 -423 16043 -367
rect 16059 -423 16114 -367
rect 16114 -423 16123 -367
rect 15979 -427 16043 -423
rect 16059 -427 16123 -423
<< metal4 >>
rect 2856 7694 16536 7695
rect 2856 7630 2857 7694
rect 2921 7630 2937 7694
rect 3001 7630 16391 7694
rect 16455 7630 16471 7694
rect 16535 7630 16536 7694
rect 2856 7629 16536 7630
rect 1675 -363 16124 -362
rect 1675 -427 1676 -363
rect 1740 -427 1756 -363
rect 1820 -427 15979 -363
rect 16043 -427 16059 -363
rect 16123 -427 16124 -363
rect 1675 -428 16124 -427
use sky130_fd_io__gpiov2_amux_ctl_inv_1  sky130_fd_io__gpiov2_amux_ctl_inv_1_0
timestamp 1666464484
transform -1 0 14983 0 1 494
box -19 -49 346 715
use sky130_fd_io__gpiov2_amux_ctl_inv_1  sky130_fd_io__gpiov2_amux_ctl_inv_1_1
timestamp 1666464484
transform -1 0 15292 0 1 494
box -19 -49 346 715
use sky130_fd_io__gpiov2_amux_ctl_ls  sky130_fd_io__gpiov2_amux_ctl_ls_0
timestamp 1666464484
transform 1 0 14705 0 1 1344
box 53 10 2203 1486
use sky130_fd_io__gpiov2_amux_ctl_lshv2hv2  sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0
timestamp 1666464484
transform 1 0 748 0 1 13628
box 172 529 4053 3493
use sky130_fd_io__gpiov2_amux_ctl_lshv2hv  sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0
timestamp 1666464484
transform -1 0 8787 0 1 10523
box 3486 559 6918 1429
use sky130_fd_io__tap_1  sky130_fd_io__tap_1_0
timestamp 1666464484
transform -1 0 14675 0 1 494
box -38 -49 134 715
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808586  sky130_fd_pr__model__nfet_highvoltage__example_55959141808586_0
timestamp 1666464484
transform -1 0 1459 0 -1 11410
box -1 0 121 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808421  sky130_fd_pr__model__pfet_highvoltage__example_55959141808421_0
timestamp 1666464484
transform 1 0 1286 0 -1 10835
box -1 0 297 1
<< labels >>
flabel metal1 s 15194 813 15222 841 3 FreeSans 280 0 0 0 ANALOG_EN
port 1 nsew
flabel metal1 s 16373 1799 16401 1827 3 FreeSans 520 0 0 0 HLD_I_H
port 2 nsew
flabel metal1 s 15578 1751 15606 1779 3 FreeSans 520 0 0 0 HLD_I_H_N
port 3 nsew
flabel metal1 s 15349 2685 15377 2713 3 FreeSans 520 0 0 0 VDDIO_Q
port 4 nsew
flabel metal1 s 2265 11538 2293 11566 3 FreeSans 520 0 0 0 VSWITCH
port 5 nsew
flabel metal1 s 3072 11397 3100 11425 3 FreeSans 520 0 0 0 AMUX_EN_VSWITCH_H
port 6 nsew
flabel metal1 s 1460 15212 1488 15240 3 FreeSans 520 0 0 0 AMUX_EN_VDDA_H_N
port 7 nsew
flabel metal1 s 1716 15162 1744 15190 3 FreeSans 520 0 0 0 VSSA
port 8 nsew
flabel metal1 s 3420 11239 3448 11267 3 FreeSans 520 0 0 0 AMUX_EN_VSWITCH_H_N
port 9 nsew
flabel metal1 s 4098 11099 4126 11127 3 FreeSans 520 0 0 0 ENABLE_VSWITCH_H
port 10 nsew
flabel metal1 s 2088 14941 2116 14969 3 FreeSans 520 0 0 0 AMUX_EN_VDDIO_H_N
port 11 nsew
flabel metal1 s 1266 14942 1294 14970 3 FreeSans 520 0 0 0 AMUX_EN_VDDIO_H
port 12 nsew
flabel metal1 s 1388 10863 1416 10891 3 FreeSans 520 0 0 0 VSWITCH
port 5 nsew
flabel metal1 s 1772 15295 1800 15323 3 FreeSans 520 0 0 0 AMUX_EN_VDDA_H
port 13 nsew
flabel metal1 s 3884 11473 3912 11501 3 FreeSans 520 0 0 0 VSSA
port 8 nsew
flabel metal1 s 2414 14295 2442 14323 3 FreeSans 520 0 0 0 VSSA
port 8 nsew
flabel metal1 s 2378 14938 2406 14966 3 FreeSans 520 0 0 0 ENABLE_VDDA_H
port 14 nsew
flabel metal1 s 1689 16916 1717 16944 3 FreeSans 520 0 0 0 VDDA
port 15 nsew
flabel metal1 s 1719 11339 1747 11367 3 FreeSans 520 0 0 0 VSSA
port 8 nsew
flabel metal1 s 15661 1459 15689 1487 3 FreeSans 280 180 0 0 VSSD
port 16 nsew
flabel metal1 s 1176 15213 1204 15241 3 FreeSans 520 0 0 0 VSSA
port 8 nsew
flabel metal1 s 16316 2358 16344 2386 3 FreeSans 280 180 0 0 VCCD
port 17 nsew
flabel metal1 s 14816 486 14844 514 3 FreeSans 280 0 0 0 VSSD
port 16 nsew
flabel metal1 s 14955 1155 14983 1183 3 FreeSans 280 0 0 0 VCCD
port 17 nsew
<< properties >>
string GDS_END 43861080
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43835424
<< end >>
