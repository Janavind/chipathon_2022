magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1471 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 487 47 517 177
rect 682 47 712 177
rect 775 47 805 177
rect 859 47 889 177
rect 963 47 993 177
rect 1082 47 1112 177
rect 1183 47 1213 177
rect 1270 47 1300 177
rect 1359 47 1389 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 651 297 681 497
rect 736 297 766 497
rect 822 297 852 497
rect 923 297 953 497
rect 1111 297 1141 497
rect 1195 297 1225 497
rect 1279 297 1309 497
rect 1363 297 1393 497
<< ndiff >>
rect 27 101 79 177
rect 27 67 35 101
rect 69 67 79 101
rect 27 47 79 67
rect 109 169 163 177
rect 109 135 119 169
rect 153 135 163 169
rect 109 47 163 135
rect 193 93 247 177
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 47 331 177
rect 361 169 415 177
rect 361 135 371 169
rect 405 135 415 169
rect 361 47 415 135
rect 445 47 487 177
rect 517 93 569 177
rect 517 59 527 93
rect 561 59 569 93
rect 517 47 569 59
rect 630 93 682 177
rect 630 59 638 93
rect 672 59 682 93
rect 630 47 682 59
rect 712 169 775 177
rect 712 135 731 169
rect 765 135 775 169
rect 712 101 775 135
rect 712 67 731 101
rect 765 67 775 101
rect 712 47 775 67
rect 805 93 859 177
rect 805 59 815 93
rect 849 59 859 93
rect 805 47 859 59
rect 889 169 963 177
rect 889 135 909 169
rect 943 135 963 169
rect 889 101 963 135
rect 889 67 909 101
rect 943 67 963 101
rect 889 47 963 67
rect 993 93 1082 177
rect 993 59 1013 93
rect 1047 59 1082 93
rect 993 47 1082 59
rect 1112 101 1183 177
rect 1112 67 1139 101
rect 1173 67 1183 101
rect 1112 47 1183 67
rect 1213 89 1270 177
rect 1213 55 1225 89
rect 1259 55 1270 89
rect 1213 47 1270 55
rect 1300 101 1359 177
rect 1300 67 1311 101
rect 1345 67 1359 101
rect 1300 47 1359 67
rect 1389 93 1445 177
rect 1389 59 1399 93
rect 1433 59 1445 93
rect 1389 47 1445 59
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 297 163 451
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 409 247 443
rect 193 375 203 409
rect 237 375 247 409
rect 193 297 247 375
rect 277 489 331 497
rect 277 455 287 489
rect 321 455 331 489
rect 277 297 331 455
rect 361 477 415 497
rect 361 443 371 477
rect 405 443 415 477
rect 361 297 415 443
rect 445 489 499 497
rect 445 455 455 489
rect 489 455 499 489
rect 445 297 499 455
rect 529 477 651 497
rect 529 443 539 477
rect 573 443 607 477
rect 641 443 651 477
rect 529 409 651 443
rect 529 375 607 409
rect 641 375 651 409
rect 529 297 651 375
rect 681 297 736 497
rect 766 489 822 497
rect 766 455 777 489
rect 811 455 822 489
rect 766 297 822 455
rect 852 297 923 497
rect 953 477 1005 497
rect 953 443 963 477
rect 997 443 1005 477
rect 953 409 1005 443
rect 953 375 963 409
rect 997 375 1005 409
rect 953 297 1005 375
rect 1059 485 1111 497
rect 1059 451 1067 485
rect 1101 451 1111 485
rect 1059 297 1111 451
rect 1141 477 1195 497
rect 1141 443 1151 477
rect 1185 443 1195 477
rect 1141 409 1195 443
rect 1141 375 1151 409
rect 1185 375 1195 409
rect 1141 297 1195 375
rect 1225 485 1279 497
rect 1225 451 1235 485
rect 1269 451 1279 485
rect 1225 417 1279 451
rect 1225 383 1235 417
rect 1269 383 1279 417
rect 1225 297 1279 383
rect 1309 477 1363 497
rect 1309 443 1319 477
rect 1353 443 1363 477
rect 1309 409 1363 443
rect 1309 375 1319 409
rect 1353 375 1363 409
rect 1309 297 1363 375
rect 1393 485 1445 497
rect 1393 451 1403 485
rect 1437 451 1445 485
rect 1393 417 1445 451
rect 1393 383 1403 417
rect 1437 383 1445 417
rect 1393 297 1445 383
<< ndiffc >>
rect 35 67 69 101
rect 119 135 153 169
rect 203 59 237 93
rect 371 135 405 169
rect 527 59 561 93
rect 638 59 672 93
rect 731 135 765 169
rect 731 67 765 101
rect 815 59 849 93
rect 909 135 943 169
rect 909 67 943 101
rect 1013 59 1047 93
rect 1139 67 1173 101
rect 1225 55 1259 89
rect 1311 67 1345 101
rect 1399 59 1433 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 451 153 485
rect 203 443 237 477
rect 203 375 237 409
rect 287 455 321 489
rect 371 443 405 477
rect 455 455 489 489
rect 539 443 573 477
rect 607 443 641 477
rect 607 375 641 409
rect 777 455 811 489
rect 963 443 997 477
rect 963 375 997 409
rect 1067 451 1101 485
rect 1151 443 1185 477
rect 1151 375 1185 409
rect 1235 451 1269 485
rect 1235 383 1269 417
rect 1319 443 1353 477
rect 1319 375 1353 409
rect 1403 451 1437 485
rect 1403 383 1437 417
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 651 497 681 523
rect 736 497 766 523
rect 822 497 852 523
rect 923 497 953 523
rect 1111 497 1141 523
rect 1195 497 1225 523
rect 1279 497 1309 523
rect 1363 497 1393 523
rect 79 265 109 297
rect 24 259 109 265
rect 163 259 193 297
rect 247 265 277 297
rect 24 249 193 259
rect 24 215 34 249
rect 68 215 193 249
rect 24 205 193 215
rect 24 199 109 205
rect 79 177 109 199
rect 163 177 193 205
rect 235 249 289 265
rect 235 215 245 249
rect 279 215 289 249
rect 235 199 289 215
rect 331 259 361 297
rect 415 259 445 297
rect 499 261 529 297
rect 499 259 564 261
rect 651 259 681 297
rect 736 282 766 297
rect 822 282 852 297
rect 331 249 445 259
rect 331 215 371 249
rect 405 215 445 249
rect 331 205 445 215
rect 247 177 277 199
rect 331 177 361 205
rect 415 177 445 205
rect 487 249 564 259
rect 487 215 514 249
rect 548 215 564 249
rect 487 203 564 215
rect 627 249 693 259
rect 736 258 852 282
rect 747 251 852 258
rect 923 281 953 297
rect 923 259 961 281
rect 1111 259 1141 297
rect 1195 259 1225 297
rect 1279 259 1309 297
rect 1363 259 1393 297
rect 923 252 997 259
rect 627 215 643 249
rect 677 220 693 249
rect 775 249 852 251
rect 677 215 712 220
rect 627 205 712 215
rect 487 177 517 203
rect 629 192 712 205
rect 682 177 712 192
rect 775 215 794 249
rect 828 227 852 249
rect 931 249 997 252
rect 828 215 889 227
rect 775 197 889 215
rect 931 215 947 249
rect 981 215 997 249
rect 931 205 997 215
rect 1082 249 1393 259
rect 1082 215 1098 249
rect 1132 215 1166 249
rect 1200 215 1234 249
rect 1268 215 1302 249
rect 1336 215 1393 249
rect 1082 205 1393 215
rect 775 177 805 197
rect 859 177 889 197
rect 963 177 993 205
rect 1082 177 1112 205
rect 1183 177 1213 205
rect 1270 177 1300 205
rect 1359 177 1389 205
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 487 21 517 47
rect 682 21 712 47
rect 775 21 805 47
rect 859 21 889 47
rect 963 21 993 47
rect 1082 21 1112 47
rect 1183 21 1213 47
rect 1270 21 1300 47
rect 1359 21 1389 47
<< polycont >>
rect 34 215 68 249
rect 245 215 279 249
rect 371 215 405 249
rect 514 215 548 249
rect 643 215 677 249
rect 794 215 828 249
rect 947 215 981 249
rect 1098 215 1132 249
rect 1166 215 1200 249
rect 1234 215 1268 249
rect 1302 215 1336 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 18 477 69 493
rect 18 443 35 477
rect 18 409 69 443
rect 103 485 169 527
rect 103 451 119 485
rect 153 451 169 485
rect 103 435 169 451
rect 203 477 246 493
rect 237 443 246 477
rect 18 375 35 409
rect 203 409 246 443
rect 280 489 325 527
rect 280 455 287 489
rect 321 455 325 489
rect 280 435 325 455
rect 359 477 405 493
rect 359 443 371 477
rect 69 375 203 401
rect 237 401 246 409
rect 359 401 405 443
rect 439 489 505 527
rect 439 455 455 489
rect 489 455 505 489
rect 439 435 505 455
rect 539 477 657 493
rect 573 443 607 477
rect 641 443 657 477
rect 539 409 657 443
rect 761 489 827 527
rect 761 455 777 489
rect 811 455 827 489
rect 761 436 827 455
rect 955 477 1013 493
rect 955 443 963 477
rect 997 443 1013 477
rect 539 401 607 409
rect 237 375 607 401
rect 641 401 657 409
rect 955 409 1013 443
rect 1049 485 1117 527
rect 1049 451 1067 485
rect 1101 451 1117 485
rect 1049 434 1117 451
rect 1151 477 1185 493
rect 955 401 963 409
rect 641 375 963 401
rect 997 400 1013 409
rect 1151 409 1185 443
rect 997 375 1110 400
rect 18 367 1110 375
rect 103 366 1110 367
rect 24 249 68 331
rect 24 215 34 249
rect 24 199 68 215
rect 103 169 172 366
rect 230 298 532 332
rect 230 249 279 298
rect 489 264 532 298
rect 661 298 965 332
rect 661 264 720 298
rect 931 264 965 298
rect 1076 264 1110 366
rect 1151 333 1185 375
rect 1219 485 1283 527
rect 1219 451 1235 485
rect 1269 451 1283 485
rect 1219 417 1283 451
rect 1219 383 1235 417
rect 1269 383 1283 417
rect 1219 367 1283 383
rect 1317 477 1355 493
rect 1317 443 1319 477
rect 1353 443 1355 477
rect 1317 409 1355 443
rect 1317 375 1319 409
rect 1353 375 1355 409
rect 1317 333 1355 375
rect 1389 485 1454 527
rect 1389 451 1403 485
rect 1437 451 1454 485
rect 1389 417 1454 451
rect 1389 383 1403 417
rect 1437 383 1454 417
rect 1389 367 1454 383
rect 1151 299 1455 333
rect 230 215 245 249
rect 355 249 443 264
rect 355 215 371 249
rect 405 215 443 249
rect 489 249 564 264
rect 629 249 720 264
rect 826 249 897 264
rect 489 216 514 249
rect 498 215 514 216
rect 548 215 564 249
rect 627 215 643 249
rect 677 215 720 249
rect 778 215 794 249
rect 828 215 897 249
rect 931 249 997 264
rect 931 215 947 249
rect 981 215 997 249
rect 1076 249 1352 264
rect 1076 215 1098 249
rect 1132 215 1166 249
rect 1200 215 1234 249
rect 1268 215 1302 249
rect 1336 215 1352 249
rect 230 199 279 215
rect 20 101 69 165
rect 103 135 119 169
rect 153 135 172 169
rect 103 131 172 135
rect 344 169 959 177
rect 1401 173 1455 299
rect 344 135 371 169
rect 405 135 731 169
rect 765 135 909 169
rect 943 135 959 169
rect 344 131 959 135
rect 20 67 35 101
rect 722 101 765 131
rect 69 93 588 97
rect 69 67 203 93
rect 20 59 203 67
rect 237 59 527 93
rect 561 59 588 93
rect 20 51 588 59
rect 622 93 688 97
rect 622 59 638 93
rect 672 59 688 93
rect 622 17 688 59
rect 722 67 731 101
rect 907 101 959 131
rect 1130 139 1455 173
rect 722 51 765 67
rect 799 93 873 97
rect 799 59 815 93
rect 849 59 873 93
rect 799 17 873 59
rect 907 67 909 101
rect 943 67 959 101
rect 907 51 959 67
rect 1007 93 1060 109
rect 1007 59 1013 93
rect 1047 59 1060 93
rect 1007 17 1060 59
rect 1130 101 1175 139
rect 1130 67 1139 101
rect 1173 67 1175 101
rect 1130 51 1175 67
rect 1215 89 1275 105
rect 1215 55 1225 89
rect 1259 55 1275 89
rect 1215 17 1275 55
rect 1309 101 1349 139
rect 1309 67 1311 101
rect 1345 67 1349 101
rect 1309 51 1349 67
rect 1383 93 1455 105
rect 1383 59 1399 93
rect 1433 59 1455 93
rect 1383 17 1455 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel locali s 1409 153 1443 187 0 FreeSans 400 0 0 0 X
port 10 nsew signal output
flabel locali s 1409 221 1443 255 0 FreeSans 400 0 0 0 X
port 10 nsew signal output
flabel locali s 1409 289 1443 323 0 FreeSans 400 0 0 0 X
port 10 nsew signal output
flabel locali s 857 221 891 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 D1
port 5 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 o2111a_4
rlabel metal1 s 0 -48 1472 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1472 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_END 945004
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 934078
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 7.360 0.000 
<< end >>
