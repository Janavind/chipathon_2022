magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect 95 503 1333 1103
<< pwell >>
rect 135 141 1293 333
<< mvnmos >>
rect 214 167 334 307
rect 390 167 510 307
rect 566 167 686 307
rect 742 167 862 307
rect 918 167 1038 307
rect 1094 167 1214 307
<< mvpmos >>
rect 214 837 334 1037
rect 390 837 510 1037
rect 566 837 686 1037
rect 742 837 862 1037
rect 918 837 1038 1037
rect 1094 837 1214 1037
rect 214 569 334 769
rect 390 569 510 769
rect 566 569 686 769
rect 742 569 862 769
rect 918 569 1038 769
rect 1094 569 1214 769
<< mvndiff >>
rect 161 281 214 307
rect 161 247 169 281
rect 203 247 214 281
rect 161 213 214 247
rect 161 179 169 213
rect 203 179 214 213
rect 161 167 214 179
rect 334 281 390 307
rect 334 247 345 281
rect 379 247 390 281
rect 334 213 390 247
rect 334 179 345 213
rect 379 179 390 213
rect 334 167 390 179
rect 510 281 566 307
rect 510 247 521 281
rect 555 247 566 281
rect 510 213 566 247
rect 510 179 521 213
rect 555 179 566 213
rect 510 167 566 179
rect 686 281 742 307
rect 686 247 697 281
rect 731 247 742 281
rect 686 213 742 247
rect 686 179 697 213
rect 731 179 742 213
rect 686 167 742 179
rect 862 281 918 307
rect 862 247 873 281
rect 907 247 918 281
rect 862 213 918 247
rect 862 179 873 213
rect 907 179 918 213
rect 862 167 918 179
rect 1038 281 1094 307
rect 1038 247 1049 281
rect 1083 247 1094 281
rect 1038 213 1094 247
rect 1038 179 1049 213
rect 1083 179 1094 213
rect 1038 167 1094 179
rect 1214 281 1267 307
rect 1214 247 1225 281
rect 1259 247 1267 281
rect 1214 213 1267 247
rect 1214 179 1225 213
rect 1259 179 1267 213
rect 1214 167 1267 179
<< mvpdiff >>
rect 161 1019 214 1037
rect 161 985 169 1019
rect 203 985 214 1019
rect 161 951 214 985
rect 161 917 169 951
rect 203 917 214 951
rect 161 883 214 917
rect 161 849 169 883
rect 203 849 214 883
rect 161 837 214 849
rect 334 1019 390 1037
rect 334 985 345 1019
rect 379 985 390 1019
rect 334 951 390 985
rect 334 917 345 951
rect 379 917 390 951
rect 334 883 390 917
rect 334 849 345 883
rect 379 849 390 883
rect 334 837 390 849
rect 510 1019 566 1037
rect 510 985 521 1019
rect 555 985 566 1019
rect 510 951 566 985
rect 510 917 521 951
rect 555 917 566 951
rect 510 883 566 917
rect 510 849 521 883
rect 555 849 566 883
rect 510 837 566 849
rect 686 1019 742 1037
rect 686 985 697 1019
rect 731 985 742 1019
rect 686 951 742 985
rect 686 917 697 951
rect 731 917 742 951
rect 686 883 742 917
rect 686 849 697 883
rect 731 849 742 883
rect 686 837 742 849
rect 862 1019 918 1037
rect 862 985 873 1019
rect 907 985 918 1019
rect 862 951 918 985
rect 862 917 873 951
rect 907 917 918 951
rect 862 883 918 917
rect 862 849 873 883
rect 907 849 918 883
rect 862 837 918 849
rect 1038 1019 1094 1037
rect 1038 985 1049 1019
rect 1083 985 1094 1019
rect 1038 951 1094 985
rect 1038 917 1049 951
rect 1083 917 1094 951
rect 1038 883 1094 917
rect 1038 849 1049 883
rect 1083 849 1094 883
rect 1038 837 1094 849
rect 1214 1019 1267 1037
rect 1214 985 1225 1019
rect 1259 985 1267 1019
rect 1214 951 1267 985
rect 1214 917 1225 951
rect 1259 917 1267 951
rect 1214 883 1267 917
rect 1214 849 1225 883
rect 1259 849 1267 883
rect 1214 837 1267 849
rect 161 751 214 769
rect 161 717 169 751
rect 203 717 214 751
rect 161 683 214 717
rect 161 649 169 683
rect 203 649 214 683
rect 161 615 214 649
rect 161 581 169 615
rect 203 581 214 615
rect 161 569 214 581
rect 334 751 390 769
rect 334 717 345 751
rect 379 717 390 751
rect 334 683 390 717
rect 334 649 345 683
rect 379 649 390 683
rect 334 615 390 649
rect 334 581 345 615
rect 379 581 390 615
rect 334 569 390 581
rect 510 751 566 769
rect 510 717 521 751
rect 555 717 566 751
rect 510 683 566 717
rect 510 649 521 683
rect 555 649 566 683
rect 510 615 566 649
rect 510 581 521 615
rect 555 581 566 615
rect 510 569 566 581
rect 686 751 742 769
rect 686 717 697 751
rect 731 717 742 751
rect 686 683 742 717
rect 686 649 697 683
rect 731 649 742 683
rect 686 615 742 649
rect 686 581 697 615
rect 731 581 742 615
rect 686 569 742 581
rect 862 751 918 769
rect 862 717 873 751
rect 907 717 918 751
rect 862 683 918 717
rect 862 649 873 683
rect 907 649 918 683
rect 862 615 918 649
rect 862 581 873 615
rect 907 581 918 615
rect 862 569 918 581
rect 1038 751 1094 769
rect 1038 717 1049 751
rect 1083 717 1094 751
rect 1038 683 1094 717
rect 1038 649 1049 683
rect 1083 649 1094 683
rect 1038 615 1094 649
rect 1038 581 1049 615
rect 1083 581 1094 615
rect 1038 569 1094 581
rect 1214 751 1267 769
rect 1214 717 1225 751
rect 1259 717 1267 751
rect 1214 683 1267 717
rect 1214 649 1225 683
rect 1259 649 1267 683
rect 1214 615 1267 649
rect 1214 581 1225 615
rect 1259 581 1267 615
rect 1214 569 1267 581
<< mvndiffc >>
rect 169 247 203 281
rect 169 179 203 213
rect 345 247 379 281
rect 345 179 379 213
rect 521 247 555 281
rect 521 179 555 213
rect 697 247 731 281
rect 697 179 731 213
rect 873 247 907 281
rect 873 179 907 213
rect 1049 247 1083 281
rect 1049 179 1083 213
rect 1225 247 1259 281
rect 1225 179 1259 213
<< mvpdiffc >>
rect 169 985 203 1019
rect 169 917 203 951
rect 169 849 203 883
rect 345 985 379 1019
rect 345 917 379 951
rect 345 849 379 883
rect 521 985 555 1019
rect 521 917 555 951
rect 521 849 555 883
rect 697 985 731 1019
rect 697 917 731 951
rect 697 849 731 883
rect 873 985 907 1019
rect 873 917 907 951
rect 873 849 907 883
rect 1049 985 1083 1019
rect 1049 917 1083 951
rect 1049 849 1083 883
rect 1225 985 1259 1019
rect 1225 917 1259 951
rect 1225 849 1259 883
rect 169 717 203 751
rect 169 649 203 683
rect 169 581 203 615
rect 345 717 379 751
rect 345 649 379 683
rect 345 581 379 615
rect 521 717 555 751
rect 521 649 555 683
rect 521 581 555 615
rect 697 717 731 751
rect 697 649 731 683
rect 697 581 731 615
rect 873 717 907 751
rect 873 649 907 683
rect 873 581 907 615
rect 1049 717 1083 751
rect 1049 649 1083 683
rect 1049 581 1083 615
rect 1225 717 1259 751
rect 1225 649 1259 683
rect 1225 581 1259 615
<< poly >>
rect 214 1119 510 1135
rect 214 1085 230 1119
rect 264 1085 307 1119
rect 341 1085 384 1119
rect 418 1085 460 1119
rect 494 1085 510 1119
rect 214 1069 510 1085
rect 734 1119 868 1135
rect 734 1085 750 1119
rect 784 1085 818 1119
rect 852 1085 868 1119
rect 734 1069 868 1085
rect 918 1119 1214 1135
rect 918 1085 934 1119
rect 968 1085 1011 1119
rect 1045 1085 1088 1119
rect 1122 1085 1164 1119
rect 1198 1085 1214 1119
rect 918 1069 1214 1085
rect 214 1037 334 1069
rect 390 1037 510 1069
rect 566 1037 686 1069
rect 742 1037 862 1069
rect 918 1037 1038 1069
rect 1094 1037 1214 1069
rect 214 769 334 837
rect 390 769 510 837
rect 566 769 686 837
rect 742 769 862 837
rect 918 769 1038 837
rect 1094 769 1214 837
rect 214 307 334 569
rect 390 307 510 569
rect 566 511 686 569
rect 566 477 608 511
rect 642 477 686 511
rect 566 443 686 477
rect 742 495 862 569
rect 918 537 1038 569
rect 742 456 1038 495
rect 566 409 608 443
rect 642 414 686 443
rect 642 409 862 414
rect 566 375 862 409
rect 566 307 686 333
rect 742 307 862 375
rect 918 307 1038 456
rect 1094 307 1214 569
rect 214 141 334 167
rect 390 141 510 167
rect 566 141 686 167
rect 742 141 862 167
rect 918 141 1038 167
rect 1094 141 1214 167
rect 214 125 510 141
rect 214 91 230 125
rect 264 91 307 125
rect 341 91 384 125
rect 418 91 460 125
rect 494 91 510 125
rect 214 75 510 91
rect 558 125 692 141
rect 558 91 574 125
rect 608 91 642 125
rect 676 91 692 125
rect 558 75 692 91
rect 1086 125 1220 141
rect 1086 91 1102 125
rect 1136 91 1170 125
rect 1204 91 1220 125
rect 1086 75 1220 91
<< polycont >>
rect 230 1085 264 1119
rect 307 1085 341 1119
rect 384 1085 418 1119
rect 460 1085 494 1119
rect 750 1085 784 1119
rect 818 1085 852 1119
rect 934 1085 968 1119
rect 1011 1085 1045 1119
rect 1088 1085 1122 1119
rect 1164 1085 1198 1119
rect 608 477 642 511
rect 608 409 642 443
rect 230 91 264 125
rect 307 91 341 125
rect 384 91 418 125
rect 460 91 494 125
rect 574 91 608 125
rect 642 91 676 125
rect 1102 91 1136 125
rect 1170 91 1204 125
<< locali >>
rect 214 1085 230 1119
rect 264 1085 307 1119
rect 341 1085 384 1119
rect 418 1085 460 1119
rect 494 1085 510 1119
rect 734 1085 750 1119
rect 784 1085 818 1119
rect 852 1085 868 1119
rect 918 1085 934 1119
rect 968 1085 1011 1119
rect 1045 1085 1088 1119
rect 1122 1085 1164 1119
rect 1198 1085 1214 1119
rect 169 1019 203 1035
rect 169 951 203 985
rect 169 883 203 917
rect 169 751 203 849
rect 169 683 203 717
rect 169 615 203 649
rect 169 518 203 581
rect 345 1025 379 1035
rect 345 953 379 985
rect 345 883 379 917
rect 345 751 379 849
rect 345 683 379 717
rect 345 615 379 649
rect 345 565 379 581
rect 203 484 241 518
rect 169 281 203 484
rect 169 213 203 247
rect 169 163 203 179
rect 345 293 379 297
rect 345 221 379 247
rect 345 163 379 179
rect 413 125 487 1085
rect 521 1019 555 1035
rect 521 951 555 985
rect 521 883 555 917
rect 521 751 555 849
rect 521 683 555 717
rect 521 615 555 649
rect 521 565 555 581
rect 697 1019 731 1035
rect 697 951 731 985
rect 697 883 731 917
rect 697 751 731 849
rect 697 683 731 717
rect 697 615 731 649
rect 608 511 642 527
rect 608 443 642 477
rect 591 409 608 441
rect 591 407 629 409
rect 608 393 642 407
rect 521 281 555 297
rect 521 213 555 247
rect 521 163 555 179
rect 697 281 731 581
rect 765 518 839 1085
rect 873 1019 907 1035
rect 873 951 907 985
rect 873 883 907 917
rect 873 751 907 849
rect 873 683 907 717
rect 873 615 907 649
rect 873 565 907 581
rect 799 484 837 518
rect 765 482 839 484
rect 697 213 731 247
rect 697 163 731 179
rect 873 281 907 297
rect 873 213 907 247
rect 873 163 907 179
rect 941 125 1015 1085
rect 1049 1025 1083 1035
rect 1049 953 1083 985
rect 1049 883 1083 917
rect 1049 751 1083 849
rect 1049 683 1083 717
rect 1049 615 1083 649
rect 1049 565 1083 581
rect 1225 1019 1259 1035
rect 1225 951 1259 985
rect 1225 883 1259 917
rect 1225 751 1259 849
rect 1225 683 1259 717
rect 1225 615 1259 649
rect 1225 441 1259 581
rect 1187 407 1225 441
rect 1049 293 1083 297
rect 1049 221 1083 247
rect 1049 163 1083 179
rect 1225 281 1259 407
rect 1225 213 1259 247
rect 1225 163 1259 179
rect 214 91 230 125
rect 264 91 307 125
rect 341 91 384 125
rect 418 91 460 125
rect 494 91 510 125
rect 558 91 574 125
rect 608 91 642 125
rect 676 91 1102 125
rect 1136 91 1170 125
rect 1204 91 1220 125
<< viali >>
rect 345 1019 379 1025
rect 345 991 379 1019
rect 345 951 379 953
rect 345 919 379 951
rect 169 484 203 518
rect 241 484 275 518
rect 345 281 379 293
rect 345 259 379 281
rect 345 213 379 221
rect 345 187 379 213
rect 557 407 591 441
rect 629 409 642 441
rect 642 409 663 441
rect 629 407 663 409
rect 765 484 799 518
rect 837 484 871 518
rect 1049 1019 1083 1025
rect 1049 991 1083 1019
rect 1049 951 1083 953
rect 1049 919 1083 951
rect 1153 407 1187 441
rect 1225 407 1259 441
rect 1049 281 1083 293
rect 1049 259 1083 281
rect 1049 213 1083 221
rect 1049 187 1083 213
<< metal1 >>
rect 339 1025 1089 1037
rect 339 991 345 1025
rect 379 991 1049 1025
rect 1083 991 1089 1025
rect 339 953 1089 991
rect 339 919 345 953
rect 379 919 1049 953
rect 1083 919 1089 953
rect 339 907 1089 919
rect 157 518 883 524
rect 157 484 169 518
rect 203 484 241 518
rect 275 484 765 518
rect 799 484 837 518
rect 871 484 883 518
rect 157 478 883 484
rect 545 441 1271 447
rect 545 407 557 441
rect 591 407 629 441
rect 663 407 1153 441
rect 1187 407 1225 441
rect 1259 407 1271 441
rect 545 401 1271 407
rect 339 293 1089 305
rect 339 259 345 293
rect 379 259 1049 293
rect 1083 259 1089 293
rect 339 221 1089 259
rect 339 187 345 221
rect 379 187 1049 221
rect 1083 187 1089 221
rect 339 175 1089 187
use sky130_fd_pr__nfet_01v8__example_55959141808417  sky130_fd_pr__nfet_01v8__example_55959141808417_0
timestamp 1666199351
transform -1 0 862 0 1 167
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808417  sky130_fd_pr__nfet_01v8__example_55959141808417_1
timestamp 1666199351
transform -1 0 1038 0 1 167
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808417  sky130_fd_pr__nfet_01v8__example_55959141808417_2
timestamp 1666199351
transform -1 0 334 0 1 167
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808417  sky130_fd_pr__nfet_01v8__example_55959141808417_3
timestamp 1666199351
transform 1 0 390 0 1 167
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808417  sky130_fd_pr__nfet_01v8__example_55959141808417_4
timestamp 1666199351
transform 1 0 1094 0 1 167
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808417  sky130_fd_pr__nfet_01v8__example_55959141808417_5
timestamp 1666199351
transform 1 0 566 0 1 167
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808416  sky130_fd_pr__pfet_01v8__example_55959141808416_0
timestamp 1666199351
transform -1 0 334 0 1 837
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808416  sky130_fd_pr__pfet_01v8__example_55959141808416_1
timestamp 1666199351
transform 1 0 566 0 1 837
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808416  sky130_fd_pr__pfet_01v8__example_55959141808416_2
timestamp 1666199351
transform -1 0 1038 0 1 837
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808416  sky130_fd_pr__pfet_01v8__example_55959141808416_3
timestamp 1666199351
transform 1 0 1094 0 1 569
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808416  sky130_fd_pr__pfet_01v8__example_55959141808416_4
timestamp 1666199351
transform -1 0 862 0 1 569
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808416  sky130_fd_pr__pfet_01v8__example_55959141808416_5
timestamp 1666199351
transform 1 0 390 0 1 569
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808416  sky130_fd_pr__pfet_01v8__example_55959141808416_6
timestamp 1666199351
transform -1 0 1038 0 1 569
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808416  sky130_fd_pr__pfet_01v8__example_55959141808416_7
timestamp 1666199351
transform -1 0 334 0 1 569
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808416  sky130_fd_pr__pfet_01v8__example_55959141808416_8
timestamp 1666199351
transform 1 0 566 0 1 569
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808416  sky130_fd_pr__pfet_01v8__example_55959141808416_9
timestamp 1666199351
transform 1 0 1094 0 1 837
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808416  sky130_fd_pr__pfet_01v8__example_55959141808416_10
timestamp 1666199351
transform -1 0 862 0 1 837
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808416  sky130_fd_pr__pfet_01v8__example_55959141808416_11
timestamp 1666199351
transform 1 0 390 0 1 837
box -1 0 121 1
<< labels >>
flabel metal1 s 570 951 802 1004 3 FreeSans 520 0 0 0 VPWR
port 1 nsew
flabel metal1 s 511 205 863 276 3 FreeSans 520 0 0 0 VGND
port 2 nsew
flabel locali s 294 92 346 125 3 FreeSans 520 0 0 0 IN0
port 3 nsew
flabel locali s 960 97 1012 149 3 FreeSans 520 0 0 0 IN1
port 4 nsew
flabel locali s 697 250 731 302 3 FreeSans 520 90 0 0 OUT
port 5 nsew
<< properties >>
string GDS_END 33676056
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 33667382
<< end >>
