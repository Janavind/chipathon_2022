magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 2890 582
<< pwell >>
rect 37 157 1011 203
rect 37 21 2834 157
rect 37 17 64 21
rect 30 -17 64 17
rect 1041 -17 1075 21
<< scnmos >>
rect 117 47 147 177
rect 311 47 341 177
rect 395 47 425 177
rect 479 47 509 177
rect 563 47 593 177
rect 647 47 677 177
rect 731 47 761 177
rect 815 47 845 177
rect 899 47 929 177
rect 1092 47 1122 131
rect 1178 47 1208 131
rect 1264 47 1294 131
rect 1350 47 1380 131
rect 1436 47 1466 131
rect 1522 47 1552 131
rect 1608 47 1638 131
rect 1694 47 1724 131
rect 1780 47 1810 131
rect 1866 47 1896 131
rect 1952 47 1982 131
rect 2038 47 2068 131
rect 2123 47 2153 131
rect 2209 47 2239 131
rect 2295 47 2325 131
rect 2381 47 2411 131
rect 2467 47 2497 131
rect 2553 47 2583 131
rect 2639 47 2669 131
rect 2725 47 2755 131
<< scpmoshvt >>
rect 117 297 147 497
rect 311 297 341 497
rect 395 297 425 497
rect 479 297 509 497
rect 563 297 593 497
rect 647 297 677 497
rect 731 297 761 497
rect 815 297 845 497
rect 899 297 929 497
rect 1092 297 1122 497
rect 1178 297 1208 497
rect 1264 297 1294 497
rect 1350 297 1380 497
rect 1436 297 1466 497
rect 1522 297 1552 497
rect 1608 297 1638 497
rect 1694 297 1724 497
rect 1780 297 1810 497
rect 1866 297 1896 497
rect 1952 297 1982 497
rect 2038 297 2068 497
rect 2123 297 2153 497
rect 2209 297 2239 497
rect 2295 297 2325 497
rect 2381 297 2411 497
rect 2467 297 2497 497
rect 2553 297 2583 497
rect 2639 297 2669 497
rect 2725 297 2755 497
<< ndiff >>
rect 63 163 117 177
rect 63 129 73 163
rect 107 129 117 163
rect 63 95 117 129
rect 63 61 73 95
rect 107 61 117 95
rect 63 47 117 61
rect 147 163 203 177
rect 147 129 157 163
rect 191 129 203 163
rect 147 95 203 129
rect 147 61 157 95
rect 191 61 203 95
rect 147 47 203 61
rect 259 163 311 177
rect 259 129 267 163
rect 301 129 311 163
rect 259 95 311 129
rect 259 61 267 95
rect 301 61 311 95
rect 259 47 311 61
rect 341 163 395 177
rect 341 129 351 163
rect 385 129 395 163
rect 341 95 395 129
rect 341 61 351 95
rect 385 61 395 95
rect 341 47 395 61
rect 425 95 479 177
rect 425 61 435 95
rect 469 61 479 95
rect 425 47 479 61
rect 509 163 563 177
rect 509 129 519 163
rect 553 129 563 163
rect 509 95 563 129
rect 509 61 519 95
rect 553 61 563 95
rect 509 47 563 61
rect 593 95 647 177
rect 593 61 603 95
rect 637 61 647 95
rect 593 47 647 61
rect 677 163 731 177
rect 677 129 687 163
rect 721 129 731 163
rect 677 95 731 129
rect 677 61 687 95
rect 721 61 731 95
rect 677 47 731 61
rect 761 95 815 177
rect 761 61 771 95
rect 805 61 815 95
rect 761 47 815 61
rect 845 163 899 177
rect 845 129 855 163
rect 889 129 899 163
rect 845 95 899 129
rect 845 61 855 95
rect 889 61 899 95
rect 845 47 899 61
rect 929 163 985 177
rect 929 129 939 163
rect 973 129 985 163
rect 929 95 985 129
rect 929 61 939 95
rect 973 61 985 95
rect 929 47 985 61
rect 1039 93 1092 131
rect 1039 59 1047 93
rect 1081 59 1092 93
rect 1039 47 1092 59
rect 1122 106 1178 131
rect 1122 72 1133 106
rect 1167 72 1178 106
rect 1122 47 1178 72
rect 1208 106 1264 131
rect 1208 72 1219 106
rect 1253 72 1264 106
rect 1208 47 1264 72
rect 1294 106 1350 131
rect 1294 72 1305 106
rect 1339 72 1350 106
rect 1294 47 1350 72
rect 1380 106 1436 131
rect 1380 72 1391 106
rect 1425 72 1436 106
rect 1380 47 1436 72
rect 1466 106 1522 131
rect 1466 72 1477 106
rect 1511 72 1522 106
rect 1466 47 1522 72
rect 1552 97 1608 131
rect 1552 63 1563 97
rect 1597 63 1608 97
rect 1552 47 1608 63
rect 1638 106 1694 131
rect 1638 72 1649 106
rect 1683 72 1694 106
rect 1638 47 1694 72
rect 1724 97 1780 131
rect 1724 63 1735 97
rect 1769 63 1780 97
rect 1724 47 1780 63
rect 1810 106 1866 131
rect 1810 72 1821 106
rect 1855 72 1866 106
rect 1810 47 1866 72
rect 1896 97 1952 131
rect 1896 63 1907 97
rect 1941 63 1952 97
rect 1896 47 1952 63
rect 1982 106 2038 131
rect 1982 72 1993 106
rect 2027 72 2038 106
rect 1982 47 2038 72
rect 2068 97 2123 131
rect 2068 63 2079 97
rect 2113 63 2123 97
rect 2068 47 2123 63
rect 2153 106 2209 131
rect 2153 72 2164 106
rect 2198 72 2209 106
rect 2153 47 2209 72
rect 2239 97 2295 131
rect 2239 63 2250 97
rect 2284 63 2295 97
rect 2239 47 2295 63
rect 2325 106 2381 131
rect 2325 72 2336 106
rect 2370 72 2381 106
rect 2325 47 2381 72
rect 2411 97 2467 131
rect 2411 63 2422 97
rect 2456 63 2467 97
rect 2411 47 2467 63
rect 2497 106 2553 131
rect 2497 72 2508 106
rect 2542 72 2553 106
rect 2497 47 2553 72
rect 2583 97 2639 131
rect 2583 63 2594 97
rect 2628 63 2639 97
rect 2583 47 2639 63
rect 2669 106 2725 131
rect 2669 72 2680 106
rect 2714 72 2725 106
rect 2669 47 2725 72
rect 2755 97 2808 131
rect 2755 63 2766 97
rect 2800 63 2808 97
rect 2755 47 2808 63
<< pdiff >>
rect 61 485 117 497
rect 61 451 73 485
rect 107 451 117 485
rect 61 417 117 451
rect 61 383 73 417
rect 107 383 117 417
rect 61 349 117 383
rect 61 315 73 349
rect 107 315 117 349
rect 61 297 117 315
rect 147 485 201 497
rect 147 451 157 485
rect 191 451 201 485
rect 147 417 201 451
rect 147 383 157 417
rect 191 383 201 417
rect 147 349 201 383
rect 147 315 157 349
rect 191 315 201 349
rect 147 297 201 315
rect 255 485 311 497
rect 255 451 267 485
rect 301 451 311 485
rect 255 417 311 451
rect 255 383 267 417
rect 301 383 311 417
rect 255 349 311 383
rect 255 315 267 349
rect 301 315 311 349
rect 255 297 311 315
rect 341 409 395 497
rect 341 375 351 409
rect 385 375 395 409
rect 341 341 395 375
rect 341 307 351 341
rect 385 307 395 341
rect 341 297 395 307
rect 425 489 479 497
rect 425 455 435 489
rect 469 455 479 489
rect 425 421 479 455
rect 425 387 435 421
rect 469 387 479 421
rect 425 297 479 387
rect 509 409 563 497
rect 509 375 519 409
rect 553 375 563 409
rect 509 341 563 375
rect 509 307 519 341
rect 553 307 563 341
rect 509 297 563 307
rect 593 485 647 497
rect 593 451 603 485
rect 637 451 647 485
rect 593 417 647 451
rect 593 383 603 417
rect 637 383 647 417
rect 593 341 647 383
rect 593 307 603 341
rect 637 307 647 341
rect 593 297 647 307
rect 677 485 731 497
rect 677 451 687 485
rect 721 451 731 485
rect 677 417 731 451
rect 677 383 687 417
rect 721 383 731 417
rect 677 297 731 383
rect 761 477 815 497
rect 761 443 771 477
rect 805 443 815 477
rect 761 409 815 443
rect 761 375 771 409
rect 805 375 815 409
rect 761 341 815 375
rect 761 307 771 341
rect 805 307 815 341
rect 761 297 815 307
rect 845 485 899 497
rect 845 451 855 485
rect 889 451 899 485
rect 845 417 899 451
rect 845 383 855 417
rect 889 383 899 417
rect 845 297 899 383
rect 929 477 985 497
rect 929 443 939 477
rect 973 443 985 477
rect 929 409 985 443
rect 929 375 939 409
rect 973 375 985 409
rect 929 341 985 375
rect 929 307 939 341
rect 973 307 985 341
rect 929 297 985 307
rect 1039 485 1092 497
rect 1039 451 1047 485
rect 1081 451 1092 485
rect 1039 417 1092 451
rect 1039 383 1047 417
rect 1081 383 1092 417
rect 1039 349 1092 383
rect 1039 315 1047 349
rect 1081 315 1092 349
rect 1039 297 1092 315
rect 1122 477 1178 497
rect 1122 443 1133 477
rect 1167 443 1178 477
rect 1122 409 1178 443
rect 1122 375 1133 409
rect 1167 375 1178 409
rect 1122 341 1178 375
rect 1122 307 1133 341
rect 1167 307 1178 341
rect 1122 297 1178 307
rect 1208 485 1264 497
rect 1208 451 1219 485
rect 1253 451 1264 485
rect 1208 417 1264 451
rect 1208 383 1219 417
rect 1253 383 1264 417
rect 1208 349 1264 383
rect 1208 315 1219 349
rect 1253 315 1264 349
rect 1208 297 1264 315
rect 1294 476 1350 497
rect 1294 442 1305 476
rect 1339 442 1350 476
rect 1294 408 1350 442
rect 1294 374 1305 408
rect 1339 374 1350 408
rect 1294 340 1350 374
rect 1294 306 1305 340
rect 1339 306 1350 340
rect 1294 297 1350 306
rect 1380 485 1436 497
rect 1380 451 1391 485
rect 1425 451 1436 485
rect 1380 417 1436 451
rect 1380 383 1391 417
rect 1425 383 1436 417
rect 1380 349 1436 383
rect 1380 315 1391 349
rect 1425 315 1436 349
rect 1380 297 1436 315
rect 1466 476 1522 497
rect 1466 442 1477 476
rect 1511 442 1522 476
rect 1466 355 1522 442
rect 1466 321 1477 355
rect 1511 321 1522 355
rect 1466 297 1522 321
rect 1552 461 1608 497
rect 1552 427 1563 461
rect 1597 427 1608 461
rect 1552 297 1608 427
rect 1638 476 1694 497
rect 1638 442 1649 476
rect 1683 442 1694 476
rect 1638 355 1694 442
rect 1638 321 1649 355
rect 1683 321 1694 355
rect 1638 297 1694 321
rect 1724 461 1780 497
rect 1724 427 1735 461
rect 1769 427 1780 461
rect 1724 297 1780 427
rect 1810 476 1866 497
rect 1810 442 1821 476
rect 1855 442 1866 476
rect 1810 355 1866 442
rect 1810 321 1821 355
rect 1855 321 1866 355
rect 1810 297 1866 321
rect 1896 461 1952 497
rect 1896 427 1907 461
rect 1941 427 1952 461
rect 1896 297 1952 427
rect 1982 476 2038 497
rect 1982 442 1993 476
rect 2027 442 2038 476
rect 1982 355 2038 442
rect 1982 321 1993 355
rect 2027 321 2038 355
rect 1982 297 2038 321
rect 2068 461 2123 497
rect 2068 427 2079 461
rect 2113 427 2123 461
rect 2068 297 2123 427
rect 2153 476 2209 497
rect 2153 442 2164 476
rect 2198 442 2209 476
rect 2153 355 2209 442
rect 2153 321 2164 355
rect 2198 321 2209 355
rect 2153 297 2209 321
rect 2239 461 2295 497
rect 2239 427 2250 461
rect 2284 427 2295 461
rect 2239 297 2295 427
rect 2325 476 2381 497
rect 2325 442 2336 476
rect 2370 442 2381 476
rect 2325 355 2381 442
rect 2325 321 2336 355
rect 2370 321 2381 355
rect 2325 297 2381 321
rect 2411 461 2467 497
rect 2411 427 2422 461
rect 2456 427 2467 461
rect 2411 297 2467 427
rect 2497 476 2553 497
rect 2497 442 2508 476
rect 2542 442 2553 476
rect 2497 355 2553 442
rect 2497 321 2508 355
rect 2542 321 2553 355
rect 2497 297 2553 321
rect 2583 461 2639 497
rect 2583 427 2594 461
rect 2628 427 2639 461
rect 2583 297 2639 427
rect 2669 476 2725 497
rect 2669 442 2680 476
rect 2714 442 2725 476
rect 2669 355 2725 442
rect 2669 321 2680 355
rect 2714 321 2725 355
rect 2669 297 2725 321
rect 2755 461 2808 497
rect 2755 427 2766 461
rect 2800 427 2808 461
rect 2755 297 2808 427
<< ndiffc >>
rect 73 129 107 163
rect 73 61 107 95
rect 157 129 191 163
rect 157 61 191 95
rect 267 129 301 163
rect 267 61 301 95
rect 351 129 385 163
rect 351 61 385 95
rect 435 61 469 95
rect 519 129 553 163
rect 519 61 553 95
rect 603 61 637 95
rect 687 129 721 163
rect 687 61 721 95
rect 771 61 805 95
rect 855 129 889 163
rect 855 61 889 95
rect 939 129 973 163
rect 939 61 973 95
rect 1047 59 1081 93
rect 1133 72 1167 106
rect 1219 72 1253 106
rect 1305 72 1339 106
rect 1391 72 1425 106
rect 1477 72 1511 106
rect 1563 63 1597 97
rect 1649 72 1683 106
rect 1735 63 1769 97
rect 1821 72 1855 106
rect 1907 63 1941 97
rect 1993 72 2027 106
rect 2079 63 2113 97
rect 2164 72 2198 106
rect 2250 63 2284 97
rect 2336 72 2370 106
rect 2422 63 2456 97
rect 2508 72 2542 106
rect 2594 63 2628 97
rect 2680 72 2714 106
rect 2766 63 2800 97
<< pdiffc >>
rect 73 451 107 485
rect 73 383 107 417
rect 73 315 107 349
rect 157 451 191 485
rect 157 383 191 417
rect 157 315 191 349
rect 267 451 301 485
rect 267 383 301 417
rect 267 315 301 349
rect 351 375 385 409
rect 351 307 385 341
rect 435 455 469 489
rect 435 387 469 421
rect 519 375 553 409
rect 519 307 553 341
rect 603 451 637 485
rect 603 383 637 417
rect 603 307 637 341
rect 687 451 721 485
rect 687 383 721 417
rect 771 443 805 477
rect 771 375 805 409
rect 771 307 805 341
rect 855 451 889 485
rect 855 383 889 417
rect 939 443 973 477
rect 939 375 973 409
rect 939 307 973 341
rect 1047 451 1081 485
rect 1047 383 1081 417
rect 1047 315 1081 349
rect 1133 443 1167 477
rect 1133 375 1167 409
rect 1133 307 1167 341
rect 1219 451 1253 485
rect 1219 383 1253 417
rect 1219 315 1253 349
rect 1305 442 1339 476
rect 1305 374 1339 408
rect 1305 306 1339 340
rect 1391 451 1425 485
rect 1391 383 1425 417
rect 1391 315 1425 349
rect 1477 442 1511 476
rect 1477 321 1511 355
rect 1563 427 1597 461
rect 1649 442 1683 476
rect 1649 321 1683 355
rect 1735 427 1769 461
rect 1821 442 1855 476
rect 1821 321 1855 355
rect 1907 427 1941 461
rect 1993 442 2027 476
rect 1993 321 2027 355
rect 2079 427 2113 461
rect 2164 442 2198 476
rect 2164 321 2198 355
rect 2250 427 2284 461
rect 2336 442 2370 476
rect 2336 321 2370 355
rect 2422 427 2456 461
rect 2508 442 2542 476
rect 2508 321 2542 355
rect 2594 427 2628 461
rect 2680 442 2714 476
rect 2680 321 2714 355
rect 2766 427 2800 461
<< poly >>
rect 117 497 147 523
rect 311 497 341 523
rect 395 497 425 523
rect 479 497 509 523
rect 563 497 593 523
rect 647 497 677 523
rect 731 497 761 523
rect 815 497 845 523
rect 899 497 929 523
rect 1092 497 1122 523
rect 1178 497 1208 523
rect 1264 497 1294 523
rect 1350 497 1380 523
rect 1436 497 1466 523
rect 1522 497 1552 523
rect 1608 497 1638 523
rect 1694 497 1724 523
rect 1780 497 1810 523
rect 1866 497 1896 523
rect 1952 497 1982 523
rect 2038 497 2068 523
rect 2123 497 2153 523
rect 2209 497 2239 523
rect 2295 497 2325 523
rect 2381 497 2411 523
rect 2467 497 2497 523
rect 2553 497 2583 523
rect 2639 497 2669 523
rect 2725 497 2755 523
rect 117 265 147 297
rect 311 265 341 297
rect 395 265 425 297
rect 479 265 509 297
rect 563 265 593 297
rect 57 249 147 265
rect 57 215 73 249
rect 107 215 147 249
rect 57 199 147 215
rect 189 249 593 265
rect 189 215 199 249
rect 233 215 267 249
rect 301 215 335 249
rect 369 215 403 249
rect 437 215 593 249
rect 189 199 593 215
rect 117 177 147 199
rect 311 177 341 199
rect 395 177 425 199
rect 479 177 509 199
rect 563 177 593 199
rect 647 265 677 297
rect 731 265 761 297
rect 815 265 845 297
rect 899 265 929 297
rect 1092 282 1122 297
rect 1178 282 1208 297
rect 1264 282 1294 297
rect 1350 282 1380 297
rect 647 249 929 265
rect 647 215 671 249
rect 705 215 739 249
rect 773 215 807 249
rect 841 215 875 249
rect 909 215 929 249
rect 647 199 929 215
rect 647 177 677 199
rect 731 177 761 199
rect 815 177 845 199
rect 899 177 929 199
rect 1033 249 1380 282
rect 1033 215 1049 249
rect 1083 215 1380 249
rect 1033 180 1380 215
rect 1092 131 1122 180
rect 1178 131 1208 180
rect 1264 131 1294 180
rect 1350 131 1380 180
rect 1436 265 1466 297
rect 1522 265 1552 297
rect 1608 265 1638 297
rect 1694 265 1724 297
rect 1780 265 1810 297
rect 1866 265 1896 297
rect 1952 265 1982 297
rect 2038 265 2068 297
rect 2123 265 2153 297
rect 2209 265 2239 297
rect 2295 265 2325 297
rect 2381 265 2411 297
rect 2467 265 2497 297
rect 2553 265 2583 297
rect 2639 265 2669 297
rect 2725 265 2755 297
rect 1436 249 2755 265
rect 1436 215 1476 249
rect 1510 215 1544 249
rect 1578 215 1612 249
rect 1646 215 1680 249
rect 1714 215 1748 249
rect 1782 215 1816 249
rect 1850 215 1884 249
rect 1918 215 1952 249
rect 1986 215 2020 249
rect 2054 215 2088 249
rect 2122 215 2156 249
rect 2190 215 2224 249
rect 2258 215 2292 249
rect 2326 215 2360 249
rect 2394 215 2428 249
rect 2462 215 2496 249
rect 2530 215 2755 249
rect 1436 190 2755 215
rect 1436 131 1466 190
rect 1522 131 1552 190
rect 1608 131 1638 190
rect 1694 131 1724 190
rect 1780 131 1810 190
rect 1866 131 1896 190
rect 1952 131 1982 190
rect 2038 131 2068 190
rect 2123 131 2153 190
rect 2209 131 2239 190
rect 2295 131 2325 190
rect 2381 131 2411 190
rect 2467 131 2497 190
rect 2553 131 2583 190
rect 2639 131 2669 190
rect 2725 131 2755 190
rect 117 21 147 47
rect 311 21 341 47
rect 395 21 425 47
rect 479 21 509 47
rect 563 21 593 47
rect 647 21 677 47
rect 731 21 761 47
rect 815 21 845 47
rect 899 21 929 47
rect 1092 21 1122 47
rect 1178 21 1208 47
rect 1264 21 1294 47
rect 1350 21 1380 47
rect 1436 21 1466 47
rect 1522 21 1552 47
rect 1608 21 1638 47
rect 1694 21 1724 47
rect 1780 21 1810 47
rect 1866 21 1896 47
rect 1952 21 1982 47
rect 2038 21 2068 47
rect 2123 21 2153 47
rect 2209 21 2239 47
rect 2295 21 2325 47
rect 2381 21 2411 47
rect 2467 21 2497 47
rect 2553 21 2583 47
rect 2639 21 2669 47
rect 2725 21 2755 47
<< polycont >>
rect 73 215 107 249
rect 199 215 233 249
rect 267 215 301 249
rect 335 215 369 249
rect 403 215 437 249
rect 671 215 705 249
rect 739 215 773 249
rect 807 215 841 249
rect 875 215 909 249
rect 1049 215 1083 249
rect 1476 215 1510 249
rect 1544 215 1578 249
rect 1612 215 1646 249
rect 1680 215 1714 249
rect 1748 215 1782 249
rect 1816 215 1850 249
rect 1884 215 1918 249
rect 1952 215 1986 249
rect 2020 215 2054 249
rect 2088 215 2122 249
rect 2156 215 2190 249
rect 2224 215 2258 249
rect 2292 215 2326 249
rect 2360 215 2394 249
rect 2428 215 2462 249
rect 2496 215 2530 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 26 485 107 527
rect 26 451 73 485
rect 26 417 107 451
rect 26 383 73 417
rect 26 349 107 383
rect 26 315 73 349
rect 141 485 207 493
rect 141 451 157 485
rect 191 451 207 485
rect 141 417 207 451
rect 141 383 157 417
rect 191 383 207 417
rect 141 349 207 383
rect 141 315 157 349
rect 191 315 207 349
rect 241 489 653 493
rect 241 485 435 489
rect 241 451 267 485
rect 301 459 435 485
rect 301 451 317 459
rect 241 417 317 451
rect 419 455 435 459
rect 469 485 653 489
rect 469 459 603 485
rect 469 455 485 459
rect 241 383 267 417
rect 301 383 317 417
rect 241 349 317 383
rect 241 315 267 349
rect 301 315 317 349
rect 351 409 385 425
rect 419 421 485 455
rect 587 451 603 459
rect 637 451 653 485
rect 419 387 435 421
rect 469 387 485 421
rect 519 409 553 425
rect 351 349 385 375
rect 519 349 553 375
rect 351 341 553 349
rect 26 299 107 315
rect 17 249 123 264
rect 17 215 73 249
rect 107 215 123 249
rect 157 255 207 315
rect 385 307 519 341
rect 351 289 553 307
rect 587 417 653 451
rect 587 383 603 417
rect 637 383 653 417
rect 587 341 653 383
rect 687 485 737 527
rect 721 451 737 485
rect 687 417 737 451
rect 721 383 737 417
rect 687 367 737 383
rect 771 477 805 493
rect 771 409 805 443
rect 587 307 603 341
rect 637 333 653 341
rect 771 341 805 375
rect 839 485 905 527
rect 839 451 855 485
rect 889 451 905 485
rect 839 417 905 451
rect 839 383 855 417
rect 889 383 905 417
rect 839 367 905 383
rect 939 477 995 493
rect 973 443 995 477
rect 939 409 995 443
rect 973 375 995 409
rect 637 307 771 333
rect 939 341 995 375
rect 805 307 939 333
rect 973 307 995 341
rect 587 291 995 307
rect 1031 485 1097 493
rect 1031 425 1047 485
rect 1081 425 1097 485
rect 1031 417 1097 425
rect 1031 383 1047 417
rect 1081 383 1097 417
rect 1031 349 1097 383
rect 1031 315 1047 349
rect 1081 315 1097 349
rect 1031 299 1097 315
rect 1131 477 1169 493
rect 1131 443 1133 477
rect 1167 443 1169 477
rect 1131 409 1169 443
rect 1131 375 1133 409
rect 1167 375 1169 409
rect 1131 341 1169 375
rect 1131 307 1133 341
rect 1167 307 1169 341
rect 157 249 453 255
rect 157 215 199 249
rect 233 215 267 249
rect 301 215 335 249
rect 369 215 403 249
rect 437 215 453 249
rect 49 163 107 181
rect 157 163 207 215
rect 487 193 553 289
rect 1131 265 1169 307
rect 1203 485 1269 493
rect 1203 425 1219 485
rect 1253 425 1269 485
rect 1203 417 1269 425
rect 1203 383 1219 417
rect 1253 383 1269 417
rect 1203 349 1269 383
rect 1203 315 1219 349
rect 1253 315 1269 349
rect 1203 299 1269 315
rect 1303 476 1341 492
rect 1303 442 1305 476
rect 1339 442 1341 476
rect 1303 408 1341 442
rect 1303 374 1305 408
rect 1339 374 1341 408
rect 1303 340 1341 374
rect 1303 306 1305 340
rect 1339 306 1341 340
rect 1303 265 1341 306
rect 1375 485 1441 493
rect 1375 459 1391 485
rect 1375 425 1390 459
rect 1425 451 1441 485
rect 1424 425 1441 451
rect 1375 417 1441 425
rect 1375 383 1391 417
rect 1425 383 1441 417
rect 1375 349 1441 383
rect 1375 315 1391 349
rect 1425 315 1441 349
rect 1375 299 1441 315
rect 1475 476 1520 492
rect 1475 442 1477 476
rect 1511 442 1520 476
rect 1475 355 1520 442
rect 1554 461 1606 493
rect 1554 459 1563 461
rect 1554 425 1560 459
rect 1597 427 1606 461
rect 1594 425 1606 427
rect 1554 381 1606 425
rect 1640 476 1692 492
rect 1640 442 1649 476
rect 1683 442 1692 476
rect 1475 321 1477 355
rect 1511 347 1520 355
rect 1640 355 1692 442
rect 1726 461 1778 493
rect 1726 427 1735 461
rect 1769 459 1778 461
rect 1726 425 1736 427
rect 1770 425 1778 459
rect 1726 381 1778 425
rect 1812 476 1864 492
rect 1812 442 1821 476
rect 1855 442 1864 476
rect 1640 347 1649 355
rect 1511 321 1649 347
rect 1683 347 1692 355
rect 1812 355 1864 442
rect 1898 461 1950 493
rect 1898 427 1907 461
rect 1941 459 1950 461
rect 1898 425 1908 427
rect 1942 425 1950 459
rect 1898 381 1950 425
rect 1984 476 2036 492
rect 1984 442 1993 476
rect 2027 442 2036 476
rect 1812 347 1821 355
rect 1683 321 1821 347
rect 1855 347 1864 355
rect 1984 355 2036 442
rect 2070 461 2119 493
rect 2070 425 2079 461
rect 2113 425 2119 461
rect 2070 381 2119 425
rect 2153 476 2205 492
rect 2153 442 2164 476
rect 2198 442 2205 476
rect 1984 347 1993 355
rect 1855 321 1993 347
rect 2027 347 2036 355
rect 2153 355 2205 442
rect 2242 461 2291 493
rect 2242 427 2250 461
rect 2284 459 2291 461
rect 2242 425 2251 427
rect 2285 425 2291 459
rect 2242 381 2291 425
rect 2325 476 2377 492
rect 2325 442 2336 476
rect 2370 442 2377 476
rect 2153 347 2164 355
rect 2027 321 2164 347
rect 2198 347 2205 355
rect 2325 355 2377 442
rect 2414 461 2463 493
rect 2414 425 2422 461
rect 2456 425 2463 461
rect 2414 381 2463 425
rect 2497 476 2549 492
rect 2497 442 2508 476
rect 2542 442 2549 476
rect 2325 347 2336 355
rect 2198 321 2336 347
rect 2370 347 2377 355
rect 2497 355 2549 442
rect 2586 461 2637 493
rect 2586 459 2594 461
rect 2586 425 2592 459
rect 2628 427 2637 461
rect 2626 425 2637 427
rect 2586 381 2637 425
rect 2671 476 2729 492
rect 2671 442 2680 476
rect 2714 442 2729 476
rect 2497 347 2508 355
rect 2370 321 2508 347
rect 2542 344 2549 355
rect 2671 355 2729 442
rect 2763 461 2817 493
rect 2763 427 2766 461
rect 2800 459 2817 461
rect 2763 425 2768 427
rect 2802 425 2817 459
rect 2763 378 2817 425
rect 2671 344 2680 355
rect 2542 321 2680 344
rect 2714 344 2729 355
rect 2714 321 2817 344
rect 1475 299 2817 321
rect 652 249 940 255
rect 652 215 671 249
rect 705 215 739 249
rect 773 215 807 249
rect 841 215 875 249
rect 909 215 940 249
rect 1029 249 1092 265
rect 1029 215 1049 249
rect 1083 215 1092 249
rect 487 187 619 193
rect 487 181 505 187
rect 49 129 73 163
rect 49 95 107 129
rect 49 61 73 95
rect 49 17 107 61
rect 141 129 157 163
rect 191 129 207 163
rect 141 95 207 129
rect 141 61 157 95
rect 191 61 207 95
rect 141 51 207 61
rect 243 163 301 181
rect 243 129 267 163
rect 243 95 301 129
rect 243 61 267 95
rect 243 17 301 61
rect 335 163 505 181
rect 539 163 577 187
rect 335 129 351 163
rect 385 153 505 163
rect 553 153 577 163
rect 611 181 619 187
rect 1029 187 1092 215
rect 611 163 905 181
rect 611 153 687 163
rect 385 145 519 153
rect 385 129 401 145
rect 335 95 401 129
rect 503 129 519 145
rect 553 145 687 153
rect 553 129 569 145
rect 335 61 351 95
rect 385 61 401 95
rect 335 51 401 61
rect 435 95 469 111
rect 435 17 469 61
rect 503 95 569 129
rect 671 129 687 145
rect 721 145 855 163
rect 721 129 737 145
rect 503 61 519 95
rect 553 61 569 95
rect 503 51 569 61
rect 603 95 637 111
rect 603 17 637 61
rect 671 95 737 129
rect 839 129 855 145
rect 889 129 905 163
rect 671 61 687 95
rect 721 61 737 95
rect 671 51 737 61
rect 771 95 805 111
rect 771 17 805 61
rect 839 95 905 129
rect 839 61 855 95
rect 889 61 905 95
rect 839 51 905 61
rect 939 163 995 181
rect 973 129 995 163
rect 1029 153 1042 187
rect 1076 153 1092 187
rect 1029 147 1092 153
rect 1131 249 2550 265
rect 1131 215 1476 249
rect 1510 215 1544 249
rect 1578 215 1612 249
rect 1646 215 1680 249
rect 1714 215 1748 249
rect 1782 215 1816 249
rect 1850 215 1884 249
rect 1918 215 1952 249
rect 1986 215 2020 249
rect 2054 215 2088 249
rect 2122 215 2156 249
rect 2190 215 2224 249
rect 2258 215 2292 249
rect 2326 215 2360 249
rect 2394 215 2428 249
rect 2462 215 2496 249
rect 2530 215 2550 249
rect 939 113 995 129
rect 939 95 1090 113
rect 973 93 1090 95
rect 973 61 1047 93
rect 939 59 1047 61
rect 1081 59 1090 93
rect 939 17 1090 59
rect 1131 106 1176 215
rect 1131 72 1133 106
rect 1167 72 1176 106
rect 1131 53 1176 72
rect 1210 106 1262 122
rect 1210 72 1219 106
rect 1253 72 1262 106
rect 1210 17 1262 72
rect 1298 106 1348 215
rect 2584 181 2817 299
rect 1468 147 2817 181
rect 1298 72 1305 106
rect 1339 72 1348 106
rect 1298 53 1348 72
rect 1382 106 1434 129
rect 1382 72 1391 106
rect 1425 72 1434 106
rect 1382 17 1434 72
rect 1468 106 1520 147
rect 1468 72 1477 106
rect 1511 72 1520 106
rect 1468 56 1520 72
rect 1554 97 1606 113
rect 1554 63 1563 97
rect 1597 63 1606 97
rect 1554 17 1606 63
rect 1640 106 1692 147
rect 1640 72 1649 106
rect 1683 72 1692 106
rect 1640 56 1692 72
rect 1726 97 1778 113
rect 1726 63 1735 97
rect 1769 63 1778 97
rect 1726 17 1778 63
rect 1812 106 1864 147
rect 1812 72 1821 106
rect 1855 72 1864 106
rect 1812 56 1864 72
rect 1898 97 1947 113
rect 1898 63 1907 97
rect 1941 63 1947 97
rect 1898 17 1947 63
rect 1981 106 2036 147
rect 1981 72 1993 106
rect 2027 72 2036 106
rect 1981 56 2036 72
rect 2070 97 2119 113
rect 2070 63 2079 97
rect 2113 63 2119 97
rect 2070 17 2119 63
rect 2153 106 2205 147
rect 2153 72 2164 106
rect 2198 72 2205 106
rect 2153 56 2205 72
rect 2241 97 2291 113
rect 2241 63 2250 97
rect 2284 63 2291 97
rect 2241 17 2291 63
rect 2325 106 2377 147
rect 2325 72 2336 106
rect 2370 72 2377 106
rect 2325 56 2377 72
rect 2413 97 2463 113
rect 2413 63 2422 97
rect 2456 63 2463 97
rect 2413 17 2463 63
rect 2497 106 2549 147
rect 2497 72 2508 106
rect 2542 72 2549 106
rect 2497 56 2549 72
rect 2585 97 2637 113
rect 2585 63 2594 97
rect 2628 63 2637 97
rect 2585 17 2637 63
rect 2671 106 2723 147
rect 2671 72 2680 106
rect 2714 72 2723 106
rect 2671 56 2723 72
rect 2757 97 2817 113
rect 2757 63 2766 97
rect 2800 63 2817 97
rect 2757 17 2817 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 1047 451 1081 459
rect 1047 425 1081 451
rect 1219 451 1253 459
rect 1219 425 1253 451
rect 1390 451 1391 459
rect 1391 451 1424 459
rect 1390 425 1424 451
rect 1560 427 1563 459
rect 1563 427 1594 459
rect 1560 425 1594 427
rect 1736 427 1769 459
rect 1769 427 1770 459
rect 1736 425 1770 427
rect 1908 427 1941 459
rect 1941 427 1942 459
rect 1908 425 1942 427
rect 2079 427 2113 459
rect 2079 425 2113 427
rect 2251 427 2284 459
rect 2284 427 2285 459
rect 2251 425 2285 427
rect 2422 427 2456 459
rect 2422 425 2456 427
rect 2592 427 2594 459
rect 2594 427 2626 459
rect 2592 425 2626 427
rect 2768 427 2800 459
rect 2800 427 2802 459
rect 2768 425 2802 427
rect 505 163 539 187
rect 505 153 519 163
rect 519 153 539 163
rect 577 153 611 187
rect 1042 153 1076 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
<< metal1 >>
rect 0 561 2852 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 0 496 2852 527
rect 14 459 2838 468
rect 14 428 1047 459
rect 1035 425 1047 428
rect 1081 428 1219 459
rect 1081 425 1093 428
rect 1035 416 1093 425
rect 1207 425 1219 428
rect 1253 428 1390 459
rect 1253 425 1265 428
rect 1207 416 1265 425
rect 1378 425 1390 428
rect 1424 428 1560 459
rect 1424 425 1436 428
rect 1378 416 1436 425
rect 1548 425 1560 428
rect 1594 428 1736 459
rect 1594 425 1606 428
rect 1548 416 1606 425
rect 1724 425 1736 428
rect 1770 428 1908 459
rect 1770 425 1782 428
rect 1724 416 1782 425
rect 1896 425 1908 428
rect 1942 428 2079 459
rect 1942 425 1954 428
rect 1896 416 1954 425
rect 2067 425 2079 428
rect 2113 428 2251 459
rect 2113 425 2125 428
rect 2067 416 2125 425
rect 2239 425 2251 428
rect 2285 428 2422 459
rect 2285 425 2297 428
rect 2239 416 2297 425
rect 2410 425 2422 428
rect 2456 428 2592 459
rect 2456 425 2468 428
rect 2410 416 2468 425
rect 2580 425 2592 428
rect 2626 428 2768 459
rect 2626 425 2638 428
rect 2580 416 2638 425
rect 2756 425 2768 428
rect 2802 428 2838 459
rect 2802 425 2814 428
rect 2756 416 2814 425
rect 493 187 623 193
rect 493 153 505 187
rect 539 153 577 187
rect 611 184 623 187
rect 1030 187 1088 193
rect 1030 184 1042 187
rect 611 156 1042 184
rect 611 153 623 156
rect 493 147 623 153
rect 1030 153 1042 156
rect 1076 153 1088 187
rect 1030 147 1088 153
rect 0 17 2852 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
rect 0 -48 2852 -17
<< labels >>
flabel locali s 2697 153 2731 187 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 2605 153 2639 187 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 2605 221 2639 255 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 2697 221 2731 255 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 2697 289 2731 323 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 2605 289 2639 323 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 50 221 84 255 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 856 221 890 255 0 FreeSans 200 180 0 0 SLEEP
port 2 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel pwell s 1041 -17 1075 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel pwell s 1058 0 1058 0 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 1041 527 1075 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 1058 544 1058 544 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 26 428 75 468 0 FreeSans 200 0 0 0 KAPWR
port 3 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 lpflow_isobufsrckapwr_16
rlabel locali s 2242 381 2291 493 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 2414 381 2463 493 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 2586 381 2637 493 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 2763 378 2817 493 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1031 299 1097 493 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1203 299 1269 493 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1375 299 1441 493 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1554 381 1606 493 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1726 381 1778 493 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1898 381 1950 493 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 2756 416 2814 428 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 2580 416 2638 428 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 2410 416 2468 428 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 2239 416 2297 428 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 2067 416 2125 428 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1896 416 1954 428 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1724 416 1782 428 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1548 416 1606 428 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1378 416 1436 428 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1207 416 1265 428 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1035 416 1093 428 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 14 428 2838 468 1 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 -48 2852 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2852 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2852 544
string GDS_END 2444532
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2422616
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 71.300 0.000 
<< end >>
