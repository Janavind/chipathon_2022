magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -36 538 404 1177
<< locali >>
rect 0 1103 368 1137
rect 64 508 98 574
rect 179 524 213 558
rect 0 -17 368 17
use pinv  pinv_0
timestamp 1666464484
transform 1 0 0 0 1 0
box -36 -17 404 1177
<< labels >>
rlabel locali s 196 541 196 541 4 Z
port 2 nsew
rlabel locali s 81 541 81 541 4 A
port 1 nsew
rlabel locali s 184 1120 184 1120 4 vdd
port 3 nsew
rlabel locali s 184 0 184 0 4 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 368 1120
string GDS_END 32706
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 31870
<< end >>
