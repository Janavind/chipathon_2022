magic
tech sky130B
magscale 1 2
timestamp 1666199351
use sky130_fd_pr__dfl1sd__example_55959141808123  sky130_fd_pr__dfl1sd__example_55959141808123_0
timestamp 1666199351
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808123  sky130_fd_pr__dfl1sd__example_55959141808123_1
timestamp 1666199351
transform 1 0 400 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 48942506
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48941456
<< end >>
