magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 1 21 1339 203
rect 29 -17 63 21
<< scnmos >>
rect 110 47 140 177
rect 216 47 246 177
rect 302 47 332 177
rect 388 47 418 177
rect 474 47 504 177
rect 628 47 658 177
rect 714 47 744 177
rect 800 47 830 177
rect 886 47 916 177
rect 972 47 1002 177
rect 1058 47 1088 177
rect 1144 47 1174 177
rect 1230 47 1260 177
<< scpmoshvt >>
rect 86 297 116 497
rect 276 297 306 497
rect 362 297 392 497
rect 448 297 478 497
rect 534 297 564 497
rect 626 297 656 497
rect 714 297 744 497
rect 800 297 830 497
rect 886 297 916 497
rect 972 297 1002 497
rect 1058 297 1088 497
rect 1144 297 1174 497
rect 1230 297 1260 497
<< ndiff >>
rect 27 157 110 177
rect 27 123 39 157
rect 73 123 110 157
rect 27 89 110 123
rect 27 55 39 89
rect 73 55 110 89
rect 27 47 110 55
rect 140 89 216 177
rect 140 55 163 89
rect 197 55 216 89
rect 140 47 216 55
rect 246 124 302 177
rect 246 90 257 124
rect 291 90 302 124
rect 246 47 302 90
rect 332 89 388 177
rect 332 55 343 89
rect 377 55 388 89
rect 332 47 388 55
rect 418 169 474 177
rect 418 135 429 169
rect 463 135 474 169
rect 418 101 474 135
rect 418 67 429 101
rect 463 67 474 101
rect 418 47 474 67
rect 504 89 628 177
rect 504 55 515 89
rect 549 55 583 89
rect 617 55 628 89
rect 504 47 628 55
rect 658 101 714 177
rect 658 67 669 101
rect 703 67 714 101
rect 658 47 714 67
rect 744 169 800 177
rect 744 135 755 169
rect 789 135 800 169
rect 744 47 800 135
rect 830 101 886 177
rect 830 67 841 101
rect 875 67 886 101
rect 830 47 886 67
rect 916 169 972 177
rect 916 135 927 169
rect 961 135 972 169
rect 916 47 972 135
rect 1002 157 1058 177
rect 1002 123 1013 157
rect 1047 123 1058 157
rect 1002 89 1058 123
rect 1002 55 1013 89
rect 1047 55 1058 89
rect 1002 47 1058 55
rect 1088 97 1144 177
rect 1088 63 1099 97
rect 1133 63 1144 97
rect 1088 47 1144 63
rect 1174 164 1230 177
rect 1174 130 1185 164
rect 1219 130 1230 164
rect 1174 96 1230 130
rect 1174 62 1185 96
rect 1219 62 1230 96
rect 1174 47 1230 62
rect 1260 161 1313 177
rect 1260 127 1271 161
rect 1305 127 1313 161
rect 1260 93 1313 127
rect 1260 59 1271 93
rect 1305 59 1313 93
rect 1260 47 1313 59
<< pdiff >>
rect 33 485 86 497
rect 33 451 41 485
rect 75 451 86 485
rect 33 417 86 451
rect 33 383 41 417
rect 75 383 86 417
rect 33 297 86 383
rect 116 485 169 497
rect 116 451 127 485
rect 161 451 169 485
rect 116 297 169 451
rect 223 477 276 497
rect 223 443 232 477
rect 266 443 276 477
rect 223 409 276 443
rect 223 375 232 409
rect 266 375 276 409
rect 223 297 276 375
rect 306 387 362 497
rect 306 353 317 387
rect 351 353 362 387
rect 306 297 362 353
rect 392 489 448 497
rect 392 455 403 489
rect 437 455 448 489
rect 392 297 448 455
rect 478 395 534 497
rect 478 361 489 395
rect 523 361 534 395
rect 478 297 534 361
rect 564 477 626 497
rect 564 443 581 477
rect 615 443 626 477
rect 564 297 626 443
rect 656 489 714 497
rect 656 455 669 489
rect 703 455 714 489
rect 656 297 714 455
rect 744 415 800 497
rect 744 381 755 415
rect 789 381 800 415
rect 744 297 800 381
rect 830 489 886 497
rect 830 455 841 489
rect 875 455 886 489
rect 830 297 886 455
rect 916 477 972 497
rect 916 443 927 477
rect 961 443 972 477
rect 916 409 972 443
rect 916 375 927 409
rect 961 375 972 409
rect 916 297 972 375
rect 1002 489 1058 497
rect 1002 455 1013 489
rect 1047 455 1058 489
rect 1002 297 1058 455
rect 1088 477 1144 497
rect 1088 443 1099 477
rect 1133 443 1144 477
rect 1088 297 1144 443
rect 1174 489 1230 497
rect 1174 455 1185 489
rect 1219 455 1230 489
rect 1174 297 1230 455
rect 1260 477 1313 497
rect 1260 443 1271 477
rect 1305 443 1313 477
rect 1260 409 1313 443
rect 1260 375 1271 409
rect 1305 375 1313 409
rect 1260 297 1313 375
<< ndiffc >>
rect 39 123 73 157
rect 39 55 73 89
rect 163 55 197 89
rect 257 90 291 124
rect 343 55 377 89
rect 429 135 463 169
rect 429 67 463 101
rect 515 55 549 89
rect 583 55 617 89
rect 669 67 703 101
rect 755 135 789 169
rect 841 67 875 101
rect 927 135 961 169
rect 1013 123 1047 157
rect 1013 55 1047 89
rect 1099 63 1133 97
rect 1185 130 1219 164
rect 1185 62 1219 96
rect 1271 127 1305 161
rect 1271 59 1305 93
<< pdiffc >>
rect 41 451 75 485
rect 41 383 75 417
rect 127 451 161 485
rect 232 443 266 477
rect 232 375 266 409
rect 317 353 351 387
rect 403 455 437 489
rect 489 361 523 395
rect 581 443 615 477
rect 669 455 703 489
rect 755 381 789 415
rect 841 455 875 489
rect 927 443 961 477
rect 927 375 961 409
rect 1013 455 1047 489
rect 1099 443 1133 477
rect 1185 455 1219 489
rect 1271 443 1305 477
rect 1271 375 1305 409
<< poly >>
rect 86 497 116 523
rect 276 497 306 523
rect 362 497 392 523
rect 448 497 478 523
rect 534 497 564 523
rect 626 497 656 523
rect 714 497 744 523
rect 800 497 830 523
rect 886 497 916 523
rect 972 497 1002 523
rect 1058 497 1088 523
rect 1144 497 1174 523
rect 1230 497 1260 523
rect 86 265 116 297
rect 276 265 306 297
rect 362 265 392 297
rect 448 265 478 297
rect 534 265 564 297
rect 626 265 656 297
rect 86 249 140 265
rect 86 215 96 249
rect 130 215 140 249
rect 86 199 140 215
rect 110 177 140 199
rect 216 249 564 265
rect 216 215 226 249
rect 260 215 294 249
rect 328 215 362 249
rect 396 215 430 249
rect 464 215 564 249
rect 216 199 564 215
rect 606 249 672 265
rect 606 215 622 249
rect 656 215 672 249
rect 606 199 672 215
rect 714 259 744 297
rect 800 259 830 297
rect 886 259 916 297
rect 972 259 1002 297
rect 714 249 1002 259
rect 714 215 738 249
rect 772 215 806 249
rect 840 215 874 249
rect 908 215 942 249
rect 976 215 1002 249
rect 216 177 246 199
rect 302 177 332 199
rect 388 177 418 199
rect 474 177 504 199
rect 628 177 658 199
rect 714 198 1002 215
rect 714 177 744 198
rect 800 177 830 198
rect 886 177 916 198
rect 972 177 1002 198
rect 1058 265 1088 297
rect 1144 265 1174 297
rect 1230 265 1260 297
rect 1058 249 1284 265
rect 1058 215 1104 249
rect 1138 215 1172 249
rect 1206 215 1240 249
rect 1274 215 1284 249
rect 1058 199 1284 215
rect 1058 177 1088 199
rect 1144 177 1174 199
rect 1230 177 1260 199
rect 110 21 140 47
rect 216 21 246 47
rect 302 21 332 47
rect 388 21 418 47
rect 474 21 504 47
rect 628 21 658 47
rect 714 21 744 47
rect 800 21 830 47
rect 886 21 916 47
rect 972 21 1002 47
rect 1058 21 1088 47
rect 1144 21 1174 47
rect 1230 21 1260 47
<< polycont >>
rect 96 215 130 249
rect 226 215 260 249
rect 294 215 328 249
rect 362 215 396 249
rect 430 215 464 249
rect 622 215 656 249
rect 738 215 772 249
rect 806 215 840 249
rect 874 215 908 249
rect 942 215 976 249
rect 1104 215 1138 249
rect 1172 215 1206 249
rect 1240 215 1274 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 25 485 91 493
rect 25 451 41 485
rect 75 451 91 485
rect 25 417 91 451
rect 125 485 177 527
rect 125 451 127 485
rect 161 451 177 485
rect 125 435 177 451
rect 232 489 619 493
rect 232 477 403 489
rect 266 455 403 477
rect 437 477 619 489
rect 437 455 581 477
rect 266 443 581 455
rect 615 443 619 477
rect 653 489 719 527
rect 653 455 669 489
rect 703 455 719 489
rect 825 489 891 527
rect 825 455 841 489
rect 875 455 891 489
rect 925 477 963 493
rect 25 383 41 417
rect 75 401 91 417
rect 232 409 271 443
rect 387 441 619 443
rect 75 383 198 401
rect 25 357 198 383
rect 266 375 271 409
rect 579 421 619 441
rect 925 443 927 477
rect 961 443 963 477
rect 997 489 1063 527
rect 997 455 1013 489
rect 1047 455 1063 489
rect 1097 477 1133 493
rect 925 421 963 443
rect 1097 443 1099 477
rect 1169 489 1235 527
rect 1169 455 1185 489
rect 1219 455 1235 489
rect 1269 477 1321 493
rect 1097 421 1133 443
rect 1269 443 1271 477
rect 1305 443 1321 477
rect 1269 421 1321 443
rect 579 415 1321 421
rect 232 359 271 375
rect 312 395 545 407
rect 312 387 489 395
rect 29 249 130 323
rect 29 215 96 249
rect 96 199 130 215
rect 164 269 198 357
rect 312 353 317 387
rect 351 361 489 387
rect 523 361 545 395
rect 579 381 755 415
rect 789 409 1321 415
rect 789 381 927 409
rect 579 375 927 381
rect 961 375 1271 409
rect 1305 375 1321 409
rect 351 353 545 361
rect 312 341 545 353
rect 312 317 572 341
rect 164 249 480 269
rect 164 215 226 249
rect 260 215 294 249
rect 328 215 362 249
rect 396 215 430 249
rect 464 215 480 249
rect 164 207 480 215
rect 164 159 221 207
rect 514 179 572 317
rect 606 296 1290 341
rect 606 249 675 296
rect 606 215 622 249
rect 656 215 675 249
rect 606 213 675 215
rect 709 249 994 262
rect 709 215 738 249
rect 772 215 806 249
rect 840 215 874 249
rect 908 215 942 249
rect 976 215 994 249
rect 1041 249 1290 296
rect 1041 215 1104 249
rect 1138 215 1172 249
rect 1206 215 1240 249
rect 1274 215 1290 249
rect 709 213 994 215
rect 514 173 977 179
rect 18 157 221 159
rect 18 123 39 157
rect 73 123 221 157
rect 255 169 977 173
rect 255 135 429 169
rect 463 139 755 169
rect 463 135 465 139
rect 651 135 755 139
rect 789 135 927 169
rect 961 135 977 169
rect 1011 164 1235 181
rect 1011 157 1185 164
rect 255 124 465 135
rect 18 89 89 123
rect 255 90 257 124
rect 291 123 465 124
rect 291 90 293 123
rect 18 55 39 89
rect 73 55 89 89
rect 18 51 89 55
rect 144 55 163 89
rect 197 55 221 89
rect 255 74 293 90
rect 427 101 465 123
rect 1011 123 1013 157
rect 1047 147 1185 157
rect 1047 123 1063 147
rect 144 17 221 55
rect 327 55 343 89
rect 377 55 393 89
rect 327 17 393 55
rect 427 67 429 101
rect 463 67 465 101
rect 427 51 465 67
rect 499 89 617 105
rect 1011 101 1063 123
rect 1169 130 1185 147
rect 1219 130 1235 164
rect 499 55 515 89
rect 549 55 583 89
rect 499 17 617 55
rect 653 67 669 101
rect 703 67 841 101
rect 875 89 1063 101
rect 875 67 1013 89
rect 653 55 1013 67
rect 1047 55 1063 89
rect 653 51 1063 55
rect 1097 97 1135 113
rect 1097 63 1099 97
rect 1133 63 1135 97
rect 1097 17 1135 63
rect 1169 96 1235 130
rect 1169 62 1185 96
rect 1219 62 1235 96
rect 1169 51 1235 62
rect 1269 161 1321 177
rect 1269 127 1271 161
rect 1305 127 1321 161
rect 1269 93 1321 127
rect 1269 59 1271 93
rect 1305 59 1321 93
rect 1269 17 1321 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel locali s 489 357 523 391 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 949 221 983 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 1225 289 1259 323 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a21boi_4
rlabel metal1 s 0 -48 1380 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1380 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1380 544
string GDS_END 4025984
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4016552
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 34.500 0.000 
<< end >>
